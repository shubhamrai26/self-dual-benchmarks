module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 ;
  assign n129 = ( x17 & ~x57 ) | ( x17 & x115 ) | ( ~x57 & x115 ) ;
  assign n130 = x22 & x116 ;
  assign n131 = n130 ^ x110 ^ 1'b0 ;
  assign n132 = x115 ^ x50 ^ 1'b0 ;
  assign n133 = x96 & n132 ;
  assign n134 = n133 ^ x75 ^ x34 ;
  assign n135 = x19 & x41 ;
  assign n136 = n135 ^ x58 ^ 1'b0 ;
  assign n137 = x41 & x94 ;
  assign n138 = ~x123 & n137 ;
  assign n139 = ( x13 & x68 ) | ( x13 & ~x92 ) | ( x68 & ~x92 ) ;
  assign n140 = ( x31 & x93 ) | ( x31 & ~x99 ) | ( x93 & ~x99 ) ;
  assign n141 = n140 ^ x94 ^ 1'b0 ;
  assign n142 = x80 & n141 ;
  assign n143 = n142 ^ x110 ^ x16 ;
  assign n144 = x36 & n140 ;
  assign n145 = ~x24 & n144 ;
  assign n146 = ( x43 & ~x92 ) | ( x43 & n145 ) | ( ~x92 & n145 ) ;
  assign n147 = x114 ^ x6 ^ 1'b0 ;
  assign n148 = x8 & n147 ;
  assign n151 = x71 & x122 ;
  assign n152 = ~x16 & n151 ;
  assign n149 = x40 & x75 ;
  assign n150 = n149 ^ x76 ^ 1'b0 ;
  assign n153 = n152 ^ n150 ^ x86 ;
  assign n154 = x93 ^ x64 ^ x45 ;
  assign n155 = x122 & n140 ;
  assign n156 = ~n154 & n155 ;
  assign n157 = n156 ^ x40 ^ 1'b0 ;
  assign n159 = x104 ^ x60 ^ 1'b0 ;
  assign n160 = x85 & n159 ;
  assign n158 = ( x36 & x63 ) | ( x36 & ~x104 ) | ( x63 & ~x104 ) ;
  assign n161 = n160 ^ n158 ^ x55 ;
  assign n162 = n161 ^ n142 ^ x65 ;
  assign n163 = ~x49 & x112 ;
  assign n164 = x106 ^ x103 ^ x76 ;
  assign n165 = ( x15 & ~x72 ) | ( x15 & n164 ) | ( ~x72 & n164 ) ;
  assign n166 = x12 & ~n165 ;
  assign n167 = n166 ^ x111 ^ 1'b0 ;
  assign n168 = ( x87 & x96 ) | ( x87 & ~n140 ) | ( x96 & ~n140 ) ;
  assign n169 = ( ~x16 & x95 ) | ( ~x16 & x108 ) | ( x95 & x108 ) ;
  assign n170 = ( x71 & x76 ) | ( x71 & ~n169 ) | ( x76 & ~n169 ) ;
  assign n171 = x122 & n133 ;
  assign n172 = n171 ^ x35 ^ 1'b0 ;
  assign n173 = ( x2 & n136 ) | ( x2 & n172 ) | ( n136 & n172 ) ;
  assign n174 = x25 & x43 ;
  assign n175 = n174 ^ n152 ^ 1'b0 ;
  assign n176 = x1 & x25 ;
  assign n177 = ~x103 & n176 ;
  assign n178 = ( ~n136 & n175 ) | ( ~n136 & n177 ) | ( n175 & n177 ) ;
  assign n179 = x0 & n178 ;
  assign n180 = n173 & n179 ;
  assign n181 = ( x0 & ~x59 ) | ( x0 & x83 ) | ( ~x59 & x83 ) ;
  assign n182 = x70 ^ x16 ^ 1'b0 ;
  assign n183 = n169 ^ x54 ^ 1'b0 ;
  assign n184 = x70 & n183 ;
  assign n185 = x127 & n140 ;
  assign n186 = n185 ^ x65 ^ 1'b0 ;
  assign n187 = x57 | n186 ;
  assign n188 = x86 & n187 ;
  assign n189 = ~x90 & n188 ;
  assign n190 = ( x52 & n153 ) | ( x52 & ~n178 ) | ( n153 & ~n178 ) ;
  assign n191 = x80 ^ x34 ^ 1'b0 ;
  assign n192 = n190 ^ x82 ^ 1'b0 ;
  assign n193 = x21 & ~n192 ;
  assign n194 = x47 ^ x28 ^ 1'b0 ;
  assign n195 = x62 & n194 ;
  assign n196 = n195 ^ x86 ^ x3 ;
  assign n197 = ( x39 & x58 ) | ( x39 & ~n187 ) | ( x58 & ~n187 ) ;
  assign n198 = x121 ^ x87 ^ 1'b0 ;
  assign n199 = x62 & n198 ;
  assign n200 = x72 & x108 ;
  assign n201 = ~x41 & n200 ;
  assign n202 = x62 & ~n201 ;
  assign n203 = ~n194 & n202 ;
  assign n204 = n190 | n203 ;
  assign n205 = x124 | n204 ;
  assign n206 = x120 & n205 ;
  assign n207 = ( ~x8 & x52 ) | ( ~x8 & x126 ) | ( x52 & x126 ) ;
  assign n208 = n207 ^ x21 ^ 1'b0 ;
  assign n209 = x33 & n208 ;
  assign n210 = n165 ^ n148 ^ x50 ;
  assign n211 = n210 ^ n206 ^ x118 ;
  assign n212 = ( x28 & ~x29 ) | ( x28 & x124 ) | ( ~x29 & x124 ) ;
  assign n213 = x61 & x65 ;
  assign n214 = ~x66 & n213 ;
  assign n215 = x63 & ~n214 ;
  assign n216 = ~n212 & n215 ;
  assign n218 = n165 ^ x93 ^ x33 ;
  assign n217 = x1 & x92 ;
  assign n219 = n218 ^ n217 ^ 1'b0 ;
  assign n220 = ( ~x7 & x104 ) | ( ~x7 & n219 ) | ( x104 & n219 ) ;
  assign n221 = ( x124 & n194 ) | ( x124 & n214 ) | ( n194 & n214 ) ;
  assign n222 = n221 ^ n205 ^ 1'b0 ;
  assign n223 = ( ~x31 & x65 ) | ( ~x31 & n219 ) | ( x65 & n219 ) ;
  assign n224 = x100 ^ x68 ^ 1'b0 ;
  assign n225 = x18 & n224 ;
  assign n226 = x88 & n225 ;
  assign n227 = ~x90 & n226 ;
  assign n228 = x26 & x36 ;
  assign n229 = n228 ^ n206 ^ 1'b0 ;
  assign n230 = x76 & x126 ;
  assign n231 = ~x86 & n230 ;
  assign n232 = n231 ^ x56 ^ x48 ;
  assign n233 = ( ~x51 & x72 ) | ( ~x51 & x120 ) | ( x72 & x120 ) ;
  assign n234 = x110 & ~n233 ;
  assign n235 = x110 ^ x64 ^ 1'b0 ;
  assign n236 = n148 & n235 ;
  assign n237 = x101 & n236 ;
  assign n238 = ~x42 & n237 ;
  assign n241 = n134 ^ x105 ^ 1'b0 ;
  assign n242 = x67 & ~n241 ;
  assign n239 = x31 & ~n164 ;
  assign n240 = ~x108 & n239 ;
  assign n243 = n242 ^ n240 ^ x61 ;
  assign n244 = n187 ^ n148 ^ 1'b0 ;
  assign n245 = x118 & n244 ;
  assign n246 = n245 ^ x49 ^ 1'b0 ;
  assign n247 = n211 ^ n191 ^ x50 ;
  assign n248 = ( ~x91 & n197 ) | ( ~x91 & n247 ) | ( n197 & n247 ) ;
  assign n249 = ( ~x120 & x127 ) | ( ~x120 & n248 ) | ( x127 & n248 ) ;
  assign n250 = n249 ^ x103 ^ 1'b0 ;
  assign n257 = x127 ^ x42 ^ x31 ;
  assign n256 = ( x4 & x36 ) | ( x4 & ~x55 ) | ( x36 & ~x55 ) ;
  assign n258 = n257 ^ n256 ^ x11 ;
  assign n259 = ~n209 & n258 ;
  assign n251 = n184 ^ x124 ^ 1'b0 ;
  assign n252 = n143 ^ n133 ^ x81 ;
  assign n253 = n252 ^ x40 ^ 1'b0 ;
  assign n254 = n251 & n253 ;
  assign n255 = x86 & n254 ;
  assign n260 = n259 ^ n255 ^ 1'b0 ;
  assign n263 = x23 & x84 ;
  assign n264 = ~x58 & n263 ;
  assign n261 = n214 ^ x112 ^ x90 ;
  assign n262 = x9 & n261 ;
  assign n265 = n264 ^ n262 ^ 1'b0 ;
  assign n266 = x17 & x113 ;
  assign n267 = x67 & ~n266 ;
  assign n268 = x97 & n160 ;
  assign n269 = n268 ^ x12 ^ 1'b0 ;
  assign n270 = n242 & ~n269 ;
  assign n271 = ~n196 & n270 ;
  assign n272 = x120 & n271 ;
  assign n273 = x68 & ~n173 ;
  assign n274 = ~x123 & n273 ;
  assign n275 = n222 ^ x93 ^ 1'b0 ;
  assign n276 = ~n274 & n275 ;
  assign n277 = n276 ^ x55 ^ 1'b0 ;
  assign n278 = x75 & n277 ;
  assign n279 = ~x77 & n160 ;
  assign n283 = x12 & ~n214 ;
  assign n284 = n283 ^ x74 ^ 1'b0 ;
  assign n280 = x37 & ~n231 ;
  assign n281 = n280 ^ x2 ^ 1'b0 ;
  assign n282 = n170 & ~n281 ;
  assign n285 = n284 ^ n282 ^ 1'b0 ;
  assign n286 = ( x44 & ~x127 ) | ( x44 & n285 ) | ( ~x127 & n285 ) ;
  assign n287 = x42 & n142 ;
  assign n288 = n287 ^ n225 ^ 1'b0 ;
  assign n289 = ( ~x109 & n158 ) | ( ~x109 & n169 ) | ( n158 & n169 ) ;
  assign n290 = n173 ^ x88 ^ x47 ;
  assign n291 = x58 & x83 ;
  assign n292 = n291 ^ n281 ^ 1'b0 ;
  assign n293 = n292 ^ n234 ^ 1'b0 ;
  assign n294 = x71 & x111 ;
  assign n295 = n294 ^ x81 ^ 1'b0 ;
  assign n296 = ( n220 & n274 ) | ( n220 & ~n295 ) | ( n274 & ~n295 ) ;
  assign n297 = x2 & n133 ;
  assign n298 = ~x97 & n297 ;
  assign n299 = n177 & ~n298 ;
  assign n300 = n299 ^ x0 ^ 1'b0 ;
  assign n301 = x69 ^ x50 ^ 1'b0 ;
  assign n302 = x61 & n301 ;
  assign n303 = n302 ^ n259 ^ x65 ;
  assign n304 = n214 ^ x106 ^ x103 ;
  assign n305 = n304 ^ n222 ^ 1'b0 ;
  assign n306 = x37 & x51 ;
  assign n307 = n306 ^ n173 ^ 1'b0 ;
  assign n308 = n307 ^ x57 ^ 1'b0 ;
  assign n309 = n308 ^ n276 ^ 1'b0 ;
  assign n310 = n139 ^ n131 ^ x2 ;
  assign n311 = n219 ^ n180 ^ 1'b0 ;
  assign n312 = x9 & n311 ;
  assign n317 = x98 ^ x14 ^ 1'b0 ;
  assign n318 = ~n269 & n317 ;
  assign n313 = n138 ^ x114 ^ x36 ;
  assign n314 = ( x78 & n134 ) | ( x78 & n158 ) | ( n134 & n158 ) ;
  assign n315 = n314 ^ x72 ^ 1'b0 ;
  assign n316 = n313 & n315 ;
  assign n319 = n318 ^ n316 ^ n261 ;
  assign n320 = n206 & ~n267 ;
  assign n323 = n199 ^ x115 ^ x56 ;
  assign n321 = x64 & x73 ;
  assign n322 = n321 ^ x80 ^ 1'b0 ;
  assign n324 = n323 ^ n322 ^ n172 ;
  assign n325 = n324 ^ n251 ^ 1'b0 ;
  assign n326 = x123 ^ x72 ^ 1'b0 ;
  assign n327 = x94 & n326 ;
  assign n328 = x119 & n327 ;
  assign n329 = x117 ^ x10 ^ 1'b0 ;
  assign n330 = x25 & n329 ;
  assign n331 = ( n145 & n168 ) | ( n145 & ~n330 ) | ( n168 & ~n330 ) ;
  assign n332 = x45 ^ x7 ^ 1'b0 ;
  assign n333 = n302 ^ x99 ^ 1'b0 ;
  assign n334 = x120 & n333 ;
  assign n335 = n324 ^ n285 ^ n180 ;
  assign n340 = ( ~x60 & x105 ) | ( ~x60 & n257 ) | ( x105 & n257 ) ;
  assign n336 = x45 & ~n152 ;
  assign n337 = n336 ^ n269 ^ 1'b0 ;
  assign n338 = x47 & n337 ;
  assign n339 = n338 ^ x10 ^ 1'b0 ;
  assign n341 = n340 ^ n339 ^ n178 ;
  assign n352 = x110 & n209 ;
  assign n353 = ~n258 & n352 ;
  assign n351 = n134 ^ x106 ^ 1'b0 ;
  assign n343 = n158 ^ x108 ^ 1'b0 ;
  assign n342 = ~n186 & n256 ;
  assign n344 = n343 ^ n342 ^ 1'b0 ;
  assign n345 = n343 ^ x30 ^ 1'b0 ;
  assign n346 = n278 & n345 ;
  assign n347 = n346 ^ x48 ^ 1'b0 ;
  assign n348 = n257 | n347 ;
  assign n349 = n348 ^ x103 ^ 1'b0 ;
  assign n350 = n344 & n349 ;
  assign n354 = n353 ^ n351 ^ n350 ;
  assign n355 = n209 ^ n129 ^ x82 ;
  assign n356 = x12 ^ x2 ^ 1'b0 ;
  assign n357 = n356 ^ n175 ^ x16 ;
  assign n358 = ( n284 & ~n355 ) | ( n284 & n357 ) | ( ~n355 & n357 ) ;
  assign n359 = x110 & ~n357 ;
  assign n360 = ~x46 & n359 ;
  assign n361 = n142 ^ x26 ^ x4 ;
  assign n362 = x24 & n361 ;
  assign n363 = n271 | n362 ;
  assign n365 = x96 ^ x65 ^ x3 ;
  assign n364 = x44 & ~n351 ;
  assign n366 = n365 ^ n364 ^ 1'b0 ;
  assign n367 = n324 ^ n172 ^ x113 ;
  assign n371 = x33 & x105 ;
  assign n372 = n371 ^ x66 ^ 1'b0 ;
  assign n376 = x102 ^ x90 ^ 1'b0 ;
  assign n377 = ~n372 & n376 ;
  assign n378 = n377 ^ x89 ^ 1'b0 ;
  assign n368 = x67 ^ x35 ^ 1'b0 ;
  assign n369 = n368 ^ n203 ^ 1'b0 ;
  assign n370 = n164 | n369 ;
  assign n373 = n214 | n372 ;
  assign n374 = n370 & ~n373 ;
  assign n375 = n320 & ~n374 ;
  assign n379 = n378 ^ n375 ^ 1'b0 ;
  assign n380 = n138 | n231 ;
  assign n381 = ( x10 & ~n146 ) | ( x10 & n380 ) | ( ~n146 & n380 ) ;
  assign n382 = ( x93 & ~n152 ) | ( x93 & n203 ) | ( ~n152 & n203 ) ;
  assign n383 = n216 ^ x104 ^ 1'b0 ;
  assign n384 = ( ~n290 & n382 ) | ( ~n290 & n383 ) | ( n382 & n383 ) ;
  assign n385 = x77 & ~n370 ;
  assign n386 = ~n155 & n385 ;
  assign n390 = ( ~x111 & n142 ) | ( ~x111 & n313 ) | ( n142 & n313 ) ;
  assign n387 = x121 & ~n134 ;
  assign n388 = n387 ^ n247 ^ 1'b0 ;
  assign n389 = x42 & n388 ;
  assign n391 = n390 ^ n389 ^ 1'b0 ;
  assign n392 = x97 & n246 ;
  assign n393 = ~x118 & n392 ;
  assign n400 = x115 ^ x7 ^ 1'b0 ;
  assign n401 = x73 & n400 ;
  assign n394 = x23 & x88 ;
  assign n395 = ~x76 & n394 ;
  assign n396 = n154 | n370 ;
  assign n397 = n395 & ~n396 ;
  assign n398 = ( ~x22 & n256 ) | ( ~x22 & n397 ) | ( n256 & n397 ) ;
  assign n399 = n398 ^ x107 ^ x35 ;
  assign n402 = n401 ^ n399 ^ 1'b0 ;
  assign n403 = n153 ^ x91 ^ 1'b0 ;
  assign n404 = ( x115 & n157 ) | ( x115 & n403 ) | ( n157 & n403 ) ;
  assign n405 = x48 & x80 ;
  assign n406 = ~x40 & n405 ;
  assign n407 = n303 ^ n157 ^ 1'b0 ;
  assign n408 = x103 & n407 ;
  assign n409 = x86 & x116 ;
  assign n410 = ~n408 & n409 ;
  assign n411 = n175 ^ n139 ^ x0 ;
  assign n412 = x127 ^ x96 ^ x43 ;
  assign n413 = n412 ^ n195 ^ x99 ;
  assign n414 = n411 & n413 ;
  assign n415 = n414 ^ n148 ^ 1'b0 ;
  assign n416 = x84 ^ x62 ^ 1'b0 ;
  assign n417 = n186 | n295 ;
  assign n418 = n417 ^ x19 ^ 1'b0 ;
  assign n419 = ( n189 & n378 ) | ( n189 & n418 ) | ( n378 & n418 ) ;
  assign n420 = ( x36 & x55 ) | ( x36 & ~x122 ) | ( x55 & ~x122 ) ;
  assign n421 = ( ~x25 & x38 ) | ( ~x25 & n264 ) | ( x38 & n264 ) ;
  assign n422 = n136 ^ x49 ^ x5 ;
  assign n423 = ~x121 & n422 ;
  assign n424 = ( n420 & n421 ) | ( n420 & ~n423 ) | ( n421 & ~n423 ) ;
  assign n425 = n187 ^ n181 ^ x62 ;
  assign n426 = x6 & x64 ;
  assign n427 = ~x74 & n426 ;
  assign n428 = n343 & ~n427 ;
  assign n429 = n190 & n428 ;
  assign n430 = x113 | n429 ;
  assign n431 = n175 & n430 ;
  assign n432 = ( ~x46 & x49 ) | ( ~x46 & x73 ) | ( x49 & x73 ) ;
  assign n433 = n290 & ~n331 ;
  assign n434 = x113 ^ x31 ^ 1'b0 ;
  assign n435 = n209 ^ x84 ^ 1'b0 ;
  assign n436 = x95 & n435 ;
  assign n437 = x18 & x86 ;
  assign n438 = n437 ^ x7 ^ 1'b0 ;
  assign n439 = n438 ^ n160 ^ 1'b0 ;
  assign n440 = n295 | n439 ;
  assign n441 = n440 ^ n337 ^ n153 ;
  assign n442 = ( ~n415 & n436 ) | ( ~n415 & n441 ) | ( n436 & n441 ) ;
  assign n443 = n390 ^ n383 ^ n218 ;
  assign n444 = ( ~x104 & n432 ) | ( ~x104 & n443 ) | ( n432 & n443 ) ;
  assign n445 = ( x22 & ~x80 ) | ( x22 & n343 ) | ( ~x80 & n343 ) ;
  assign n446 = n445 ^ x31 ^ 1'b0 ;
  assign n447 = n212 & n446 ;
  assign n448 = n447 ^ n216 ^ x34 ;
  assign n449 = n340 ^ x84 ^ 1'b0 ;
  assign n450 = n190 ^ x57 ^ 1'b0 ;
  assign n451 = n449 | n450 ;
  assign n452 = n212 ^ x61 ^ 1'b0 ;
  assign n453 = n452 ^ n261 ^ 1'b0 ;
  assign n455 = x108 & ~n150 ;
  assign n456 = ~x60 & n455 ;
  assign n457 = x107 & ~n201 ;
  assign n458 = n456 & n457 ;
  assign n454 = n181 & ~n231 ;
  assign n459 = n458 ^ n454 ^ 1'b0 ;
  assign n460 = x95 & n236 ;
  assign n461 = n460 ^ x106 ^ 1'b0 ;
  assign n462 = ( x72 & ~n459 ) | ( x72 & n461 ) | ( ~n459 & n461 ) ;
  assign n463 = n456 ^ n377 ^ x57 ;
  assign n469 = x80 | n257 ;
  assign n464 = x15 & ~n134 ;
  assign n465 = ~x91 & n464 ;
  assign n466 = x100 ^ x53 ^ 1'b0 ;
  assign n467 = x26 & n466 ;
  assign n468 = ~n465 & n467 ;
  assign n470 = n469 ^ n468 ^ 1'b0 ;
  assign n471 = x122 | n470 ;
  assign n472 = x49 & ~n344 ;
  assign n473 = n472 ^ x24 ^ 1'b0 ;
  assign n477 = ~x2 & x73 ;
  assign n474 = n269 ^ n143 ^ x10 ;
  assign n475 = n474 ^ n214 ^ x20 ;
  assign n476 = n186 | n475 ;
  assign n478 = n477 ^ n476 ^ 1'b0 ;
  assign n479 = ~n325 & n478 ;
  assign n480 = n473 & n479 ;
  assign n481 = ~n164 & n304 ;
  assign n482 = ~n431 & n481 ;
  assign n485 = x123 ^ x60 ^ 1'b0 ;
  assign n483 = x31 & x44 ;
  assign n484 = n483 ^ x84 ^ 1'b0 ;
  assign n486 = n485 ^ n484 ^ 1'b0 ;
  assign n487 = x111 & ~n486 ;
  assign n488 = n261 & ~n386 ;
  assign n489 = ~n139 & n488 ;
  assign n490 = n341 ^ n142 ^ x114 ;
  assign n491 = n490 ^ n259 ^ n249 ;
  assign n492 = n184 ^ x32 ^ 1'b0 ;
  assign n493 = x94 & n492 ;
  assign n494 = x102 & ~n493 ;
  assign n495 = n438 ^ n169 ^ 1'b0 ;
  assign n496 = n218 & ~n495 ;
  assign n497 = ( x54 & ~n327 ) | ( x54 & n421 ) | ( ~n327 & n421 ) ;
  assign n498 = n497 ^ n434 ^ 1'b0 ;
  assign n499 = ~n279 & n498 ;
  assign n500 = n497 ^ x16 ^ 1'b0 ;
  assign n501 = x110 & ~n500 ;
  assign n502 = n441 ^ n349 ^ x6 ;
  assign n503 = x49 & n389 ;
  assign n504 = ~n502 & n503 ;
  assign n505 = x120 & ~n441 ;
  assign n506 = n505 ^ n401 ^ 1'b0 ;
  assign n507 = n471 & ~n506 ;
  assign n508 = n507 ^ n381 ^ 1'b0 ;
  assign n509 = n347 ^ n288 ^ x77 ;
  assign n510 = x34 & n186 ;
  assign n511 = n510 ^ n456 ^ n452 ;
  assign n513 = x127 & ~n231 ;
  assign n514 = n227 & n513 ;
  assign n512 = n232 ^ x97 ^ 1'b0 ;
  assign n515 = n514 ^ n512 ^ n216 ;
  assign n516 = n131 | n231 ;
  assign n517 = x16 | n516 ;
  assign n518 = n517 ^ n372 ^ x82 ;
  assign n519 = n518 ^ n332 ^ 1'b0 ;
  assign n520 = x75 & n519 ;
  assign n521 = x126 ^ x4 ^ 1'b0 ;
  assign n522 = ( n193 & ~n281 ) | ( n193 & n340 ) | ( ~n281 & n340 ) ;
  assign n523 = x87 & ~x119 ;
  assign n524 = x15 & n523 ;
  assign n525 = n524 ^ x20 ^ 1'b0 ;
  assign n526 = n525 ^ n370 ^ x106 ;
  assign n527 = n290 & ~n458 ;
  assign n528 = n527 ^ n227 ^ 1'b0 ;
  assign n529 = ( ~n522 & n526 ) | ( ~n522 & n528 ) | ( n526 & n528 ) ;
  assign n530 = n438 ^ x65 ^ x43 ;
  assign n531 = n530 ^ n487 ^ x125 ;
  assign n532 = x24 & n158 ;
  assign n533 = n532 ^ x52 ^ 1'b0 ;
  assign n534 = n272 & ~n533 ;
  assign n535 = n534 ^ n316 ^ 1'b0 ;
  assign n536 = ( x66 & ~n140 ) | ( x66 & n281 ) | ( ~n140 & n281 ) ;
  assign n537 = n536 ^ n289 ^ n205 ;
  assign n539 = x77 & n318 ;
  assign n540 = n539 ^ x35 ^ 1'b0 ;
  assign n541 = n540 ^ n252 ^ x116 ;
  assign n538 = x17 & n436 ;
  assign n542 = n541 ^ n538 ^ 1'b0 ;
  assign n543 = x116 | n542 ;
  assign n544 = n138 ^ x47 ^ 1'b0 ;
  assign n545 = x94 & ~n544 ;
  assign n546 = x2 & n545 ;
  assign n547 = n272 & n546 ;
  assign n548 = n547 ^ n420 ^ 1'b0 ;
  assign n549 = x54 ^ x12 ^ 1'b0 ;
  assign n550 = n207 & n549 ;
  assign n551 = ( x71 & n303 ) | ( x71 & ~n550 ) | ( n303 & ~n550 ) ;
  assign n552 = n216 | n551 ;
  assign n553 = n552 ^ x96 ^ 1'b0 ;
  assign n554 = n379 ^ x117 ^ 1'b0 ;
  assign n555 = ( x49 & ~x56 ) | ( x49 & n554 ) | ( ~x56 & n554 ) ;
  assign n556 = n233 & ~n473 ;
  assign n557 = ~n304 & n556 ;
  assign n559 = n165 ^ x35 ^ 1'b0 ;
  assign n560 = x52 & ~n559 ;
  assign n558 = n162 & n276 ;
  assign n561 = n560 ^ n558 ^ 1'b0 ;
  assign n562 = n561 ^ n528 ^ n207 ;
  assign n563 = ( ~x18 & x24 ) | ( ~x18 & x45 ) | ( x24 & x45 ) ;
  assign n564 = n563 ^ x77 ^ 1'b0 ;
  assign n565 = ~n190 & n564 ;
  assign n566 = n195 ^ x58 ^ 1'b0 ;
  assign n567 = n566 ^ n474 ^ 1'b0 ;
  assign n568 = n533 | n567 ;
  assign n569 = n140 ^ x0 ^ 1'b0 ;
  assign n571 = ~n157 & n296 ;
  assign n570 = x115 & n245 ;
  assign n572 = n571 ^ n570 ^ 1'b0 ;
  assign n573 = n536 ^ n154 ^ n138 ;
  assign n574 = n129 & n258 ;
  assign n575 = ~x119 & n574 ;
  assign n576 = ( n158 & n573 ) | ( n158 & n575 ) | ( n573 & n575 ) ;
  assign n577 = n222 & ~n451 ;
  assign n578 = ~n576 & n577 ;
  assign n579 = ( n136 & n365 ) | ( n136 & ~n578 ) | ( n365 & ~n578 ) ;
  assign n580 = n499 ^ n415 ^ n320 ;
  assign n581 = ~n331 & n522 ;
  assign n582 = n484 & n581 ;
  assign n583 = n463 & ~n582 ;
  assign n584 = n583 ^ x11 ^ 1'b0 ;
  assign n585 = n526 ^ x35 ^ 1'b0 ;
  assign n586 = n582 ^ x45 ^ x5 ;
  assign n587 = n207 ^ n164 ^ 1'b0 ;
  assign n588 = n434 ^ x75 ^ 1'b0 ;
  assign n589 = n588 ^ n384 ^ n365 ;
  assign n590 = n168 & n413 ;
  assign n591 = n590 ^ x81 ^ 1'b0 ;
  assign n592 = n589 & ~n591 ;
  assign n593 = ~x26 & n592 ;
  assign n594 = n234 ^ n219 ^ x46 ;
  assign n595 = ( ~x112 & n196 ) | ( ~x112 & n594 ) | ( n196 & n594 ) ;
  assign n596 = x18 & ~n595 ;
  assign n597 = n596 ^ x15 ^ 1'b0 ;
  assign n598 = n360 | n597 ;
  assign n599 = n139 | n598 ;
  assign n600 = n521 ^ x77 ^ x18 ;
  assign n601 = n211 & n232 ;
  assign n605 = x28 & ~n134 ;
  assign n606 = ~x33 & n605 ;
  assign n602 = x120 & n324 ;
  assign n603 = n281 & n602 ;
  assign n604 = n484 | n603 ;
  assign n607 = n606 ^ n604 ^ 1'b0 ;
  assign n608 = n350 ^ n298 ^ n206 ;
  assign n609 = n608 ^ n292 ^ n133 ;
  assign n610 = n142 & n609 ;
  assign n611 = n607 & n610 ;
  assign n612 = n601 | n611 ;
  assign n613 = n600 & ~n612 ;
  assign n614 = n355 | n475 ;
  assign n615 = n614 ^ n266 ^ 1'b0 ;
  assign n616 = x98 & ~n615 ;
  assign n617 = n207 ^ x11 ^ 1'b0 ;
  assign n618 = ( n161 & ~n257 ) | ( n161 & n617 ) | ( ~n257 & n617 ) ;
  assign n619 = n271 & ~n618 ;
  assign n620 = n619 ^ x125 ^ 1'b0 ;
  assign n621 = n620 ^ n452 ^ 1'b0 ;
  assign n622 = ( x59 & ~n616 ) | ( x59 & n621 ) | ( ~n616 & n621 ) ;
  assign n623 = x49 & n424 ;
  assign n624 = n623 ^ x114 ^ 1'b0 ;
  assign n625 = ( ~n343 & n413 ) | ( ~n343 & n545 ) | ( n413 & n545 ) ;
  assign n626 = n165 ^ x112 ^ 1'b0 ;
  assign n627 = n626 ^ n164 ^ x87 ;
  assign n628 = n299 ^ x125 ^ 1'b0 ;
  assign n629 = n627 & ~n628 ;
  assign n630 = ~x86 & n629 ;
  assign n631 = n586 ^ n256 ^ x6 ;
  assign n632 = n161 ^ x96 ^ 1'b0 ;
  assign n633 = n415 ^ n350 ^ 1'b0 ;
  assign n634 = n632 & n633 ;
  assign n635 = x93 | n154 ;
  assign n636 = x119 ^ x53 ^ 1'b0 ;
  assign n637 = n401 & n636 ;
  assign n638 = n637 ^ n425 ^ 1'b0 ;
  assign n639 = x87 & ~n638 ;
  assign n640 = ~n380 & n639 ;
  assign n641 = n640 ^ n389 ^ 1'b0 ;
  assign n642 = x50 & ~n641 ;
  assign n643 = ~n635 & n642 ;
  assign n644 = ( x67 & n393 ) | ( x67 & ~n643 ) | ( n393 & ~n643 ) ;
  assign n645 = x119 & n313 ;
  assign n646 = n645 ^ x40 ^ 1'b0 ;
  assign n650 = n134 ^ x81 ^ x68 ;
  assign n647 = n419 & n566 ;
  assign n648 = ~n404 & n647 ;
  assign n649 = ( x27 & ~n309 ) | ( x27 & n648 ) | ( ~n309 & n648 ) ;
  assign n651 = n650 ^ n649 ^ 1'b0 ;
  assign n652 = n643 | n651 ;
  assign n653 = n349 ^ n157 ^ x80 ;
  assign n654 = n606 ^ n496 ^ x49 ;
  assign n656 = n606 ^ n541 ^ 1'b0 ;
  assign n657 = x118 & ~n656 ;
  assign n655 = n167 | n614 ;
  assign n658 = n657 ^ n655 ^ 1'b0 ;
  assign n659 = ~n643 & n658 ;
  assign n660 = n659 ^ n356 ^ 1'b0 ;
  assign n663 = x72 ^ x51 ^ 1'b0 ;
  assign n661 = ~n421 & n525 ;
  assign n662 = x73 & ~n661 ;
  assign n664 = n663 ^ n662 ^ 1'b0 ;
  assign n665 = n403 ^ n368 ^ x85 ;
  assign n666 = x116 & ~n514 ;
  assign n667 = n666 ^ n289 ^ 1'b0 ;
  assign n668 = ~n665 & n667 ;
  assign n669 = n668 ^ x121 ^ 1'b0 ;
  assign n670 = n225 & ~n669 ;
  assign n671 = ~n161 & n206 ;
  assign n672 = ~x18 & n671 ;
  assign n673 = n672 ^ n143 ^ 1'b0 ;
  assign n683 = n314 ^ n139 ^ 1'b0 ;
  assign n684 = x3 & n683 ;
  assign n674 = n186 ^ n184 ^ 1'b0 ;
  assign n675 = x37 & ~n674 ;
  assign n676 = n675 ^ x30 ^ 1'b0 ;
  assign n677 = x25 & n676 ;
  assign n678 = x91 ^ x4 ^ 1'b0 ;
  assign n679 = x118 & n678 ;
  assign n680 = ~n150 & n679 ;
  assign n681 = ~n677 & n680 ;
  assign n682 = n485 & ~n681 ;
  assign n685 = n684 ^ n682 ^ 1'b0 ;
  assign n686 = n626 ^ n252 ^ n164 ;
  assign n687 = n686 ^ n624 ^ 1'b0 ;
  assign n688 = n292 & ~n687 ;
  assign n689 = ~n138 & n622 ;
  assign n690 = n504 & n689 ;
  assign n691 = x38 & x120 ;
  assign n692 = ~n635 & n691 ;
  assign n693 = n514 & ~n692 ;
  assign n694 = n323 ^ x27 ^ 1'b0 ;
  assign n695 = ~x106 & n286 ;
  assign n696 = ~n477 & n695 ;
  assign n697 = n250 | n696 ;
  assign n698 = n307 & ~n412 ;
  assign n699 = ~n276 & n698 ;
  assign n700 = ( ~x31 & x81 ) | ( ~x31 & n699 ) | ( x81 & n699 ) ;
  assign n701 = n467 ^ n266 ^ x108 ;
  assign n703 = x87 & n158 ;
  assign n704 = n703 ^ n313 ^ 1'b0 ;
  assign n702 = x42 & x127 ;
  assign n705 = n704 ^ n702 ^ 1'b0 ;
  assign n706 = n240 | n256 ;
  assign n707 = ~n579 & n706 ;
  assign n708 = ~n139 & n707 ;
  assign n709 = ( n652 & n705 ) | ( n652 & ~n708 ) | ( n705 & ~n708 ) ;
  assign n710 = n169 ^ n146 ^ x65 ;
  assign n711 = n710 ^ n582 ^ 1'b0 ;
  assign n712 = n146 & ~n167 ;
  assign n713 = x47 & n377 ;
  assign n714 = n713 ^ n627 ^ 1'b0 ;
  assign n716 = ( ~x72 & x87 ) | ( ~x72 & n168 ) | ( x87 & n168 ) ;
  assign n715 = n398 ^ n358 ^ n216 ;
  assign n717 = n716 ^ n715 ^ 1'b0 ;
  assign n718 = x110 & n717 ;
  assign n719 = n718 ^ n349 ^ 1'b0 ;
  assign n720 = n563 ^ x37 ^ 1'b0 ;
  assign n721 = x94 & n720 ;
  assign n722 = n721 ^ n459 ^ 1'b0 ;
  assign n723 = ~n227 & n722 ;
  assign n724 = x36 & n723 ;
  assign n725 = ~x108 & n724 ;
  assign n726 = n725 ^ n575 ^ n528 ;
  assign n727 = n139 & ~n679 ;
  assign n728 = x91 & ~n595 ;
  assign n729 = n728 ^ x102 ^ 1'b0 ;
  assign n730 = n289 & ~n641 ;
  assign n731 = n474 & n730 ;
  assign n732 = ( x79 & n355 ) | ( x79 & ~n731 ) | ( n355 & ~n731 ) ;
  assign n733 = x13 & n401 ;
  assign n734 = n372 & n733 ;
  assign n735 = n422 ^ n290 ^ 1'b0 ;
  assign n736 = ( n398 & n734 ) | ( n398 & n735 ) | ( n734 & n735 ) ;
  assign n737 = ( x17 & n523 ) | ( x17 & n736 ) | ( n523 & n736 ) ;
  assign n738 = n737 ^ x45 ^ 1'b0 ;
  assign n739 = n444 & n738 ;
  assign n740 = n138 ^ x93 ^ x20 ;
  assign n741 = ( x122 & n203 ) | ( x122 & n740 ) | ( n203 & n740 ) ;
  assign n742 = n225 ^ x49 ^ 1'b0 ;
  assign n743 = n742 ^ n160 ^ 1'b0 ;
  assign n744 = n741 & n743 ;
  assign n745 = x51 & x80 ;
  assign n746 = n745 ^ n175 ^ 1'b0 ;
  assign n747 = n620 | n664 ;
  assign n748 = n594 ^ n272 ^ n207 ;
  assign n749 = n413 & ~n748 ;
  assign n750 = ~n374 & n749 ;
  assign n751 = ~n424 & n750 ;
  assign n752 = n332 & n337 ;
  assign n753 = n752 ^ n288 ^ 1'b0 ;
  assign n759 = n362 | n449 ;
  assign n754 = x3 & x10 ;
  assign n755 = n754 ^ n368 ^ 1'b0 ;
  assign n756 = n218 & ~n755 ;
  assign n760 = n759 ^ n756 ^ 1'b0 ;
  assign n757 = x125 & n756 ;
  assign n758 = n757 ^ n430 ^ 1'b0 ;
  assign n761 = n760 ^ n758 ^ n293 ;
  assign n762 = n227 | n761 ;
  assign n763 = n762 ^ n573 ^ 1'b0 ;
  assign n764 = x61 & n233 ;
  assign n765 = n764 ^ n456 ^ 1'b0 ;
  assign n766 = x115 ^ x23 ^ 1'b0 ;
  assign n767 = n155 & n766 ;
  assign n768 = ( n433 & ~n765 ) | ( n433 & n767 ) | ( ~n765 & n767 ) ;
  assign n769 = n768 ^ n709 ^ 1'b0 ;
  assign n770 = ~n694 & n769 ;
  assign n771 = n393 ^ n142 ^ 1'b0 ;
  assign n772 = n771 ^ n250 ^ 1'b0 ;
  assign n773 = n205 & ~n772 ;
  assign n774 = x68 ^ x10 ^ 1'b0 ;
  assign n775 = n723 & n774 ;
  assign n776 = x81 | n267 ;
  assign n777 = ~n361 & n776 ;
  assign n778 = ~n775 & n777 ;
  assign n779 = n444 ^ n233 ^ x40 ;
  assign n780 = n334 & ~n779 ;
  assign n781 = n780 ^ n474 ^ 1'b0 ;
  assign n782 = n608 & n781 ;
  assign n783 = x34 & ~n189 ;
  assign n784 = n783 ^ x43 ^ 1'b0 ;
  assign n785 = n784 ^ n553 ^ n531 ;
  assign n786 = n328 | n548 ;
  assign n787 = x77 & ~n133 ;
  assign n788 = n787 ^ n173 ^ 1'b0 ;
  assign n789 = n442 ^ n167 ^ 1'b0 ;
  assign n790 = n776 & ~n789 ;
  assign n791 = n303 ^ x55 ^ x19 ;
  assign n792 = n744 ^ x86 ^ 1'b0 ;
  assign n793 = n791 & n792 ;
  assign n794 = n335 | n624 ;
  assign n795 = n413 ^ x109 ^ 1'b0 ;
  assign n796 = n522 & n741 ;
  assign n797 = ~n207 & n354 ;
  assign n798 = n797 ^ n343 ^ n221 ;
  assign n799 = ( x109 & n797 ) | ( x109 & n798 ) | ( n797 & n798 ) ;
  assign n800 = n443 ^ n247 ^ x105 ;
  assign n801 = n236 & n800 ;
  assign n802 = ( x12 & x43 ) | ( x12 & n322 ) | ( x43 & n322 ) ;
  assign n803 = n802 ^ n746 ^ n686 ;
  assign n804 = ( n240 & n517 ) | ( n240 & n560 ) | ( n517 & n560 ) ;
  assign n805 = ( n304 & ~n313 ) | ( n304 & n804 ) | ( ~n313 & n804 ) ;
  assign n806 = n723 & n781 ;
  assign n807 = ~n737 & n806 ;
  assign n808 = n210 & n807 ;
  assign n809 = ~n526 & n585 ;
  assign n811 = ( x8 & ~n163 ) | ( x8 & n355 ) | ( ~n163 & n355 ) ;
  assign n810 = ~x107 & n252 ;
  assign n812 = n811 ^ n810 ^ n779 ;
  assign n819 = n248 ^ n162 ^ 1'b0 ;
  assign n820 = n649 ^ n461 ^ x13 ;
  assign n821 = n819 & ~n820 ;
  assign n822 = n821 ^ n194 ^ 1'b0 ;
  assign n814 = x110 ^ x1 ^ 1'b0 ;
  assign n815 = x30 & n814 ;
  assign n816 = n815 ^ n517 ^ x71 ;
  assign n817 = n816 ^ n389 ^ n285 ;
  assign n813 = ~x33 & x110 ;
  assign n818 = n817 ^ n813 ^ 1'b0 ;
  assign n823 = n822 ^ n818 ^ n541 ;
  assign n824 = ( x101 & ~n162 ) | ( x101 & n603 ) | ( ~n162 & n603 ) ;
  assign n825 = n286 ^ x109 ^ 1'b0 ;
  assign n826 = ~n824 & n825 ;
  assign n827 = ~n621 & n826 ;
  assign n828 = ( x60 & x81 ) | ( x60 & ~x94 ) | ( x81 & ~x94 ) ;
  assign n829 = ( x108 & ~n247 ) | ( x108 & n828 ) | ( ~n247 & n828 ) ;
  assign n830 = n168 & n829 ;
  assign n831 = ~x49 & n830 ;
  assign n832 = n831 ^ n462 ^ x14 ;
  assign n833 = n211 ^ x23 ^ 1'b0 ;
  assign n834 = n833 ^ x76 ^ x25 ;
  assign n835 = x27 & x65 ;
  assign n836 = ~x41 & n835 ;
  assign n837 = n134 | n836 ;
  assign n838 = n837 ^ n180 ^ 1'b0 ;
  assign n839 = ~x25 & n637 ;
  assign n840 = n838 | n839 ;
  assign n841 = n840 ^ n458 ^ 1'b0 ;
  assign n842 = n209 & ~n494 ;
  assign n843 = ~x20 & n842 ;
  assign n844 = n843 ^ n677 ^ 1'b0 ;
  assign n845 = n543 ^ n170 ^ 1'b0 ;
  assign n846 = n542 ^ n430 ^ 1'b0 ;
  assign n847 = n391 | n846 ;
  assign n848 = n644 ^ n195 ^ 1'b0 ;
  assign n849 = n631 & n663 ;
  assign n850 = n210 ^ n177 ^ x6 ;
  assign n851 = x101 ^ x33 ^ 1'b0 ;
  assign n852 = x16 & n851 ;
  assign n853 = ~n692 & n852 ;
  assign n854 = n853 ^ n309 ^ 1'b0 ;
  assign n855 = n850 & n854 ;
  assign n856 = n855 ^ n701 ^ 1'b0 ;
  assign n857 = ~n849 & n856 ;
  assign n858 = n361 ^ n341 ^ x43 ;
  assign n859 = x24 | n858 ;
  assign n860 = n706 ^ n694 ^ 1'b0 ;
  assign n861 = n184 & ~n353 ;
  assign n862 = ~n401 & n861 ;
  assign n864 = n334 & ~n617 ;
  assign n865 = n864 ^ n370 ^ 1'b0 ;
  assign n863 = x106 | n186 ;
  assign n866 = n865 ^ n863 ^ 1'b0 ;
  assign n867 = n173 | n866 ;
  assign n868 = n867 ^ n787 ^ n214 ;
  assign n869 = n862 | n868 ;
  assign n870 = x64 | n869 ;
  assign n871 = n723 ^ x94 ^ 1'b0 ;
  assign n872 = n562 & n871 ;
  assign n873 = x79 ^ x24 ^ 1'b0 ;
  assign n874 = n245 & n873 ;
  assign n875 = ~n154 & n874 ;
  assign n876 = n875 ^ n608 ^ 1'b0 ;
  assign n877 = ~x65 & n876 ;
  assign n878 = n181 & ~n209 ;
  assign n879 = n878 ^ n672 ^ n588 ;
  assign n880 = n748 ^ n418 ^ 1'b0 ;
  assign n881 = n363 & n880 ;
  assign n882 = ( x108 & n657 ) | ( x108 & ~n881 ) | ( n657 & ~n881 ) ;
  assign n883 = ( ~x26 & x71 ) | ( ~x26 & x73 ) | ( x71 & x73 ) ;
  assign n884 = n741 & n883 ;
  assign n885 = n384 & n884 ;
  assign n886 = ~n219 & n264 ;
  assign n887 = n886 ^ n178 ^ 1'b0 ;
  assign n892 = n279 ^ x59 ^ 1'b0 ;
  assign n893 = n271 & n892 ;
  assign n894 = n232 & n251 ;
  assign n895 = ~x31 & n894 ;
  assign n896 = n221 ^ x112 ^ 1'b0 ;
  assign n897 = x115 & n896 ;
  assign n898 = n897 ^ n585 ^ 1'b0 ;
  assign n899 = n895 | n898 ;
  assign n900 = n893 & ~n899 ;
  assign n889 = n177 ^ x65 ^ 1'b0 ;
  assign n890 = n264 | n889 ;
  assign n891 = n829 | n890 ;
  assign n888 = n712 ^ n704 ^ x83 ;
  assign n901 = n900 ^ n891 ^ n888 ;
  assign n902 = n368 & ~n890 ;
  assign n903 = n902 ^ x30 ^ 1'b0 ;
  assign n904 = ( ~x48 & n337 ) | ( ~x48 & n903 ) | ( n337 & n903 ) ;
  assign n905 = n146 & ~n212 ;
  assign n906 = n692 | n905 ;
  assign n907 = x84 & x113 ;
  assign n908 = n907 ^ n787 ^ 1'b0 ;
  assign n909 = n908 ^ n850 ^ n256 ;
  assign n912 = n550 ^ n469 ^ 1'b0 ;
  assign n913 = ~n452 & n912 ;
  assign n910 = n390 & ~n708 ;
  assign n911 = n910 ^ n776 ^ 1'b0 ;
  assign n914 = n913 ^ n911 ^ n456 ;
  assign n915 = n632 ^ n351 ^ x101 ;
  assign n916 = n153 ^ x44 ^ 1'b0 ;
  assign n917 = n916 ^ x23 ^ 1'b0 ;
  assign n918 = n917 ^ n650 ^ n611 ;
  assign n919 = ~n551 & n918 ;
  assign n920 = n919 ^ n145 ^ 1'b0 ;
  assign n921 = n723 ^ n284 ^ 1'b0 ;
  assign n922 = n415 | n921 ;
  assign n923 = ( n915 & ~n920 ) | ( n915 & n922 ) | ( ~n920 & n922 ) ;
  assign n924 = ~n161 & n828 ;
  assign n925 = n924 ^ n382 ^ 1'b0 ;
  assign n926 = x15 & n271 ;
  assign n927 = n925 & n926 ;
  assign n928 = n927 ^ n816 ^ 1'b0 ;
  assign n930 = n514 | n606 ;
  assign n931 = n930 ^ n276 ^ 1'b0 ;
  assign n929 = n199 ^ x20 ^ 1'b0 ;
  assign n932 = n931 ^ n929 ^ 1'b0 ;
  assign n933 = x122 & ~n932 ;
  assign n934 = x67 & ~n933 ;
  assign n935 = n415 ^ x11 ^ 1'b0 ;
  assign n936 = n935 ^ n748 ^ 1'b0 ;
  assign n937 = n747 ^ n675 ^ 1'b0 ;
  assign n945 = n579 ^ n530 ^ 1'b0 ;
  assign n946 = n945 ^ n561 ^ x97 ;
  assign n940 = x126 ^ x70 ^ 1'b0 ;
  assign n938 = x70 & ~n716 ;
  assign n939 = x56 & ~n938 ;
  assign n941 = n940 ^ n939 ^ 1'b0 ;
  assign n942 = ~n514 & n771 ;
  assign n943 = n942 ^ n641 ^ 1'b0 ;
  assign n944 = n941 | n943 ;
  assign n947 = n946 ^ n944 ^ 1'b0 ;
  assign n948 = ( ~x88 & n418 ) | ( ~x88 & n441 ) | ( n418 & n441 ) ;
  assign n949 = n948 ^ n441 ^ 1'b0 ;
  assign n950 = ~n545 & n949 ;
  assign n951 = n950 ^ n386 ^ n362 ;
  assign n952 = n148 & n706 ;
  assign n953 = ~n951 & n952 ;
  assign n954 = n942 ^ n843 ^ x82 ;
  assign n955 = n314 & ~n423 ;
  assign n956 = n955 ^ x18 ^ 1'b0 ;
  assign n957 = n956 ^ x5 ^ 1'b0 ;
  assign n958 = n251 & ~n957 ;
  assign n959 = n730 & n958 ;
  assign n960 = n959 ^ n891 ^ 1'b0 ;
  assign n967 = ~n238 & n643 ;
  assign n968 = n967 ^ x79 ^ 1'b0 ;
  assign n969 = x86 & ~n968 ;
  assign n961 = n712 ^ x75 ^ 1'b0 ;
  assign n962 = n471 & n961 ;
  assign n963 = n606 ^ n560 ^ n447 ;
  assign n964 = ( x75 & ~n334 ) | ( x75 & n963 ) | ( ~n334 & n963 ) ;
  assign n965 = n964 ^ n849 ^ n561 ;
  assign n966 = n962 & ~n965 ;
  assign n970 = n969 ^ n966 ^ 1'b0 ;
  assign n971 = n607 ^ n292 ^ x14 ;
  assign n972 = n971 ^ n358 ^ 1'b0 ;
  assign n973 = x118 ^ x62 ^ 1'b0 ;
  assign n974 = n459 & n973 ;
  assign n975 = n157 & n184 ;
  assign n976 = n975 ^ n293 ^ 1'b0 ;
  assign n977 = n974 & n976 ;
  assign n983 = n575 ^ n514 ^ n372 ;
  assign n984 = n983 ^ n925 ^ n663 ;
  assign n978 = n199 & n543 ;
  assign n979 = n978 ^ n478 ^ 1'b0 ;
  assign n980 = n828 ^ x40 ^ x18 ;
  assign n981 = n980 ^ n242 ^ 1'b0 ;
  assign n982 = n979 | n981 ;
  assign n985 = n984 ^ n982 ^ 1'b0 ;
  assign n986 = ( n972 & n977 ) | ( n972 & n985 ) | ( n977 & n985 ) ;
  assign n989 = x76 & ~n209 ;
  assign n990 = n293 & n989 ;
  assign n991 = n335 & ~n990 ;
  assign n992 = n211 & n991 ;
  assign n987 = x70 & n485 ;
  assign n988 = ( ~x74 & n330 ) | ( ~x74 & n987 ) | ( n330 & n987 ) ;
  assign n993 = n992 ^ n988 ^ 1'b0 ;
  assign n994 = x40 & ~n614 ;
  assign n995 = ~x9 & n994 ;
  assign n996 = n419 & ~n995 ;
  assign n997 = n996 ^ n931 ^ 1'b0 ;
  assign n998 = ( x74 & n828 ) | ( x74 & n997 ) | ( n828 & n997 ) ;
  assign n999 = n998 ^ n632 ^ 1'b0 ;
  assign n1000 = ~n993 & n999 ;
  assign n1001 = x124 & n225 ;
  assign n1002 = ~n1000 & n1001 ;
  assign n1003 = n249 & n345 ;
  assign n1004 = ( n276 & n810 ) | ( n276 & n1003 ) | ( n810 & n1003 ) ;
  assign n1005 = n229 ^ x10 ^ 1'b0 ;
  assign n1006 = n458 | n1005 ;
  assign n1007 = n535 ^ n430 ^ 1'b0 ;
  assign n1008 = n1006 | n1007 ;
  assign n1009 = n1008 ^ n811 ^ 1'b0 ;
  assign n1010 = n331 | n1009 ;
  assign n1011 = ( n778 & n833 ) | ( n778 & ~n1010 ) | ( n833 & ~n1010 ) ;
  assign n1012 = x96 & n415 ;
  assign n1013 = n751 ^ n573 ^ 1'b0 ;
  assign n1014 = n131 | n1013 ;
  assign n1015 = ~n1012 & n1014 ;
  assign n1016 = n660 | n898 ;
  assign n1017 = n514 & ~n1016 ;
  assign n1018 = n883 ^ n470 ^ n445 ;
  assign n1019 = x86 & ~n820 ;
  assign n1020 = n1019 ^ n663 ^ 1'b0 ;
  assign n1021 = n189 | n608 ;
  assign n1022 = n550 | n1021 ;
  assign n1023 = n1022 ^ n401 ^ x29 ;
  assign n1024 = x102 & n270 ;
  assign n1025 = ~x70 & n1024 ;
  assign n1026 = n169 & n563 ;
  assign n1027 = n1026 ^ x79 ^ 1'b0 ;
  assign n1028 = n1027 ^ x116 ^ 1'b0 ;
  assign n1029 = n1025 | n1028 ;
  assign n1030 = n1023 | n1029 ;
  assign n1031 = n1020 | n1030 ;
  assign n1032 = n813 ^ n276 ^ 1'b0 ;
  assign n1033 = ~n551 & n1032 ;
  assign n1034 = n657 ^ n533 ^ 1'b0 ;
  assign n1035 = n1034 ^ n232 ^ 1'b0 ;
  assign n1036 = ~n372 & n1035 ;
  assign n1037 = ~n288 & n427 ;
  assign n1038 = n1037 ^ n347 ^ 1'b0 ;
  assign n1039 = x18 & ~n1038 ;
  assign n1040 = n403 ^ x126 ^ x75 ;
  assign n1041 = n1040 ^ n327 ^ n153 ;
  assign n1042 = ( n181 & ~n900 ) | ( n181 & n1041 ) | ( ~n900 & n1041 ) ;
  assign n1043 = x61 & n563 ;
  assign n1044 = n525 ^ n136 ^ 1'b0 ;
  assign n1045 = n1043 & n1044 ;
  assign n1046 = ~n737 & n1045 ;
  assign n1047 = n447 | n1046 ;
  assign n1048 = ~n295 & n328 ;
  assign n1049 = ~n290 & n1048 ;
  assign n1050 = n278 & ~n595 ;
  assign n1051 = n1050 ^ n677 ^ 1'b0 ;
  assign n1052 = n300 | n1051 ;
  assign n1053 = n497 & ~n1052 ;
  assign n1054 = ( n307 & n1049 ) | ( n307 & n1053 ) | ( n1049 & n1053 ) ;
  assign n1055 = n138 | n1054 ;
  assign n1056 = n314 ^ x45 ^ 1'b0 ;
  assign n1057 = x90 & n1056 ;
  assign n1058 = n1057 ^ n849 ^ 1'b0 ;
  assign n1059 = n1058 ^ n491 ^ 1'b0 ;
  assign n1060 = n478 & ~n1059 ;
  assign n1061 = n850 ^ x115 ^ x83 ;
  assign n1062 = n1061 ^ n639 ^ n469 ;
  assign n1063 = n399 & n1062 ;
  assign n1064 = n1063 ^ n129 ^ 1'b0 ;
  assign n1065 = n916 ^ n588 ^ n427 ;
  assign n1066 = x90 & ~n510 ;
  assign n1067 = x17 & n1066 ;
  assign n1068 = x26 & ~n1067 ;
  assign n1070 = n473 ^ x12 ^ 1'b0 ;
  assign n1071 = n320 & ~n1070 ;
  assign n1072 = ~n216 & n1071 ;
  assign n1073 = n711 & n1072 ;
  assign n1069 = n307 | n325 ;
  assign n1074 = n1073 ^ n1069 ^ n667 ;
  assign n1075 = ~n307 & n490 ;
  assign n1076 = ( n218 & n412 ) | ( n218 & n1075 ) | ( n412 & n1075 ) ;
  assign n1077 = n622 ^ n550 ^ 1'b0 ;
  assign n1078 = n1076 & n1077 ;
  assign n1079 = n419 ^ n356 ^ 1'b0 ;
  assign n1080 = ( ~n309 & n314 ) | ( ~n309 & n1006 ) | ( n314 & n1006 ) ;
  assign n1081 = n948 ^ x108 ^ 1'b0 ;
  assign n1082 = n443 & ~n1081 ;
  assign n1083 = ( n617 & ~n953 ) | ( n617 & n1082 ) | ( ~n953 & n1082 ) ;
  assign n1084 = ( x20 & x24 ) | ( x20 & ~n247 ) | ( x24 & ~n247 ) ;
  assign n1085 = n760 & n1084 ;
  assign n1086 = n1085 ^ n848 ^ 1'b0 ;
  assign n1087 = n715 ^ n443 ^ 1'b0 ;
  assign n1088 = x2 & n1087 ;
  assign n1089 = n429 & n1088 ;
  assign n1090 = n811 & ~n1089 ;
  assign n1091 = ( n339 & n542 ) | ( n339 & n964 ) | ( n542 & n964 ) ;
  assign n1092 = ( x30 & ~n433 ) | ( x30 & n1091 ) | ( ~n433 & n1091 ) ;
  assign n1093 = n429 & n478 ;
  assign n1094 = n1093 ^ n196 ^ x81 ;
  assign n1095 = n874 ^ n831 ^ 1'b0 ;
  assign n1096 = n1094 | n1095 ;
  assign n1097 = n1092 | n1096 ;
  assign n1098 = x2 | n1097 ;
  assign n1099 = n163 | n845 ;
  assign n1100 = n828 ^ n679 ^ 1'b0 ;
  assign n1101 = ~n281 & n510 ;
  assign n1102 = ( n730 & n935 ) | ( n730 & n1101 ) | ( n935 & n1101 ) ;
  assign n1103 = n1100 & n1102 ;
  assign n1104 = ~n634 & n1103 ;
  assign n1109 = n209 ^ x103 ^ 1'b0 ;
  assign n1110 = n260 | n1109 ;
  assign n1111 = n1110 ^ n210 ^ 1'b0 ;
  assign n1112 = x4 & ~n1111 ;
  assign n1113 = n1112 ^ n508 ^ 1'b0 ;
  assign n1105 = ~n229 & n381 ;
  assign n1106 = n1105 ^ x43 ^ 1'b0 ;
  assign n1107 = ( ~n441 & n618 ) | ( ~n441 & n1106 ) | ( n618 & n1106 ) ;
  assign n1108 = n1107 ^ n927 ^ n467 ;
  assign n1114 = n1113 ^ n1108 ^ 1'b0 ;
  assign n1116 = ( x127 & n432 ) | ( x127 & ~n718 ) | ( n432 & ~n718 ) ;
  assign n1117 = n345 & ~n734 ;
  assign n1118 = ~n1116 & n1117 ;
  assign n1119 = n569 | n1118 ;
  assign n1120 = n1119 ^ n331 ^ 1'b0 ;
  assign n1115 = n278 & n697 ;
  assign n1121 = n1120 ^ n1115 ^ 1'b0 ;
  assign n1122 = n354 ^ n300 ^ 1'b0 ;
  assign n1123 = n461 | n1122 ;
  assign n1124 = n1042 & ~n1123 ;
  assign n1125 = ( ~n323 & n853 ) | ( ~n323 & n927 ) | ( n853 & n927 ) ;
  assign n1126 = n781 & ~n1125 ;
  assign n1127 = x28 & n1126 ;
  assign n1128 = n550 & ~n603 ;
  assign n1129 = n134 & n1128 ;
  assign n1130 = ( n285 & n561 ) | ( n285 & n611 ) | ( n561 & n611 ) ;
  assign n1131 = ( x31 & ~n1129 ) | ( x31 & n1130 ) | ( ~n1129 & n1130 ) ;
  assign n1132 = ( n572 & n586 ) | ( n572 & n679 ) | ( n586 & n679 ) ;
  assign n1133 = ( n172 & n270 ) | ( n172 & ~n1132 ) | ( n270 & ~n1132 ) ;
  assign n1136 = ( x47 & ~n471 ) | ( x47 & n704 ) | ( ~n471 & n704 ) ;
  assign n1137 = n1136 ^ n404 ^ 1'b0 ;
  assign n1134 = x12 & n975 ;
  assign n1135 = ~n675 & n1134 ;
  assign n1138 = n1137 ^ n1135 ^ 1'b0 ;
  assign n1140 = n948 ^ n365 ^ x12 ;
  assign n1139 = n668 ^ n608 ^ 1'b0 ;
  assign n1141 = n1140 ^ n1139 ^ n609 ;
  assign n1142 = n828 & ~n1141 ;
  assign n1143 = n1142 ^ n770 ^ 1'b0 ;
  assign n1144 = x17 & n537 ;
  assign n1145 = n510 & n1144 ;
  assign n1146 = n1145 ^ n425 ^ 1'b0 ;
  assign n1152 = n627 ^ x19 ^ 1'b0 ;
  assign n1147 = x87 ^ x60 ^ 1'b0 ;
  assign n1148 = n438 | n566 ;
  assign n1149 = n1148 ^ n508 ^ 1'b0 ;
  assign n1150 = n1147 | n1149 ;
  assign n1151 = n419 & ~n1150 ;
  assign n1153 = n1152 ^ n1151 ^ 1'b0 ;
  assign n1154 = n609 ^ n199 ^ 1'b0 ;
  assign n1155 = x3 & ~n1154 ;
  assign n1156 = n1155 ^ n220 ^ 1'b0 ;
  assign n1157 = n1156 ^ n824 ^ n453 ;
  assign n1158 = n735 ^ n684 ^ 1'b0 ;
  assign n1159 = n1158 ^ n569 ^ n475 ;
  assign n1160 = n390 | n1159 ;
  assign n1165 = n413 ^ n380 ^ n195 ;
  assign n1164 = n232 ^ n209 ^ x116 ;
  assign n1161 = n214 | n938 ;
  assign n1162 = n1161 ^ n357 ^ 1'b0 ;
  assign n1163 = n1162 ^ n1075 ^ n487 ;
  assign n1166 = n1165 ^ n1164 ^ n1163 ;
  assign n1167 = ( n629 & n1160 ) | ( n629 & ~n1166 ) | ( n1160 & ~n1166 ) ;
  assign n1168 = x122 ^ x108 ^ 1'b0 ;
  assign n1169 = x18 & x101 ;
  assign n1170 = ~x37 & n1169 ;
  assign n1171 = n1170 ^ n214 ^ n211 ;
  assign n1172 = n987 ^ x99 ^ 1'b0 ;
  assign n1173 = ~n154 & n1172 ;
  assign n1174 = n231 | n575 ;
  assign n1175 = n1173 | n1174 ;
  assign n1176 = n988 ^ n456 ^ n223 ;
  assign n1177 = ( n1171 & n1175 ) | ( n1171 & n1176 ) | ( n1175 & n1176 ) ;
  assign n1178 = n1177 ^ n270 ^ 1'b0 ;
  assign n1179 = n1168 & n1178 ;
  assign n1180 = n1124 ^ x16 ^ 1'b0 ;
  assign n1181 = n706 & n1180 ;
  assign n1182 = x15 & x17 ;
  assign n1183 = n347 & n1182 ;
  assign n1184 = n1183 ^ n1076 ^ n650 ;
  assign n1185 = n693 ^ n650 ^ 1'b0 ;
  assign n1186 = n285 ^ x1 ^ 1'b0 ;
  assign n1187 = n1035 & n1186 ;
  assign n1188 = ~n356 & n1187 ;
  assign n1191 = n365 | n465 ;
  assign n1192 = n684 | n1191 ;
  assign n1189 = n979 ^ n506 ^ 1'b0 ;
  assign n1190 = n310 & n1189 ;
  assign n1193 = n1192 ^ n1190 ^ 1'b0 ;
  assign n1194 = ~n374 & n1193 ;
  assign n1195 = n589 ^ n211 ^ 1'b0 ;
  assign n1196 = ~n585 & n1195 ;
  assign n1197 = n1196 ^ n1175 ^ 1'b0 ;
  assign n1198 = n274 | n1197 ;
  assign n1199 = n557 & ~n944 ;
  assign n1200 = ( x0 & ~x53 ) | ( x0 & n609 ) | ( ~x53 & n609 ) ;
  assign n1201 = n1200 ^ n322 ^ x58 ;
  assign n1202 = n452 ^ x45 ^ 1'b0 ;
  assign n1203 = n1202 ^ n1010 ^ 1'b0 ;
  assign n1204 = x49 ^ x24 ^ 1'b0 ;
  assign n1205 = x39 & n1204 ;
  assign n1206 = n1205 ^ n390 ^ 1'b0 ;
  assign n1207 = n1203 & n1206 ;
  assign n1209 = ( n303 & n673 ) | ( n303 & ~n992 ) | ( n673 & ~n992 ) ;
  assign n1208 = n401 & ~n1046 ;
  assign n1210 = n1209 ^ n1208 ^ 1'b0 ;
  assign n1211 = n1210 ^ n1181 ^ 1'b0 ;
  assign n1218 = n565 ^ x82 ^ 1'b0 ;
  assign n1219 = n1218 ^ x113 ^ 1'b0 ;
  assign n1220 = ~n434 & n1219 ;
  assign n1212 = n829 ^ n637 ^ x43 ;
  assign n1213 = n846 | n938 ;
  assign n1214 = n1212 & ~n1213 ;
  assign n1215 = n673 ^ n148 ^ 1'b0 ;
  assign n1216 = ~n588 & n1215 ;
  assign n1217 = n1214 | n1216 ;
  assign n1221 = n1220 ^ n1217 ^ 1'b0 ;
  assign n1222 = n788 ^ n664 ^ x17 ;
  assign n1223 = n250 & n1222 ;
  assign n1224 = n1223 ^ n918 ^ 1'b0 ;
  assign n1225 = n187 & ~n465 ;
  assign n1226 = n196 & n1225 ;
  assign n1227 = x11 & ~n1226 ;
  assign n1228 = ~n259 & n349 ;
  assign n1229 = n1228 ^ n974 ^ 1'b0 ;
  assign n1230 = n474 | n1229 ;
  assign n1231 = x88 & n152 ;
  assign n1232 = ~n340 & n1231 ;
  assign n1233 = n1230 & n1232 ;
  assign n1234 = n1233 ^ n331 ^ 1'b0 ;
  assign n1235 = n240 | n859 ;
  assign n1236 = x99 | n1235 ;
  assign n1237 = x93 & n721 ;
  assign n1238 = ~n389 & n1237 ;
  assign n1239 = n1238 ^ x113 ^ 1'b0 ;
  assign n1240 = n415 | n1239 ;
  assign n1241 = n1240 ^ n776 ^ 1'b0 ;
  assign n1242 = n221 & ~n1241 ;
  assign n1243 = n983 ^ n353 ^ 1'b0 ;
  assign n1244 = x54 & ~n1243 ;
  assign n1250 = ~n739 & n749 ;
  assign n1247 = x53 & ~n710 ;
  assign n1248 = n1247 ^ n663 ^ 1'b0 ;
  assign n1245 = ~n449 & n1082 ;
  assign n1246 = n1245 ^ n705 ^ 1'b0 ;
  assign n1249 = n1248 ^ n1246 ^ n888 ;
  assign n1251 = n1250 ^ n1249 ^ n413 ;
  assign n1252 = ( n225 & ~n809 ) | ( n225 & n1251 ) | ( ~n809 & n1251 ) ;
  assign n1253 = ( ~n1242 & n1244 ) | ( ~n1242 & n1252 ) | ( n1244 & n1252 ) ;
  assign n1254 = n995 ^ n399 ^ x21 ;
  assign n1255 = ~n1051 & n1254 ;
  assign n1256 = ~n931 & n1255 ;
  assign n1257 = n1256 ^ n721 ^ x116 ;
  assign n1258 = ~n281 & n977 ;
  assign n1259 = n1258 ^ n1017 ^ 1'b0 ;
  assign n1261 = ~n164 & n431 ;
  assign n1260 = n289 & ~n865 ;
  assign n1262 = n1261 ^ n1260 ^ n234 ;
  assign n1263 = n272 & ~n860 ;
  assign n1264 = ~n1262 & n1263 ;
  assign n1265 = n920 ^ x127 ^ 1'b0 ;
  assign n1266 = ~n1264 & n1265 ;
  assign n1267 = n1266 ^ n593 ^ 1'b0 ;
  assign n1268 = n881 & ~n1267 ;
  assign n1269 = n992 ^ x6 ^ 1'b0 ;
  assign n1270 = n207 & ~n1269 ;
  assign n1271 = ~n560 & n1270 ;
  assign n1272 = n843 ^ n618 ^ 1'b0 ;
  assign n1273 = ~n269 & n1272 ;
  assign n1274 = ( x123 & ~n1272 ) | ( x123 & n1273 ) | ( ~n1272 & n1273 ) ;
  assign n1278 = n675 & ~n1110 ;
  assign n1279 = n1278 ^ n404 ^ 1'b0 ;
  assign n1280 = n497 | n1279 ;
  assign n1275 = x86 & ~n614 ;
  assign n1276 = ~n635 & n1275 ;
  assign n1277 = n799 & ~n1276 ;
  assign n1281 = n1280 ^ n1277 ^ 1'b0 ;
  assign n1282 = ( n196 & ~n416 ) | ( n196 & n641 ) | ( ~n416 & n641 ) ;
  assign n1283 = n1282 ^ x36 ^ 1'b0 ;
  assign n1284 = n155 & ~n210 ;
  assign n1285 = n1057 ^ n892 ^ n327 ;
  assign n1286 = n1078 & n1285 ;
  assign n1287 = n1284 & n1286 ;
  assign n1288 = ~n1283 & n1287 ;
  assign n1289 = n531 | n761 ;
  assign n1290 = n1283 & ~n1289 ;
  assign n1291 = n1290 ^ n1060 ^ 1'b0 ;
  assign n1292 = n796 ^ n453 ^ 1'b0 ;
  assign n1293 = n627 ^ n162 ^ 1'b0 ;
  assign n1294 = x30 & n1293 ;
  assign n1295 = n1294 ^ n1283 ^ x105 ;
  assign n1296 = x45 & n1295 ;
  assign n1297 = ~n571 & n1296 ;
  assign n1298 = ( x25 & x90 ) | ( x25 & ~n381 ) | ( x90 & ~n381 ) ;
  assign n1299 = n1298 ^ n1273 ^ n307 ;
  assign n1300 = x53 & ~n1040 ;
  assign n1301 = ~n572 & n1300 ;
  assign n1302 = n1301 ^ n129 ^ 1'b0 ;
  assign n1303 = n456 ^ n199 ^ 1'b0 ;
  assign n1304 = n626 & ~n1303 ;
  assign n1305 = ~n453 & n1304 ;
  assign n1306 = n485 & ~n940 ;
  assign n1307 = x34 & ~n1306 ;
  assign n1308 = n543 & n1307 ;
  assign n1309 = n1308 ^ n1276 ^ n1135 ;
  assign n1313 = n419 ^ n155 ^ 1'b0 ;
  assign n1311 = ( x78 & n184 ) | ( x78 & ~n663 ) | ( n184 & ~n663 ) ;
  assign n1310 = n1020 ^ n874 ^ n211 ;
  assign n1312 = n1311 ^ n1310 ^ 1'b0 ;
  assign n1314 = n1313 ^ n1312 ^ x13 ;
  assign n1315 = x9 & x51 ;
  assign n1316 = ~n644 & n1315 ;
  assign n1317 = n1061 ^ n259 ^ 1'b0 ;
  assign n1318 = ( n657 & n686 ) | ( n657 & n1317 ) | ( n686 & n1317 ) ;
  assign n1319 = n697 & n977 ;
  assign n1320 = n1319 ^ n195 ^ 1'b0 ;
  assign n1321 = n139 & n420 ;
  assign n1322 = n1321 ^ n1280 ^ 1'b0 ;
  assign n1330 = n1290 ^ n946 ^ n916 ;
  assign n1331 = n1330 ^ n1269 ^ x75 ;
  assign n1323 = n548 ^ n245 ^ n196 ;
  assign n1324 = n146 & n1323 ;
  assign n1325 = ~n221 & n616 ;
  assign n1326 = n1325 ^ x5 ^ 1'b0 ;
  assign n1327 = ( x126 & ~n225 ) | ( x126 & n1326 ) | ( ~n225 & n1326 ) ;
  assign n1328 = n1327 ^ n681 ^ 1'b0 ;
  assign n1329 = ~n1324 & n1328 ;
  assign n1332 = n1331 ^ n1329 ^ n913 ;
  assign n1333 = n496 ^ n404 ^ 1'b0 ;
  assign n1334 = n918 & n1333 ;
  assign n1335 = ( ~x9 & n838 ) | ( ~x9 & n1334 ) | ( n838 & n1334 ) ;
  assign n1336 = n167 & ~n269 ;
  assign n1337 = x68 & n1336 ;
  assign n1338 = ~x97 & n1337 ;
  assign n1339 = ~n885 & n1058 ;
  assign n1340 = ~n1069 & n1339 ;
  assign n1341 = n331 & ~n1340 ;
  assign n1342 = n365 & ~n927 ;
  assign n1343 = ~n1104 & n1342 ;
  assign n1346 = x92 & ~n725 ;
  assign n1347 = ~n459 & n1346 ;
  assign n1344 = x93 & ~n1280 ;
  assign n1345 = n1344 ^ n349 ^ 1'b0 ;
  assign n1348 = n1347 ^ n1345 ^ n522 ;
  assign n1349 = ~n1320 & n1348 ;
  assign n1350 = n514 ^ x117 ^ x112 ;
  assign n1351 = ( x55 & n1064 ) | ( x55 & n1350 ) | ( n1064 & n1350 ) ;
  assign n1352 = n1298 ^ n716 ^ 1'b0 ;
  assign n1353 = n429 ^ x10 ^ 1'b0 ;
  assign n1355 = n699 | n983 ;
  assign n1354 = ~n221 & n354 ;
  assign n1356 = n1355 ^ n1354 ^ n214 ;
  assign n1357 = x59 & ~n1356 ;
  assign n1358 = n1353 & n1357 ;
  assign n1359 = n1352 | n1358 ;
  assign n1360 = n328 | n1359 ;
  assign n1361 = n1165 ^ n886 ^ 1'b0 ;
  assign n1362 = n535 | n1361 ;
  assign n1363 = n1360 & n1362 ;
  assign n1364 = n1238 ^ n411 ^ 1'b0 ;
  assign n1365 = x120 & ~n1364 ;
  assign n1366 = n803 ^ n196 ^ 1'b0 ;
  assign n1367 = n138 | n1366 ;
  assign n1368 = n1367 ^ n948 ^ 1'b0 ;
  assign n1369 = n463 ^ n445 ^ n395 ;
  assign n1370 = n1369 ^ n1092 ^ 1'b0 ;
  assign n1371 = n1370 ^ n1240 ^ 1'b0 ;
  assign n1372 = n1371 ^ n561 ^ 1'b0 ;
  assign n1373 = x87 & ~n1372 ;
  assign n1374 = n1373 ^ n303 ^ 1'b0 ;
  assign n1375 = n613 | n1000 ;
  assign n1376 = ( n434 & ~n551 ) | ( n434 & n1375 ) | ( ~n551 & n1375 ) ;
  assign n1377 = n663 & ~n795 ;
  assign n1378 = ~x93 & n1377 ;
  assign n1379 = n1378 ^ n349 ^ 1'b0 ;
  assign n1380 = x39 & n968 ;
  assign n1381 = n1379 & n1380 ;
  assign n1382 = ( n381 & ~n1003 ) | ( n381 & n1378 ) | ( ~n1003 & n1378 ) ;
  assign n1383 = ( n229 & n353 ) | ( n229 & ~n1382 ) | ( n353 & ~n1382 ) ;
  assign n1384 = n1101 ^ n393 ^ 1'b0 ;
  assign n1385 = n182 ^ x56 ^ 1'b0 ;
  assign n1386 = x31 & ~n1385 ;
  assign n1387 = ~n465 & n1259 ;
  assign n1388 = ~n1386 & n1387 ;
  assign n1389 = ~n153 & n421 ;
  assign n1390 = ~n380 & n1389 ;
  assign n1391 = ~n165 & n1390 ;
  assign n1392 = n1388 & n1391 ;
  assign n1393 = n1012 ^ n903 ^ 1'b0 ;
  assign n1394 = n1393 ^ n489 ^ n209 ;
  assign n1395 = n726 | n761 ;
  assign n1396 = n1373 | n1395 ;
  assign n1397 = x52 & ~n988 ;
  assign n1398 = n222 & n1397 ;
  assign n1399 = n649 | n1398 ;
  assign n1400 = n1399 ^ n609 ^ 1'b0 ;
  assign n1401 = n712 & n1400 ;
  assign n1402 = n1401 ^ n541 ^ 1'b0 ;
  assign n1403 = ~n1196 & n1402 ;
  assign n1404 = x120 ^ x73 ^ 1'b0 ;
  assign n1405 = n227 | n1404 ;
  assign n1406 = n1405 ^ n1002 ^ 1'b0 ;
  assign n1407 = x67 & n432 ;
  assign n1408 = ~n791 & n1407 ;
  assign n1409 = n1329 & ~n1408 ;
  assign n1410 = n1406 & n1409 ;
  assign n1411 = n1284 ^ n589 ^ 1'b0 ;
  assign n1412 = n261 & ~n1411 ;
  assign n1413 = x98 & n1412 ;
  assign n1414 = n614 & n1413 ;
  assign n1415 = n1414 ^ x107 ^ x75 ;
  assign n1416 = n1415 ^ n588 ^ 1'b0 ;
  assign n1417 = x67 & ~n1416 ;
  assign n1418 = n696 & n1417 ;
  assign n1419 = x104 & n860 ;
  assign n1420 = n933 | n1419 ;
  assign n1425 = n184 ^ x2 ^ 1'b0 ;
  assign n1426 = n398 | n1347 ;
  assign n1427 = n1425 | n1426 ;
  assign n1421 = n178 & n232 ;
  assign n1422 = n1421 ^ x75 ^ 1'b0 ;
  assign n1423 = ( n203 & n250 ) | ( n203 & n1422 ) | ( n250 & n1422 ) ;
  assign n1424 = ( n660 & n773 ) | ( n660 & n1423 ) | ( n773 & n1423 ) ;
  assign n1428 = n1427 ^ n1424 ^ 1'b0 ;
  assign n1429 = n145 | n916 ;
  assign n1430 = n509 & ~n1429 ;
  assign n1431 = ( ~x34 & x46 ) | ( ~x34 & x84 ) | ( x46 & x84 ) ;
  assign n1432 = n1431 ^ n1312 ^ 1'b0 ;
  assign n1433 = n1430 | n1432 ;
  assign n1434 = n1424 ^ x6 ^ 1'b0 ;
  assign n1435 = ~n1244 & n1262 ;
  assign n1437 = n463 & ~n748 ;
  assign n1438 = n1437 ^ n393 ^ 1'b0 ;
  assign n1436 = n344 ^ x107 ^ 1'b0 ;
  assign n1439 = n1438 ^ n1436 ^ 1'b0 ;
  assign n1440 = ~n1074 & n1439 ;
  assign n1441 = n1192 ^ n521 ^ 1'b0 ;
  assign n1442 = n462 ^ x21 ^ 1'b0 ;
  assign n1444 = n650 ^ n410 ^ n286 ;
  assign n1445 = ( ~n181 & n1170 ) | ( ~n181 & n1444 ) | ( n1170 & n1444 ) ;
  assign n1446 = x3 & n271 ;
  assign n1447 = n1445 & n1446 ;
  assign n1443 = ~n164 & n650 ;
  assign n1448 = n1447 ^ n1443 ^ 1'b0 ;
  assign n1449 = n1078 ^ n909 ^ 1'b0 ;
  assign n1455 = n430 & ~n715 ;
  assign n1450 = n967 ^ n285 ^ 1'b0 ;
  assign n1451 = n1216 ^ n828 ^ 1'b0 ;
  assign n1452 = ( n756 & n1450 ) | ( n756 & ~n1451 ) | ( n1450 & ~n1451 ) ;
  assign n1453 = n1285 & n1452 ;
  assign n1454 = ~n469 & n1453 ;
  assign n1456 = n1455 ^ n1454 ^ 1'b0 ;
  assign n1459 = n233 ^ x13 ^ x7 ;
  assign n1457 = n756 & n816 ;
  assign n1458 = n1457 ^ n1129 ^ 1'b0 ;
  assign n1460 = n1459 ^ n1458 ^ n218 ;
  assign n1461 = n298 | n1460 ;
  assign n1462 = ( n941 & n1456 ) | ( n941 & n1461 ) | ( n1456 & n1461 ) ;
  assign n1463 = n1027 ^ n776 ^ 1'b0 ;
  assign n1464 = n1463 ^ n614 ^ 1'b0 ;
  assign n1465 = n935 & n1464 ;
  assign n1466 = n1288 ^ n880 ^ n381 ;
  assign n1467 = n1466 ^ n844 ^ n469 ;
  assign n1468 = x88 & x127 ;
  assign n1469 = n1468 ^ n723 ^ 1'b0 ;
  assign n1470 = ( n184 & ~n258 ) | ( n184 & n1469 ) | ( ~n258 & n1469 ) ;
  assign n1471 = n1470 ^ x17 ^ 1'b0 ;
  assign n1472 = n1012 | n1471 ;
  assign n1475 = n1457 ^ n531 ^ n387 ;
  assign n1473 = ~n1222 & n1417 ;
  assign n1474 = n1436 & n1473 ;
  assign n1476 = n1475 ^ n1474 ^ 1'b0 ;
  assign n1477 = ( x33 & ~x42 ) | ( x33 & n1244 ) | ( ~x42 & n1244 ) ;
  assign n1478 = n1477 ^ n1252 ^ n879 ;
  assign n1479 = x29 & ~n1478 ;
  assign n1480 = n1479 ^ n1051 ^ 1'b0 ;
  assign n1481 = n1023 ^ n134 ^ 1'b0 ;
  assign n1482 = ~n664 & n713 ;
  assign n1483 = ~n418 & n1482 ;
  assign n1484 = n1483 ^ x33 ^ 1'b0 ;
  assign n1485 = n807 | n1484 ;
  assign n1486 = n447 & ~n603 ;
  assign n1487 = ~n205 & n1486 ;
  assign n1488 = n1036 & ~n1487 ;
  assign n1489 = ~n1129 & n1488 ;
  assign n1490 = n1370 ^ n328 ^ 1'b0 ;
  assign n1491 = ~n1284 & n1490 ;
  assign n1492 = n134 | n1459 ;
  assign n1493 = n1492 ^ n330 ^ 1'b0 ;
  assign n1494 = x80 & ~n1256 ;
  assign n1495 = ~n1493 & n1494 ;
  assign n1496 = n1252 | n1495 ;
  assign n1497 = n383 ^ x80 ^ 1'b0 ;
  assign n1498 = n995 | n1497 ;
  assign n1499 = n668 ^ n281 ^ x104 ;
  assign n1500 = n731 | n1499 ;
  assign n1501 = n307 | n1500 ;
  assign n1502 = n1501 ^ x91 ^ 1'b0 ;
  assign n1503 = n1502 ^ n229 ^ 1'b0 ;
  assign n1504 = ~n223 & n825 ;
  assign n1505 = n1504 ^ n847 ^ 1'b0 ;
  assign n1506 = n1505 ^ n746 ^ 1'b0 ;
  assign n1507 = ~n1036 & n1152 ;
  assign n1511 = n1183 | n1226 ;
  assign n1512 = ( x75 & n646 ) | ( x75 & n1511 ) | ( n646 & n1511 ) ;
  assign n1508 = ~n186 & n725 ;
  assign n1509 = n1508 ^ n997 ^ 1'b0 ;
  assign n1510 = n852 & ~n1509 ;
  assign n1513 = n1512 ^ n1510 ^ 1'b0 ;
  assign n1514 = n469 ^ n362 ^ x91 ;
  assign n1515 = n1419 | n1514 ;
  assign n1516 = x92 & ~n146 ;
  assign n1517 = n319 | n1516 ;
  assign n1518 = n1517 ^ n267 ^ x42 ;
  assign n1519 = n286 | n1120 ;
  assign n1520 = x76 & x103 ;
  assign n1521 = n393 & n1520 ;
  assign n1522 = n1521 ^ n867 ^ 1'b0 ;
  assign n1523 = ( n802 & n1120 ) | ( n802 & ~n1522 ) | ( n1120 & ~n1522 ) ;
  assign n1524 = n1523 ^ n1502 ^ n1403 ;
  assign n1525 = n1020 ^ x85 ^ 1'b0 ;
  assign n1526 = n746 ^ n305 ^ 1'b0 ;
  assign n1527 = n465 | n1526 ;
  assign n1528 = n843 ^ n491 ^ 1'b0 ;
  assign n1529 = n1304 ^ n307 ^ 1'b0 ;
  assign n1534 = n1087 ^ n489 ^ x26 ;
  assign n1530 = n744 & ~n886 ;
  assign n1531 = n1530 ^ n1371 ^ 1'b0 ;
  assign n1532 = n1298 ^ n744 ^ 1'b0 ;
  assign n1533 = n1531 | n1532 ;
  assign n1535 = n1534 ^ n1533 ^ 1'b0 ;
  assign n1536 = n533 | n1306 ;
  assign n1537 = n271 & ~n1536 ;
  assign n1541 = n663 & n1173 ;
  assign n1542 = n380 & n1541 ;
  assign n1538 = n1022 | n1240 ;
  assign n1539 = ~n415 & n787 ;
  assign n1540 = n1538 & ~n1539 ;
  assign n1543 = n1542 ^ n1540 ^ 1'b0 ;
  assign n1544 = n670 | n779 ;
  assign n1545 = ( n161 & n1123 ) | ( n161 & n1534 ) | ( n1123 & n1534 ) ;
  assign n1546 = n1545 ^ x116 ^ 1'b0 ;
  assign n1547 = n704 | n1546 ;
  assign n1548 = n281 & ~n1547 ;
  assign n1549 = n608 | n1451 ;
  assign n1550 = n1549 ^ x16 ^ 1'b0 ;
  assign n1551 = ~n1548 & n1550 ;
  assign n1552 = ~n1544 & n1551 ;
  assign n1553 = n614 ^ n510 ^ 1'b0 ;
  assign n1554 = n1552 | n1553 ;
  assign n1555 = n1488 ^ n463 ^ x91 ;
  assign n1557 = n536 ^ n168 ^ 1'b0 ;
  assign n1558 = n254 & ~n1557 ;
  assign n1559 = n735 & n1558 ;
  assign n1560 = n725 & n1559 ;
  assign n1556 = n1170 ^ n1116 ^ 1'b0 ;
  assign n1561 = n1560 ^ n1556 ^ n510 ;
  assign n1562 = n1272 ^ n357 ^ 1'b0 ;
  assign n1563 = n1369 & ~n1562 ;
  assign n1564 = n401 & n1563 ;
  assign n1565 = n1564 ^ n1061 ^ n1036 ;
  assign n1566 = n424 ^ n390 ^ 1'b0 ;
  assign n1567 = n1565 & n1566 ;
  assign n1568 = n1440 ^ n340 ^ 1'b0 ;
  assign n1569 = n1567 & ~n1568 ;
  assign n1570 = ~n1410 & n1569 ;
  assign n1571 = ~x84 & n1570 ;
  assign n1572 = n271 & ~n1358 ;
  assign n1573 = ~n1420 & n1572 ;
  assign n1574 = n456 | n551 ;
  assign n1575 = n1574 ^ n701 ^ 1'b0 ;
  assign n1576 = n1575 ^ n343 ^ x62 ;
  assign n1577 = n1576 ^ n157 ^ 1'b0 ;
  assign n1586 = ( n201 & n248 ) | ( n201 & ~n897 ) | ( n248 & ~n897 ) ;
  assign n1587 = n874 & n1586 ;
  assign n1579 = x117 & ~n535 ;
  assign n1580 = n1579 ^ n1445 ^ 1'b0 ;
  assign n1581 = n337 & ~n1580 ;
  assign n1582 = n1581 ^ n1256 ^ n508 ;
  assign n1583 = n493 & ~n1582 ;
  assign n1584 = ~n1194 & n1583 ;
  assign n1585 = n1584 ^ n866 ^ n303 ;
  assign n1588 = n1587 ^ n1585 ^ 1'b0 ;
  assign n1578 = ~n843 & n877 ;
  assign n1589 = n1588 ^ n1578 ^ 1'b0 ;
  assign n1590 = n1034 ^ x49 ^ 1'b0 ;
  assign n1591 = n298 | n1590 ;
  assign n1592 = x69 & n377 ;
  assign n1593 = ~n688 & n1592 ;
  assign n1594 = ( ~n136 & n494 ) | ( ~n136 & n1593 ) | ( n494 & n1593 ) ;
  assign n1595 = ( x3 & ~n1228 ) | ( x3 & n1594 ) | ( ~n1228 & n1594 ) ;
  assign n1596 = n1591 | n1595 ;
  assign n1597 = n571 & ~n967 ;
  assign n1598 = n1597 ^ n1108 ^ 1'b0 ;
  assign n1599 = ~n406 & n1598 ;
  assign n1600 = ~n573 & n1599 ;
  assign n1601 = n398 ^ n267 ^ 1'b0 ;
  assign n1602 = ~n190 & n1601 ;
  assign n1603 = n653 ^ x113 ^ 1'b0 ;
  assign n1604 = ~n397 & n855 ;
  assign n1605 = n1604 ^ n1029 ^ 1'b0 ;
  assign n1608 = n613 ^ n600 ^ 1'b0 ;
  assign n1606 = n1170 | n1282 ;
  assign n1607 = n1606 ^ n260 ^ 1'b0 ;
  assign n1609 = n1608 ^ n1607 ^ 1'b0 ;
  assign n1610 = n606 | n1609 ;
  assign n1611 = n1610 ^ n1057 ^ 1'b0 ;
  assign n1612 = n1611 ^ n1473 ^ x63 ;
  assign n1613 = n1312 ^ n1010 ^ 1'b0 ;
  assign n1614 = ( n915 & n1135 ) | ( n915 & n1552 ) | ( n1135 & n1552 ) ;
  assign n1615 = x6 & n173 ;
  assign n1616 = n1615 ^ n711 ^ 1'b0 ;
  assign n1617 = n1262 & n1616 ;
  assign n1618 = ~n1284 & n1596 ;
  assign n1619 = n1489 ^ n888 ^ 1'b0 ;
  assign n1620 = n1475 ^ n491 ^ 1'b0 ;
  assign n1621 = x61 & n1620 ;
  assign n1622 = n1621 ^ n881 ^ 1'b0 ;
  assign n1623 = n264 | n563 ;
  assign n1624 = n1467 ^ n778 ^ 1'b0 ;
  assign n1625 = n1623 | n1624 ;
  assign n1626 = ~n1483 & n1625 ;
  assign n1627 = x39 & n1438 ;
  assign n1628 = n308 & n1627 ;
  assign n1629 = n1628 ^ n805 ^ 1'b0 ;
  assign n1630 = n584 ^ n214 ^ 1'b0 ;
  assign n1631 = n399 & n1630 ;
  assign n1632 = n1045 & ~n1631 ;
  assign n1633 = ( ~x35 & x114 ) | ( ~x35 & n261 ) | ( x114 & n261 ) ;
  assign n1634 = n1633 ^ n1331 ^ 1'b0 ;
  assign n1635 = n1376 ^ n530 ^ 1'b0 ;
  assign n1636 = ~n1393 & n1635 ;
  assign n1637 = ( n986 & n1102 ) | ( n986 & ~n1322 ) | ( n1102 & ~n1322 ) ;
  assign n1638 = n143 | n1637 ;
  assign n1639 = n1638 ^ n319 ^ 1'b0 ;
  assign n1640 = n347 ^ x118 ^ 1'b0 ;
  assign n1641 = n631 | n1640 ;
  assign n1642 = n1641 ^ n366 ^ 1'b0 ;
  assign n1643 = n710 ^ n629 ^ n413 ;
  assign n1644 = n1643 ^ n261 ^ 1'b0 ;
  assign n1645 = n1644 ^ n1284 ^ n134 ;
  assign n1650 = n345 & n791 ;
  assign n1651 = n1327 & n1650 ;
  assign n1646 = n515 ^ n154 ^ 1'b0 ;
  assign n1647 = n246 & n1646 ;
  assign n1648 = ( n850 & n911 ) | ( n850 & n1647 ) | ( n911 & n1647 ) ;
  assign n1649 = ( n380 & n990 ) | ( n380 & n1648 ) | ( n990 & n1648 ) ;
  assign n1652 = n1651 ^ n1649 ^ n672 ;
  assign n1655 = n737 ^ x66 ^ 1'b0 ;
  assign n1653 = ~x2 & x125 ;
  assign n1654 = n1653 ^ x109 ^ 1'b0 ;
  assign n1656 = n1655 ^ n1654 ^ n721 ;
  assign n1657 = n1457 ^ n540 ^ 1'b0 ;
  assign n1658 = n971 ^ n316 ^ 1'b0 ;
  assign n1659 = n201 & ~n447 ;
  assign n1660 = n1659 ^ n194 ^ 1'b0 ;
  assign n1661 = n1425 & ~n1660 ;
  assign n1662 = n1661 ^ n782 ^ 1'b0 ;
  assign n1663 = n620 | n1662 ;
  assign n1664 = n1663 ^ n1392 ^ n1257 ;
  assign n1665 = n1292 ^ n850 ^ 1'b0 ;
  assign n1666 = n1665 ^ n1168 ^ n805 ;
  assign n1667 = n1666 ^ n1091 ^ 1'b0 ;
  assign n1668 = n803 ^ x19 ^ 1'b0 ;
  assign n1669 = n931 & ~n1668 ;
  assign n1670 = x23 & ~n1512 ;
  assign n1671 = ~n1669 & n1670 ;
  assign n1672 = x116 & ~n760 ;
  assign n1673 = x0 & n1672 ;
  assign n1674 = n836 ^ n196 ^ x46 ;
  assign n1675 = ~n296 & n580 ;
  assign n1676 = n1675 ^ n1209 ^ 1'b0 ;
  assign n1677 = n1517 & n1676 ;
  assign n1678 = n1674 | n1677 ;
  assign n1679 = n1666 ^ n536 ^ n473 ;
  assign n1680 = n1027 ^ n771 ^ 1'b0 ;
  assign n1681 = ~n421 & n1633 ;
  assign n1682 = n285 & n1681 ;
  assign n1683 = n250 ^ x33 ^ 1'b0 ;
  assign n1684 = ( n811 & n990 ) | ( n811 & ~n1683 ) | ( n990 & ~n1683 ) ;
  assign n1685 = ~n1682 & n1684 ;
  assign n1686 = n573 ^ n372 ^ 1'b0 ;
  assign n1687 = x64 & n1686 ;
  assign n1688 = n1687 ^ n1106 ^ 1'b0 ;
  assign n1689 = ~n510 & n1688 ;
  assign n1690 = ( n554 & ~n793 ) | ( n554 & n1148 ) | ( ~n793 & n1148 ) ;
  assign n1691 = x93 & ~n335 ;
  assign n1692 = n1691 ^ n1615 ^ 1'b0 ;
  assign n1693 = n477 ^ n295 ^ 1'b0 ;
  assign n1694 = n205 & ~n1693 ;
  assign n1695 = n221 & ~n1694 ;
  assign n1696 = ( n677 & n1629 ) | ( n677 & ~n1695 ) | ( n1629 & ~n1695 ) ;
  assign n1697 = ( ~n834 & n882 ) | ( ~n834 & n1290 ) | ( n882 & n1290 ) ;
  assign n1700 = n1027 ^ n824 ^ n169 ;
  assign n1698 = x29 & n142 ;
  assign n1699 = n1698 ^ n1212 ^ 1'b0 ;
  assign n1701 = n1700 ^ n1699 ^ 1'b0 ;
  assign n1702 = x70 & n1701 ;
  assign n1703 = n1528 ^ n770 ^ n550 ;
  assign n1704 = ( n531 & n744 ) | ( n531 & n1510 ) | ( n744 & n1510 ) ;
  assign n1708 = n603 ^ n201 ^ x87 ;
  assign n1709 = n1708 ^ n560 ^ x74 ;
  assign n1705 = n1008 | n1290 ;
  assign n1706 = n1705 ^ n1154 ^ 1'b0 ;
  assign n1707 = x78 & ~n1706 ;
  assign n1710 = n1709 ^ n1707 ^ 1'b0 ;
  assign n1711 = n1689 ^ x102 ^ 1'b0 ;
  assign n1712 = n278 & n1711 ;
  assign n1713 = n1712 ^ n1696 ^ n1375 ;
  assign n1714 = n1295 ^ n893 ^ n804 ;
  assign n1715 = n591 & n1714 ;
  assign n1716 = n323 ^ x64 ^ 1'b0 ;
  assign n1717 = ~n1459 & n1716 ;
  assign n1718 = ~n1715 & n1717 ;
  assign n1720 = ( ~n627 & n684 ) | ( ~n627 & n1579 ) | ( n684 & n1579 ) ;
  assign n1719 = ~x10 & n1058 ;
  assign n1721 = n1720 ^ n1719 ^ 1'b0 ;
  assign n1722 = n923 | n1721 ;
  assign n1723 = n1326 | n1431 ;
  assign n1724 = n716 ^ x55 ^ 1'b0 ;
  assign n1725 = n1723 & n1724 ;
  assign n1726 = n1722 & ~n1725 ;
  assign n1727 = ( n387 & n704 ) | ( n387 & n916 ) | ( n704 & n916 ) ;
  assign n1728 = n995 ^ n214 ^ 1'b0 ;
  assign n1729 = n1107 ^ x78 ^ 1'b0 ;
  assign n1730 = n1729 ^ n1051 ^ 1'b0 ;
  assign n1731 = n1728 & n1730 ;
  assign n1732 = n1556 ^ n1348 ^ n278 ;
  assign n1733 = n517 ^ n322 ^ n257 ;
  assign n1734 = n625 & n1733 ;
  assign n1735 = n1334 & n1734 ;
  assign n1736 = ~n232 & n1735 ;
  assign n1737 = n974 & ~n1736 ;
  assign n1738 = n1737 ^ n901 ^ 1'b0 ;
  assign n1739 = n1738 ^ n1295 ^ n493 ;
  assign n1740 = n1571 ^ n1268 ^ x105 ;
  assign n1742 = x113 & n390 ;
  assign n1743 = n1742 ^ n430 ^ 1'b0 ;
  assign n1744 = n459 & ~n1743 ;
  assign n1745 = n1744 ^ n960 ^ 1'b0 ;
  assign n1746 = n254 & n1745 ;
  assign n1747 = n1310 & n1746 ;
  assign n1741 = n456 & ~n1323 ;
  assign n1748 = n1747 ^ n1741 ^ 1'b0 ;
  assign n1749 = n357 | n922 ;
  assign n1750 = n1749 ^ n1613 ^ 1'b0 ;
  assign n1751 = n1748 | n1750 ;
  assign n1752 = ( n740 & n1242 ) | ( n740 & ~n1751 ) | ( n1242 & ~n1751 ) ;
  assign n1753 = ~n617 & n697 ;
  assign n1754 = n1162 & n1753 ;
  assign n1755 = n1754 ^ n341 ^ 1'b0 ;
  assign n1756 = ~n982 & n1755 ;
  assign n1757 = ~n1424 & n1756 ;
  assign n1758 = n1757 ^ n431 ^ 1'b0 ;
  assign n1759 = n1324 ^ n805 ^ n541 ;
  assign n1760 = x51 & ~n148 ;
  assign n1761 = x68 & n1760 ;
  assign n1762 = n1761 ^ n490 ^ 1'b0 ;
  assign n1763 = n205 & ~n1762 ;
  assign n1764 = n1763 ^ n411 ^ n207 ;
  assign n1765 = n1163 | n1764 ;
  assign n1766 = n515 & ~n1765 ;
  assign n1767 = n1766 ^ n1221 ^ 1'b0 ;
  assign n1770 = ( x0 & n456 ) | ( x0 & n1425 ) | ( n456 & n1425 ) ;
  assign n1768 = x39 & n1445 ;
  assign n1769 = x86 & n1768 ;
  assign n1771 = n1770 ^ n1769 ^ 1'b0 ;
  assign n1772 = ~n1354 & n1771 ;
  assign n1773 = n1186 ^ n967 ^ 1'b0 ;
  assign n1774 = n758 ^ x2 ^ 1'b0 ;
  assign n1775 = n1220 ^ n997 ^ 1'b0 ;
  assign n1776 = n1774 | n1775 ;
  assign n1777 = n310 & n1776 ;
  assign n1778 = n1057 & ~n1457 ;
  assign n1779 = ( n298 & ~n467 ) | ( n298 & n487 ) | ( ~n467 & n487 ) ;
  assign n1780 = n1778 & ~n1779 ;
  assign n1781 = n1777 & n1780 ;
  assign n1785 = n370 ^ x4 ^ 1'b0 ;
  assign n1786 = x1 | n1785 ;
  assign n1787 = n390 | n1786 ;
  assign n1782 = n152 & ~n672 ;
  assign n1783 = n1014 ^ n937 ^ n485 ;
  assign n1784 = n1782 & n1783 ;
  assign n1788 = n1787 ^ n1784 ^ x2 ;
  assign n1789 = n998 ^ n606 ^ n560 ;
  assign n1790 = n419 & ~n423 ;
  assign n1791 = ~n1789 & n1790 ;
  assign n1793 = n1297 ^ n1201 ^ 1'b0 ;
  assign n1792 = n236 | n557 ;
  assign n1794 = n1793 ^ n1792 ^ 1'b0 ;
  assign n1795 = n232 | n1053 ;
  assign n1796 = ( n250 & n925 ) | ( n250 & ~n1499 ) | ( n925 & ~n1499 ) ;
  assign n1797 = n1796 ^ n1610 ^ 1'b0 ;
  assign n1798 = n1550 ^ x61 ^ 1'b0 ;
  assign n1800 = ( ~x70 & n798 ) | ( ~x70 & n815 ) | ( n798 & n815 ) ;
  assign n1799 = ( ~n480 & n525 ) | ( ~n480 & n1254 ) | ( n525 & n1254 ) ;
  assign n1801 = n1800 ^ n1799 ^ 1'b0 ;
  assign n1802 = n1798 & n1801 ;
  assign n1803 = ( n155 & ~n285 ) | ( n155 & n415 ) | ( ~n285 & n415 ) ;
  assign n1804 = n1306 & ~n1803 ;
  assign n1805 = n1804 ^ n1203 ^ 1'b0 ;
  assign n1806 = n1805 ^ n1259 ^ 1'b0 ;
  assign n1807 = n449 | n836 ;
  assign n1808 = n1807 ^ n1256 ^ 1'b0 ;
  assign n1809 = ( n1027 & ~n1469 ) | ( n1027 & n1808 ) | ( ~n1469 & n1808 ) ;
  assign n1810 = n672 ^ n403 ^ 1'b0 ;
  assign n1813 = ~n293 & n1004 ;
  assign n1814 = ~n242 & n1813 ;
  assign n1815 = n1814 ^ n960 ^ n415 ;
  assign n1811 = n855 ^ n546 ^ 1'b0 ;
  assign n1812 = ( n591 & n1071 ) | ( n591 & ~n1811 ) | ( n1071 & ~n1811 ) ;
  assign n1816 = n1815 ^ n1812 ^ 1'b0 ;
  assign n1817 = n1810 | n1816 ;
  assign n1818 = ( ~n843 & n1809 ) | ( ~n843 & n1817 ) | ( n1809 & n1817 ) ;
  assign n1819 = n931 ^ n898 ^ 1'b0 ;
  assign n1820 = ~n1659 & n1819 ;
  assign n1821 = n243 ^ n133 ^ 1'b0 ;
  assign n1822 = ~n606 & n1821 ;
  assign n1823 = n456 | n917 ;
  assign n1824 = n1822 & n1823 ;
  assign n1825 = n1824 ^ n882 ^ 1'b0 ;
  assign n1826 = ( n1055 & n1490 ) | ( n1055 & ~n1825 ) | ( n1490 & ~n1825 ) ;
  assign n1827 = ~n1107 & n1826 ;
  assign n1828 = ~n1473 & n1827 ;
  assign n1829 = ( n163 & n657 ) | ( n163 & n867 ) | ( n657 & n867 ) ;
  assign n1830 = n337 & n530 ;
  assign n1831 = n331 & n1830 ;
  assign n1832 = n1831 ^ n1605 ^ n879 ;
  assign n1833 = n1130 ^ n825 ^ 1'b0 ;
  assign n1834 = ~n1613 & n1833 ;
  assign n1835 = n330 & n1331 ;
  assign n1836 = n1835 ^ n1470 ^ 1'b0 ;
  assign n1837 = n986 & n1798 ;
  assign n1838 = n918 & n1313 ;
  assign n1839 = ~n920 & n1838 ;
  assign n1840 = n1254 & n1839 ;
  assign n1841 = n1840 ^ n1729 ^ x39 ;
  assign n1842 = n1841 ^ n234 ^ 1'b0 ;
  assign n1843 = ( ~x116 & n419 ) | ( ~x116 & n808 ) | ( n419 & n808 ) ;
  assign n1846 = ~n152 & n1525 ;
  assign n1844 = n553 & ~n859 ;
  assign n1845 = n1844 ^ n1831 ^ 1'b0 ;
  assign n1847 = n1846 ^ n1845 ^ 1'b0 ;
  assign n1848 = ~n1843 & n1847 ;
  assign n1849 = n1487 ^ n1388 ^ 1'b0 ;
  assign n1850 = n194 & n1849 ;
  assign n1851 = n1425 ^ n458 ^ 1'b0 ;
  assign n1852 = n1851 ^ n232 ^ 1'b0 ;
  assign n1853 = n154 | n1852 ;
  assign n1854 = n1853 ^ n517 ^ x88 ;
  assign n1855 = n1854 ^ n1510 ^ 1'b0 ;
  assign n1856 = n1608 ^ n1396 ^ 1'b0 ;
  assign n1857 = n573 & ~n1249 ;
  assign n1858 = n214 & n1857 ;
  assign n1859 = n391 | n1858 ;
  assign n1860 = n1856 | n1859 ;
  assign n1861 = ~x10 & n1756 ;
  assign n1862 = ~x52 & n382 ;
  assign n1863 = n1862 ^ n822 ^ 1'b0 ;
  assign n1865 = n1008 ^ n343 ^ 1'b0 ;
  assign n1864 = n357 ^ n269 ^ n152 ;
  assign n1866 = n1865 ^ n1864 ^ 1'b0 ;
  assign n1867 = n201 | n1866 ;
  assign n1868 = n709 & ~n1311 ;
  assign n1869 = n1868 ^ n732 ^ 1'b0 ;
  assign n1870 = n730 & n1869 ;
  assign n1871 = n1867 & n1870 ;
  assign n1872 = n1376 ^ n715 ^ 1'b0 ;
  assign n1873 = ~n1871 & n1872 ;
  assign n1874 = ~n386 & n1216 ;
  assign n1875 = n1874 ^ x1 ^ 1'b0 ;
  assign n1876 = n1525 & ~n1875 ;
  assign n1877 = n1075 & n1876 ;
  assign n1878 = ~x94 & n1877 ;
  assign n1881 = n1564 ^ n529 ^ 1'b0 ;
  assign n1879 = ~n434 & n501 ;
  assign n1880 = n1879 ^ n1325 ^ 1'b0 ;
  assign n1882 = n1881 ^ n1880 ^ 1'b0 ;
  assign n1883 = n1412 & ~n1882 ;
  assign n1884 = ~n1465 & n1883 ;
  assign n1886 = ~n421 & n905 ;
  assign n1887 = ~n723 & n1886 ;
  assign n1885 = x21 & ~n1531 ;
  assign n1888 = n1887 ^ n1885 ^ 1'b0 ;
  assign n1889 = x120 & n522 ;
  assign n1890 = ~n1888 & n1889 ;
  assign n1891 = n1408 ^ x67 ^ 1'b0 ;
  assign n1892 = n1284 | n1891 ;
  assign n1893 = n1808 ^ n410 ^ x29 ;
  assign n1894 = n1893 ^ n1079 ^ n911 ;
  assign n1895 = ( n575 & n677 ) | ( n575 & ~n1894 ) | ( n677 & ~n1894 ) ;
  assign n1898 = ( ~n471 & n582 ) | ( ~n471 & n1071 ) | ( n582 & n1071 ) ;
  assign n1896 = n536 ^ n307 ^ 1'b0 ;
  assign n1897 = n1412 & ~n1896 ;
  assign n1899 = n1898 ^ n1897 ^ n413 ;
  assign n1900 = n1899 ^ n1679 ^ n461 ;
  assign n1901 = x13 | n358 ;
  assign n1902 = n1901 ^ n663 ^ 1'b0 ;
  assign n1903 = n451 ^ n368 ^ n334 ;
  assign n1904 = n1903 ^ n688 ^ 1'b0 ;
  assign n1905 = n1904 ^ n1538 ^ n1525 ;
  assign n1906 = ( ~n1165 & n1902 ) | ( ~n1165 & n1905 ) | ( n1902 & n1905 ) ;
  assign n1907 = n178 ^ x30 ^ 1'b0 ;
  assign n1908 = n227 & ~n1843 ;
  assign n1909 = n1907 & ~n1908 ;
  assign n1910 = n1909 ^ x109 ^ 1'b0 ;
  assign n1911 = n1020 ^ x91 ^ 1'b0 ;
  assign n1912 = n1911 ^ n1093 ^ 1'b0 ;
  assign n1913 = x3 & n1912 ;
  assign n1914 = n1913 ^ n971 ^ n630 ;
  assign n1915 = n1254 | n1584 ;
  assign n1916 = n1915 ^ n522 ^ 1'b0 ;
  assign n1917 = n1914 & n1916 ;
  assign n1918 = n1582 ^ n936 ^ 1'b0 ;
  assign n1919 = n1918 ^ n934 ^ 1'b0 ;
  assign n1920 = x103 & n771 ;
  assign n1921 = ( n368 & n1733 ) | ( n368 & ~n1815 ) | ( n1733 & ~n1815 ) ;
  assign n1922 = n726 ^ x121 ^ 1'b0 ;
  assign n1923 = n1660 | n1922 ;
  assign n1924 = n1923 ^ n938 ^ n768 ;
  assign n1925 = n1921 & n1924 ;
  assign n1926 = x95 & ~n554 ;
  assign n1927 = n1926 ^ n742 ^ 1'b0 ;
  assign n1928 = n1927 ^ n1714 ^ n240 ;
  assign n1929 = n390 & n1118 ;
  assign n1930 = n1929 ^ n1865 ^ n1524 ;
  assign n1935 = n751 & ~n1107 ;
  assign n1936 = n1935 ^ n1268 ^ n322 ;
  assign n1933 = ( n475 & n723 ) | ( n475 & ~n1785 ) | ( n723 & ~n1785 ) ;
  assign n1934 = ~n1040 & n1933 ;
  assign n1931 = n1839 ^ n622 ^ 1'b0 ;
  assign n1932 = n1931 ^ n1199 ^ 1'b0 ;
  assign n1937 = n1936 ^ n1934 ^ n1932 ;
  assign n1938 = n1937 ^ n1340 ^ x86 ;
  assign n1939 = n295 ^ x19 ^ 1'b0 ;
  assign n1942 = n425 & n770 ;
  assign n1940 = ( n868 & n1065 ) | ( n868 & ~n1087 ) | ( n1065 & ~n1087 ) ;
  assign n1941 = n246 & ~n1940 ;
  assign n1943 = n1942 ^ n1941 ^ 1'b0 ;
  assign n1950 = ~n175 & n546 ;
  assign n1951 = n1950 ^ n1427 ^ 1'b0 ;
  assign n1952 = n836 | n1951 ;
  assign n1945 = n350 | n693 ;
  assign n1946 = n597 & ~n1945 ;
  assign n1944 = n823 & n1076 ;
  assign n1947 = n1946 ^ n1944 ^ 1'b0 ;
  assign n1948 = n1947 ^ n914 ^ 1'b0 ;
  assign n1949 = x103 & ~n1948 ;
  assign n1953 = n1952 ^ n1949 ^ n260 ;
  assign n1957 = n210 & n793 ;
  assign n1958 = n1487 & n1957 ;
  assign n1954 = n361 | n1331 ;
  assign n1955 = n1954 ^ n182 ^ 1'b0 ;
  assign n1956 = n1955 ^ n384 ^ n340 ;
  assign n1959 = n1958 ^ n1956 ^ 1'b0 ;
  assign n1960 = ( n307 & n608 ) | ( n307 & ~n749 ) | ( n608 & ~n749 ) ;
  assign n1961 = n1960 ^ n1280 ^ 1'b0 ;
  assign n1962 = n1588 & n1961 ;
  assign n1971 = n363 | n731 ;
  assign n1972 = n484 | n1971 ;
  assign n1973 = ( n611 & n1694 ) | ( n611 & ~n1972 ) | ( n1694 & ~n1972 ) ;
  assign n1963 = n1743 ^ n803 ^ 1'b0 ;
  assign n1964 = ~n1183 & n1963 ;
  assign n1965 = ( ~n201 & n704 ) | ( ~n201 & n1913 ) | ( n704 & n1913 ) ;
  assign n1966 = n1964 & ~n1965 ;
  assign n1967 = ~n1218 & n1966 ;
  assign n1968 = n1967 ^ n1376 ^ 1'b0 ;
  assign n1969 = n1511 | n1968 ;
  assign n1970 = ( ~n872 & n1205 ) | ( ~n872 & n1969 ) | ( n1205 & n1969 ) ;
  assign n1974 = n1973 ^ n1970 ^ n888 ;
  assign n1976 = n786 ^ x93 ^ x59 ;
  assign n1977 = n1669 & ~n1976 ;
  assign n1975 = n1595 & ~n1840 ;
  assign n1978 = n1977 ^ n1975 ^ 1'b0 ;
  assign n1979 = ( n1011 & ~n1406 ) | ( n1011 & n1978 ) | ( ~n1406 & n1978 ) ;
  assign n1980 = n923 | n1923 ;
  assign n1981 = n1980 ^ n903 ^ 1'b0 ;
  assign n1982 = n917 | n1188 ;
  assign n1983 = ~n1629 & n1982 ;
  assign n1984 = n191 & ~n1475 ;
  assign n1985 = n756 ^ n293 ^ n219 ;
  assign n1986 = n1985 ^ n298 ^ 1'b0 ;
  assign n1987 = n1986 ^ n1836 ^ 1'b0 ;
  assign n1988 = n1244 & n1987 ;
  assign n1992 = n1240 | n1398 ;
  assign n1989 = x101 & n562 ;
  assign n1990 = n1989 ^ x122 ^ 1'b0 ;
  assign n1991 = n1637 | n1990 ;
  assign n1993 = n1992 ^ n1991 ^ 1'b0 ;
  assign n1995 = ( x44 & n303 ) | ( x44 & n555 ) | ( n303 & n555 ) ;
  assign n1994 = n1280 ^ n494 ^ n339 ;
  assign n1996 = n1995 ^ n1994 ^ n1691 ;
  assign n2004 = n278 ^ x104 ^ 1'b0 ;
  assign n2005 = x76 & n2004 ;
  assign n2006 = n2005 ^ n1809 ^ 1'b0 ;
  assign n1998 = n740 ^ n447 ^ x1 ;
  assign n1997 = n1238 ^ n393 ^ 1'b0 ;
  assign n1999 = n1998 ^ n1997 ^ 1'b0 ;
  assign n2000 = n569 & ~n822 ;
  assign n2001 = n433 ^ n177 ^ 1'b0 ;
  assign n2002 = n2000 | n2001 ;
  assign n2003 = n1999 | n2002 ;
  assign n2007 = n2006 ^ n2003 ^ 1'b0 ;
  assign n2008 = ~n257 & n1756 ;
  assign n2009 = n1284 ^ n420 ^ n281 ;
  assign n2010 = n378 & ~n1307 ;
  assign n2011 = ~n1020 & n2010 ;
  assign n2012 = n1539 ^ n1336 ^ 1'b0 ;
  assign n2013 = n478 & n2012 ;
  assign n2014 = n2013 ^ n1461 ^ 1'b0 ;
  assign n2015 = n1146 ^ x46 ^ 1'b0 ;
  assign n2016 = n2014 | n2015 ;
  assign n2017 = n1469 | n2016 ;
  assign n2024 = n504 | n578 ;
  assign n2025 = n2024 ^ n429 ^ 1'b0 ;
  assign n2018 = n1475 ^ n1053 ^ 1'b0 ;
  assign n2019 = n172 ^ n161 ^ 1'b0 ;
  assign n2020 = n285 & n2019 ;
  assign n2021 = n2020 ^ n1135 ^ 1'b0 ;
  assign n2022 = n1131 & n2021 ;
  assign n2023 = ~n2018 & n2022 ;
  assign n2026 = n2025 ^ n2023 ^ 1'b0 ;
  assign n2031 = n1262 ^ n817 ^ n413 ;
  assign n2027 = n129 & ~n1615 ;
  assign n2028 = ~n781 & n2027 ;
  assign n2029 = n1843 ^ n1090 ^ 1'b0 ;
  assign n2030 = ( n425 & ~n2028 ) | ( n425 & n2029 ) | ( ~n2028 & n2029 ) ;
  assign n2032 = n2031 ^ n2030 ^ n254 ;
  assign n2037 = n886 ^ x60 ^ 1'b0 ;
  assign n2038 = n1116 & ~n2037 ;
  assign n2039 = n2038 ^ n1903 ^ n1311 ;
  assign n2033 = x53 & ~n833 ;
  assign n2034 = n2033 ^ n1997 ^ 1'b0 ;
  assign n2035 = ~n1542 & n2034 ;
  assign n2036 = n2035 ^ n1449 ^ 1'b0 ;
  assign n2040 = n2039 ^ n2036 ^ n853 ;
  assign n2041 = n422 & n1428 ;
  assign n2042 = n979 ^ n833 ^ 1'b0 ;
  assign n2043 = n512 & ~n2042 ;
  assign n2044 = n2043 ^ n1754 ^ 1'b0 ;
  assign n2045 = ~n1248 & n2044 ;
  assign n2046 = n2045 ^ n625 ^ 1'b0 ;
  assign n2047 = ( n614 & n629 ) | ( n614 & n1397 ) | ( n629 & n1397 ) ;
  assign n2048 = n1584 ^ n983 ^ 1'b0 ;
  assign n2049 = x39 | n347 ;
  assign n2050 = x115 & ~n696 ;
  assign n2051 = n1282 & n2050 ;
  assign n2052 = n2051 ^ n1027 ^ 1'b0 ;
  assign n2053 = n2049 & n2052 ;
  assign n2054 = ( n1837 & n1996 ) | ( n1837 & ~n2053 ) | ( n1996 & ~n2053 ) ;
  assign n2055 = n730 ^ n379 ^ n225 ;
  assign n2056 = ~n1647 & n2055 ;
  assign n2057 = n1227 ^ n190 ^ 1'b0 ;
  assign n2058 = n1810 | n2057 ;
  assign n2059 = ( n1470 & ~n2056 ) | ( n1470 & n2058 ) | ( ~n2056 & n2058 ) ;
  assign n2060 = n1334 & ~n1378 ;
  assign n2061 = n685 & ~n736 ;
  assign n2062 = n2061 ^ n741 ^ 1'b0 ;
  assign n2063 = n1675 ^ n1036 ^ n186 ;
  assign n2064 = ~x53 & n160 ;
  assign n2065 = n1116 & ~n1513 ;
  assign n2066 = ~n937 & n2065 ;
  assign n2067 = x65 & ~n1976 ;
  assign n2068 = n2067 ^ x49 ^ 1'b0 ;
  assign n2069 = ( n950 & n1976 ) | ( n950 & ~n2068 ) | ( n1976 & ~n2068 ) ;
  assign n2070 = n1626 ^ n1006 ^ n715 ;
  assign n2071 = n143 | n412 ;
  assign n2072 = n1774 & ~n2071 ;
  assign n2073 = n1294 & ~n2072 ;
  assign n2074 = n2073 ^ x6 ^ 1'b0 ;
  assign n2075 = n1096 ^ n327 ^ 1'b0 ;
  assign n2076 = n1231 & ~n2075 ;
  assign n2077 = n1065 & n2076 ;
  assign n2078 = ( ~n696 & n1260 ) | ( ~n696 & n2077 ) | ( n1260 & n2077 ) ;
  assign n2079 = ( ~n944 & n1455 ) | ( ~n944 & n1942 ) | ( n1455 & n1942 ) ;
  assign n2080 = n925 | n1469 ;
  assign n2081 = n2079 & ~n2080 ;
  assign n2082 = n2081 ^ n1545 ^ 1'b0 ;
  assign n2083 = n2082 ^ n363 ^ 1'b0 ;
  assign n2084 = ( n700 & ~n1370 ) | ( n700 & n2083 ) | ( ~n1370 & n2083 ) ;
  assign n2085 = n609 | n1523 ;
  assign n2086 = ( n597 & n1667 ) | ( n597 & n2085 ) | ( n1667 & n2085 ) ;
  assign n2087 = n541 ^ x105 ^ 1'b0 ;
  assign n2090 = n391 & ~n945 ;
  assign n2091 = ~n1785 & n2090 ;
  assign n2092 = ~x22 & n2091 ;
  assign n2093 = n350 | n2092 ;
  assign n2094 = n2093 ^ n1714 ^ 1'b0 ;
  assign n2088 = n660 | n681 ;
  assign n2089 = n2088 ^ x126 ^ 1'b0 ;
  assign n2095 = n2094 ^ n2089 ^ n1046 ;
  assign n2096 = n2095 ^ n1873 ^ 1'b0 ;
  assign n2097 = n2087 | n2096 ;
  assign n2098 = x61 & ~n1018 ;
  assign n2099 = ( n386 & ~n1452 ) | ( n386 & n2098 ) | ( ~n1452 & n2098 ) ;
  assign n2100 = n1560 ^ n1306 ^ n211 ;
  assign n2101 = n2099 & ~n2100 ;
  assign n2107 = n418 & n885 ;
  assign n2102 = n573 ^ n305 ^ x69 ;
  assign n2103 = n473 ^ x119 ^ 1'b0 ;
  assign n2104 = n900 | n2103 ;
  assign n2105 = n2104 ^ n947 ^ x64 ;
  assign n2106 = n2102 & n2105 ;
  assign n2108 = n2107 ^ n2106 ^ 1'b0 ;
  assign n2109 = n1955 ^ n770 ^ 1'b0 ;
  assign n2110 = n2109 ^ n296 ^ 1'b0 ;
  assign n2111 = ~n279 & n839 ;
  assign n2112 = n2111 ^ n1841 ^ 1'b0 ;
  assign n2113 = n1192 & n2112 ;
  assign n2114 = n2113 ^ n1338 ^ 1'b0 ;
  assign n2115 = n913 & ~n2114 ;
  assign n2116 = n471 ^ n220 ^ 1'b0 ;
  assign n2117 = n568 | n2116 ;
  assign n2118 = n2117 ^ n980 ^ 1'b0 ;
  assign n2119 = x97 & n2118 ;
  assign n2120 = ~n828 & n2119 ;
  assign n2122 = n1903 ^ n546 ^ n152 ;
  assign n2121 = n1582 ^ n1454 ^ n673 ;
  assign n2123 = n2122 ^ n2121 ^ 1'b0 ;
  assign n2124 = n362 | n2123 ;
  assign n2128 = n337 ^ n155 ^ 1'b0 ;
  assign n2125 = n711 ^ n278 ^ 1'b0 ;
  assign n2126 = ( n353 & ~n1648 ) | ( n353 & n2125 ) | ( ~n1648 & n2125 ) ;
  assign n2127 = n2126 ^ n272 ^ 1'b0 ;
  assign n2129 = n2128 ^ n2127 ^ 1'b0 ;
  assign n2130 = n755 ^ n641 ^ 1'b0 ;
  assign n2131 = n1475 ^ n1164 ^ 1'b0 ;
  assign n2132 = n330 & ~n1457 ;
  assign n2133 = ~n302 & n2132 ;
  assign n2134 = n325 | n2133 ;
  assign n2135 = n284 | n341 ;
  assign n2136 = n447 | n2135 ;
  assign n2137 = n278 | n1524 ;
  assign n2138 = ~n2136 & n2137 ;
  assign n2139 = n412 & n1440 ;
  assign n2146 = n833 ^ n701 ^ 1'b0 ;
  assign n2140 = n1573 & n2018 ;
  assign n2141 = ( n462 & n877 ) | ( n462 & ~n893 ) | ( n877 & ~n893 ) ;
  assign n2142 = n1266 ^ x113 ^ 1'b0 ;
  assign n2143 = ~n1654 & n2142 ;
  assign n2144 = ( n1613 & n2141 ) | ( n1613 & ~n2143 ) | ( n2141 & ~n2143 ) ;
  assign n2145 = ( n251 & n2140 ) | ( n251 & ~n2144 ) | ( n2140 & ~n2144 ) ;
  assign n2147 = n2146 ^ n2145 ^ 1'b0 ;
  assign n2148 = n962 & ~n2147 ;
  assign n2149 = n189 | n672 ;
  assign n2150 = n2149 ^ n1074 ^ n942 ;
  assign n2151 = n2150 ^ n1127 ^ 1'b0 ;
  assign n2155 = n341 & ~n603 ;
  assign n2156 = ( n1294 & n1323 ) | ( n1294 & ~n2155 ) | ( n1323 & ~n2155 ) ;
  assign n2152 = x54 ^ x27 ^ 1'b0 ;
  assign n2153 = ~n847 & n2152 ;
  assign n2154 = x79 & n2153 ;
  assign n2157 = n2156 ^ n2154 ^ 1'b0 ;
  assign n2158 = n739 ^ x79 ^ 1'b0 ;
  assign n2159 = ~n2157 & n2158 ;
  assign n2160 = x108 & n523 ;
  assign n2161 = ~n234 & n2160 ;
  assign n2162 = n411 | n1682 ;
  assign n2163 = n2161 & ~n2162 ;
  assign n2164 = ~n779 & n878 ;
  assign n2165 = n822 & n2164 ;
  assign n2166 = n1990 | n2165 ;
  assign n2167 = n2163 & ~n2166 ;
  assign n2168 = x127 & n1168 ;
  assign n2169 = n2168 ^ n195 ^ 1'b0 ;
  assign n2170 = n622 & ~n859 ;
  assign n2171 = n2170 ^ n2092 ^ 1'b0 ;
  assign n2172 = ~n785 & n2171 ;
  assign n2173 = ( x24 & n2169 ) | ( x24 & ~n2172 ) | ( n2169 & ~n2172 ) ;
  assign n2174 = n289 & ~n712 ;
  assign n2175 = n2173 | n2174 ;
  assign n2176 = n2175 ^ n1659 ^ 1'b0 ;
  assign n2177 = n685 ^ n429 ^ 1'b0 ;
  assign n2178 = n2177 ^ n904 ^ n247 ;
  assign n2179 = n2178 ^ n563 ^ n175 ;
  assign n2180 = n1130 ^ x42 ^ 1'b0 ;
  assign n2181 = n238 | n2180 ;
  assign n2182 = n1800 ^ x54 ^ 1'b0 ;
  assign n2183 = n2182 ^ n1532 ^ 1'b0 ;
  assign n2184 = n175 & n190 ;
  assign n2185 = ~n1575 & n2184 ;
  assign n2186 = n2185 ^ n367 ^ 1'b0 ;
  assign n2187 = n1680 & ~n2186 ;
  assign n2188 = ( n449 & n848 ) | ( n449 & n1881 ) | ( n848 & n1881 ) ;
  assign n2189 = n2188 ^ n1459 ^ 1'b0 ;
  assign n2192 = n173 | n704 ;
  assign n2193 = n2192 ^ x3 ^ 1'b0 ;
  assign n2190 = ~n506 & n1220 ;
  assign n2191 = n795 & n2190 ;
  assign n2194 = n2193 ^ n2191 ^ 1'b0 ;
  assign n2195 = n2189 & n2194 ;
  assign n2196 = n2068 ^ n1020 ^ n970 ;
  assign n2197 = n2196 ^ n2179 ^ n187 ;
  assign n2198 = n963 & n1459 ;
  assign n2199 = ~n2126 & n2198 ;
  assign n2200 = n384 & n2199 ;
  assign n2201 = n2200 ^ n134 ^ 1'b0 ;
  assign n2202 = n1876 ^ n1689 ^ n883 ;
  assign n2203 = n1022 ^ n982 ^ 1'b0 ;
  assign n2204 = ( n1152 & n1379 ) | ( n1152 & n2203 ) | ( n1379 & n2203 ) ;
  assign n2205 = n588 ^ n165 ^ 1'b0 ;
  assign n2206 = ~n2204 & n2205 ;
  assign n2207 = n857 | n1126 ;
  assign n2208 = n1743 ^ n522 ^ 1'b0 ;
  assign n2209 = n2207 & ~n2208 ;
  assign n2210 = n1266 ^ n992 ^ 1'b0 ;
  assign n2211 = n2209 & ~n2210 ;
  assign n2212 = n2211 ^ n684 ^ n540 ;
  assign n2213 = n2206 & n2212 ;
  assign n2214 = x100 ^ x35 ^ 1'b0 ;
  assign n2215 = n1067 & n2214 ;
  assign n2216 = n1918 ^ n1110 ^ n672 ;
  assign n2217 = n1490 & ~n2216 ;
  assign n2218 = ( n568 & n1675 ) | ( n568 & ~n2182 ) | ( n1675 & ~n2182 ) ;
  assign n2219 = n1750 ^ x47 ^ 1'b0 ;
  assign n2220 = n2090 ^ n231 ^ 1'b0 ;
  assign n2221 = n1090 & ~n2220 ;
  assign n2222 = n2221 ^ n1058 ^ 1'b0 ;
  assign n2223 = n155 & n918 ;
  assign n2224 = ~n1683 & n2223 ;
  assign n2225 = n2224 ^ n1695 ^ 1'b0 ;
  assign n2226 = n1931 & n2225 ;
  assign n2227 = n2226 ^ n787 ^ 1'b0 ;
  assign n2228 = n1356 | n2227 ;
  assign n2229 = n1906 ^ n1744 ^ 1'b0 ;
  assign n2230 = n1272 & n1298 ;
  assign n2231 = n2229 & n2230 ;
  assign n2232 = x40 & x80 ;
  assign n2233 = n1485 & n2232 ;
  assign n2234 = n1956 ^ n1101 ^ 1'b0 ;
  assign n2235 = n2233 | n2234 ;
  assign n2238 = ( ~n146 & n250 ) | ( ~n146 & n1536 ) | ( n250 & n1536 ) ;
  assign n2236 = n1694 & n1774 ;
  assign n2237 = n2236 ^ n1728 ^ 1'b0 ;
  assign n2239 = n2238 ^ n2237 ^ n1545 ;
  assign n2241 = n2028 ^ n1818 ^ 1'b0 ;
  assign n2242 = n2241 ^ n523 ^ 1'b0 ;
  assign n2240 = ~n1992 & n2034 ;
  assign n2243 = n2242 ^ n2240 ^ 1'b0 ;
  assign n2246 = ~x13 & n730 ;
  assign n2244 = n1902 ^ n685 ^ 1'b0 ;
  assign n2245 = n303 | n2244 ;
  assign n2247 = n2246 ^ n2245 ^ 1'b0 ;
  assign n2248 = n2082 | n2247 ;
  assign n2249 = x13 & n1535 ;
  assign n2250 = n2248 & n2249 ;
  assign n2251 = n1826 ^ n1655 ^ 1'b0 ;
  assign n2252 = ( n131 & ~n1271 ) | ( n131 & n1764 ) | ( ~n1271 & n1764 ) ;
  assign n2253 = n2252 ^ n1510 ^ 1'b0 ;
  assign n2254 = n2253 ^ n1375 ^ n1101 ;
  assign n2255 = n2251 & n2254 ;
  assign n2256 = n2250 & n2255 ;
  assign n2263 = n312 & ~n1023 ;
  assign n2264 = n2263 ^ n459 ^ 1'b0 ;
  assign n2260 = ( n360 & n496 ) | ( n360 & ~n1647 ) | ( n496 & ~n1647 ) ;
  assign n2261 = ~n391 & n2260 ;
  assign n2262 = n2261 ^ n1143 ^ 1'b0 ;
  assign n2257 = n463 ^ x2 ^ 1'b0 ;
  assign n2258 = x20 & n2257 ;
  assign n2259 = ( n203 & n1348 ) | ( n203 & n2258 ) | ( n1348 & n2258 ) ;
  assign n2265 = n2264 ^ n2262 ^ n2259 ;
  assign n2266 = n2265 ^ n927 ^ 1'b0 ;
  assign n2267 = n1035 & n2266 ;
  assign n2268 = n1587 ^ n901 ^ x28 ;
  assign n2269 = ( n1181 & n1648 ) | ( n1181 & n2268 ) | ( n1648 & n2268 ) ;
  assign n2272 = ~n211 & n1998 ;
  assign n2270 = ( x75 & ~n788 ) | ( x75 & n1534 ) | ( ~n788 & n1534 ) ;
  assign n2271 = ~n1170 & n2270 ;
  assign n2273 = n2272 ^ n2271 ^ 1'b0 ;
  assign n2274 = ~n1141 & n2273 ;
  assign n2275 = ~x8 & n2274 ;
  assign n2276 = n931 & n2268 ;
  assign n2277 = n1035 ^ n936 ^ 1'b0 ;
  assign n2278 = ~n438 & n2277 ;
  assign n2279 = n2278 ^ n1708 ^ 1'b0 ;
  assign n2280 = ( ~n1104 & n1982 ) | ( ~n1104 & n2279 ) | ( n1982 & n2279 ) ;
  assign n2281 = n1067 ^ n207 ^ 1'b0 ;
  assign n2282 = n744 & n2281 ;
  assign n2283 = ( n1715 & ~n1937 ) | ( n1715 & n2188 ) | ( ~n1937 & n2188 ) ;
  assign n2284 = ~n661 & n1709 ;
  assign n2285 = ~n335 & n2284 ;
  assign n2286 = n2282 ^ n1798 ^ 1'b0 ;
  assign n2287 = n521 & n1756 ;
  assign n2288 = n1529 & n2287 ;
  assign n2289 = x113 & n1175 ;
  assign n2290 = n2289 ^ n709 ^ 1'b0 ;
  assign n2291 = n2290 ^ x97 ^ 1'b0 ;
  assign n2295 = n377 & ~n1140 ;
  assign n2296 = n461 & n2295 ;
  assign n2297 = ( ~n729 & n936 ) | ( ~n729 & n2296 ) | ( n936 & n2296 ) ;
  assign n2292 = n704 ^ n201 ^ 1'b0 ;
  assign n2293 = n603 | n2292 ;
  assign n2294 = n1057 & ~n2293 ;
  assign n2298 = n2297 ^ n2294 ^ 1'b0 ;
  assign n2299 = n2291 & ~n2298 ;
  assign n2307 = n849 & n1617 ;
  assign n2308 = n2307 ^ n438 ^ 1'b0 ;
  assign n2300 = n881 ^ n741 ^ 1'b0 ;
  assign n2301 = x95 & n247 ;
  assign n2302 = n1478 ^ x96 ^ 1'b0 ;
  assign n2303 = n2301 & ~n2302 ;
  assign n2304 = n1761 ^ n1758 ^ 1'b0 ;
  assign n2305 = n2303 & n2304 ;
  assign n2306 = ~n2300 & n2305 ;
  assign n2309 = n2308 ^ n2306 ^ 1'b0 ;
  assign n2310 = n2299 | n2309 ;
  assign n2314 = n1810 | n2042 ;
  assign n2315 = n473 & ~n2314 ;
  assign n2311 = n1911 ^ n1094 ^ 1'b0 ;
  assign n2312 = ~n648 & n2311 ;
  assign n2313 = n1505 & n2312 ;
  assign n2316 = n2315 ^ n2313 ^ 1'b0 ;
  assign n2317 = n1876 & ~n2042 ;
  assign n2318 = ~n2316 & n2317 ;
  assign n2319 = n2318 ^ n802 ^ 1'b0 ;
  assign n2320 = n404 & ~n2319 ;
  assign n2321 = n408 & n2097 ;
  assign n2323 = n427 & ~n1141 ;
  assign n2322 = n1563 ^ x0 ^ 1'b0 ;
  assign n2324 = n2323 ^ n2322 ^ n1309 ;
  assign n2325 = n1495 | n1965 ;
  assign n2326 = n2325 ^ n259 ^ 1'b0 ;
  assign n2327 = n1973 ^ n591 ^ 1'b0 ;
  assign n2328 = ~n665 & n2327 ;
  assign n2329 = n506 & n1371 ;
  assign n2330 = n2329 ^ n988 ^ 1'b0 ;
  assign n2331 = n2328 & ~n2330 ;
  assign n2332 = n2331 ^ n309 ^ 1'b0 ;
  assign n2333 = n1554 ^ n933 ^ 1'b0 ;
  assign n2335 = n2169 ^ n1003 ^ 1'b0 ;
  assign n2334 = ( n557 & n1006 ) | ( n557 & ~n1868 ) | ( n1006 & ~n1868 ) ;
  assign n2336 = n2335 ^ n2334 ^ 1'b0 ;
  assign n2337 = n732 & n2336 ;
  assign n2338 = n2337 ^ n161 ^ 1'b0 ;
  assign n2339 = n347 | n2338 ;
  assign n2340 = n2333 & ~n2339 ;
  assign n2342 = ( x116 & n436 ) | ( x116 & ~n739 ) | ( n436 & ~n739 ) ;
  assign n2343 = ~n1923 & n2342 ;
  assign n2344 = n2343 ^ n1561 ^ 1'b0 ;
  assign n2345 = n2344 ^ n1434 ^ 1'b0 ;
  assign n2341 = n1589 ^ n522 ^ 1'b0 ;
  assign n2346 = n2345 ^ n2341 ^ 1'b0 ;
  assign n2347 = n1370 | n2346 ;
  assign n2348 = x55 & n178 ;
  assign n2349 = ~n511 & n2348 ;
  assign n2350 = ~n661 & n2349 ;
  assign n2351 = n254 & ~n932 ;
  assign n2352 = n2350 & n2351 ;
  assign n2353 = ( n384 & n397 ) | ( n384 & ~n2352 ) | ( n397 & ~n2352 ) ;
  assign n2354 = ~n281 & n1294 ;
  assign n2355 = ~n791 & n2354 ;
  assign n2356 = n788 & ~n2355 ;
  assign n2357 = n2353 & n2356 ;
  assign n2358 = ( n805 & ~n831 ) | ( n805 & n2357 ) | ( ~n831 & n2357 ) ;
  assign n2359 = ( ~n1972 & n1999 ) | ( ~n1972 & n2358 ) | ( n1999 & n2358 ) ;
  assign n2363 = n362 ^ n201 ^ 1'b0 ;
  assign n2364 = ( n932 & n2315 ) | ( n932 & n2363 ) | ( n2315 & n2363 ) ;
  assign n2360 = n572 ^ n293 ^ 1'b0 ;
  assign n2361 = ~n506 & n2360 ;
  assign n2362 = ~n227 & n2361 ;
  assign n2365 = n2364 ^ n2362 ^ 1'b0 ;
  assign n2366 = n1373 | n1976 ;
  assign n2367 = n2366 ^ n1726 ^ 1'b0 ;
  assign n2368 = n2365 & n2367 ;
  assign n2369 = n1291 ^ n320 ^ 1'b0 ;
  assign n2370 = ~n227 & n2369 ;
  assign n2371 = ( ~x17 & n1761 ) | ( ~x17 & n2370 ) | ( n1761 & n2370 ) ;
  assign n2372 = n2371 ^ n2229 ^ 1'b0 ;
  assign n2373 = n568 | n1079 ;
  assign n2374 = n748 & ~n2373 ;
  assign n2375 = n1246 ^ n420 ^ 1'b0 ;
  assign n2376 = n1435 ^ n381 ^ 1'b0 ;
  assign n2377 = x27 & n2376 ;
  assign n2378 = n216 | n2377 ;
  assign n2379 = n905 ^ n672 ^ 1'b0 ;
  assign n2380 = n2379 ^ n1579 ^ n563 ;
  assign n2381 = n2378 | n2380 ;
  assign n2382 = n850 ^ n245 ^ x114 ;
  assign n2383 = ( ~n584 & n1459 ) | ( ~n584 & n2382 ) | ( n1459 & n2382 ) ;
  assign n2384 = n2383 ^ n403 ^ 1'b0 ;
  assign n2385 = n668 | n2384 ;
  assign n2386 = n2385 ^ n1259 ^ 1'b0 ;
  assign n2387 = ( n465 & n2365 ) | ( n465 & n2386 ) | ( n2365 & n2386 ) ;
  assign n2388 = n730 | n1403 ;
  assign n2389 = ( n506 & ~n641 ) | ( n506 & n1853 ) | ( ~n641 & n1853 ) ;
  assign n2390 = n1513 ^ n540 ^ 1'b0 ;
  assign n2391 = ( n227 & ~n381 ) | ( n227 & n1037 ) | ( ~n381 & n1037 ) ;
  assign n2392 = n1422 | n2391 ;
  assign n2393 = n2390 & ~n2392 ;
  assign n2394 = n915 ^ n561 ^ 1'b0 ;
  assign n2395 = x20 & ~n2394 ;
  assign n2396 = n324 & n697 ;
  assign n2397 = ~n270 & n2396 ;
  assign n2398 = n1057 ^ x99 ^ 1'b0 ;
  assign n2399 = ~n2397 & n2398 ;
  assign n2400 = ( n493 & ~n528 ) | ( n493 & n1006 ) | ( ~n528 & n1006 ) ;
  assign n2401 = x99 & n421 ;
  assign n2402 = ( ~n1402 & n2400 ) | ( ~n1402 & n2401 ) | ( n2400 & n2401 ) ;
  assign n2403 = ~n1332 & n2402 ;
  assign n2404 = n2248 & n2403 ;
  assign n2405 = n641 | n690 ;
  assign n2406 = n2405 ^ x70 ^ 1'b0 ;
  assign n2407 = n421 & n1060 ;
  assign n2408 = n2407 ^ n903 ^ 1'b0 ;
  assign n2409 = x7 & n267 ;
  assign n2410 = x101 & n935 ;
  assign n2411 = n2410 ^ x1 ^ 1'b0 ;
  assign n2412 = n2239 & ~n2411 ;
  assign n2413 = n2409 & n2412 ;
  assign n2414 = x35 & ~n579 ;
  assign n2415 = n2414 ^ n1252 ^ 1'b0 ;
  assign n2416 = n1826 | n2233 ;
  assign n2424 = n970 | n1283 ;
  assign n2425 = n2424 ^ n1342 ^ 1'b0 ;
  assign n2426 = ~n180 & n2425 ;
  assign n2417 = n1483 ^ n797 ^ 1'b0 ;
  assign n2418 = ( n1132 & n1949 ) | ( n1132 & ~n2417 ) | ( n1949 & ~n2417 ) ;
  assign n2419 = n2418 ^ n1202 ^ n649 ;
  assign n2420 = n1156 ^ n847 ^ x78 ;
  assign n2421 = n848 & n2420 ;
  assign n2422 = ~n2312 & n2421 ;
  assign n2423 = ( n1929 & n2419 ) | ( n1929 & n2422 ) | ( n2419 & n2422 ) ;
  assign n2427 = n2426 ^ n2423 ^ 1'b0 ;
  assign n2436 = ~n298 & n436 ;
  assign n2437 = n2436 ^ n535 ^ 1'b0 ;
  assign n2433 = n1933 ^ n266 ^ 1'b0 ;
  assign n2434 = n155 & n2433 ;
  assign n2435 = ( x80 & ~n378 ) | ( x80 & n2434 ) | ( ~n378 & n2434 ) ;
  assign n2428 = n557 ^ x34 ^ 1'b0 ;
  assign n2429 = n2428 ^ n1660 ^ 1'b0 ;
  assign n2430 = ~n1470 & n2429 ;
  assign n2431 = n2430 ^ n1623 ^ 1'b0 ;
  assign n2432 = n2431 ^ n555 ^ 1'b0 ;
  assign n2438 = n2437 ^ n2435 ^ n2432 ;
  assign n2439 = n1881 ^ n140 ^ 1'b0 ;
  assign n2440 = n714 & n2439 ;
  assign n2441 = ~n1280 & n2440 ;
  assign n2442 = n565 ^ n206 ^ 1'b0 ;
  assign n2443 = n520 & n2442 ;
  assign n2444 = n242 & n2443 ;
  assign n2445 = n796 & ~n1695 ;
  assign n2446 = n2445 ^ n1729 ^ 1'b0 ;
  assign n2447 = n904 | n2446 ;
  assign n2448 = n2141 ^ n1943 ^ 1'b0 ;
  assign n2449 = n956 ^ n187 ^ 1'b0 ;
  assign n2450 = ~n1282 & n2449 ;
  assign n2451 = n390 & n767 ;
  assign n2452 = n1023 ^ n408 ^ 1'b0 ;
  assign n2453 = n2452 ^ n1976 ^ 1'b0 ;
  assign n2454 = n261 & n2453 ;
  assign n2455 = ( ~n254 & n2451 ) | ( ~n254 & n2454 ) | ( n2451 & n2454 ) ;
  assign n2456 = n2434 ^ n942 ^ 1'b0 ;
  assign n2457 = n2456 ^ n1555 ^ n1165 ;
  assign n2458 = n657 ^ x33 ^ 1'b0 ;
  assign n2459 = ~n318 & n1078 ;
  assign n2460 = ( n1713 & n2458 ) | ( n1713 & n2459 ) | ( n2458 & n2459 ) ;
  assign n2461 = n2457 & ~n2460 ;
  assign n2462 = n2461 ^ n170 ^ 1'b0 ;
  assign n2463 = n395 ^ n233 ^ 1'b0 ;
  assign n2464 = n432 & ~n2463 ;
  assign n2465 = n1438 ^ n1139 ^ 1'b0 ;
  assign n2466 = n2464 & ~n2465 ;
  assign n2467 = n512 & ~n2466 ;
  assign n2468 = n834 & n1988 ;
  assign n2469 = n578 & n2468 ;
  assign n2470 = ~n2467 & n2469 ;
  assign n2471 = n175 & ~n1414 ;
  assign n2472 = ( n970 & n1672 ) | ( n970 & ~n2169 ) | ( n1672 & ~n2169 ) ;
  assign n2473 = ( x119 & n761 ) | ( x119 & n816 ) | ( n761 & n816 ) ;
  assign n2474 = n2473 ^ n1441 ^ 1'b0 ;
  assign n2475 = n2472 | n2474 ;
  assign n2476 = n2475 ^ n1613 ^ 1'b0 ;
  assign n2477 = n1283 | n2476 ;
  assign n2478 = n1102 ^ n906 ^ 1'b0 ;
  assign n2479 = n2477 ^ n206 ^ 1'b0 ;
  assign n2480 = n2102 ^ n1459 ^ 1'b0 ;
  assign n2481 = n874 & ~n2480 ;
  assign n2482 = n1000 & n2481 ;
  assign n2483 = n2482 ^ n1459 ^ 1'b0 ;
  assign n2484 = n739 & ~n2483 ;
  assign n2485 = n1946 ^ n511 ^ 1'b0 ;
  assign n2486 = n2484 | n2485 ;
  assign n2487 = n2280 ^ n785 ^ 1'b0 ;
  assign n2488 = ~n279 & n2406 ;
  assign n2490 = n781 & ~n893 ;
  assign n2491 = n618 & n2490 ;
  assign n2489 = n1145 ^ n256 ^ n165 ;
  assign n2492 = n2491 ^ n2489 ^ n458 ;
  assign n2493 = n1677 & n1998 ;
  assign n2494 = n2493 ^ x91 ^ x50 ;
  assign n2495 = n340 ^ n154 ^ 1'b0 ;
  assign n2496 = ~n1154 & n2495 ;
  assign n2497 = n1200 ^ n597 ^ n525 ;
  assign n2498 = ~n569 & n1306 ;
  assign n2499 = ( n2496 & n2497 ) | ( n2496 & n2498 ) | ( n2497 & n2498 ) ;
  assign n2500 = n1502 ^ n1340 ^ n129 ;
  assign n2501 = ( n580 & n800 ) | ( n580 & ~n1658 ) | ( n800 & ~n1658 ) ;
  assign n2502 = n161 & ~n267 ;
  assign n2503 = n2502 ^ n160 ^ 1'b0 ;
  assign n2504 = n563 & ~n2503 ;
  assign n2505 = n2504 ^ x44 ^ 1'b0 ;
  assign n2506 = ~n1923 & n2505 ;
  assign n2507 = n553 & ~n1558 ;
  assign n2508 = n2507 ^ n2236 ^ 1'b0 ;
  assign n2509 = n2055 ^ n940 ^ 1'b0 ;
  assign n2510 = n1669 & n2509 ;
  assign n2511 = ( ~n1856 & n1931 ) | ( ~n1856 & n2510 ) | ( n1931 & n2510 ) ;
  assign n2512 = n499 & n1445 ;
  assign n2513 = ( ~n1349 & n2243 ) | ( ~n1349 & n2512 ) | ( n2243 & n2512 ) ;
  assign n2514 = ( x75 & x113 ) | ( x75 & n2513 ) | ( x113 & n2513 ) ;
  assign n2515 = ~n254 & n1648 ;
  assign n2516 = n2432 & ~n2515 ;
  assign n2517 = x89 | n1325 ;
  assign n2524 = n1054 ^ n378 ^ n366 ;
  assign n2518 = n578 | n1674 ;
  assign n2519 = x121 | n2518 ;
  assign n2520 = ( n1558 & n1560 ) | ( n1558 & n2329 ) | ( n1560 & n2329 ) ;
  assign n2521 = ( n1363 & n2519 ) | ( n1363 & ~n2520 ) | ( n2519 & ~n2520 ) ;
  assign n2522 = n1788 ^ n1162 ^ 1'b0 ;
  assign n2523 = n2521 & n2522 ;
  assign n2525 = n2524 ^ n2523 ^ 1'b0 ;
  assign n2526 = n2517 & n2525 ;
  assign n2527 = n152 | n190 ;
  assign n2533 = n1516 & ~n2452 ;
  assign n2534 = n2533 ^ n1029 ^ 1'b0 ;
  assign n2535 = n2534 ^ n512 ^ 1'b0 ;
  assign n2530 = n622 ^ n575 ^ 1'b0 ;
  assign n2528 = n314 & ~n509 ;
  assign n2529 = n829 & n2528 ;
  assign n2531 = n2530 ^ n2529 ^ 1'b0 ;
  assign n2532 = ( n932 & ~n1587 ) | ( n932 & n2531 ) | ( ~n1587 & n2531 ) ;
  assign n2536 = n2535 ^ n2532 ^ n1658 ;
  assign n2537 = n1106 ^ n917 ^ 1'b0 ;
  assign n2538 = n451 | n2537 ;
  assign n2539 = n307 & n1306 ;
  assign n2540 = n299 & n2539 ;
  assign n2541 = n2540 ^ n1777 ^ 1'b0 ;
  assign n2542 = ~n2538 & n2541 ;
  assign n2543 = n1168 & n1463 ;
  assign n2544 = n2543 ^ n2278 ^ 1'b0 ;
  assign n2546 = ( n319 & n444 ) | ( n319 & ~n1135 ) | ( n444 & ~n1135 ) ;
  assign n2545 = n1351 & n2018 ;
  assign n2547 = n2546 ^ n2545 ^ 1'b0 ;
  assign n2548 = n928 & ~n1682 ;
  assign n2549 = ~n1647 & n2548 ;
  assign n2550 = n1240 | n1406 ;
  assign n2551 = n2549 & ~n2550 ;
  assign n2558 = n469 & ~n771 ;
  assign n2559 = n2558 ^ n363 ^ 1'b0 ;
  assign n2556 = n697 & n775 ;
  assign n2557 = n2556 ^ n236 ^ 1'b0 ;
  assign n2560 = n2559 ^ n2557 ^ n412 ;
  assign n2561 = n293 & n2049 ;
  assign n2562 = ~n2560 & n2561 ;
  assign n2553 = n843 ^ n723 ^ 1'b0 ;
  assign n2554 = n2553 ^ n1544 ^ n1176 ;
  assign n2555 = n2554 ^ n1365 ^ n1209 ;
  assign n2552 = n639 ^ n586 ^ 1'b0 ;
  assign n2563 = n2562 ^ n2555 ^ n2552 ;
  assign n2564 = n560 & ~n1269 ;
  assign n2565 = n785 & n2564 ;
  assign n2566 = n2565 ^ n1648 ^ 1'b0 ;
  assign n2573 = n1228 ^ x25 ^ 1'b0 ;
  assign n2567 = n1419 ^ n1290 ^ 1'b0 ;
  assign n2568 = n1720 ^ n925 ^ 1'b0 ;
  assign n2569 = n2568 ^ n934 ^ 1'b0 ;
  assign n2570 = n2569 ^ n850 ^ 1'b0 ;
  assign n2571 = n2570 ^ n824 ^ 1'b0 ;
  assign n2572 = n2567 | n2571 ;
  assign n2574 = n2573 ^ n2572 ^ 1'b0 ;
  assign n2575 = n270 & ~n2161 ;
  assign n2576 = ~n530 & n2182 ;
  assign n2577 = ( n1613 & ~n2575 ) | ( n1613 & n2576 ) | ( ~n2575 & n2576 ) ;
  assign n2578 = n1138 ^ n557 ^ 1'b0 ;
  assign n2579 = ( n220 & ~n1290 ) | ( n220 & n2578 ) | ( ~n1290 & n2578 ) ;
  assign n2580 = n2579 ^ n2007 ^ n1215 ;
  assign n2581 = n758 ^ n424 ^ n146 ;
  assign n2582 = n2581 ^ n2283 ^ 1'b0 ;
  assign n2583 = n2246 ^ n1721 ^ 1'b0 ;
  assign n2584 = n2254 & ~n2583 ;
  assign n2585 = n729 ^ n390 ^ 1'b0 ;
  assign n2586 = n168 & ~n2585 ;
  assign n2587 = x96 & ~n1221 ;
  assign n2588 = n2587 ^ n946 ^ n833 ;
  assign n2589 = ( n1311 & ~n2586 ) | ( n1311 & n2588 ) | ( ~n2586 & n2588 ) ;
  assign n2590 = n502 & n597 ;
  assign n2591 = ~x42 & n2019 ;
  assign n2592 = n2591 ^ n1326 ^ n1294 ;
  assign n2593 = n1853 & n2483 ;
  assign n2594 = n839 | n2574 ;
  assign n2595 = n1338 & ~n2594 ;
  assign n2596 = ~n1246 & n2359 ;
  assign n2597 = n1430 ^ n936 ^ n734 ;
  assign n2598 = n1825 ^ n1352 ^ n172 ;
  assign n2599 = n1020 ^ n800 ^ n740 ;
  assign n2605 = n1430 ^ n249 ^ 1'b0 ;
  assign n2606 = n499 & ~n2605 ;
  assign n2602 = ( n335 & n543 ) | ( n335 & ~n2128 ) | ( n543 & ~n2128 ) ;
  assign n2603 = n1159 ^ n541 ^ 1'b0 ;
  assign n2604 = n2602 & ~n2603 ;
  assign n2600 = ~n618 & n1313 ;
  assign n2601 = n2600 ^ n820 ^ 1'b0 ;
  assign n2607 = n2606 ^ n2604 ^ n2601 ;
  assign n2608 = n2607 ^ n1202 ^ 1'b0 ;
  assign n2609 = n2599 & n2608 ;
  assign n2610 = n1984 ^ n718 ^ 1'b0 ;
  assign n2611 = n865 & n2610 ;
  assign n2612 = ( ~n1373 & n1820 ) | ( ~n1373 & n1836 ) | ( n1820 & n1836 ) ;
  assign n2613 = x106 & n257 ;
  assign n2614 = n2613 ^ n2012 ^ n626 ;
  assign n2615 = n692 | n1148 ;
  assign n2616 = n838 & n2615 ;
  assign n2617 = n718 ^ x24 ^ 1'b0 ;
  assign n2618 = n1729 | n2617 ;
  assign n2619 = n438 | n2618 ;
  assign n2621 = n211 & ~n970 ;
  assign n2620 = ~n1017 & n1375 ;
  assign n2622 = n2621 ^ n2620 ^ 1'b0 ;
  assign n2623 = n2622 ^ x5 ^ 1'b0 ;
  assign n2624 = n2384 | n2623 ;
  assign n2625 = n209 | n2624 ;
  assign n2626 = n1259 ^ n419 ^ 1'b0 ;
  assign n2627 = n1489 & n2626 ;
  assign n2628 = ~n2496 & n2627 ;
  assign n2629 = n2628 ^ n727 ^ 1'b0 ;
  assign n2630 = n2625 & n2629 ;
  assign n2631 = n945 | n1720 ;
  assign n2632 = n2631 ^ n1959 ^ 1'b0 ;
  assign n2633 = n2406 & ~n2632 ;
  assign n2634 = n207 & ~n836 ;
  assign n2635 = n2634 ^ n734 ^ 1'b0 ;
  assign n2636 = x114 & n2635 ;
  assign n2637 = ~n1812 & n2636 ;
  assign n2638 = ( x12 & ~n222 ) | ( x12 & n967 ) | ( ~n222 & n967 ) ;
  assign n2639 = x61 & ~n2296 ;
  assign n2640 = n2638 & n2639 ;
  assign n2641 = n2640 ^ n797 ^ 1'b0 ;
  assign n2642 = n2349 ^ x62 ^ 1'b0 ;
  assign n2643 = x63 & ~n2642 ;
  assign n2644 = ~n1653 & n2643 ;
  assign n2645 = n2644 ^ n848 ^ 1'b0 ;
  assign n2646 = n2641 | n2645 ;
  assign n2647 = n2646 ^ n2148 ^ 1'b0 ;
  assign n2648 = ( ~n1683 & n2637 ) | ( ~n1683 & n2647 ) | ( n2637 & n2647 ) ;
  assign n2650 = n763 | n1218 ;
  assign n2649 = n436 & n1355 ;
  assign n2651 = n2650 ^ n2649 ^ 1'b0 ;
  assign n2652 = n1435 ^ n1018 ^ 1'b0 ;
  assign n2653 = ~n2651 & n2652 ;
  assign n2654 = n2653 ^ n1491 ^ 1'b0 ;
  assign n2655 = ( n1495 & n1658 ) | ( n1495 & n2654 ) | ( n1658 & n2654 ) ;
  assign n2656 = x97 & n349 ;
  assign n2657 = n2656 ^ n1644 ^ 1'b0 ;
  assign n2658 = ( x94 & ~n712 ) | ( x94 & n2657 ) | ( ~n712 & n2657 ) ;
  assign n2659 = n1355 & ~n1868 ;
  assign n2660 = ~n2658 & n2659 ;
  assign n2661 = n254 & n1678 ;
  assign n2662 = ( n271 & n776 ) | ( n271 & n1308 ) | ( n776 & n1308 ) ;
  assign n2663 = n2662 ^ n866 ^ 1'b0 ;
  assign n2664 = n1532 & n2663 ;
  assign n2667 = x57 & ~n358 ;
  assign n2668 = n2667 ^ n463 ^ 1'b0 ;
  assign n2665 = n686 & n1290 ;
  assign n2666 = n1982 | n2665 ;
  assign n2669 = n2668 ^ n2666 ^ n1451 ;
  assign n2670 = n2662 & ~n2669 ;
  assign n2671 = ~n190 & n408 ;
  assign n2672 = ~n408 & n2671 ;
  assign n2673 = n704 | n2672 ;
  assign n2674 = n2672 & ~n2673 ;
  assign n2675 = n578 | n2674 ;
  assign n2676 = n1438 & ~n2675 ;
  assign n2677 = n2676 ^ n563 ^ 1'b0 ;
  assign n2680 = n370 | n1761 ;
  assign n2681 = n855 ^ x35 ^ 1'b0 ;
  assign n2682 = ~n2680 & n2681 ;
  assign n2679 = ~n425 & n1022 ;
  assign n2683 = n2682 ^ n2679 ^ 1'b0 ;
  assign n2684 = ~n2364 & n2683 ;
  assign n2678 = n923 ^ n243 ^ 1'b0 ;
  assign n2685 = n2684 ^ n2678 ^ n331 ;
  assign n2686 = n1118 & ~n2425 ;
  assign n2687 = ~n708 & n1965 ;
  assign n2688 = n390 & n404 ;
  assign n2689 = n2599 & n2688 ;
  assign n2690 = n1760 & n2689 ;
  assign n2691 = n2471 ^ x7 ^ 1'b0 ;
  assign n2692 = ~n2690 & n2691 ;
  assign n2693 = ( ~x13 & n747 ) | ( ~x13 & n2542 ) | ( n747 & n2542 ) ;
  assign n2698 = n2680 ^ n653 ^ 1'b0 ;
  assign n2696 = x123 & n737 ;
  assign n2697 = n2696 ^ n1648 ^ 1'b0 ;
  assign n2699 = n2698 ^ n2697 ^ n2363 ;
  assign n2694 = n499 & ~n1160 ;
  assign n2695 = n2694 ^ x121 ^ 1'b0 ;
  assign n2700 = n2699 ^ n2695 ^ 1'b0 ;
  assign n2701 = n833 | n898 ;
  assign n2702 = n920 | n2701 ;
  assign n2703 = n1633 & ~n2702 ;
  assign n2704 = n2524 ^ n265 ^ 1'b0 ;
  assign n2705 = n2703 & n2704 ;
  assign n2706 = n2705 ^ n1550 ^ n138 ;
  assign n2707 = ~n2587 & n2706 ;
  assign n2708 = n2707 ^ n1507 ^ 1'b0 ;
  assign n2709 = ~n1831 & n2708 ;
  assign n2710 = ( n260 & n474 ) | ( n260 & n887 ) | ( n474 & n887 ) ;
  assign n2711 = n1010 | n1136 ;
  assign n2712 = n2711 ^ n1977 ^ 1'b0 ;
  assign n2713 = ~n704 & n2712 ;
  assign n2714 = n2710 & n2713 ;
  assign n2715 = ( ~n1318 & n1534 ) | ( ~n1318 & n2248 ) | ( n1534 & n2248 ) ;
  assign n2716 = ( n811 & n2714 ) | ( n811 & n2715 ) | ( n2714 & n2715 ) ;
  assign n2717 = n2002 | n2422 ;
  assign n2718 = x21 & ~n145 ;
  assign n2719 = n2718 ^ n430 ^ 1'b0 ;
  assign n2720 = n331 | n572 ;
  assign n2721 = n2720 ^ x51 ^ 1'b0 ;
  assign n2723 = n700 & n1162 ;
  assign n2722 = ~n778 & n1331 ;
  assign n2724 = n2723 ^ n2722 ^ 1'b0 ;
  assign n2725 = n238 | n818 ;
  assign n2726 = ( ~n2721 & n2724 ) | ( ~n2721 & n2725 ) | ( n2724 & n2725 ) ;
  assign n2727 = n2726 ^ n138 ^ 1'b0 ;
  assign n2728 = n2719 | n2727 ;
  assign n2729 = x120 & n1738 ;
  assign n2730 = n1163 & n2729 ;
  assign n2731 = n2728 & ~n2730 ;
  assign n2732 = ~n452 & n819 ;
  assign n2733 = n1283 & n2732 ;
  assign n2734 = ~n1271 & n2733 ;
  assign n2735 = n870 & n2421 ;
  assign n2736 = ~n1645 & n2735 ;
  assign n2737 = ( n1358 & ~n1647 ) | ( n1358 & n1752 ) | ( ~n1647 & n1752 ) ;
  assign n2738 = n1435 ^ n1329 ^ 1'b0 ;
  assign n2739 = n1768 ^ n692 ^ 1'b0 ;
  assign n2740 = ( n1806 & n2738 ) | ( n1806 & n2739 ) | ( n2738 & n2739 ) ;
  assign n2741 = ( n1354 & ~n2031 ) | ( n1354 & n2740 ) | ( ~n2031 & n2740 ) ;
  assign n2742 = n2332 ^ n416 ^ 1'b0 ;
  assign n2743 = x67 & ~n2742 ;
  assign n2744 = ( n1497 & ~n1582 ) | ( n1497 & n1760 ) | ( ~n1582 & n1760 ) ;
  assign n2745 = n2744 ^ n980 ^ n142 ;
  assign n2746 = n1600 ^ n700 ^ n313 ;
  assign n2747 = n874 & ~n1743 ;
  assign n2748 = n2747 ^ n318 ^ 1'b0 ;
  assign n2749 = n2748 ^ n771 ^ 1'b0 ;
  assign n2750 = ~n2746 & n2749 ;
  assign n2751 = ~n1423 & n2189 ;
  assign n2752 = n2458 ^ n1539 ^ n1499 ;
  assign n2753 = ( x11 & ~x89 ) | ( x11 & n2752 ) | ( ~x89 & n2752 ) ;
  assign n2754 = ( n618 & n1084 ) | ( n618 & n2753 ) | ( n1084 & n2753 ) ;
  assign n2755 = n1689 & ~n2754 ;
  assign n2756 = n1503 | n1898 ;
  assign n2757 = n2653 ^ n1729 ^ 1'b0 ;
  assign n2758 = n2756 | n2757 ;
  assign n2759 = n1990 & n2521 ;
  assign n2760 = ( n1251 & ~n1342 ) | ( n1251 & n2641 ) | ( ~n1342 & n2641 ) ;
  assign n2761 = n1356 & ~n2760 ;
  assign n2767 = ( n140 & ~n168 ) | ( n140 & n536 ) | ( ~n168 & n536 ) ;
  assign n2766 = n295 | n2051 ;
  assign n2768 = n2767 ^ n2766 ^ 1'b0 ;
  assign n2765 = n378 & n1631 ;
  assign n2769 = n2768 ^ n2765 ^ 1'b0 ;
  assign n2762 = ~n995 & n1902 ;
  assign n2763 = ~n853 & n2762 ;
  assign n2764 = n1709 & ~n2763 ;
  assign n2770 = n2769 ^ n2764 ^ 1'b0 ;
  assign n2771 = n681 | n2770 ;
  assign n2776 = ( x110 & n1160 ) | ( x110 & n1862 ) | ( n1160 & n1862 ) ;
  assign n2777 = n2326 & n2776 ;
  assign n2778 = n2777 ^ n644 ^ 1'b0 ;
  assign n2772 = n857 ^ n184 ^ 1'b0 ;
  assign n2773 = n493 & n734 ;
  assign n2774 = ( ~n951 & n2772 ) | ( ~n951 & n2773 ) | ( n2772 & n2773 ) ;
  assign n2775 = n804 & n2774 ;
  assign n2779 = n2778 ^ n2775 ^ 1'b0 ;
  assign n2780 = n1457 ^ n303 ^ 1'b0 ;
  assign n2781 = n1539 & n2780 ;
  assign n2782 = n1702 | n2389 ;
  assign n2783 = n2384 ^ n2108 ^ x109 ;
  assign n2794 = n2238 ^ n1400 ^ 1'b0 ;
  assign n2795 = ~n1591 & n2794 ;
  assign n2796 = n456 & n2795 ;
  assign n2797 = n1544 & ~n2796 ;
  assign n2791 = n1516 ^ n1276 ^ 1'b0 ;
  assign n2784 = n1538 ^ n1231 ^ 1'b0 ;
  assign n2785 = x7 & n2784 ;
  assign n2786 = n1352 ^ n819 ^ 1'b0 ;
  assign n2787 = n2785 & ~n2786 ;
  assign n2788 = n2787 ^ n1706 ^ n416 ;
  assign n2789 = n1996 | n2788 ;
  assign n2790 = n1797 & n2789 ;
  assign n2792 = n2791 ^ n2790 ^ 1'b0 ;
  assign n2793 = n1503 | n2792 ;
  assign n2798 = n2797 ^ n2793 ^ 1'b0 ;
  assign n2799 = x63 | n172 ;
  assign n2800 = n1475 ^ n330 ^ 1'b0 ;
  assign n2801 = n427 & ~n2800 ;
  assign n2802 = n2038 ^ n225 ^ 1'b0 ;
  assign n2803 = n2557 | n2802 ;
  assign n2804 = n1728 & ~n2803 ;
  assign n2811 = n146 & ~n1485 ;
  assign n2812 = n186 | n1370 ;
  assign n2813 = n1759 | n2812 ;
  assign n2814 = n1269 ^ n809 ^ 1'b0 ;
  assign n2815 = n2813 & ~n2814 ;
  assign n2816 = ( n2031 & ~n2811 ) | ( n2031 & n2815 ) | ( ~n2811 & n2815 ) ;
  assign n2805 = n399 & ~n1014 ;
  assign n2806 = n2805 ^ n354 ^ 1'b0 ;
  assign n2807 = n1096 | n2806 ;
  assign n2808 = n2401 | n2807 ;
  assign n2809 = ~n2344 & n2808 ;
  assign n2810 = ~n1202 & n2809 ;
  assign n2817 = n2816 ^ n2810 ^ 1'b0 ;
  assign n2818 = n2004 ^ n1937 ^ 1'b0 ;
  assign n2819 = n2818 ^ x60 ^ 1'b0 ;
  assign n2820 = n1331 | n1376 ;
  assign n2821 = n1645 ^ n337 ^ 1'b0 ;
  assign n2822 = ~n1341 & n2821 ;
  assign n2825 = n1545 ^ n320 ^ 1'b0 ;
  assign n2826 = n715 & ~n2825 ;
  assign n2823 = n1087 & n1575 ;
  assign n2824 = n2823 ^ n1282 ^ n950 ;
  assign n2827 = n2826 ^ n2824 ^ 1'b0 ;
  assign n2828 = ( x16 & n389 ) | ( x16 & n1414 ) | ( n389 & n1414 ) ;
  assign n2829 = ( x62 & ~n526 ) | ( x62 & n2828 ) | ( ~n526 & n2828 ) ;
  assign n2830 = x73 & ~n293 ;
  assign n2831 = ~n2829 & n2830 ;
  assign n2832 = n868 | n2831 ;
  assign n2833 = n2832 ^ n1637 ^ 1'b0 ;
  assign n2834 = n1422 | n2833 ;
  assign n2835 = n322 | n2834 ;
  assign n2836 = ( n1651 & n1904 ) | ( n1651 & ~n2835 ) | ( n1904 & ~n2835 ) ;
  assign n2837 = ( n599 & n1228 ) | ( n599 & n2157 ) | ( n1228 & n2157 ) ;
  assign n2838 = x90 & x93 ;
  assign n2839 = n2838 ^ x87 ^ 1'b0 ;
  assign n2840 = n2039 ^ n206 ^ 1'b0 ;
  assign n2841 = n2839 | n2840 ;
  assign n2842 = ( n162 & n489 ) | ( n162 & n2841 ) | ( n489 & n2841 ) ;
  assign n2843 = n804 | n2842 ;
  assign n2844 = ( ~n1288 & n2837 ) | ( ~n1288 & n2843 ) | ( n2837 & n2843 ) ;
  assign n2845 = n1368 | n1660 ;
  assign n2846 = ( ~n1280 & n1485 ) | ( ~n1280 & n2845 ) | ( n1485 & n2845 ) ;
  assign n2847 = x13 | n784 ;
  assign n2848 = n2847 ^ x9 ^ 1'b0 ;
  assign n2849 = n2172 & ~n2848 ;
  assign n2850 = ( n131 & ~n616 ) | ( n131 & n2237 ) | ( ~n616 & n2237 ) ;
  assign n2851 = x23 & n2042 ;
  assign n2852 = n2851 ^ n1466 ^ 1'b0 ;
  assign n2853 = ~n2850 & n2852 ;
  assign n2854 = n2853 ^ n2715 ^ n410 ;
  assign n2855 = n705 | n1127 ;
  assign n2856 = n2855 ^ n1536 ^ 1'b0 ;
  assign n2857 = ( n367 & n1412 ) | ( n367 & n1586 ) | ( n1412 & n1586 ) ;
  assign n2858 = n684 & n1593 ;
  assign n2859 = n2857 & ~n2858 ;
  assign n2860 = ( ~n320 & n1227 ) | ( ~n320 & n1341 ) | ( n1227 & n1341 ) ;
  assign n2861 = n2395 & ~n2860 ;
  assign n2862 = n2767 & n2861 ;
  assign n2863 = n2179 ^ n2063 ^ 1'b0 ;
  assign n2864 = n1669 & ~n2863 ;
  assign n2865 = n2864 ^ n1240 ^ 1'b0 ;
  assign n2866 = n325 ^ n227 ^ 1'b0 ;
  assign n2867 = ~n725 & n2866 ;
  assign n2868 = n1452 ^ n1078 ^ n484 ;
  assign n2869 = n2868 ^ n323 ^ 1'b0 ;
  assign n2870 = n2867 | n2869 ;
  assign n2871 = n2870 ^ n2524 ^ 1'b0 ;
  assign n2872 = n1745 & ~n2871 ;
  assign n2873 = n1422 ^ n1124 ^ 1'b0 ;
  assign n2874 = n1593 ^ n1148 ^ n653 ;
  assign n2875 = n1114 & n2874 ;
  assign n2876 = ~n795 & n1719 ;
  assign n2877 = ~n2875 & n2876 ;
  assign n2878 = ( n565 & n2245 ) | ( n565 & ~n2877 ) | ( n2245 & ~n2877 ) ;
  assign n2879 = n2878 ^ n641 ^ 1'b0 ;
  assign n2880 = n2879 ^ n1773 ^ 1'b0 ;
  assign n2881 = n401 & ~n1327 ;
  assign n2882 = n2881 ^ n611 ^ 1'b0 ;
  assign n2883 = n2882 ^ n1268 ^ 1'b0 ;
  assign n2884 = n2449 & n2883 ;
  assign n2885 = ~n824 & n2884 ;
  assign n2886 = n1946 & n2885 ;
  assign n2887 = n677 & n1200 ;
  assign n2888 = n2886 & n2887 ;
  assign n2889 = ( ~n142 & n288 ) | ( ~n142 & n1205 ) | ( n288 & n1205 ) ;
  assign n2890 = ( n1920 & n2655 ) | ( n1920 & ~n2889 ) | ( n2655 & ~n2889 ) ;
  assign n2891 = n2660 ^ n1522 ^ n749 ;
  assign n2892 = x127 & n566 ;
  assign n2893 = n2892 ^ n2874 ^ 1'b0 ;
  assign n2894 = n2893 ^ n1244 ^ 1'b0 ;
  assign n2895 = n2894 ^ n2868 ^ n413 ;
  assign n2896 = ( n536 & ~n554 ) | ( n536 & n1785 ) | ( ~n554 & n1785 ) ;
  assign n2897 = n2323 ^ n2118 ^ n879 ;
  assign n2898 = n2897 ^ n885 ^ 1'b0 ;
  assign n2899 = ~n755 & n2038 ;
  assign n2900 = n136 & n2899 ;
  assign n2901 = n1200 & ~n1511 ;
  assign n2902 = ~n670 & n2901 ;
  assign n2903 = n2902 ^ x4 ^ 1'b0 ;
  assign n2904 = n2334 | n2903 ;
  assign n2905 = n433 ^ n284 ^ 1'b0 ;
  assign n2906 = ~n1748 & n2905 ;
  assign n2907 = n2906 ^ n880 ^ n879 ;
  assign n2908 = n221 & n715 ;
  assign n2909 = n555 & n2908 ;
  assign n2910 = ( n530 & n795 ) | ( n530 & n1869 ) | ( n795 & n1869 ) ;
  assign n2911 = n2895 ^ n1116 ^ 1'b0 ;
  assign n2912 = n2910 & n2911 ;
  assign n2913 = n705 ^ n433 ^ 1'b0 ;
  assign n2914 = n2110 ^ n654 ^ 1'b0 ;
  assign n2915 = n2913 & n2914 ;
  assign n2924 = ( n2089 & n2169 ) | ( n2089 & ~n2293 ) | ( n2169 & ~n2293 ) ;
  assign n2916 = n1011 | n1054 ;
  assign n2917 = n2916 ^ n1302 ^ 1'b0 ;
  assign n2918 = x61 & ~n1764 ;
  assign n2919 = n2918 ^ n1871 ^ 1'b0 ;
  assign n2920 = n444 & n2919 ;
  assign n2921 = n2920 ^ n209 ^ 1'b0 ;
  assign n2922 = n2921 ^ x15 ^ 1'b0 ;
  assign n2923 = n2917 | n2922 ;
  assign n2925 = n2924 ^ n2923 ^ 1'b0 ;
  assign n2926 = n2484 | n2925 ;
  assign n2927 = n1378 ^ n653 ^ n366 ;
  assign n2928 = n2927 ^ n2780 ^ n584 ;
  assign n2929 = n2349 ^ n1329 ^ n1297 ;
  assign n2930 = ( x14 & n209 ) | ( x14 & n987 ) | ( n209 & n987 ) ;
  assign n2931 = n845 ^ n285 ^ 1'b0 ;
  assign n2932 = n142 & ~n2931 ;
  assign n2933 = n2932 ^ x52 ^ 1'b0 ;
  assign n2934 = ~n536 & n2933 ;
  assign n2935 = n2930 & ~n2934 ;
  assign n2936 = n673 & ~n779 ;
  assign n2937 = n1240 & n2936 ;
  assign n2938 = n1294 & ~n2937 ;
  assign n2939 = n2938 ^ n2095 ^ 1'b0 ;
  assign n2940 = n1487 ^ n528 ^ 1'b0 ;
  assign n2941 = x61 & ~n779 ;
  assign n2942 = n1238 & n2941 ;
  assign n2943 = n1689 & n2813 ;
  assign n2944 = ~n2702 & n2943 ;
  assign n2945 = n2092 ^ n1140 ^ n593 ;
  assign n2946 = ( n313 & n1445 ) | ( n313 & ~n2945 ) | ( n1445 & ~n2945 ) ;
  assign n2952 = ( n1181 & n1985 ) | ( n1181 & n2044 ) | ( n1985 & n2044 ) ;
  assign n2953 = ~n1499 & n2952 ;
  assign n2954 = n2953 ^ n1240 ^ 1'b0 ;
  assign n2948 = ( n697 & n998 ) | ( n697 & ~n2297 ) | ( n998 & ~n2297 ) ;
  assign n2947 = n2884 ^ n2204 ^ 1'b0 ;
  assign n2949 = n2948 ^ n2947 ^ 1'b0 ;
  assign n2950 = ~x13 & n2949 ;
  assign n2951 = ~n915 & n2950 ;
  assign n2955 = n2954 ^ n2951 ^ 1'b0 ;
  assign n2956 = n2435 & ~n2955 ;
  assign n2957 = n1538 ^ n828 ^ 1'b0 ;
  assign n2958 = x83 & ~n2957 ;
  assign n2959 = ~n304 & n2958 ;
  assign n2960 = n836 & ~n2959 ;
  assign n2961 = ( n332 & ~n753 ) | ( n332 & n2960 ) | ( ~n753 & n2960 ) ;
  assign n2962 = n962 ^ n686 ^ n463 ;
  assign n2963 = n162 & n920 ;
  assign n2964 = n904 & n2963 ;
  assign n2965 = ( n370 & n571 ) | ( n370 & n808 ) | ( n571 & n808 ) ;
  assign n2966 = x17 & n571 ;
  assign n2967 = n2965 & n2966 ;
  assign n2968 = ~n2964 & n2967 ;
  assign n2969 = ( ~n1402 & n2962 ) | ( ~n1402 & n2968 ) | ( n2962 & n2968 ) ;
  assign n2970 = n1362 | n1398 ;
  assign n2971 = n2407 & ~n2970 ;
  assign n2972 = n2576 | n2971 ;
  assign n2973 = n579 | n2879 ;
  assign n2974 = n2973 ^ n1199 ^ 1'b0 ;
  assign n2975 = x33 & ~n360 ;
  assign n2976 = n2975 ^ n2125 ^ 1'b0 ;
  assign n2977 = n665 ^ n537 ^ 1'b0 ;
  assign n2978 = n1353 | n2977 ;
  assign n2979 = n1695 & ~n2978 ;
  assign n2980 = n2979 ^ n2072 ^ n424 ;
  assign n2981 = n2976 & ~n2980 ;
  assign n2982 = ( ~n694 & n893 ) | ( ~n694 & n1438 ) | ( n893 & n1438 ) ;
  assign n2983 = n1139 | n2188 ;
  assign n2984 = n2982 | n2983 ;
  assign n2988 = n2882 ^ n1542 ^ n368 ;
  assign n2985 = n1476 ^ n844 ^ n403 ;
  assign n2986 = n629 ^ n528 ^ 1'b0 ;
  assign n2987 = ~n2985 & n2986 ;
  assign n2989 = n2988 ^ n2987 ^ 1'b0 ;
  assign n2990 = n303 | n515 ;
  assign n2991 = ( n1240 & n2880 ) | ( n1240 & n2990 ) | ( n2880 & n2990 ) ;
  assign n2992 = n1888 ^ n701 ^ 1'b0 ;
  assign n2993 = n2992 ^ n985 ^ 1'b0 ;
  assign n2994 = n542 | n2972 ;
  assign n2995 = n737 | n2994 ;
  assign n2996 = n836 ^ n548 ^ 1'b0 ;
  assign n2997 = ~n1785 & n2996 ;
  assign n2998 = n2997 ^ n551 ^ 1'b0 ;
  assign n2999 = n427 | n2998 ;
  assign n3000 = n421 ^ n358 ^ 1'b0 ;
  assign n3001 = ~n2999 & n3000 ;
  assign n3002 = n1175 & ~n3001 ;
  assign n3003 = n531 | n905 ;
  assign n3004 = n2638 | n2860 ;
  assign n3005 = n1417 | n3004 ;
  assign n3006 = ( ~n2651 & n3003 ) | ( ~n2651 & n3005 ) | ( n3003 & n3005 ) ;
  assign n3007 = ~n2862 & n3006 ;
  assign n3008 = n1586 ^ n1137 ^ 1'b0 ;
  assign n3009 = ~n1483 & n3008 ;
  assign n3010 = n579 & n3009 ;
  assign n3011 = ( n1292 & n1747 ) | ( n1292 & ~n2025 ) | ( n1747 & ~n2025 ) ;
  assign n3012 = n2009 ^ n1617 ^ n246 ;
  assign n3013 = n1246 | n2375 ;
  assign n3016 = n609 | n898 ;
  assign n3014 = n494 ^ x73 ^ 1'b0 ;
  assign n3015 = n716 & ~n3014 ;
  assign n3017 = n3016 ^ n3015 ^ n510 ;
  assign n3018 = ~x0 & n1288 ;
  assign n3019 = ~n1152 & n3018 ;
  assign n3020 = n3017 | n3019 ;
  assign n3023 = ~n381 & n741 ;
  assign n3021 = n1908 ^ n1004 ^ 1'b0 ;
  assign n3022 = n2524 & ~n3021 ;
  assign n3024 = n3023 ^ n3022 ^ 1'b0 ;
  assign n3025 = n2128 | n3024 ;
  assign n3026 = ( n272 & n1124 ) | ( n272 & ~n1389 ) | ( n1124 & ~n1389 ) ;
  assign n3027 = n1911 ^ n343 ^ 1'b0 ;
  assign n3028 = n3026 & ~n3027 ;
  assign n3029 = n3028 ^ n1266 ^ 1'b0 ;
  assign n3030 = ( ~n729 & n1023 ) | ( ~n729 & n1764 ) | ( n1023 & n1764 ) ;
  assign n3031 = n3030 ^ n1329 ^ 1'b0 ;
  assign n3032 = n1489 & ~n3031 ;
  assign n3033 = n946 | n1714 ;
  assign n3034 = n1170 ^ n918 ^ x32 ;
  assign n3035 = ( n1554 & n1984 ) | ( n1554 & n3034 ) | ( n1984 & n3034 ) ;
  assign n3036 = n389 & ~n1129 ;
  assign n3037 = n797 & n3036 ;
  assign n3038 = ~n148 & n3037 ;
  assign n3039 = n1268 ^ n606 ^ 1'b0 ;
  assign n3040 = n3038 & ~n3039 ;
  assign n3041 = n3040 ^ n2891 ^ n1353 ;
  assign n3042 = n229 & n2402 ;
  assign n3043 = n3041 | n3042 ;
  assign n3044 = n2420 ^ n357 ^ 1'b0 ;
  assign n3045 = x117 & ~n931 ;
  assign n3046 = n1690 | n3045 ;
  assign n3047 = ( ~n1882 & n2827 ) | ( ~n1882 & n3046 ) | ( n2827 & n3046 ) ;
  assign n3048 = n1171 & n1248 ;
  assign n3049 = n865 & ~n3048 ;
  assign n3050 = n1012 ^ n675 ^ x84 ;
  assign n3051 = n3050 ^ x113 ^ 1'b0 ;
  assign n3052 = x1 | n3051 ;
  assign n3053 = n3052 ^ n2258 ^ 1'b0 ;
  assign n3054 = n508 ^ x113 ^ 1'b0 ;
  assign n3055 = n951 & n2457 ;
  assign n3056 = n3055 ^ n1992 ^ 1'b0 ;
  assign n3057 = ~n726 & n1298 ;
  assign n3058 = n3057 ^ n1137 ^ 1'b0 ;
  assign n3059 = n3058 ^ n575 ^ n207 ;
  assign n3060 = n1778 ^ n1521 ^ 1'b0 ;
  assign n3061 = n142 & n184 ;
  assign n3062 = ~n1177 & n3061 ;
  assign n3063 = x45 & ~n1341 ;
  assign n3064 = n2363 & n3063 ;
  assign n3065 = n3064 ^ n1445 ^ 1'b0 ;
  assign n3066 = n1713 | n3065 ;
  assign n3067 = n1093 | n1341 ;
  assign n3068 = n259 | n3067 ;
  assign n3069 = n2243 ^ n1455 ^ 1'b0 ;
  assign n3070 = n1350 & n3069 ;
  assign n3071 = ~n1523 & n2524 ;
  assign n3072 = n3071 ^ n2089 ^ 1'b0 ;
  assign n3073 = n761 | n1308 ;
  assign n3074 = n3072 & ~n3073 ;
  assign n3075 = n3074 ^ n1470 ^ 1'b0 ;
  assign n3076 = n2054 & n3075 ;
  assign n3081 = n2571 | n2833 ;
  assign n3082 = n3081 ^ n1508 ^ 1'b0 ;
  assign n3083 = n3082 ^ n911 ^ n901 ;
  assign n3077 = n1160 ^ x93 ^ x51 ;
  assign n3078 = ~n319 & n3077 ;
  assign n3079 = n3078 ^ n191 ^ 1'b0 ;
  assign n3080 = n3079 ^ n2375 ^ 1'b0 ;
  assign n3084 = n3083 ^ n3080 ^ n823 ;
  assign n3085 = x65 & ~n696 ;
  assign n3086 = ~n805 & n3085 ;
  assign n3087 = ~n410 & n1309 ;
  assign n3088 = n3086 & n3087 ;
  assign n3089 = n1702 & ~n3088 ;
  assign n3090 = n2806 & n3089 ;
  assign n3091 = n2128 & ~n3090 ;
  assign n3092 = n2029 ^ n1487 ^ n1227 ;
  assign n3095 = ( ~n350 & n716 ) | ( ~n350 & n1252 ) | ( n716 & n1252 ) ;
  assign n3096 = n3095 ^ n562 ^ x0 ;
  assign n3093 = n2431 ^ n1473 ^ n1376 ;
  assign n3094 = n1776 & n3093 ;
  assign n3097 = n3096 ^ n3094 ^ 1'b0 ;
  assign n3098 = n246 & ~n3097 ;
  assign n3099 = n995 & ~n2404 ;
  assign n3100 = n3098 & n3099 ;
  assign n3110 = n1012 | n1456 ;
  assign n3111 = n3110 ^ n1222 ^ 1'b0 ;
  assign n3112 = n2018 & n3111 ;
  assign n3113 = n3112 ^ n142 ^ 1'b0 ;
  assign n3105 = x22 & ~n2990 ;
  assign n3106 = n3105 ^ x73 ^ 1'b0 ;
  assign n3107 = n422 & n530 ;
  assign n3108 = n3106 & n3107 ;
  assign n3101 = n300 ^ n148 ^ 1'b0 ;
  assign n3102 = n843 | n3101 ;
  assign n3103 = n3102 ^ n1331 ^ 1'b0 ;
  assign n3104 = n3103 ^ n2383 ^ n1594 ;
  assign n3109 = n3108 ^ n3104 ^ n2307 ;
  assign n3114 = n3113 ^ n3109 ^ n2597 ;
  assign n3115 = n2177 & n2458 ;
  assign n3116 = n3115 ^ n1776 ^ 1'b0 ;
  assign n3117 = ~n1035 & n1543 ;
  assign n3118 = n3116 & ~n3117 ;
  assign n3119 = n2368 ^ n1538 ^ 1'b0 ;
  assign n3122 = ( n787 & ~n849 ) | ( n787 & n1430 ) | ( ~n849 & n1430 ) ;
  assign n3123 = n2111 & n3122 ;
  assign n3124 = n2064 ^ n1962 ^ 1'b0 ;
  assign n3125 = ~n3123 & n3124 ;
  assign n3120 = n345 | n704 ;
  assign n3121 = n2647 & n3120 ;
  assign n3126 = n3125 ^ n3121 ^ 1'b0 ;
  assign n3127 = n1418 ^ n1284 ^ n1168 ;
  assign n3128 = ( ~n493 & n1709 ) | ( ~n493 & n1715 ) | ( n1709 & n1715 ) ;
  assign n3129 = n2513 | n3054 ;
  assign n3130 = n1335 ^ n1012 ^ 1'b0 ;
  assign n3131 = n1129 | n2530 ;
  assign n3132 = n3131 ^ n2018 ^ 1'b0 ;
  assign n3133 = ~n1781 & n3132 ;
  assign n3134 = ~n2669 & n3133 ;
  assign n3135 = n3134 ^ n2089 ^ 1'b0 ;
  assign n3136 = n3130 & ~n3135 ;
  assign n3137 = x40 & x114 ;
  assign n3138 = ~n918 & n3137 ;
  assign n3139 = n211 | n3138 ;
  assign n3140 = ( n1047 & n2494 ) | ( n1047 & ~n2917 ) | ( n2494 & ~n2917 ) ;
  assign n3141 = n2352 ^ n1230 ^ 1'b0 ;
  assign n3142 = n2107 ^ n1791 ^ x111 ;
  assign n3143 = ( ~x59 & n266 ) | ( ~x59 & n665 ) | ( n266 & n665 ) ;
  assign n3144 = n1709 ^ n1591 ^ 1'b0 ;
  assign n3145 = n877 & n3144 ;
  assign n3146 = n3145 ^ n709 ^ 1'b0 ;
  assign n3147 = ( n292 & n3143 ) | ( n292 & ~n3146 ) | ( n3143 & ~n3146 ) ;
  assign n3148 = n2724 & n3147 ;
  assign n3149 = n3148 ^ n944 ^ 1'b0 ;
  assign n3150 = ~n138 & n827 ;
  assign n3154 = n2889 ^ n2384 ^ 1'b0 ;
  assign n3151 = n2270 & ~n2930 ;
  assign n3152 = ~n2849 & n3151 ;
  assign n3153 = n322 | n3152 ;
  assign n3155 = n3154 ^ n3153 ^ 1'b0 ;
  assign n3156 = n274 | n845 ;
  assign n3157 = n3156 ^ n160 ^ 1'b0 ;
  assign n3158 = n2929 & n3157 ;
  assign n3159 = x52 & ~x117 ;
  assign n3160 = ( ~n209 & n518 ) | ( ~n209 & n1444 ) | ( n518 & n1444 ) ;
  assign n3161 = ~n2086 & n3160 ;
  assign n3162 = n2411 & n3161 ;
  assign n3163 = n3162 ^ n2992 ^ n2976 ;
  assign n3164 = ( n1738 & n2077 ) | ( n1738 & ~n3163 ) | ( n2077 & ~n3163 ) ;
  assign n3165 = x89 & n3164 ;
  assign n3166 = n219 & n3165 ;
  assign n3167 = n1990 ^ n740 ^ 1'b0 ;
  assign n3168 = n1510 & ~n3167 ;
  assign n3169 = n3168 ^ n963 ^ 1'b0 ;
  assign n3170 = n3169 ^ n2651 ^ 1'b0 ;
  assign n3171 = n3119 & n3170 ;
  assign n3172 = ( n541 & ~n1651 ) | ( n541 & n2540 ) | ( ~n1651 & n2540 ) ;
  assign n3173 = ( n2062 & n2195 ) | ( n2062 & ~n3172 ) | ( n2195 & ~n3172 ) ;
  assign n3174 = n2905 ^ x54 ^ 1'b0 ;
  assign n3175 = n3174 ^ n2829 ^ 1'b0 ;
  assign n3176 = n1882 | n3175 ;
  assign n3177 = n2423 ^ n1280 ^ 1'b0 ;
  assign n3178 = n1697 | n3177 ;
  assign n3179 = ( x43 & ~n942 ) | ( x43 & n2519 ) | ( ~n942 & n2519 ) ;
  assign n3180 = n1089 & n3179 ;
  assign n3181 = n3180 ^ n2158 ^ n1548 ;
  assign n3182 = n1682 ^ n681 ^ 1'b0 ;
  assign n3183 = n2869 ^ n755 ^ 1'b0 ;
  assign n3184 = n3182 & n3183 ;
  assign n3185 = n2937 ^ n586 ^ 1'b0 ;
  assign n3186 = n2987 ^ n2301 ^ n168 ;
  assign n3189 = n697 & n2380 ;
  assign n3190 = n1582 | n3189 ;
  assign n3187 = n2440 ^ n1522 ^ 1'b0 ;
  assign n3188 = ~n2014 & n3187 ;
  assign n3191 = n3190 ^ n3188 ^ 1'b0 ;
  assign n3192 = n2420 ^ n630 ^ 1'b0 ;
  assign n3195 = n181 & ~n2133 ;
  assign n3193 = ( x87 & n211 ) | ( x87 & n2334 ) | ( n211 & n2334 ) ;
  assign n3194 = ~n834 & n3193 ;
  assign n3196 = n3195 ^ n3194 ^ n1718 ;
  assign n3197 = n506 | n2124 ;
  assign n3198 = n3197 ^ n1281 ^ 1'b0 ;
  assign n3201 = n2192 ^ n950 ^ 1'b0 ;
  assign n3202 = n2095 | n3201 ;
  assign n3199 = n246 & n2837 ;
  assign n3200 = n2772 & ~n3199 ;
  assign n3203 = n3202 ^ n3200 ^ 1'b0 ;
  assign n3204 = n2931 ^ n1973 ^ 1'b0 ;
  assign n3205 = n139 & ~n3204 ;
  assign n3212 = n684 & ~n1586 ;
  assign n3213 = ~n452 & n3212 ;
  assign n3214 = n3213 ^ n2927 ^ 1'b0 ;
  assign n3208 = n1078 & ~n1905 ;
  assign n3209 = n3208 ^ n563 ^ 1'b0 ;
  assign n3210 = n1379 | n3209 ;
  assign n3211 = n1644 & ~n3210 ;
  assign n3206 = n1485 ^ n1071 ^ 1'b0 ;
  assign n3207 = n2506 & ~n3206 ;
  assign n3215 = n3214 ^ n3211 ^ n3207 ;
  assign n3216 = x8 & ~n186 ;
  assign n3217 = n3216 ^ x2 ^ 1'b0 ;
  assign n3218 = n412 & ~n3217 ;
  assign n3219 = n3218 ^ n2069 ^ n1496 ;
  assign n3220 = n236 ^ n160 ^ 1'b0 ;
  assign n3221 = n3132 & n3220 ;
  assign n3222 = ( ~n1046 & n1496 ) | ( ~n1046 & n3221 ) | ( n1496 & n3221 ) ;
  assign n3223 = n1360 & ~n3222 ;
  assign n3224 = n3223 ^ n170 ^ 1'b0 ;
  assign n3225 = n2974 ^ n904 ^ 1'b0 ;
  assign n3226 = n1414 ^ n1012 ^ 1'b0 ;
  assign n3227 = x57 & n3226 ;
  assign n3228 = n3225 & ~n3227 ;
  assign n3229 = n1351 & n3228 ;
  assign n3230 = ~n686 & n3229 ;
  assign n3231 = n736 ^ n434 ^ n236 ;
  assign n3232 = n3231 ^ n1971 ^ 1'b0 ;
  assign n3233 = n677 & ~n1937 ;
  assign n3234 = n358 & n3233 ;
  assign n3235 = n1904 ^ n1723 ^ 1'b0 ;
  assign n3236 = ~n1145 & n3235 ;
  assign n3237 = n1495 ^ n410 ^ 1'b0 ;
  assign n3238 = n3090 ^ x116 ^ 1'b0 ;
  assign n3239 = n1410 ^ n866 ^ 1'b0 ;
  assign n3240 = ( n635 & ~n1888 ) | ( n635 & n2434 ) | ( ~n1888 & n2434 ) ;
  assign n3241 = n285 & ~n3240 ;
  assign n3242 = n2406 ^ n433 ^ 1'b0 ;
  assign n3244 = ~n1276 & n1908 ;
  assign n3243 = n1455 | n3242 ;
  assign n3245 = n3244 ^ n3243 ^ 1'b0 ;
  assign n3246 = n2771 ^ n2723 ^ 1'b0 ;
  assign n3247 = ( n550 & ~n2984 ) | ( n550 & n3246 ) | ( ~n2984 & n3246 ) ;
  assign n3248 = ( n3242 & n3245 ) | ( n3242 & n3247 ) | ( n3245 & n3247 ) ;
  assign n3249 = n138 | n355 ;
  assign n3250 = n3249 ^ n1280 ^ 1'b0 ;
  assign n3251 = n3023 | n3250 ;
  assign n3252 = n3189 | n3251 ;
  assign n3253 = n962 & n3252 ;
  assign n3254 = n3253 ^ n2058 ^ 1'b0 ;
  assign n3255 = n3050 ^ n2038 ^ n227 ;
  assign n3256 = n723 & n3255 ;
  assign n3257 = n3256 ^ n2122 ^ 1'b0 ;
  assign n3258 = n2741 & ~n3257 ;
  assign n3259 = n1535 ^ n372 ^ 1'b0 ;
  assign n3260 = n2923 | n3259 ;
  assign n3261 = n1576 & ~n1831 ;
  assign n3262 = n3261 ^ n751 ^ 1'b0 ;
  assign n3263 = ( n2826 & n3260 ) | ( n2826 & n3262 ) | ( n3260 & n3262 ) ;
  assign n3264 = ( ~n295 & n1150 ) | ( ~n295 & n1703 ) | ( n1150 & n1703 ) ;
  assign n3269 = n818 ^ n661 ^ 1'b0 ;
  assign n3270 = n718 & ~n3269 ;
  assign n3268 = ~n177 & n1648 ;
  assign n3271 = n3270 ^ n3268 ^ 1'b0 ;
  assign n3272 = n3271 ^ n2930 ^ n903 ;
  assign n3273 = n3272 ^ n363 ^ 1'b0 ;
  assign n3274 = n934 & n3273 ;
  assign n3265 = n1814 ^ n1538 ^ n319 ;
  assign n3266 = n2320 & ~n3265 ;
  assign n3267 = n923 & n3266 ;
  assign n3275 = n3274 ^ n3267 ^ n1925 ;
  assign n3276 = ( n734 & n1475 ) | ( n734 & n2187 ) | ( n1475 & n2187 ) ;
  assign n3277 = ( ~n829 & n1960 ) | ( ~n829 & n2342 ) | ( n1960 & n2342 ) ;
  assign n3278 = n3277 ^ n799 ^ 1'b0 ;
  assign n3279 = ( n985 & n2602 ) | ( n985 & n3278 ) | ( n2602 & n3278 ) ;
  assign n3280 = n585 & n3279 ;
  assign n3281 = ~n2930 & n3280 ;
  assign n3282 = n2753 ^ n1874 ^ n1420 ;
  assign n3283 = n1487 ^ n1100 ^ 1'b0 ;
  assign n3284 = n2968 | n3283 ;
  assign n3285 = n616 & n1460 ;
  assign n3286 = ~n258 & n3285 ;
  assign n3287 = ( n1282 & n1350 ) | ( n1282 & ~n3286 ) | ( n1350 & ~n3286 ) ;
  assign n3288 = n1846 & n3287 ;
  assign n3289 = n3288 ^ n2364 ^ 1'b0 ;
  assign n3293 = ( n145 & n2128 ) | ( n145 & n2657 ) | ( n2128 & n2657 ) ;
  assign n3290 = ~n595 & n983 ;
  assign n3291 = ~n2344 & n3290 ;
  assign n3292 = n2995 & ~n3291 ;
  assign n3294 = n3293 ^ n3292 ^ 1'b0 ;
  assign n3295 = n911 | n1282 ;
  assign n3296 = n3295 ^ n1919 ^ 1'b0 ;
  assign n3297 = n3296 ^ n535 ^ x19 ;
  assign n3298 = n2945 & ~n3297 ;
  assign n3299 = n2859 ^ n1352 ^ 1'b0 ;
  assign n3300 = ~n1199 & n3299 ;
  assign n3301 = n2472 ^ n608 ^ 1'b0 ;
  assign n3302 = n2399 & n3301 ;
  assign n3303 = n3278 ^ n778 ^ 1'b0 ;
  assign n3304 = ~n2469 & n3303 ;
  assign n3305 = n510 & n3304 ;
  assign n3306 = n1653 ^ n744 ^ 1'b0 ;
  assign n3307 = ~n2333 & n3306 ;
  assign n3308 = n3307 ^ n3302 ^ n3196 ;
  assign n3309 = n1502 & n2604 ;
  assign n3310 = n1470 & n3309 ;
  assign n3311 = ( n1015 & ~n1586 ) | ( n1015 & n3278 ) | ( ~n1586 & n3278 ) ;
  assign n3312 = ~n3310 & n3311 ;
  assign n3313 = n740 & n2851 ;
  assign n3314 = n3313 ^ x28 ^ 1'b0 ;
  assign n3315 = ( n148 & n692 ) | ( n148 & n945 ) | ( n692 & n945 ) ;
  assign n3316 = n2246 ^ n1728 ^ 1'b0 ;
  assign n3317 = n3316 ^ n1138 ^ 1'b0 ;
  assign n3318 = n3015 ^ n2643 ^ 1'b0 ;
  assign n3319 = n736 ^ n266 ^ 1'b0 ;
  assign n3320 = n3319 ^ n380 ^ 1'b0 ;
  assign n3322 = n1365 & ~n1614 ;
  assign n3323 = n3322 ^ n212 ^ 1'b0 ;
  assign n3324 = n3323 ^ n1573 ^ 1'b0 ;
  assign n3325 = n3324 ^ n953 ^ 1'b0 ;
  assign n3326 = n1491 & ~n3325 ;
  assign n3321 = ~n154 & n3009 ;
  assign n3327 = n3326 ^ n3321 ^ 1'b0 ;
  assign n3328 = ~n817 & n2724 ;
  assign n3329 = n3327 & n3328 ;
  assign n3331 = ~n438 & n742 ;
  assign n3332 = ~n714 & n3331 ;
  assign n3330 = ( ~n778 & n1083 ) | ( ~n778 & n1133 ) | ( n1083 & n1133 ) ;
  assign n3333 = n3332 ^ n3330 ^ 1'b0 ;
  assign n3334 = x36 & ~n3333 ;
  assign n3335 = n1171 ^ n798 ^ 1'b0 ;
  assign n3336 = n160 & n732 ;
  assign n3337 = n3336 ^ n1084 ^ 1'b0 ;
  assign n3338 = ( n915 & ~n1529 ) | ( n915 & n3337 ) | ( ~n1529 & n3337 ) ;
  assign n3339 = n2999 ^ n2746 ^ n1913 ;
  assign n3340 = n3339 ^ n661 ^ n419 ;
  assign n3343 = n2196 ^ n1659 ^ 1'b0 ;
  assign n3344 = n1613 & ~n3343 ;
  assign n3345 = ~n520 & n3344 ;
  assign n3346 = n1817 | n3345 ;
  assign n3347 = n2651 & ~n3346 ;
  assign n3341 = ( n134 & ~n1139 ) | ( n134 & n1744 ) | ( ~n1139 & n1744 ) ;
  assign n3342 = n3341 ^ n828 ^ n227 ;
  assign n3348 = n3347 ^ n3342 ^ n699 ;
  assign n3352 = n1795 ^ n787 ^ 1'b0 ;
  assign n3349 = n2051 ^ n672 ^ 1'b0 ;
  assign n3350 = ( n1256 & n2146 ) | ( n1256 & n3349 ) | ( n2146 & n3349 ) ;
  assign n3351 = ~n2597 & n3350 ;
  assign n3353 = n3352 ^ n3351 ^ 1'b0 ;
  assign n3355 = ~n990 & n1894 ;
  assign n3357 = n1123 ^ n586 ^ n274 ;
  assign n3358 = n3357 ^ n1458 ^ n145 ;
  assign n3356 = n1069 ^ n399 ^ 1'b0 ;
  assign n3359 = n3358 ^ n3356 ^ 1'b0 ;
  assign n3360 = n3359 ^ n1924 ^ 1'b0 ;
  assign n3361 = n3355 & ~n3360 ;
  assign n3354 = n1832 | n2345 ;
  assign n3362 = n3361 ^ n3354 ^ 1'b0 ;
  assign n3363 = ( n1384 & n2382 ) | ( n1384 & ~n2466 ) | ( n2382 & ~n2466 ) ;
  assign n3364 = n2826 & n3363 ;
  assign n3365 = n1428 | n3218 ;
  assign n3366 = n3365 ^ n1036 ^ n487 ;
  assign n3367 = ( n2174 & n2813 ) | ( n2174 & ~n3366 ) | ( n2813 & ~n3366 ) ;
  assign n3368 = n146 & ~n1534 ;
  assign n3369 = n2370 ^ n958 ^ 1'b0 ;
  assign n3370 = ~n648 & n3369 ;
  assign n3371 = n3370 ^ n1933 ^ n1462 ;
  assign n3372 = ( n3011 & n3368 ) | ( n3011 & n3371 ) | ( n3368 & n3371 ) ;
  assign n3373 = n3372 ^ n2823 ^ n330 ;
  assign n3382 = ( n143 & n1354 ) | ( n143 & ~n2053 ) | ( n1354 & ~n2053 ) ;
  assign n3383 = ( n1812 & ~n2038 ) | ( n1812 & n3382 ) | ( ~n2038 & n3382 ) ;
  assign n3374 = n1501 ^ n427 ^ 1'b0 ;
  assign n3375 = x15 & ~n3374 ;
  assign n3376 = x108 & n1233 ;
  assign n3377 = n1548 | n2680 ;
  assign n3378 = n299 & ~n3377 ;
  assign n3379 = ( n1652 & ~n3376 ) | ( n1652 & n3378 ) | ( ~n3376 & n3378 ) ;
  assign n3380 = n3375 & n3379 ;
  assign n3381 = ~x3 & n3380 ;
  assign n3384 = n3383 ^ n3381 ^ n139 ;
  assign n3385 = ~n1020 & n1719 ;
  assign n3386 = n3385 ^ n2055 ^ 1'b0 ;
  assign n3387 = n3386 ^ n2467 ^ 1'b0 ;
  assign n3388 = n3387 ^ n576 ^ 1'b0 ;
  assign n3389 = n1102 & n3388 ;
  assign n3390 = ~n3384 & n3389 ;
  assign n3391 = n2538 ^ n1324 ^ 1'b0 ;
  assign n3392 = n1972 & n3391 ;
  assign n3393 = n1455 ^ n735 ^ 1'b0 ;
  assign n3394 = n3324 & ~n3357 ;
  assign n3395 = n164 & n3394 ;
  assign n3396 = ~n1271 & n3395 ;
  assign n3397 = ~n3393 & n3396 ;
  assign n3398 = n3397 ^ n3032 ^ 1'b0 ;
  assign n3399 = n2760 ^ x12 ^ 1'b0 ;
  assign n3400 = n1853 ^ n530 ^ 1'b0 ;
  assign n3401 = n2131 | n3400 ;
  assign n3402 = n2789 ^ n2388 ^ n1493 ;
  assign n3403 = n1789 & ~n3402 ;
  assign n3404 = n3403 ^ n916 ^ 1'b0 ;
  assign n3405 = n1320 | n3315 ;
  assign n3406 = n3405 ^ n800 ^ 1'b0 ;
  assign n3407 = n2323 ^ n1376 ^ n858 ;
  assign n3408 = n3407 ^ n2650 ^ 1'b0 ;
  assign n3409 = x30 & n1897 ;
  assign n3410 = n3408 & n3409 ;
  assign n3411 = n1703 | n3410 ;
  assign n3412 = n3411 ^ n1162 ^ 1'b0 ;
  assign n3413 = n3412 ^ n2982 ^ n1069 ;
  assign n3414 = n2105 ^ n1864 ^ 1'b0 ;
  assign n3415 = n3187 & n3414 ;
  assign n3416 = ~n2928 & n3415 ;
  assign n3417 = n3404 ^ n299 ^ 1'b0 ;
  assign n3419 = n1379 | n2568 ;
  assign n3420 = n1982 | n3419 ;
  assign n3418 = n293 & ~n1784 ;
  assign n3421 = n3420 ^ n3418 ^ n1356 ;
  assign n3429 = n271 & n904 ;
  assign n3422 = ~n620 & n2128 ;
  assign n3423 = n3422 ^ n945 ^ 1'b0 ;
  assign n3424 = n1907 & n3423 ;
  assign n3425 = n3424 ^ n178 ^ 1'b0 ;
  assign n3426 = n3034 | n3425 ;
  assign n3427 = n3426 ^ n690 ^ 1'b0 ;
  assign n3428 = x103 & ~n3427 ;
  assign n3430 = n3429 ^ n3428 ^ n1118 ;
  assign n3431 = n2663 | n2767 ;
  assign n3432 = n3431 ^ n2999 ^ 1'b0 ;
  assign n3433 = n2470 | n3432 ;
  assign n3434 = n2026 ^ n229 ^ 1'b0 ;
  assign n3435 = n1890 ^ n1573 ^ 1'b0 ;
  assign n3436 = ~n2023 & n3435 ;
  assign n3437 = n3436 ^ n1331 ^ 1'b0 ;
  assign n3438 = n3434 & n3437 ;
  assign n3439 = x12 & n3438 ;
  assign n3440 = n3439 ^ n746 ^ 1'b0 ;
  assign n3441 = n3440 ^ n1342 ^ 1'b0 ;
  assign n3442 = n1389 ^ n802 ^ n607 ;
  assign n3443 = n2182 ^ n1033 ^ 1'b0 ;
  assign n3444 = n243 & n3443 ;
  assign n3445 = ( n1039 & n3442 ) | ( n1039 & ~n3444 ) | ( n3442 & ~n3444 ) ;
  assign n3446 = ( n1252 & n1552 ) | ( n1252 & n3445 ) | ( n1552 & n3445 ) ;
  assign n3447 = n2074 & n2521 ;
  assign n3448 = n3146 ^ n1843 ^ n478 ;
  assign n3449 = n3447 & ~n3448 ;
  assign n3450 = n1060 ^ n254 ^ 1'b0 ;
  assign n3451 = n3450 ^ n1795 ^ 1'b0 ;
  assign n3452 = n1673 | n3451 ;
  assign n3453 = n737 ^ x61 ^ 1'b0 ;
  assign n3454 = n322 & ~n3453 ;
  assign n3455 = ~n811 & n3454 ;
  assign n3457 = n310 ^ x86 ^ 1'b0 ;
  assign n3456 = n1259 ^ n1067 ^ 1'b0 ;
  assign n3458 = n3457 ^ n3456 ^ 1'b0 ;
  assign n3459 = n2498 & n3458 ;
  assign n3460 = ~n1340 & n1442 ;
  assign n3461 = n3460 ^ n3381 ^ 1'b0 ;
  assign n3462 = n3461 ^ n911 ^ 1'b0 ;
  assign n3463 = n697 & ~n3462 ;
  assign n3464 = ~n2976 & n3463 ;
  assign n3465 = ~n920 & n3464 ;
  assign n3466 = n3453 ^ n2256 ^ 1'b0 ;
  assign n3467 = n3452 ^ n2018 ^ 1'b0 ;
  assign n3468 = ( ~n1290 & n1535 ) | ( ~n1290 & n1952 ) | ( n1535 & n1952 ) ;
  assign n3469 = ( ~n3149 & n3291 ) | ( ~n3149 & n3468 ) | ( n3291 & n3468 ) ;
  assign n3470 = n3381 ^ n936 ^ 1'b0 ;
  assign n3471 = n1643 ^ n1091 ^ n576 ;
  assign n3472 = n963 ^ n254 ^ 1'b0 ;
  assign n3473 = ~n929 & n3472 ;
  assign n3474 = n3473 ^ n1378 ^ 1'b0 ;
  assign n3475 = n1764 ^ n403 ^ 1'b0 ;
  assign n3476 = n798 & ~n3475 ;
  assign n3477 = n3476 ^ n1854 ^ n779 ;
  assign n3478 = ( n589 & n1306 ) | ( n589 & ~n3477 ) | ( n1306 & ~n3477 ) ;
  assign n3479 = ( n1355 & n1768 ) | ( n1355 & ~n2407 ) | ( n1768 & ~n2407 ) ;
  assign n3481 = x31 & ~n1896 ;
  assign n3482 = n1674 & n3481 ;
  assign n3480 = n2171 & n2189 ;
  assign n3483 = n3482 ^ n3480 ^ 1'b0 ;
  assign n3484 = n2184 ^ n325 ^ 1'b0 ;
  assign n3485 = n639 & ~n1662 ;
  assign n3486 = n3485 ^ n1373 ^ 1'b0 ;
  assign n3487 = n2258 & n3486 ;
  assign n3488 = ~n3484 & n3487 ;
  assign n3489 = n463 & ~n1591 ;
  assign n3490 = n1997 & n3489 ;
  assign n3491 = ( ~x82 & n1066 ) | ( ~x82 & n3490 ) | ( n1066 & n3490 ) ;
  assign n3492 = ~n941 & n1744 ;
  assign n3493 = n3491 & n3492 ;
  assign n3494 = ( n1435 & n1971 ) | ( n1435 & n3425 ) | ( n1971 & n3425 ) ;
  assign n3495 = n1834 ^ n491 ^ 1'b0 ;
  assign n3496 = ~n308 & n3495 ;
  assign n3497 = n1937 | n2961 ;
  assign n3498 = n227 & ~n3497 ;
  assign n3499 = ( n389 & ~n2837 ) | ( n389 & n3498 ) | ( ~n2837 & n3498 ) ;
  assign n3500 = n3499 ^ n1622 ^ 1'b0 ;
  assign n3501 = n3106 | n3500 ;
  assign n3502 = n2364 ^ n1523 ^ 1'b0 ;
  assign n3503 = ~n1006 & n3502 ;
  assign n3504 = n3503 ^ n561 ^ 1'b0 ;
  assign n3508 = ~n1447 & n2370 ;
  assign n3505 = n432 & ~n485 ;
  assign n3506 = n397 | n1447 ;
  assign n3507 = ( ~n2174 & n3505 ) | ( ~n2174 & n3506 ) | ( n3505 & n3506 ) ;
  assign n3509 = n3508 ^ n3507 ^ x35 ;
  assign n3513 = n543 | n1788 ;
  assign n3510 = n2200 ^ n474 ^ 1'b0 ;
  assign n3511 = ~n822 & n3510 ;
  assign n3512 = ( x57 & ~n1943 ) | ( x57 & n3511 ) | ( ~n1943 & n3511 ) ;
  assign n3514 = n3513 ^ n3512 ^ 1'b0 ;
  assign n3515 = x71 & n3459 ;
  assign n3516 = n805 & ~n2824 ;
  assign n3517 = n1512 & n3516 ;
  assign n3518 = n1083 & ~n1107 ;
  assign n3519 = n3518 ^ x4 ^ 1'b0 ;
  assign n3520 = n668 ^ n172 ^ 1'b0 ;
  assign n3521 = ~n157 & n3520 ;
  assign n3522 = n3386 & ~n3521 ;
  assign n3523 = n1041 & ~n3522 ;
  assign n3524 = n3523 ^ n872 ^ n849 ;
  assign n3525 = ( ~x32 & n195 ) | ( ~x32 & n402 ) | ( n195 & n402 ) ;
  assign n3526 = n3525 ^ n2521 ^ n209 ;
  assign n3527 = n2822 & ~n3013 ;
  assign n3528 = n1320 & n3527 ;
  assign n3529 = n2066 ^ n726 ^ x55 ;
  assign n3530 = ( n712 & n1881 ) | ( n712 & ~n3529 ) | ( n1881 & ~n3529 ) ;
  assign n3536 = n1546 ^ n485 ^ 1'b0 ;
  assign n3537 = n1135 | n3536 ;
  assign n3533 = n1778 ^ n1455 ^ 1'b0 ;
  assign n3534 = n3533 ^ n162 ^ 1'b0 ;
  assign n3535 = n344 | n3534 ;
  assign n3538 = n3537 ^ n3535 ^ 1'b0 ;
  assign n3539 = n3538 ^ n1930 ^ 1'b0 ;
  assign n3531 = ~n929 & n1291 ;
  assign n3532 = n630 & n3531 ;
  assign n3540 = n3539 ^ n3532 ^ 1'b0 ;
  assign n3541 = ~n2613 & n3540 ;
  assign n3542 = ~n701 & n3240 ;
  assign n3543 = ~n1576 & n3542 ;
  assign n3544 = n992 ^ n688 ^ 1'b0 ;
  assign n3545 = n938 | n3544 ;
  assign n3546 = n3545 ^ x113 ^ 1'b0 ;
  assign n3547 = n1770 ^ n1371 ^ 1'b0 ;
  assign n3548 = ~n1575 & n3547 ;
  assign n3549 = ( ~n1386 & n1760 ) | ( ~n1386 & n2657 ) | ( n1760 & n2657 ) ;
  assign n3550 = n2680 ^ x14 ^ x13 ;
  assign n3551 = ( n334 & n3549 ) | ( n334 & n3550 ) | ( n3549 & n3550 ) ;
  assign n3552 = n785 | n1418 ;
  assign n3553 = n887 & n1234 ;
  assign n3554 = ( n554 & n726 ) | ( n554 & ~n1747 ) | ( n726 & ~n1747 ) ;
  assign n3555 = n1003 ^ n932 ^ 1'b0 ;
  assign n3556 = n1858 | n3555 ;
  assign n3557 = n3556 ^ n893 ^ 1'b0 ;
  assign n3558 = ~n822 & n3557 ;
  assign n3559 = ( n251 & n1323 ) | ( n251 & ~n3558 ) | ( n1323 & ~n3558 ) ;
  assign n3560 = ( n3553 & n3554 ) | ( n3553 & n3559 ) | ( n3554 & n3559 ) ;
  assign n3561 = n1573 | n1766 ;
  assign n3562 = n1242 ^ n133 ^ 1'b0 ;
  assign n3563 = ~n165 & n3562 ;
  assign n3566 = n2149 ^ n432 ^ 1'b0 ;
  assign n3567 = n3566 ^ n2246 ^ n356 ;
  assign n3564 = n2965 ^ n1931 ^ n219 ;
  assign n3565 = ~n693 & n3564 ;
  assign n3568 = n3567 ^ n3565 ^ x30 ;
  assign n3569 = x75 & n3568 ;
  assign n3570 = ~n3563 & n3569 ;
  assign n3571 = n247 | n1347 ;
  assign n3572 = n298 & ~n3571 ;
  assign n3573 = x52 & ~n3572 ;
  assign n3574 = n3573 ^ n995 ^ 1'b0 ;
  assign n3575 = n3574 ^ n3154 ^ 1'b0 ;
  assign n3576 = n876 & n1764 ;
  assign n3577 = n3576 ^ n2148 ^ 1'b0 ;
  assign n3578 = n1150 | n3577 ;
  assign n3580 = n212 & n1514 ;
  assign n3581 = n3580 ^ n1108 ^ 1'b0 ;
  assign n3579 = n1481 | n1684 ;
  assign n3582 = n3581 ^ n3579 ^ 1'b0 ;
  assign n3583 = n1779 & n3582 ;
  assign n3584 = n3583 ^ n1305 ^ n1298 ;
  assign n3585 = n3584 ^ n1828 ^ 1'b0 ;
  assign n3586 = n323 | n3585 ;
  assign n3587 = ( n578 & n1034 ) | ( n578 & ~n3586 ) | ( n1034 & ~n3586 ) ;
  assign n3588 = n335 & ~n1643 ;
  assign n3589 = n1290 & n3588 ;
  assign n3590 = n3589 ^ n848 ^ 1'b0 ;
  assign n3591 = n918 & ~n3590 ;
  assign n3592 = ( n184 & n1347 ) | ( n184 & n3591 ) | ( n1347 & n3591 ) ;
  assign n3593 = n3592 ^ n2049 ^ 1'b0 ;
  assign n3594 = n2475 & n3593 ;
  assign n3595 = n1170 ^ x91 ^ 1'b0 ;
  assign n3596 = n3595 ^ n339 ^ 1'b0 ;
  assign n3597 = ~n3365 & n3596 ;
  assign n3598 = n2131 & n2399 ;
  assign n3599 = ( n836 & n1789 ) | ( n836 & n3106 ) | ( n1789 & n3106 ) ;
  assign n3603 = n2875 ^ x36 ^ 1'b0 ;
  assign n3604 = ~n1545 & n3603 ;
  assign n3605 = n1784 ^ x101 ^ 1'b0 ;
  assign n3606 = n3604 & n3605 ;
  assign n3602 = n1138 & n3418 ;
  assign n3607 = n3606 ^ n3602 ^ 1'b0 ;
  assign n3600 = n285 | n903 ;
  assign n3601 = x34 & n3600 ;
  assign n3608 = n3607 ^ n3601 ^ 1'b0 ;
  assign n3609 = n3461 ^ n2450 ^ n718 ;
  assign n3610 = ( ~n489 & n1666 ) | ( ~n489 & n2748 ) | ( n1666 & n2748 ) ;
  assign n3611 = ( n146 & n3609 ) | ( n146 & n3610 ) | ( n3609 & n3610 ) ;
  assign n3612 = n2984 ^ x44 ^ 1'b0 ;
  assign n3613 = n1779 ^ n1104 ^ n920 ;
  assign n3614 = n2902 & n3613 ;
  assign n3615 = n1863 & n2767 ;
  assign n3620 = n2012 ^ n812 ^ x38 ;
  assign n3616 = n1167 ^ n299 ^ n148 ;
  assign n3617 = n307 ^ n143 ^ 1'b0 ;
  assign n3618 = ( n356 & n1470 ) | ( n356 & ~n3617 ) | ( n1470 & ~n3617 ) ;
  assign n3619 = ~n3616 & n3618 ;
  assign n3621 = n3620 ^ n3619 ^ 1'b0 ;
  assign n3622 = n2340 ^ n2081 ^ x63 ;
  assign n3623 = n1853 ^ n387 ^ 1'b0 ;
  assign n3624 = n2025 | n3623 ;
  assign n3625 = n3624 ^ n1171 ^ n221 ;
  assign n3626 = n3625 ^ n531 ^ 1'b0 ;
  assign n3627 = n563 ^ n221 ^ 1'b0 ;
  assign n3628 = ~n361 & n3627 ;
  assign n3629 = n3628 ^ n345 ^ 1'b0 ;
  assign n3642 = n478 & ~n594 ;
  assign n3643 = n1868 | n3642 ;
  assign n3644 = n3237 & ~n3643 ;
  assign n3645 = n3644 ^ n2169 ^ 1'b0 ;
  assign n3646 = n3645 ^ n870 ^ 1'b0 ;
  assign n3647 = n502 & n3646 ;
  assign n3639 = n1738 & ~n2233 ;
  assign n3640 = n3639 ^ n1078 ^ 1'b0 ;
  assign n3641 = n784 | n3640 ;
  assign n3648 = n3647 ^ n3641 ^ 1'b0 ;
  assign n3630 = ( n1034 & n1763 ) | ( n1034 & ~n2496 ) | ( n1763 & ~n2496 ) ;
  assign n3631 = n730 & n734 ;
  assign n3632 = ( n1023 & n3261 ) | ( n1023 & ~n3631 ) | ( n3261 & ~n3631 ) ;
  assign n3633 = n557 | n982 ;
  assign n3634 = x18 | n3633 ;
  assign n3635 = n1352 ^ n193 ^ 1'b0 ;
  assign n3636 = n3634 & ~n3635 ;
  assign n3637 = ( n2345 & n3116 ) | ( n2345 & n3636 ) | ( n3116 & n3636 ) ;
  assign n3638 = ( n3630 & n3632 ) | ( n3630 & ~n3637 ) | ( n3632 & ~n3637 ) ;
  assign n3649 = n3648 ^ n3638 ^ n2014 ;
  assign n3650 = x84 & ~n706 ;
  assign n3651 = ( n433 & n1025 ) | ( n433 & n1045 ) | ( n1025 & n1045 ) ;
  assign n3652 = n3650 & n3651 ;
  assign n3653 = ~n569 & n3125 ;
  assign n3654 = n3653 ^ n242 ^ 1'b0 ;
  assign n3655 = ~n355 & n732 ;
  assign n3656 = n220 | n3655 ;
  assign n3657 = x6 & ~n3656 ;
  assign n3658 = x56 & ~n3381 ;
  assign n3659 = ( n221 & n1014 ) | ( n221 & n2110 ) | ( n1014 & n2110 ) ;
  assign n3660 = n593 ^ x60 ^ 1'b0 ;
  assign n3661 = n3529 ^ n2193 ^ 1'b0 ;
  assign n3662 = n3050 & ~n3661 ;
  assign n3663 = n211 & n3662 ;
  assign n3664 = ( x76 & ~n3660 ) | ( x76 & n3663 ) | ( ~n3660 & n3663 ) ;
  assign n3665 = n2038 ^ n415 ^ 1'b0 ;
  assign n3666 = n3665 ^ n231 ^ 1'b0 ;
  assign n3667 = n589 | n1014 ;
  assign n3668 = n3667 ^ n2997 ^ 1'b0 ;
  assign n3669 = n1576 & ~n3668 ;
  assign n3670 = ~x0 & n850 ;
  assign n3671 = n3670 ^ n2006 ^ 1'b0 ;
  assign n3672 = n2680 ^ n1353 ^ 1'b0 ;
  assign n3673 = ~n2783 & n3672 ;
  assign n3674 = ~n801 & n3381 ;
  assign n3675 = n3674 ^ n1440 ^ 1'b0 ;
  assign n3676 = n1322 & ~n3675 ;
  assign n3677 = n2827 ^ n1211 ^ n509 ;
  assign n3678 = n411 & n1212 ;
  assign n3679 = ( n664 & ~n784 ) | ( n664 & n3678 ) | ( ~n784 & n3678 ) ;
  assign n3680 = n3679 ^ n3532 ^ 1'b0 ;
  assign n3681 = ~n2204 & n3680 ;
  assign n3682 = ( n553 & ~n1125 ) | ( n553 & n2581 ) | ( ~n1125 & n2581 ) ;
  assign n3683 = n2776 ^ n2478 ^ 1'b0 ;
  assign n3684 = n3682 | n3683 ;
  assign n3685 = n3684 ^ n3234 ^ 1'b0 ;
  assign n3686 = n3154 & n3685 ;
  assign n3690 = n251 & ~n2095 ;
  assign n3691 = ~n1501 & n3690 ;
  assign n3692 = n3691 ^ n2714 ^ 1'b0 ;
  assign n3693 = n1556 & n3692 ;
  assign n3687 = n2260 ^ n397 ^ 1'b0 ;
  assign n3688 = n2270 & n3687 ;
  assign n3689 = n319 | n3688 ;
  assign n3694 = n3693 ^ n3689 ^ n1714 ;
  assign n3695 = n3686 | n3694 ;
  assign n3696 = n3319 ^ n1997 ^ n154 ;
  assign n3697 = n3553 ^ n3345 ^ 1'b0 ;
  assign n3700 = n1993 & n2930 ;
  assign n3698 = ( n1069 & n1622 ) | ( n1069 & n2421 ) | ( n1622 & n2421 ) ;
  assign n3699 = n3698 ^ n2576 ^ n2211 ;
  assign n3701 = n3700 ^ n3699 ^ x70 ;
  assign n3702 = n3697 & ~n3701 ;
  assign n3703 = n3702 ^ n2486 ^ 1'b0 ;
  assign n3704 = n3703 ^ n2709 ^ n1483 ;
  assign n3705 = n2645 ^ n316 ^ 1'b0 ;
  assign n3706 = n3705 ^ n1470 ^ n425 ;
  assign n3707 = n1579 ^ n148 ^ 1'b0 ;
  assign n3708 = n727 | n1805 ;
  assign n3709 = x40 | n3708 ;
  assign n3710 = ( ~n2032 & n3707 ) | ( ~n2032 & n3709 ) | ( n3707 & n3709 ) ;
  assign n3711 = n3710 ^ n3607 ^ 1'b0 ;
  assign n3712 = n3121 ^ n2664 ^ 1'b0 ;
  assign n3713 = n510 | n3712 ;
  assign n3714 = n3194 ^ n2340 ^ 1'b0 ;
  assign n3715 = n1378 ^ n540 ^ 1'b0 ;
  assign n3716 = ~n1176 & n3715 ;
  assign n3717 = n3716 ^ n1460 ^ x36 ;
  assign n3718 = n2788 & ~n3717 ;
  assign n3719 = ~n1427 & n3718 ;
  assign n3720 = n3719 ^ x42 ^ 1'b0 ;
  assign n3722 = n2540 ^ n1087 ^ 1'b0 ;
  assign n3721 = x63 | n1591 ;
  assign n3723 = n3722 ^ n3721 ^ 1'b0 ;
  assign n3724 = n992 & n2930 ;
  assign n3725 = n3724 ^ n303 ^ 1'b0 ;
  assign n3726 = ~n3332 & n3725 ;
  assign n3729 = n2312 ^ n1719 ^ n618 ;
  assign n3727 = n1640 | n2042 ;
  assign n3728 = n3169 & ~n3727 ;
  assign n3730 = n3729 ^ n3728 ^ 1'b0 ;
  assign n3731 = n3676 ^ n3545 ^ 1'b0 ;
  assign n3732 = n2555 ^ n284 ^ 1'b0 ;
  assign n3733 = ~n1080 & n1272 ;
  assign n3734 = n3556 & n3733 ;
  assign n3735 = n3734 ^ n2666 ^ n1017 ;
  assign n3736 = n1420 & n3735 ;
  assign n3737 = ~n3254 & n3736 ;
  assign n3738 = n585 & ~n2293 ;
  assign n3739 = n3738 ^ n1455 ^ 1'b0 ;
  assign n3740 = n1958 ^ n882 ^ 1'b0 ;
  assign n3741 = n1658 | n3740 ;
  assign n3742 = n2320 & ~n3741 ;
  assign n3743 = ~n3739 & n3742 ;
  assign n3744 = n2698 ^ n2143 ^ n256 ;
  assign n3745 = ~n1341 & n3744 ;
  assign n3746 = n3745 ^ n1433 ^ 1'b0 ;
  assign n3747 = n1647 & ~n3746 ;
  assign n3748 = n2034 & ~n3747 ;
  assign n3749 = ( n470 & ~n923 ) | ( n470 & n2976 ) | ( ~n923 & n2976 ) ;
  assign n3751 = n2772 ^ n2614 ^ 1'b0 ;
  assign n3752 = n2355 | n3751 ;
  assign n3750 = n1544 & ~n3129 ;
  assign n3753 = n3752 ^ n3750 ^ 1'b0 ;
  assign n3754 = ~n3749 & n3753 ;
  assign n3755 = ~x69 & n3754 ;
  assign n3756 = ~n387 & n881 ;
  assign n3757 = n3756 ^ n922 ^ n337 ;
  assign n3758 = ( x30 & ~n318 ) | ( x30 & n3757 ) | ( ~n318 & n3757 ) ;
  assign n3759 = ~n2860 & n3758 ;
  assign n3760 = n1832 & n3759 ;
  assign n3761 = ~n3613 & n3693 ;
  assign n3762 = n3761 ^ n3643 ^ 1'b0 ;
  assign n3765 = n320 | n1210 ;
  assign n3763 = n1595 ^ x0 ^ 1'b0 ;
  assign n3764 = n386 | n3763 ;
  assign n3766 = n3765 ^ n3764 ^ 1'b0 ;
  assign n3767 = ( n221 & ~n2039 ) | ( n221 & n2371 ) | ( ~n2039 & n2371 ) ;
  assign n3768 = n2322 & n3767 ;
  assign n3769 = n350 & n3768 ;
  assign n3770 = n987 & n1869 ;
  assign n3771 = n2028 ^ n145 ^ 1'b0 ;
  assign n3772 = n2039 & n2297 ;
  assign n3773 = ( n1417 & ~n1438 ) | ( n1417 & n1631 ) | ( ~n1438 & n1631 ) ;
  assign n3774 = ~n474 & n3773 ;
  assign n3775 = n3774 ^ n3116 ^ 1'b0 ;
  assign n3776 = n3775 ^ n2919 ^ n238 ;
  assign n3777 = n3776 ^ n2645 ^ 1'b0 ;
  assign n3778 = n1710 | n3777 ;
  assign n3779 = n1656 ^ n1575 ^ n1014 ;
  assign n3780 = n697 & n2877 ;
  assign n3781 = n1625 ^ n279 ^ 1'b0 ;
  assign n3782 = n1101 ^ n843 ^ 1'b0 ;
  assign n3783 = ~n3114 & n3782 ;
  assign n3784 = n909 ^ n327 ^ 1'b0 ;
  assign n3785 = ( n1147 & ~n1623 ) | ( n1147 & n3572 ) | ( ~n1623 & n3572 ) ;
  assign n3788 = n2106 ^ n1864 ^ 1'b0 ;
  assign n3786 = n367 & ~n2285 ;
  assign n3787 = n3786 ^ n1175 ^ 1'b0 ;
  assign n3789 = n3788 ^ n3787 ^ 1'b0 ;
  assign n3790 = n511 & ~n3789 ;
  assign n3791 = n931 & n1418 ;
  assign n3793 = n1100 ^ n402 ^ 1'b0 ;
  assign n3794 = n511 & n3793 ;
  assign n3792 = ~x62 & n453 ;
  assign n3795 = n3794 ^ n3792 ^ 1'b0 ;
  assign n3796 = ( n256 & ~n3791 ) | ( n256 & n3795 ) | ( ~n3791 & n3795 ) ;
  assign n3797 = ~n2039 & n3796 ;
  assign n3798 = n831 & n3797 ;
  assign n3803 = n2496 ^ n1438 ^ x107 ;
  assign n3801 = n1985 ^ n322 ^ 1'b0 ;
  assign n3802 = ~n340 & n3801 ;
  assign n3804 = n3803 ^ n3802 ^ 1'b0 ;
  assign n3805 = n493 & ~n3804 ;
  assign n3799 = ~n2062 & n2930 ;
  assign n3800 = n3799 ^ n438 ^ 1'b0 ;
  assign n3806 = n3805 ^ n3800 ^ n2359 ;
  assign n3807 = ( ~n3790 & n3798 ) | ( ~n3790 & n3806 ) | ( n3798 & n3806 ) ;
  assign n3808 = n2930 ^ n2804 ^ 1'b0 ;
  assign n3809 = n3807 & ~n3808 ;
  assign n3810 = ~n3785 & n3809 ;
  assign n3811 = ~n332 & n3810 ;
  assign n3812 = n1084 & ~n2290 ;
  assign n3813 = n3812 ^ n153 ^ 1'b0 ;
  assign n3814 = ( n3096 & n3258 ) | ( n3096 & n3813 ) | ( n3258 & n3813 ) ;
  assign n3815 = n2584 ^ n2449 ^ n1837 ;
  assign n3816 = n1215 ^ n793 ^ 1'b0 ;
  assign n3817 = n3816 ^ n2645 ^ n2113 ;
  assign n3818 = n3817 ^ n3122 ^ 1'b0 ;
  assign n3819 = n832 | n3818 ;
  assign n3820 = n3819 ^ n2264 ^ 1'b0 ;
  assign n3821 = n2372 & ~n2800 ;
  assign n3822 = n2144 ^ n1198 ^ 1'b0 ;
  assign n3823 = n3821 & ~n3822 ;
  assign n3824 = n504 ^ n266 ^ 1'b0 ;
  assign n3825 = ~n886 & n1626 ;
  assign n3826 = ~n1869 & n3825 ;
  assign n3827 = n3785 ^ n2850 ^ n2267 ;
  assign n3828 = ( n2965 & ~n3549 ) | ( n2965 & n3827 ) | ( ~n3549 & n3827 ) ;
  assign n3829 = n3379 ^ n2338 ^ 1'b0 ;
  assign n3830 = n883 & ~n2905 ;
  assign n3831 = ( ~n2055 & n3383 ) | ( ~n2055 & n3830 ) | ( n3383 & n3830 ) ;
  assign n3832 = n3831 ^ n1511 ^ 1'b0 ;
  assign n3833 = n1045 ^ n944 ^ 1'b0 ;
  assign n3834 = n3832 & ~n3833 ;
  assign n3835 = n3829 & n3834 ;
  assign n3836 = ~n236 & n3835 ;
  assign n3837 = n914 & ~n1276 ;
  assign n3838 = n3837 ^ n322 ^ 1'b0 ;
  assign n3839 = n2515 ^ n1715 ^ n1546 ;
  assign n3840 = ( n2371 & n2855 ) | ( n2371 & ~n3839 ) | ( n2855 & ~n3839 ) ;
  assign n3841 = n2843 ^ n2297 ^ 1'b0 ;
  assign n3842 = ~n2788 & n3841 ;
  assign n3843 = ~n231 & n2258 ;
  assign n3844 = n3843 ^ n305 ^ 1'b0 ;
  assign n3845 = ( n1679 & n1862 ) | ( n1679 & ~n3050 ) | ( n1862 & ~n3050 ) ;
  assign n3846 = n568 | n3845 ;
  assign n3847 = n3844 | n3846 ;
  assign n3848 = n971 & ~n1881 ;
  assign n3849 = ~n992 & n1725 ;
  assign n3850 = n3849 ^ n232 ^ 1'b0 ;
  assign n3851 = n3850 ^ n3701 ^ n963 ;
  assign n3852 = ~n993 & n1491 ;
  assign n3853 = ( ~n395 & n1170 ) | ( ~n395 & n3852 ) | ( n1170 & n3852 ) ;
  assign n3854 = n1320 & n2221 ;
  assign n3855 = ~n1682 & n3854 ;
  assign n3856 = n248 & n1350 ;
  assign n3857 = n760 & ~n3086 ;
  assign n3858 = ~n3856 & n3857 ;
  assign n3859 = n3858 ^ n1329 ^ x48 ;
  assign n3860 = n3859 ^ x126 ^ 1'b0 ;
  assign n3861 = ~n1199 & n3860 ;
  assign n3862 = n3861 ^ n2896 ^ 1'b0 ;
  assign n3863 = ( n679 & ~n1537 ) | ( n679 & n3862 ) | ( ~n1537 & n3862 ) ;
  assign n3872 = n2038 ^ n165 ^ 1'b0 ;
  assign n3873 = n1743 | n3872 ;
  assign n3864 = n3660 ^ n1655 ^ n1160 ;
  assign n3865 = n887 ^ n693 ^ n493 ;
  assign n3866 = ( n290 & n646 ) | ( n290 & n2246 ) | ( n646 & n2246 ) ;
  assign n3867 = n3866 ^ n1743 ^ 1'b0 ;
  assign n3868 = n3865 & n3867 ;
  assign n3869 = n3868 ^ n2868 ^ 1'b0 ;
  assign n3870 = n261 & ~n3869 ;
  assign n3871 = n3864 & n3870 ;
  assign n3874 = n3873 ^ n3871 ^ 1'b0 ;
  assign n3875 = ~n2224 & n3874 ;
  assign n3876 = n1814 & n3875 ;
  assign n3877 = ( n629 & ~n775 ) | ( n629 & n779 ) | ( ~n775 & n779 ) ;
  assign n3878 = ( n211 & ~n2077 ) | ( n211 & n3877 ) | ( ~n2077 & n3877 ) ;
  assign n3879 = ~n281 & n1768 ;
  assign n3880 = n1165 & n2528 ;
  assign n3881 = ~n1511 & n3880 ;
  assign n3882 = ~n3879 & n3881 ;
  assign n3883 = n3878 & n3882 ;
  assign n3884 = ( n1177 & n1260 ) | ( n1177 & ~n1584 ) | ( n1260 & ~n1584 ) ;
  assign n3885 = ~n3467 & n3659 ;
  assign n3886 = ~n3884 & n3885 ;
  assign n3887 = n2219 ^ n2100 ^ n246 ;
  assign n3888 = n406 & ~n3887 ;
  assign n3889 = n652 | n2268 ;
  assign n3890 = n1603 & ~n3889 ;
  assign n3891 = n3752 | n3890 ;
  assign n3892 = n3891 ^ n3011 ^ 1'b0 ;
  assign n3893 = n2614 & ~n3719 ;
  assign n3894 = n3893 ^ n2837 ^ 1'b0 ;
  assign n3895 = n3045 ^ n829 ^ 1'b0 ;
  assign n3896 = n1165 & n3895 ;
  assign n3897 = n739 & ~n3682 ;
  assign n3898 = n929 & n3897 ;
  assign n3899 = ~n339 & n2118 ;
  assign n3900 = ~x31 & n3899 ;
  assign n3901 = n3900 ^ n2382 ^ 1'b0 ;
  assign n3902 = ~n3898 & n3901 ;
  assign n3903 = n3190 ^ n2435 ^ n1708 ;
  assign n3904 = n3903 ^ n3051 ^ 1'b0 ;
  assign n3905 = x92 & ~n3904 ;
  assign n3906 = n1442 ^ x66 ^ 1'b0 ;
  assign n3907 = n1894 & n3906 ;
  assign n3908 = n3907 ^ n3713 ^ 1'b0 ;
  assign n3909 = n1770 ^ n1365 ^ 1'b0 ;
  assign n3910 = x112 & n3909 ;
  assign n3911 = n3910 ^ n1107 ^ 1'b0 ;
  assign n3912 = n3911 ^ n3681 ^ n833 ;
  assign n3913 = ~n900 & n2258 ;
  assign n3914 = n3913 ^ n1281 ^ 1'b0 ;
  assign n3915 = n3914 ^ n3739 ^ 1'b0 ;
  assign n3916 = n3915 ^ n1185 ^ 1'b0 ;
  assign n3917 = n1958 ^ n1818 ^ 1'b0 ;
  assign n3918 = n3917 ^ n1082 ^ 1'b0 ;
  assign n3919 = n2278 & n3918 ;
  assign n3920 = n721 & ~n2986 ;
  assign n3921 = n2236 ^ n818 ^ 1'b0 ;
  assign n3922 = x40 ^ x19 ^ 1'b0 ;
  assign n3923 = ~n3921 & n3922 ;
  assign n3925 = n2251 & ~n2688 ;
  assign n3924 = n1809 | n3090 ;
  assign n3926 = n3925 ^ n3924 ^ 1'b0 ;
  assign n3927 = ~n1587 & n2657 ;
  assign n3928 = n3926 & n3927 ;
  assign n3929 = n3928 ^ n2835 ^ 1'b0 ;
  assign n3930 = n3016 & n3929 ;
  assign n3931 = ( ~n1556 & n3923 ) | ( ~n1556 & n3930 ) | ( n3923 & n3930 ) ;
  assign n3932 = ( n502 & n548 ) | ( n502 & ~n890 ) | ( n548 & ~n890 ) ;
  assign n3933 = ( n1022 & ~n2524 ) | ( n1022 & n3932 ) | ( ~n2524 & n3932 ) ;
  assign n3934 = n3933 ^ n3191 ^ 1'b0 ;
  assign n3935 = n2326 & n3563 ;
  assign n3936 = n1101 ^ n363 ^ 1'b0 ;
  assign n3937 = x46 & ~n3936 ;
  assign n3939 = x59 & n827 ;
  assign n3938 = n377 & ~n2047 ;
  assign n3940 = n3939 ^ n3938 ^ 1'b0 ;
  assign n3941 = n3937 & ~n3940 ;
  assign n3942 = n3920 ^ n2889 ^ n2535 ;
  assign n3943 = ( ~n963 & n1087 ) | ( ~n963 & n3552 ) | ( n1087 & n3552 ) ;
  assign n3944 = n3245 ^ n408 ^ 1'b0 ;
  assign n3945 = n3693 & ~n3944 ;
  assign n3946 = n3945 ^ n1923 ^ 1'b0 ;
  assign n3947 = n436 & ~n1435 ;
  assign n3951 = x43 & ~n3212 ;
  assign n3952 = n1853 & n2368 ;
  assign n3953 = ( x76 & n3951 ) | ( x76 & ~n3952 ) | ( n3951 & ~n3952 ) ;
  assign n3948 = n923 ^ n827 ^ 1'b0 ;
  assign n3949 = n3948 ^ n2056 ^ n424 ;
  assign n3950 = n3949 ^ n1682 ^ n349 ;
  assign n3954 = n3953 ^ n3950 ^ 1'b0 ;
  assign n3955 = n3954 ^ n3716 ^ n3242 ;
  assign n3956 = n443 ^ n258 ^ 1'b0 ;
  assign n3957 = n1699 | n3956 ;
  assign n3958 = n664 | n2397 ;
  assign n3959 = n1925 | n3958 ;
  assign n3960 = n3957 & ~n3959 ;
  assign n3961 = n512 ^ n288 ^ x86 ;
  assign n3962 = n1447 & n3961 ;
  assign n3967 = ~n194 & n3739 ;
  assign n3968 = n2831 ^ n2530 ^ 1'b0 ;
  assign n3969 = x103 | n434 ;
  assign n3970 = n3968 & n3969 ;
  assign n3971 = ~n3676 & n3970 ;
  assign n3972 = n3967 | n3971 ;
  assign n3963 = n1611 | n2165 ;
  assign n3964 = n3963 ^ n2049 ^ 1'b0 ;
  assign n3965 = n3964 ^ n708 ^ 1'b0 ;
  assign n3966 = n788 & ~n3965 ;
  assign n3973 = n3972 ^ n3966 ^ 1'b0 ;
  assign n3984 = n2337 ^ n2036 ^ 1'b0 ;
  assign n3985 = ~n412 & n1162 ;
  assign n3986 = ~n3984 & n3985 ;
  assign n3974 = ( n322 & n356 ) | ( n322 & n977 ) | ( n356 & n977 ) ;
  assign n3977 = n233 & ~n2117 ;
  assign n3978 = ~n193 & n3977 ;
  assign n3979 = n1841 ^ n1153 ^ 1'b0 ;
  assign n3980 = ~n3978 & n3979 ;
  assign n3975 = n1648 ^ n1183 ^ n761 ;
  assign n3976 = n3975 ^ n2452 ^ n1978 ;
  assign n3981 = n3980 ^ n3976 ^ 1'b0 ;
  assign n3982 = n3974 & n3981 ;
  assign n3983 = n3982 ^ n1163 ^ 1'b0 ;
  assign n3987 = n3986 ^ n3983 ^ n2138 ;
  assign n3988 = n2815 ^ n313 ^ 1'b0 ;
  assign n3989 = n3914 ^ n1818 ^ 1'b0 ;
  assign n3990 = n983 & n3976 ;
  assign n3991 = ~n512 & n3990 ;
  assign n3992 = n3884 ^ n1936 ^ 1'b0 ;
  assign n3993 = n3991 | n3992 ;
  assign n3994 = n1475 ^ n824 ^ n790 ;
  assign n3995 = n2984 ^ n152 ^ 1'b0 ;
  assign n3996 = ~n2173 & n3651 ;
  assign n3997 = ~n2416 & n3996 ;
  assign n3998 = n1386 ^ n621 ^ 1'b0 ;
  assign n3999 = n2535 & n3998 ;
  assign n4000 = n1761 & n3999 ;
  assign n4001 = ~n2555 & n4000 ;
  assign n4002 = n1066 & ~n3616 ;
  assign n4003 = ~x68 & n4002 ;
  assign n4004 = n4003 ^ n1529 ^ 1'b0 ;
  assign n4005 = ~n4001 & n4004 ;
  assign n4006 = ( n977 & ~n3962 ) | ( n977 & n4005 ) | ( ~n3962 & n4005 ) ;
  assign n4007 = ~n554 & n805 ;
  assign n4008 = ~n3250 & n4007 ;
  assign n4009 = n4008 ^ n995 ^ 1'b0 ;
  assign n4010 = n3046 ^ n1839 ^ 1'b0 ;
  assign n4011 = n234 & n2059 ;
  assign n4012 = n2712 ^ n1626 ^ n657 ;
  assign n4013 = x100 | n1512 ;
  assign n4014 = n4013 ^ n2538 ^ 1'b0 ;
  assign n4015 = ( ~n4011 & n4012 ) | ( ~n4011 & n4014 ) | ( n4012 & n4014 ) ;
  assign n4018 = ( n209 & n1690 ) | ( n209 & n3428 ) | ( n1690 & n3428 ) ;
  assign n4019 = n4018 ^ x1 ^ 1'b0 ;
  assign n4020 = ~n1651 & n4019 ;
  assign n4016 = n988 & ~n3978 ;
  assign n4017 = ~n2596 & n4016 ;
  assign n4021 = n4020 ^ n4017 ^ 1'b0 ;
  assign n4022 = n3636 ^ n304 ^ 1'b0 ;
  assign n4023 = n278 & n1655 ;
  assign n4024 = ~n2705 & n4023 ;
  assign n4025 = n4024 ^ n290 ^ 1'b0 ;
  assign n4026 = n227 | n4025 ;
  assign n4027 = ( n148 & n222 ) | ( n148 & ~n1764 ) | ( n222 & ~n1764 ) ;
  assign n4028 = n1302 & ~n3003 ;
  assign n4029 = n4027 & n4028 ;
  assign n4030 = ~n4026 & n4029 ;
  assign n4031 = ~n4022 & n4030 ;
  assign n4037 = x8 & x116 ;
  assign n4038 = n1843 ^ n1415 ^ 1'b0 ;
  assign n4039 = ~n4037 & n4038 ;
  assign n4040 = n1388 ^ n688 ^ 1'b0 ;
  assign n4041 = n4039 | n4040 ;
  assign n4032 = n1212 ^ n247 ^ x89 ;
  assign n4033 = ( n1841 & ~n2109 ) | ( n1841 & n3261 ) | ( ~n2109 & n3261 ) ;
  assign n4034 = n1249 | n4033 ;
  assign n4035 = n4032 | n4034 ;
  assign n4036 = ~n2976 & n4035 ;
  assign n4042 = n4041 ^ n4036 ^ 1'b0 ;
  assign n4043 = n1858 ^ n1727 ^ n1320 ;
  assign n4044 = n4043 ^ n1714 ^ 1'b0 ;
  assign n4045 = n2102 & ~n4044 ;
  assign n4046 = ( ~n1326 & n2218 ) | ( ~n1326 & n4045 ) | ( n2218 & n4045 ) ;
  assign n4047 = ~n841 & n2153 ;
  assign n4048 = ~n701 & n4047 ;
  assign n4049 = n668 & ~n4048 ;
  assign n4050 = n4049 ^ n3395 ^ x31 ;
  assign n4051 = ~n387 & n586 ;
  assign n4052 = n4051 ^ n1977 ^ 1'b0 ;
  assign n4053 = n2251 ^ n1025 ^ 1'b0 ;
  assign n4054 = n627 & ~n4053 ;
  assign n4055 = n4054 ^ n941 ^ x21 ;
  assign n4061 = n2245 ^ n300 ^ x19 ;
  assign n4058 = x44 & n1491 ;
  assign n4059 = n4058 ^ n3218 ^ 1'b0 ;
  assign n4060 = n1425 & n4059 ;
  assign n4062 = n4061 ^ n4060 ^ 1'b0 ;
  assign n4063 = n4062 ^ n2081 ^ n165 ;
  assign n4056 = ~n595 & n775 ;
  assign n4057 = n2425 & n4056 ;
  assign n4064 = n4063 ^ n4057 ^ 1'b0 ;
  assign n4065 = n4055 & n4064 ;
  assign n4066 = n2557 ^ n1476 ^ 1'b0 ;
  assign n4067 = n2357 ^ x107 ^ 1'b0 ;
  assign n4068 = n828 ^ n606 ^ 1'b0 ;
  assign n4069 = ( n948 & ~n1256 ) | ( n948 & n4068 ) | ( ~n1256 & n4068 ) ;
  assign n4070 = n4069 ^ n1163 ^ 1'b0 ;
  assign n4071 = n4070 ^ n2335 ^ 1'b0 ;
  assign n4072 = ( n490 & ~n942 ) | ( n490 & n1065 ) | ( ~n942 & n1065 ) ;
  assign n4073 = n4072 ^ n881 ^ 1'b0 ;
  assign n4074 = ~n4071 & n4073 ;
  assign n4078 = n3556 ^ n3033 ^ x37 ;
  assign n4075 = n3739 ^ n1741 ^ n533 ;
  assign n4076 = n2526 ^ n620 ^ 1'b0 ;
  assign n4077 = n4075 | n4076 ;
  assign n4079 = n4078 ^ n4077 ^ 1'b0 ;
  assign n4080 = n775 & ~n2310 ;
  assign n4081 = n153 & n4080 ;
  assign n4082 = n1524 | n4081 ;
  assign n4083 = n4082 ^ n1936 ^ 1'b0 ;
  assign n4084 = ( ~x30 & x37 ) | ( ~x30 & n4083 ) | ( x37 & n4083 ) ;
  assign n4085 = n1937 ^ n1802 ^ n153 ;
  assign n4086 = ~n236 & n4085 ;
  assign n4087 = n2647 ^ n2584 ^ x72 ;
  assign n4088 = ~n1195 & n2535 ;
  assign n4089 = n4038 ^ n2379 ^ 1'b0 ;
  assign n4090 = ~n2079 & n4089 ;
  assign n4091 = n1035 & n1998 ;
  assign n4092 = ~x37 & n4091 ;
  assign n4093 = n3341 & ~n3429 ;
  assign n4094 = ~n1425 & n4093 ;
  assign n4095 = ~n1445 & n4094 ;
  assign n4096 = ( x83 & n4092 ) | ( x83 & ~n4095 ) | ( n4092 & ~n4095 ) ;
  assign n4097 = n4096 ^ n3416 ^ 1'b0 ;
  assign n4102 = n1738 & n2083 ;
  assign n4099 = n1008 & ~n3864 ;
  assign n4098 = n175 & ~n950 ;
  assign n4100 = n4099 ^ n4098 ^ 1'b0 ;
  assign n4101 = n4100 ^ n2213 ^ 1'b0 ;
  assign n4103 = n4102 ^ n4101 ^ n2619 ;
  assign n4104 = n4103 ^ n3486 ^ n2221 ;
  assign n4105 = n520 & ~n1455 ;
  assign n4106 = n700 & n4105 ;
  assign n4107 = ( n1020 & n1459 ) | ( n1020 & ~n4106 ) | ( n1459 & ~n4106 ) ;
  assign n4108 = n4107 ^ n2165 ^ 1'b0 ;
  assign n4109 = n4104 & ~n4108 ;
  assign n4110 = n4109 ^ n3509 ^ 1'b0 ;
  assign n4111 = n2767 ^ n2549 ^ 1'b0 ;
  assign n4112 = ( n1639 & n3831 ) | ( n1639 & ~n4077 ) | ( n3831 & ~n4077 ) ;
  assign n4113 = ~n755 & n796 ;
  assign n4114 = n4113 ^ n1485 ^ 1'b0 ;
  assign n4115 = n4114 ^ n1335 ^ 1'b0 ;
  assign n4116 = ( n276 & n664 ) | ( n276 & ~n800 ) | ( n664 & ~n800 ) ;
  assign n4117 = n266 & ~n4116 ;
  assign n4118 = n4117 ^ n756 ^ 1'b0 ;
  assign n4119 = n4115 & ~n4118 ;
  assign n4120 = ( ~n193 & n815 ) | ( ~n193 & n890 ) | ( n815 & n890 ) ;
  assign n4121 = n4120 ^ n3565 ^ 1'b0 ;
  assign n4122 = ~n482 & n1147 ;
  assign n4123 = n313 | n1260 ;
  assign n4124 = n1930 & ~n3195 ;
  assign n4125 = ( n211 & ~n3389 ) | ( n211 & n4124 ) | ( ~n3389 & n4124 ) ;
  assign n4126 = n3607 ^ n1744 ^ 1'b0 ;
  assign n4127 = n3777 & ~n4126 ;
  assign n4128 = n4127 ^ n334 ^ 1'b0 ;
  assign n4129 = n1249 | n2104 ;
  assign n4130 = n2352 & ~n4129 ;
  assign n4131 = n2053 ^ n629 ^ n493 ;
  assign n4132 = n3117 ^ n1831 ^ 1'b0 ;
  assign n4133 = n3508 | n4132 ;
  assign n4134 = ~n860 & n925 ;
  assign n4135 = n1893 ^ n1436 ^ 1'b0 ;
  assign n4136 = n1074 | n4135 ;
  assign n4137 = n3659 | n4136 ;
  assign n4140 = n1066 & ~n1249 ;
  assign n4141 = n4140 ^ n781 ^ 1'b0 ;
  assign n4142 = n927 ^ n211 ^ 1'b0 ;
  assign n4143 = n4142 ^ n2368 ^ 1'b0 ;
  assign n4144 = n1764 ^ n433 ^ 1'b0 ;
  assign n4145 = x121 & n4144 ;
  assign n4146 = ~n4143 & n4145 ;
  assign n4147 = n4141 & ~n4146 ;
  assign n4148 = n4147 ^ n1812 ^ n867 ;
  assign n4138 = ~n1299 & n3466 ;
  assign n4139 = n4138 ^ n2706 ^ 1'b0 ;
  assign n4149 = n4148 ^ n4139 ^ 1'b0 ;
  assign n4155 = n3244 ^ n2047 ^ 1'b0 ;
  assign n4150 = ( x13 & ~x85 ) | ( x13 & n3172 ) | ( ~x85 & n3172 ) ;
  assign n4151 = n4150 ^ n229 ^ 1'b0 ;
  assign n4152 = n1335 | n4151 ;
  assign n4153 = n1893 | n4152 ;
  assign n4154 = n4153 ^ n4062 ^ 1'b0 ;
  assign n4156 = n4155 ^ n4154 ^ n2705 ;
  assign n4157 = n1971 ^ n1964 ^ 1'b0 ;
  assign n4158 = n1719 & n4157 ;
  assign n4159 = n360 ^ n201 ^ 1'b0 ;
  assign n4160 = n2544 ^ n958 ^ n300 ;
  assign n4161 = n4160 ^ n3593 ^ n1536 ;
  assign n4162 = n4159 & ~n4161 ;
  assign n4163 = ~n4158 & n4162 ;
  assign n4164 = ( ~n1184 & n1218 ) | ( ~n1184 & n1543 ) | ( n1218 & n1543 ) ;
  assign n4165 = n1490 & n4164 ;
  assign n4166 = ~n4143 & n4165 ;
  assign n4167 = n4166 ^ n1475 ^ x57 ;
  assign n4168 = n1190 ^ n756 ^ 1'b0 ;
  assign n4169 = ~n2617 & n4168 ;
  assign n4170 = n4169 ^ n1797 ^ n846 ;
  assign n4171 = n4170 ^ n2846 ^ 1'b0 ;
  assign n4172 = n2726 & n4171 ;
  assign n4173 = n979 ^ n713 ^ 1'b0 ;
  assign n4174 = n4173 ^ n2889 ^ 1'b0 ;
  assign n4175 = n4014 ^ n2070 ^ 1'b0 ;
  assign n4176 = n2012 ^ n1334 ^ 1'b0 ;
  assign n4177 = n1515 & n4176 ;
  assign n4178 = ~n403 & n4177 ;
  assign n4179 = ( ~n963 & n1605 ) | ( ~n963 & n4178 ) | ( n1605 & n4178 ) ;
  assign n4180 = ~n1382 & n1619 ;
  assign n4181 = n4180 ^ n2880 ^ 1'b0 ;
  assign n4184 = n1398 ^ n1350 ^ 1'b0 ;
  assign n4183 = n1422 ^ x52 ^ 1'b0 ;
  assign n4182 = n813 ^ n485 ^ 1'b0 ;
  assign n4185 = n4184 ^ n4183 ^ n4182 ;
  assign n4186 = ( n2231 & n2726 ) | ( n2231 & ~n3507 ) | ( n2726 & ~n3507 ) ;
  assign n4187 = n1587 | n4186 ;
  assign n4188 = n4187 ^ n1865 ^ n1126 ;
  assign n4189 = ~n2340 & n3513 ;
  assign n4190 = ~n2201 & n4189 ;
  assign n4191 = ( n285 & n411 ) | ( n285 & ~n4190 ) | ( n411 & ~n4190 ) ;
  assign n4192 = n1318 & ~n1445 ;
  assign n4193 = n4191 & n4192 ;
  assign n4194 = ~n911 & n4059 ;
  assign n4195 = n4194 ^ n595 ^ 1'b0 ;
  assign n4196 = n2391 ^ n613 ^ 1'b0 ;
  assign n4197 = x29 & n4196 ;
  assign n4198 = n4197 ^ n956 ^ 1'b0 ;
  assign n4199 = n4092 | n4198 ;
  assign n4200 = n3317 | n4199 ;
  assign n4201 = n2971 & n4200 ;
  assign n4203 = n2155 ^ n1175 ^ 1'b0 ;
  assign n4202 = n1947 ^ n882 ^ 1'b0 ;
  assign n4204 = n4203 ^ n4202 ^ n2018 ;
  assign n4205 = n916 | n1146 ;
  assign n4206 = n349 | n4205 ;
  assign n4207 = n4206 ^ n874 ^ 1'b0 ;
  assign n4208 = ( ~x7 & n3293 ) | ( ~x7 & n4207 ) | ( n3293 & n4207 ) ;
  assign n4214 = n2008 ^ x96 ^ 1'b0 ;
  assign n4209 = n2617 ^ n1537 ^ 1'b0 ;
  assign n4210 = ( ~x57 & n1854 ) | ( ~x57 & n4209 ) | ( n1854 & n4209 ) ;
  assign n4211 = n362 & n4210 ;
  assign n4212 = n1608 & ~n4211 ;
  assign n4213 = n953 & n4212 ;
  assign n4215 = n4214 ^ n4213 ^ 1'b0 ;
  assign n4216 = n2951 & ~n4215 ;
  assign n4217 = ( n1548 & n1860 ) | ( n1548 & n2430 ) | ( n1860 & n2430 ) ;
  assign n4218 = n2332 ^ n247 ^ 1'b0 ;
  assign n4219 = n4218 ^ n2929 ^ 1'b0 ;
  assign n4220 = n477 & n4219 ;
  assign n4221 = n4220 ^ n3672 ^ n1025 ;
  assign n4222 = ~n134 & n1071 ;
  assign n4223 = ~n1261 & n4222 ;
  assign n4224 = n4223 ^ n3878 ^ 1'b0 ;
  assign n4225 = n4224 ^ x74 ^ 1'b0 ;
  assign n4226 = n575 | n4225 ;
  assign n4227 = ( ~n289 & n408 ) | ( ~n289 & n667 ) | ( n408 & n667 ) ;
  assign n4228 = n796 & ~n2349 ;
  assign n4229 = n4227 & n4228 ;
  assign n4230 = ( n1555 & n3326 ) | ( n1555 & n4229 ) | ( n3326 & n4229 ) ;
  assign n4231 = ~n2235 & n4230 ;
  assign n4232 = x104 & n1907 ;
  assign n4233 = n900 & n4232 ;
  assign n4234 = n4233 ^ n4211 ^ 1'b0 ;
  assign n4235 = n3890 | n4234 ;
  assign n4236 = n940 & ~n4235 ;
  assign n4237 = ~n979 & n4236 ;
  assign n4238 = ~n3604 & n4237 ;
  assign n4239 = n191 & n2231 ;
  assign n4240 = n3108 ^ n747 ^ n660 ;
  assign n4241 = n4240 ^ n3272 ^ 1'b0 ;
  assign n4242 = ~n1881 & n4241 ;
  assign n4243 = n4242 ^ n2124 ^ n194 ;
  assign n4244 = n725 | n4243 ;
  assign n4245 = n4244 ^ n2357 ^ 1'b0 ;
  assign n4246 = n4245 ^ n2997 ^ 1'b0 ;
  assign n4247 = n4246 ^ n2290 ^ n1305 ;
  assign n4248 = n2038 ^ n1921 ^ n1314 ;
  assign n4249 = n3429 & n3693 ;
  assign n4250 = n225 | n391 ;
  assign n4251 = n4250 ^ n2207 ^ 1'b0 ;
  assign n4252 = n4249 | n4251 ;
  assign n4253 = n4248 & n4252 ;
  assign n4256 = n4048 ^ n2262 ^ 1'b0 ;
  assign n4254 = x5 & n3375 ;
  assign n4255 = n3643 & n4254 ;
  assign n4257 = n4256 ^ n4255 ^ n3705 ;
  assign n4258 = n1992 | n2076 ;
  assign n4259 = n384 & ~n4258 ;
  assign n4260 = n1931 ^ x73 ^ 1'b0 ;
  assign n4261 = ~n4259 & n4260 ;
  assign n4277 = ~x23 & n3272 ;
  assign n4278 = ~n1049 & n4277 ;
  assign n4279 = n4278 ^ x75 ^ 1'b0 ;
  assign n4280 = n1214 | n1686 ;
  assign n4281 = n613 & ~n4280 ;
  assign n4282 = n521 & ~n4281 ;
  assign n4283 = n4279 & n4282 ;
  assign n4262 = n2161 | n4233 ;
  assign n4263 = n4262 ^ n1379 ^ 1'b0 ;
  assign n4264 = n2905 | n4263 ;
  assign n4265 = n1665 & ~n4264 ;
  assign n4266 = x21 & x69 ;
  assign n4267 = n2157 & n4266 ;
  assign n4268 = n3341 ^ n1764 ^ 1'b0 ;
  assign n4269 = n611 | n4268 ;
  assign n4270 = n833 | n4269 ;
  assign n4271 = n4270 ^ n4016 ^ 1'b0 ;
  assign n4272 = ~n219 & n4271 ;
  assign n4273 = n4267 & n4272 ;
  assign n4274 = ( n3088 & n4265 ) | ( n3088 & ~n4273 ) | ( n4265 & ~n4273 ) ;
  assign n4275 = n1184 & ~n2500 ;
  assign n4276 = ~n4274 & n4275 ;
  assign n4284 = n4283 ^ n4276 ^ 1'b0 ;
  assign n4285 = x4 & n594 ;
  assign n4286 = n4285 ^ n2298 ^ 1'b0 ;
  assign n4287 = ( n1012 & n2640 ) | ( n1012 & ~n3839 ) | ( n2640 & ~n3839 ) ;
  assign n4288 = ( ~n3420 & n4286 ) | ( ~n3420 & n4287 ) | ( n4286 & n4287 ) ;
  assign n4289 = n3431 ^ n1958 ^ 1'b0 ;
  assign n4290 = n3697 ^ n2303 ^ 1'b0 ;
  assign n4291 = n4290 ^ n3950 ^ 1'b0 ;
  assign n4292 = ~n4289 & n4291 ;
  assign n4293 = n404 ^ x20 ^ 1'b0 ;
  assign n4294 = ~n2604 & n4293 ;
  assign n4295 = n4024 ^ n2546 ^ 1'b0 ;
  assign n4296 = n4294 & n4295 ;
  assign n4297 = n1615 ^ n212 ^ 1'b0 ;
  assign n4298 = n2534 & ~n4297 ;
  assign n4299 = ~n1055 & n2312 ;
  assign n4300 = ~n3255 & n4299 ;
  assign n4301 = n3270 & n4300 ;
  assign n4302 = n2031 ^ n1201 ^ 1'b0 ;
  assign n4303 = ( ~n927 & n4301 ) | ( ~n927 & n4302 ) | ( n4301 & n4302 ) ;
  assign n4304 = n1750 ^ n557 ^ 1'b0 ;
  assign n4305 = n1913 & ~n3704 ;
  assign n4306 = ~n4304 & n4305 ;
  assign n4307 = n954 & ~n2062 ;
  assign n4308 = ( n1098 & n1818 ) | ( n1098 & ~n4307 ) | ( n1818 & ~n4307 ) ;
  assign n4323 = ( n2174 & n2215 ) | ( n2174 & ~n3393 ) | ( n2215 & ~n3393 ) ;
  assign n4310 = n514 | n536 ;
  assign n4311 = x105 & n537 ;
  assign n4312 = n4310 & n4311 ;
  assign n4313 = n4312 ^ n980 ^ 1'b0 ;
  assign n4309 = ~n2285 & n3964 ;
  assign n4314 = n4313 ^ n4309 ^ 1'b0 ;
  assign n4315 = n4314 ^ n1336 ^ 1'b0 ;
  assign n4316 = n573 & ~n4315 ;
  assign n4317 = n2070 ^ n445 ^ 1'b0 ;
  assign n4318 = n2426 & n4317 ;
  assign n4319 = n2641 | n4318 ;
  assign n4320 = n1240 & ~n4319 ;
  assign n4321 = n4320 ^ n3515 ^ 1'b0 ;
  assign n4322 = n4316 & n4321 ;
  assign n4324 = n4323 ^ n4322 ^ 1'b0 ;
  assign n4325 = n1921 & ~n2145 ;
  assign n4326 = n4325 ^ n1970 ^ 1'b0 ;
  assign n4327 = n1697 ^ n1408 ^ 1'b0 ;
  assign n4328 = n4326 & n4327 ;
  assign n4329 = ( n1042 & n2430 ) | ( n1042 & n2699 ) | ( n2430 & n2699 ) ;
  assign n4330 = n2499 & n4329 ;
  assign n4331 = x117 & ~n1107 ;
  assign n4332 = ~n670 & n2008 ;
  assign n4333 = ( n1106 & n4028 ) | ( n1106 & n4332 ) | ( n4028 & n4332 ) ;
  assign n4334 = ( ~n1199 & n4331 ) | ( ~n1199 & n4333 ) | ( n4331 & n4333 ) ;
  assign n4335 = x126 & n3182 ;
  assign n4336 = n410 & n4335 ;
  assign n4337 = n4336 ^ n2337 ^ 1'b0 ;
  assign n4338 = ~n1240 & n3534 ;
  assign n4339 = n2124 | n3871 ;
  assign n4340 = n4339 ^ n2549 ^ 1'b0 ;
  assign n4341 = ~n2297 & n4248 ;
  assign n4342 = ( n663 & n4340 ) | ( n663 & n4341 ) | ( n4340 & n4341 ) ;
  assign n4343 = n4342 ^ n1649 ^ 1'b0 ;
  assign n4344 = n3227 ^ n1836 ^ 1'b0 ;
  assign n4345 = n3017 ^ n2990 ^ x37 ;
  assign n4346 = ( n2431 & ~n3117 ) | ( n2431 & n4345 ) | ( ~n3117 & n4345 ) ;
  assign n4347 = x32 & ~n1084 ;
  assign n4348 = n4346 | n4347 ;
  assign n4349 = n4344 | n4348 ;
  assign n4350 = ~x47 & n4349 ;
  assign n4351 = n3388 ^ n1689 ^ 1'b0 ;
  assign n4352 = n3914 | n4351 ;
  assign n4353 = n4352 ^ n4116 ^ 1'b0 ;
  assign n4354 = ~n535 & n4353 ;
  assign n4355 = n2514 ^ n922 ^ 1'b0 ;
  assign n4356 = ~n1996 & n3757 ;
  assign n4357 = n4356 ^ n1612 ^ n1042 ;
  assign n4358 = ( n1969 & n3718 ) | ( n1969 & n4357 ) | ( n3718 & n4357 ) ;
  assign n4359 = ~n299 & n2516 ;
  assign n4360 = n4359 ^ n3997 ^ 1'b0 ;
  assign n4361 = n4071 ^ n746 ^ 1'b0 ;
  assign n4368 = ~n1663 & n2070 ;
  assign n4369 = n4368 ^ n2758 ^ 1'b0 ;
  assign n4362 = n1475 ^ n1469 ^ n485 ;
  assign n4363 = n798 & ~n1878 ;
  assign n4364 = n4362 & n4363 ;
  assign n4365 = ( n195 & n1312 ) | ( n195 & n4364 ) | ( n1312 & n4364 ) ;
  assign n4366 = n2531 & ~n4365 ;
  assign n4367 = ~n3241 & n4366 ;
  assign n4370 = n4369 ^ n4367 ^ n3160 ;
  assign n4371 = n915 & ~n4175 ;
  assign n4372 = ~n3080 & n4371 ;
  assign n4373 = n3713 ^ n1699 ^ 1'b0 ;
  assign n4374 = ( ~n708 & n932 ) | ( ~n708 & n3873 ) | ( n932 & n3873 ) ;
  assign n4375 = n4374 ^ n2540 ^ n850 ;
  assign n4376 = n4375 ^ n1403 ^ 1'b0 ;
  assign n4377 = n4376 ^ n4086 ^ 1'b0 ;
  assign n4378 = x31 & ~n4377 ;
  assign n4379 = n2303 ^ n1211 ^ 1'b0 ;
  assign n4380 = n3227 & ~n4379 ;
  assign n4381 = n1995 ^ n510 ^ 1'b0 ;
  assign n4382 = n3476 & n4381 ;
  assign n4383 = n3364 ^ n1347 ^ 1'b0 ;
  assign n4384 = n3988 ^ n3686 ^ n1785 ;
  assign n4387 = ~n332 & n1972 ;
  assign n4385 = n1410 | n1660 ;
  assign n4386 = n372 | n4385 ;
  assign n4388 = n4387 ^ n4386 ^ 1'b0 ;
  assign n4389 = ( ~n561 & n2767 ) | ( ~n561 & n3707 ) | ( n2767 & n3707 ) ;
  assign n4402 = n3504 ^ n2475 ^ n927 ;
  assign n4399 = n673 & ~n1982 ;
  assign n4391 = n1784 & ~n4281 ;
  assign n4392 = ~n2102 & n4391 ;
  assign n4393 = ( ~n705 & n971 ) | ( ~n705 & n1430 ) | ( n971 & n1430 ) ;
  assign n4394 = ( ~n186 & n848 ) | ( ~n186 & n4393 ) | ( n848 & n4393 ) ;
  assign n4395 = n4394 ^ n2306 ^ 1'b0 ;
  assign n4396 = n4392 | n4395 ;
  assign n4390 = n951 & ~n1340 ;
  assign n4397 = n4396 ^ n4390 ^ 1'b0 ;
  assign n4398 = n4397 ^ n2012 ^ n947 ;
  assign n4400 = n4399 ^ n4398 ^ 1'b0 ;
  assign n4401 = x24 & ~n4400 ;
  assign n4403 = n4402 ^ n4401 ^ n761 ;
  assign n4404 = ( n1992 & n1995 ) | ( n1992 & n4403 ) | ( n1995 & n4403 ) ;
  assign n4405 = ~n517 & n2947 ;
  assign n4406 = n876 & n3503 ;
  assign n4407 = n1284 & n4406 ;
  assign n4408 = ( x106 & n1340 ) | ( x106 & ~n4407 ) | ( n1340 & ~n4407 ) ;
  assign n4409 = n4405 | n4408 ;
  assign n4410 = n3186 ^ n964 ^ 1'b0 ;
  assign n4411 = n4409 | n4410 ;
  assign n4412 = n1819 | n2236 ;
  assign n4413 = n1715 | n4412 ;
  assign n4414 = x27 & n3678 ;
  assign n4415 = n3178 ^ n2836 ^ 1'b0 ;
  assign n4416 = n4099 ^ n3964 ^ 1'b0 ;
  assign n4417 = n4416 ^ n4086 ^ 1'b0 ;
  assign n4420 = n3548 ^ n3001 ^ 1'b0 ;
  assign n4418 = n4132 ^ n3616 ^ 1'b0 ;
  assign n4419 = n4418 ^ n3340 ^ 1'b0 ;
  assign n4421 = n4420 ^ n4419 ^ 1'b0 ;
  assign n4422 = n1269 | n4421 ;
  assign n4425 = n2124 | n2264 ;
  assign n4423 = n1997 ^ n799 ^ 1'b0 ;
  assign n4424 = n599 & ~n4423 ;
  assign n4426 = n4425 ^ n4424 ^ 1'b0 ;
  assign n4427 = n3677 ^ n1116 ^ 1'b0 ;
  assign n4428 = ~n4250 & n4427 ;
  assign n4429 = n3261 ^ n1082 ^ 1'b0 ;
  assign n4430 = ( n1652 & n2030 ) | ( n1652 & ~n4429 ) | ( n2030 & ~n4429 ) ;
  assign n4433 = n3553 ^ n3016 ^ 1'b0 ;
  assign n4431 = ( n1460 & ~n2826 ) | ( n1460 & n3925 ) | ( ~n2826 & n3925 ) ;
  assign n4432 = n4431 ^ n3287 ^ 1'b0 ;
  assign n4434 = n4433 ^ n4432 ^ n299 ;
  assign n4439 = n467 & n2609 ;
  assign n4440 = n4439 ^ n1356 ^ 1'b0 ;
  assign n4435 = ~n1234 & n3001 ;
  assign n4436 = n4435 ^ n1012 ^ 1'b0 ;
  assign n4437 = ( x0 & n420 ) | ( x0 & n4436 ) | ( n420 & n4436 ) ;
  assign n4438 = ~n474 & n4437 ;
  assign n4441 = n4440 ^ n4438 ^ 1'b0 ;
  assign n4442 = n1738 ^ n1481 ^ n1306 ;
  assign n4443 = n4442 ^ n4085 ^ n1491 ;
  assign n4444 = n1506 ^ n866 ^ 1'b0 ;
  assign n4445 = ( x68 & n1330 ) | ( x68 & ~n4444 ) | ( n1330 & ~n4444 ) ;
  assign n4446 = n4445 ^ x54 ^ 1'b0 ;
  assign n4447 = n3181 ^ n1626 ^ 1'b0 ;
  assign n4448 = n2931 & n3999 ;
  assign n4449 = n2614 & n4448 ;
  assign n4450 = n4434 ^ n3735 ^ n825 ;
  assign n4451 = n211 & ~n4264 ;
  assign n4452 = n4451 ^ n1739 ^ x53 ;
  assign n4453 = n2196 & ~n4259 ;
  assign n4454 = n4453 ^ n1956 ^ 1'b0 ;
  assign n4455 = ( n998 & n1552 ) | ( n998 & n4454 ) | ( n1552 & n4454 ) ;
  assign n4456 = n608 ^ n607 ^ n378 ;
  assign n4457 = n2059 ^ n447 ^ 1'b0 ;
  assign n4458 = n1718 | n4457 ;
  assign n4459 = ( n313 & n4456 ) | ( n313 & ~n4458 ) | ( n4456 & ~n4458 ) ;
  assign n4460 = n4343 ^ n4334 ^ 1'b0 ;
  assign n4461 = n4459 & n4460 ;
  assign n4462 = ~n218 & n3999 ;
  assign n4463 = ~n1076 & n3356 ;
  assign n4464 = n4462 | n4463 ;
  assign n4465 = n2565 & ~n4464 ;
  assign n4466 = ~n578 & n2712 ;
  assign n4467 = n4466 ^ n1308 ^ 1'b0 ;
  assign n4468 = n4467 ^ n2440 ^ n2303 ;
  assign n4469 = ( x88 & ~n248 ) | ( x88 & n1138 ) | ( ~n248 & n1138 ) ;
  assign n4470 = ~n2791 & n4469 ;
  assign n4471 = ~n911 & n1311 ;
  assign n4472 = n4470 & n4471 ;
  assign n4473 = n307 & ~n4472 ;
  assign n4474 = ~n3560 & n4473 ;
  assign n4475 = n4474 ^ n3378 ^ 1'b0 ;
  assign n4476 = n4475 ^ n3485 ^ n3180 ;
  assign n4477 = n1430 | n4095 ;
  assign n4478 = n1083 | n4477 ;
  assign n4479 = n1233 ^ n711 ^ 1'b0 ;
  assign n4480 = n1154 & n4326 ;
  assign n4481 = n1525 & n1759 ;
  assign n4482 = n1379 & n4481 ;
  assign n4483 = n2349 | n4269 ;
  assign n4484 = n3710 ^ n2204 ^ n1622 ;
  assign n4485 = ( x52 & ~n1389 ) | ( x52 & n4062 ) | ( ~n1389 & n4062 ) ;
  assign n4486 = ( n540 & n1120 ) | ( n540 & n4485 ) | ( n1120 & n4485 ) ;
  assign n4487 = n4486 ^ n2695 ^ n1211 ;
  assign n4488 = n1939 ^ n1903 ^ 1'b0 ;
  assign n4489 = ( x92 & ~n337 ) | ( x92 & n1727 ) | ( ~n337 & n1727 ) ;
  assign n4490 = ( n860 & n4488 ) | ( n860 & n4489 ) | ( n4488 & n4489 ) ;
  assign n4492 = n2105 | n2893 ;
  assign n4491 = n429 & ~n3329 ;
  assign n4493 = n4492 ^ n4491 ^ 1'b0 ;
  assign n4494 = n1644 | n4493 ;
  assign n4495 = n2913 ^ n634 ^ 1'b0 ;
  assign n4496 = n3631 ^ n719 ^ 1'b0 ;
  assign n4497 = n4495 & n4496 ;
  assign n4498 = n4199 ^ n990 ^ 1'b0 ;
  assign n4499 = n3185 ^ n1674 ^ 1'b0 ;
  assign n4500 = n1745 ^ x37 ^ 1'b0 ;
  assign n4501 = ~n3572 & n4500 ;
  assign n4502 = n741 & n2772 ;
  assign n4503 = ~n1288 & n4502 ;
  assign n4504 = n4503 ^ n456 ^ x68 ;
  assign n4505 = n3212 ^ n557 ^ n181 ;
  assign n4506 = ~n4048 & n4505 ;
  assign n4507 = ~n206 & n4506 ;
  assign n4508 = ( n838 & ~n1249 ) | ( n838 & n4507 ) | ( ~n1249 & n4507 ) ;
  assign n4509 = n2236 | n4508 ;
  assign n4510 = n4509 ^ n1454 ^ 1'b0 ;
  assign n4511 = x0 | n1725 ;
  assign n4512 = n4511 ^ n2523 ^ 1'b0 ;
  assign n4513 = n4083 ^ n2131 ^ n1324 ;
  assign n4514 = n3513 ^ n796 ^ 1'b0 ;
  assign n4515 = n251 & n4514 ;
  assign n4516 = ~n2282 & n4515 ;
  assign n4517 = n4516 ^ n3262 ^ 1'b0 ;
  assign n4518 = n860 | n4259 ;
  assign n4519 = n4518 ^ n1162 ^ 1'b0 ;
  assign n4520 = n298 ^ x117 ^ 1'b0 ;
  assign n4521 = x39 & ~n4520 ;
  assign n4522 = n1292 | n1980 ;
  assign n4523 = n4522 ^ n1680 ^ 1'b0 ;
  assign n4524 = ( n3951 & n4521 ) | ( n3951 & ~n4523 ) | ( n4521 & ~n4523 ) ;
  assign n4525 = n2819 ^ n2809 ^ n2693 ;
  assign n4526 = ( n726 & n1327 ) | ( n726 & ~n3748 ) | ( n1327 & ~n3748 ) ;
  assign n4527 = ( x31 & ~n4214 ) | ( x31 & n4320 ) | ( ~n4214 & n4320 ) ;
  assign n4537 = n713 & n2721 ;
  assign n4538 = n4537 ^ n477 ^ 1'b0 ;
  assign n4539 = n4538 ^ n2770 ^ n169 ;
  assign n4540 = ~x123 & n2954 ;
  assign n4541 = n4539 & n4540 ;
  assign n4528 = n2575 ^ n1803 ^ 1'b0 ;
  assign n4529 = n1713 | n4528 ;
  assign n4530 = n2530 & ~n4529 ;
  assign n4531 = n3043 & ~n4530 ;
  assign n4532 = ~n236 & n4531 ;
  assign n4533 = ( ~n1373 & n1799 ) | ( ~n1373 & n2622 ) | ( n1799 & n2622 ) ;
  assign n4534 = n1584 | n4533 ;
  assign n4535 = n4532 & ~n4534 ;
  assign n4536 = n679 & ~n4535 ;
  assign n4542 = n4541 ^ n4536 ^ 1'b0 ;
  assign n4543 = n4373 ^ n1986 ^ 1'b0 ;
  assign n4544 = n521 & ~n4376 ;
  assign n4545 = n1784 ^ n1408 ^ 1'b0 ;
  assign n4546 = n4393 | n4545 ;
  assign n4549 = n1608 ^ n1595 ^ n739 ;
  assign n4547 = n494 | n3323 ;
  assign n4548 = n877 | n4547 ;
  assign n4550 = n4549 ^ n4548 ^ 1'b0 ;
  assign n4551 = ~n4546 & n4550 ;
  assign n4552 = n4551 ^ n1977 ^ 1'b0 ;
  assign n4553 = n4013 ^ n2619 ^ n2355 ;
  assign n4554 = n573 & n694 ;
  assign n4555 = ( n2552 & n2751 ) | ( n2552 & n4554 ) | ( n2751 & n4554 ) ;
  assign n4556 = ( n980 & n1302 ) | ( n980 & n2444 ) | ( n1302 & n2444 ) ;
  assign n4557 = n2478 | n4556 ;
  assign n4558 = n1306 & ~n3019 ;
  assign n4559 = n4558 ^ n1971 ^ 1'b0 ;
  assign n4560 = n493 & ~n3576 ;
  assign n4561 = n1555 & n4560 ;
  assign n4562 = n2785 & n4561 ;
  assign n4570 = ( ~n1550 & n1633 ) | ( ~n1550 & n2272 ) | ( n1633 & n2272 ) ;
  assign n4571 = ( n827 & n1918 ) | ( n827 & ~n4570 ) | ( n1918 & ~n4570 ) ;
  assign n4565 = n1228 | n1591 ;
  assign n4566 = n4565 ^ n2637 ^ 1'b0 ;
  assign n4567 = n3045 & ~n4566 ;
  assign n4568 = n2481 & n4567 ;
  assign n4569 = n747 & n4568 ;
  assign n4563 = n1362 ^ x123 ^ 1'b0 ;
  assign n4564 = n3522 & ~n4563 ;
  assign n4572 = n4571 ^ n4569 ^ n4564 ;
  assign n4573 = n1164 | n1342 ;
  assign n4574 = n1874 | n4573 ;
  assign n4575 = n233 & n4574 ;
  assign n4576 = n4575 ^ n4172 ^ 1'b0 ;
  assign n4577 = n589 & n1502 ;
  assign n4578 = n4577 ^ n663 ^ 1'b0 ;
  assign n4579 = n2499 & ~n4578 ;
  assign n4580 = n4579 ^ n690 ^ 1'b0 ;
  assign n4581 = n4393 ^ n877 ^ x45 ;
  assign n4582 = n1046 & n2089 ;
  assign n4583 = ~n4581 & n4582 ;
  assign n4584 = ( n2169 & n2663 ) | ( n2169 & n4583 ) | ( n2663 & n4583 ) ;
  assign n4585 = ~n506 & n1745 ;
  assign n4586 = ( ~n2470 & n4584 ) | ( ~n2470 & n4585 ) | ( n4584 & n4585 ) ;
  assign n4587 = n4586 ^ n2280 ^ 1'b0 ;
  assign n4588 = ~n3615 & n4587 ;
  assign n4589 = n521 | n4213 ;
  assign n4590 = n4589 ^ n1336 ^ 1'b0 ;
  assign n4591 = n1567 & ~n4392 ;
  assign n4592 = n4591 ^ n927 ^ n686 ;
  assign n4593 = n1967 ^ n1617 ^ 1'b0 ;
  assign n4594 = n4592 & ~n4593 ;
  assign n4597 = n2917 ^ n2643 ^ n1198 ;
  assign n4595 = ~n1895 & n2128 ;
  assign n4596 = n4595 ^ n1833 ^ 1'b0 ;
  assign n4598 = n4597 ^ n4596 ^ n410 ;
  assign n4599 = n3939 ^ n3376 ^ n2767 ;
  assign n4600 = n4599 ^ n3672 ^ 1'b0 ;
  assign n4605 = ( ~x49 & n537 ) | ( ~x49 & n582 ) | ( n537 & n582 ) ;
  assign n4606 = n922 ^ n256 ^ 1'b0 ;
  assign n4607 = n4605 & ~n4606 ;
  assign n4601 = n1156 & ~n1476 ;
  assign n4602 = n920 & n4601 ;
  assign n4603 = n4602 ^ n1669 ^ 1'b0 ;
  assign n4604 = n2133 | n4603 ;
  assign n4608 = n4607 ^ n4604 ^ 1'b0 ;
  assign n4609 = ( n753 & ~n2386 ) | ( n753 & n2878 ) | ( ~n2386 & n2878 ) ;
  assign n4610 = ~n1090 & n2038 ;
  assign n4611 = n4609 & n4610 ;
  assign n4612 = n4611 ^ n499 ^ 1'b0 ;
  assign n4613 = n1147 | n3665 ;
  assign n4614 = n4613 ^ n3539 ^ 1'b0 ;
  assign n4615 = n530 | n4614 ;
  assign n4616 = x53 & n2042 ;
  assign n4617 = ( n520 & n1603 ) | ( n520 & n2042 ) | ( n1603 & n2042 ) ;
  assign n4618 = n3926 ^ n1214 ^ x81 ;
  assign n4619 = ~n4617 & n4618 ;
  assign n4620 = n4574 ^ n2361 ^ 1'b0 ;
  assign n4621 = ( ~n2146 & n4619 ) | ( ~n2146 & n4620 ) | ( n4619 & n4620 ) ;
  assign n4622 = n4621 ^ n2555 ^ 1'b0 ;
  assign n4623 = n4616 & n4622 ;
  assign n4624 = n4623 ^ n2085 ^ 1'b0 ;
  assign n4625 = n1890 & n4624 ;
  assign n4630 = n201 & n2724 ;
  assign n4631 = ~n178 & n4630 ;
  assign n4629 = n1833 & n2795 ;
  assign n4632 = n4631 ^ n4629 ^ 1'b0 ;
  assign n4626 = n2816 & n3688 ;
  assign n4627 = n3024 & n4626 ;
  assign n4628 = n4539 & ~n4627 ;
  assign n4633 = n4632 ^ n4628 ^ n803 ;
  assign n4634 = ( ~n165 & n221 ) | ( ~n165 & n992 ) | ( n221 & n992 ) ;
  assign n4635 = n3187 ^ n2460 ^ 1'b0 ;
  assign n4636 = n4634 & ~n4635 ;
  assign n4640 = n2557 ^ n988 ^ 1'b0 ;
  assign n4641 = n2698 | n4640 ;
  assign n4637 = n562 ^ n290 ^ 1'b0 ;
  assign n4638 = x18 & ~n4637 ;
  assign n4639 = ( ~n521 & n2499 ) | ( ~n521 & n4638 ) | ( n2499 & n4638 ) ;
  assign n4642 = n4641 ^ n4639 ^ n212 ;
  assign n4643 = n4636 & ~n4642 ;
  assign n4644 = n4633 & n4643 ;
  assign n4645 = n2760 ^ n1080 ^ 1'b0 ;
  assign n4646 = n1436 & ~n4645 ;
  assign n4647 = ( x91 & n3252 ) | ( x91 & ~n4646 ) | ( n3252 & ~n4646 ) ;
  assign n4648 = n3926 ^ n3859 ^ 1'b0 ;
  assign n4649 = n4394 & ~n4648 ;
  assign n4650 = ( n618 & n2443 ) | ( n618 & n3134 ) | ( n2443 & n3134 ) ;
  assign n4651 = n367 & n3307 ;
  assign n4652 = n4651 ^ n247 ^ 1'b0 ;
  assign n4653 = n4652 ^ n4169 ^ n2800 ;
  assign n4654 = n958 | n1196 ;
  assign n4655 = n3819 ^ n1067 ^ 1'b0 ;
  assign n4656 = n2658 & ~n4655 ;
  assign n4657 = ~n4654 & n4656 ;
  assign n4658 = ~n1166 & n1819 ;
  assign n4659 = n4289 ^ n339 ^ 1'b0 ;
  assign n4660 = n4658 & n4659 ;
  assign n4661 = ( n979 & n2304 ) | ( n979 & ~n4610 ) | ( n2304 & ~n4610 ) ;
  assign n4662 = n3512 ^ n2584 ^ n1515 ;
  assign n4663 = n819 & n2136 ;
  assign n4664 = ( n1106 & ~n1545 ) | ( n1106 & n4663 ) | ( ~n1545 & n4663 ) ;
  assign n4665 = x98 | n4664 ;
  assign n4666 = n270 | n1841 ;
  assign n4667 = n3999 | n4666 ;
  assign n4668 = ~n4665 & n4667 ;
  assign n4669 = n1871 & n4668 ;
  assign n4670 = n2638 | n4669 ;
  assign n4671 = ~n3388 & n4670 ;
  assign n4672 = n3084 ^ n2097 ^ 1'b0 ;
  assign n4673 = n4078 & ~n4672 ;
  assign n4675 = n3948 ^ n839 ^ x64 ;
  assign n4676 = n339 & n908 ;
  assign n4677 = ~n1887 & n4676 ;
  assign n4678 = ~n4675 & n4677 ;
  assign n4674 = n3236 ^ n1427 ^ n511 ;
  assign n4679 = n4678 ^ n4674 ^ n1955 ;
  assign n4680 = n1633 & n2063 ;
  assign n4681 = n2304 ^ n626 ^ 1'b0 ;
  assign n4684 = n1617 & n2212 ;
  assign n4685 = n816 & n4684 ;
  assign n4686 = n4685 ^ n1953 ^ n1485 ;
  assign n4682 = n1914 ^ n214 ^ x117 ;
  assign n4683 = x64 & n4682 ;
  assign n4687 = n4686 ^ n4683 ^ 1'b0 ;
  assign n4688 = n251 | n2203 ;
  assign n4693 = n265 & ~n1896 ;
  assign n4694 = n4693 ^ n3968 ^ 1'b0 ;
  assign n4689 = n3655 ^ n1162 ^ n704 ;
  assign n4690 = n163 | n196 ;
  assign n4691 = n4690 ^ n3144 ^ 1'b0 ;
  assign n4692 = ~n4689 & n4691 ;
  assign n4695 = n4694 ^ n4692 ^ 1'b0 ;
  assign n4696 = ~n4688 & n4695 ;
  assign n4697 = n1501 & n4077 ;
  assign n4698 = ( n293 & ~n803 ) | ( n293 & n4062 ) | ( ~n803 & n4062 ) ;
  assign n4699 = n4698 ^ n4154 ^ 1'b0 ;
  assign n4700 = n1748 | n4699 ;
  assign n4701 = n221 & ~n2507 ;
  assign n4702 = x45 & x111 ;
  assign n4703 = n4702 ^ n2846 ^ 1'b0 ;
  assign n4704 = n4701 & ~n4703 ;
  assign n4705 = n203 | n274 ;
  assign n4706 = n4705 ^ n4658 ^ 1'b0 ;
  assign n4707 = n4706 ^ n1882 ^ n246 ;
  assign n4709 = n2964 ^ n2072 ^ n2034 ;
  assign n4708 = ~n1078 & n4277 ;
  assign n4710 = n4709 ^ n4708 ^ n2772 ;
  assign n4711 = x25 & n580 ;
  assign n4712 = n4711 ^ n730 ^ 1'b0 ;
  assign n4713 = n4712 ^ n3933 ^ n2844 ;
  assign n4714 = n4402 ^ n4252 ^ 1'b0 ;
  assign n4715 = n2125 & ~n2844 ;
  assign n4716 = n449 & n4715 ;
  assign n4717 = n4091 ^ n2651 ^ n986 ;
  assign n4718 = n4717 ^ n4592 ^ 1'b0 ;
  assign n4719 = n2372 & n4247 ;
  assign n4720 = n4719 ^ n1660 ^ 1'b0 ;
  assign n4723 = ( n378 & n1803 ) | ( n378 & ~n3485 ) | ( n1803 & ~n3485 ) ;
  assign n4721 = n1165 ^ n167 ^ 1'b0 ;
  assign n4722 = n4664 & ~n4721 ;
  assign n4724 = n4723 ^ n4722 ^ 1'b0 ;
  assign n4725 = ~n2976 & n4383 ;
  assign n4726 = ~n4209 & n4725 ;
  assign n4727 = n2471 ^ n1550 ^ 1'b0 ;
  assign n4728 = ~n771 & n4727 ;
  assign n4729 = n290 & ~n578 ;
  assign n4730 = n4729 ^ n3356 ^ 1'b0 ;
  assign n4731 = n4730 ^ n2868 ^ n927 ;
  assign n4732 = x88 & n4731 ;
  assign n4733 = n4732 ^ n3914 ^ 1'b0 ;
  assign n4734 = ( n225 & n618 ) | ( n225 & n2680 ) | ( n618 & n2680 ) ;
  assign n4735 = ( n1895 & n3844 ) | ( n1895 & ~n4734 ) | ( n3844 & ~n4734 ) ;
  assign n4736 = n1680 & n4735 ;
  assign n4737 = n3549 & n4736 ;
  assign n4738 = ( n535 & n1000 ) | ( n535 & n4392 ) | ( n1000 & n4392 ) ;
  assign n4739 = n4738 ^ n1666 ^ n427 ;
  assign n4740 = n4737 | n4739 ;
  assign n4741 = n4740 ^ n2497 ^ 1'b0 ;
  assign n4742 = n3072 ^ n2575 ^ x67 ;
  assign n4743 = n4742 ^ n2046 ^ 1'b0 ;
  assign n4744 = n3886 ^ x64 ^ 1'b0 ;
  assign n4745 = n1767 | n4744 ;
  assign n4746 = ~n578 & n820 ;
  assign n4747 = n653 & n4746 ;
  assign n4748 = n2710 & n4747 ;
  assign n4752 = n2418 ^ n1631 ^ 1'b0 ;
  assign n4753 = n511 & n4752 ;
  assign n4749 = ~n234 & n2138 ;
  assign n4750 = x11 & x54 ;
  assign n4751 = n4749 & n4750 ;
  assign n4754 = n4753 ^ n4751 ^ n739 ;
  assign n4755 = n1297 ^ n618 ^ 1'b0 ;
  assign n4756 = ~n1205 & n4755 ;
  assign n4757 = n3506 | n4544 ;
  assign n4758 = n675 ^ x108 ^ 1'b0 ;
  assign n4759 = n760 & ~n1093 ;
  assign n4760 = n4758 & n4759 ;
  assign n4761 = n2328 & n4760 ;
  assign n4762 = n4761 ^ n2939 ^ n890 ;
  assign n4766 = n1694 ^ n726 ^ 1'b0 ;
  assign n4767 = x50 & ~n4766 ;
  assign n4764 = ( ~x100 & n796 ) | ( ~x100 & n1318 ) | ( n796 & n1318 ) ;
  assign n4763 = ~n731 & n4467 ;
  assign n4765 = n4764 ^ n4763 ^ 1'b0 ;
  assign n4768 = n4767 ^ n4765 ^ n1116 ;
  assign n4769 = n4739 ^ n2919 ^ 1'b0 ;
  assign n4770 = n1195 & ~n4769 ;
  assign n4771 = n2624 | n4392 ;
  assign n4772 = n2364 & ~n4771 ;
  assign n4773 = ~n2894 & n3045 ;
  assign n4774 = ~n4676 & n4773 ;
  assign n4775 = n518 & ~n4774 ;
  assign n4776 = n4775 ^ n1949 ^ 1'b0 ;
  assign n4777 = n4776 ^ n1972 ^ 1'b0 ;
  assign n4778 = n4306 ^ n3297 ^ 1'b0 ;
  assign n4779 = n2094 ^ n1370 ^ n223 ;
  assign n4780 = x85 & n936 ;
  assign n4781 = n4780 ^ n1643 ^ 1'b0 ;
  assign n4782 = ~n4779 & n4781 ;
  assign n4783 = n4782 ^ n3958 ^ 1'b0 ;
  assign n4784 = n1499 | n2770 ;
  assign n4785 = n2601 | n4784 ;
  assign n4786 = n356 & n1242 ;
  assign n4787 = ~n1311 & n4786 ;
  assign n4788 = ( n1683 & ~n2171 ) | ( n1683 & n4787 ) | ( ~n2171 & n4787 ) ;
  assign n4789 = n4788 ^ n3796 ^ 1'b0 ;
  assign n4790 = n3747 ^ n787 ^ 1'b0 ;
  assign n4793 = n3262 ^ n2413 ^ n859 ;
  assign n4791 = n1503 | n2352 ;
  assign n4792 = n4791 ^ n1893 ^ 1'b0 ;
  assign n4794 = n4793 ^ n4792 ^ n1923 ;
  assign n4795 = n2574 ^ n2141 ^ n746 ;
  assign n4796 = n2834 | n4795 ;
  assign n4797 = n1478 | n4796 ;
  assign n4798 = n3491 ^ n1307 ^ n381 ;
  assign n4799 = n2517 & n3098 ;
  assign n4800 = n4798 & n4799 ;
  assign n4801 = n4800 ^ n4147 ^ n639 ;
  assign n4802 = ( n1150 & n3163 ) | ( n1150 & ~n4737 ) | ( n3163 & ~n4737 ) ;
  assign n4803 = n4802 ^ n1435 ^ 1'b0 ;
  assign n4804 = ~n699 & n2743 ;
  assign n4805 = n4804 ^ n3093 ^ 1'b0 ;
  assign n4806 = n4805 ^ n2390 ^ 1'b0 ;
  assign n4807 = ~n480 & n4806 ;
  assign n4808 = ~n746 & n4807 ;
  assign n4809 = ( ~n157 & n485 ) | ( ~n157 & n2106 ) | ( n485 & n2106 ) ;
  assign n4810 = n2031 & ~n4809 ;
  assign n4811 = n4248 ^ n3524 ^ 1'b0 ;
  assign n4812 = n979 ^ x8 ^ 1'b0 ;
  assign n4813 = n2688 & ~n4812 ;
  assign n4814 = ( n2449 & n4243 ) | ( n2449 & n4813 ) | ( n4243 & n4813 ) ;
  assign n4815 = n1967 ^ n1441 ^ 1'b0 ;
  assign n4816 = n1179 & ~n1725 ;
  assign n4817 = ( n3798 & ~n4815 ) | ( n3798 & n4816 ) | ( ~n4815 & n4816 ) ;
  assign n4818 = n4714 & ~n4817 ;
  assign n4819 = ~n4814 & n4818 ;
  assign n4821 = n3190 ^ n2349 ^ 1'b0 ;
  assign n4820 = ( n705 & n1481 ) | ( n705 & n2328 ) | ( n1481 & n2328 ) ;
  assign n4822 = n4821 ^ n4820 ^ n3027 ;
  assign n4823 = n2192 | n2719 ;
  assign n4824 = n983 | n4823 ;
  assign n4825 = x90 & n4824 ;
  assign n4826 = n4825 ^ n1822 ^ 1'b0 ;
  assign n4827 = n3440 & n3831 ;
  assign n4828 = ( ~n3338 & n4826 ) | ( ~n3338 & n4827 ) | ( n4826 & n4827 ) ;
  assign n4829 = n4570 ^ n2180 ^ 1'b0 ;
  assign n4830 = ( ~n825 & n4495 ) | ( ~n825 & n4829 ) | ( n4495 & n4829 ) ;
  assign n4831 = n1305 & ~n3971 ;
  assign n4832 = n4830 & n4831 ;
  assign n4833 = n3877 ^ n1074 ^ n478 ;
  assign n4834 = n4833 ^ n4567 ^ n2945 ;
  assign n4835 = n4834 ^ n2816 ^ 1'b0 ;
  assign n4838 = x20 & n2456 ;
  assign n4839 = n4838 ^ n984 ^ 1'b0 ;
  assign n4836 = n701 | n3587 ;
  assign n4837 = n4836 ^ n2481 ^ 1'b0 ;
  assign n4840 = n4839 ^ n4837 ^ 1'b0 ;
  assign n4841 = ( n502 & ~n553 ) | ( n502 & n2122 ) | ( ~n553 & n2122 ) ;
  assign n4842 = n2705 & n4841 ;
  assign n4843 = n4840 & n4842 ;
  assign n4846 = n327 & n3017 ;
  assign n4847 = n4846 ^ n2682 ^ 1'b0 ;
  assign n4844 = n2344 ^ n1692 ^ 1'b0 ;
  assign n4845 = n1822 & n4844 ;
  assign n4848 = n4847 ^ n4845 ^ 1'b0 ;
  assign n4849 = ~n2261 & n4848 ;
  assign n4850 = n2799 ^ n157 ^ 1'b0 ;
  assign n4851 = n1982 | n2771 ;
  assign n4852 = n4851 ^ x23 ^ 1'b0 ;
  assign n4856 = n2182 ^ x3 ^ 1'b0 ;
  assign n4857 = ~n3693 & n4856 ;
  assign n4853 = n594 & n2382 ;
  assign n4854 = ( n1216 & n1798 ) | ( n1216 & ~n2117 ) | ( n1798 & ~n2117 ) ;
  assign n4855 = ( ~n247 & n4853 ) | ( ~n247 & n4854 ) | ( n4853 & n4854 ) ;
  assign n4858 = n4857 ^ n4855 ^ n1515 ;
  assign n4859 = n4858 ^ n451 ^ 1'b0 ;
  assign n4860 = n2508 ^ n1292 ^ 1'b0 ;
  assign n4861 = n3651 ^ n2202 ^ 1'b0 ;
  assign n4867 = n4271 ^ n3871 ^ 1'b0 ;
  assign n4863 = n1378 ^ n827 ^ n420 ;
  assign n4862 = n4521 ^ n1528 ^ n1094 ;
  assign n4864 = n4863 ^ n4862 ^ 1'b0 ;
  assign n4865 = n3693 & n4864 ;
  assign n4866 = ( ~n367 & n3119 ) | ( ~n367 & n4865 ) | ( n3119 & n4865 ) ;
  assign n4868 = n4867 ^ n4866 ^ 1'b0 ;
  assign n4869 = n546 & n1656 ;
  assign n4870 = n4869 ^ n4191 ^ 1'b0 ;
  assign n4872 = n2278 ^ n2041 ^ 1'b0 ;
  assign n4871 = n3092 ^ n1810 ^ n1317 ;
  assign n4873 = n4872 ^ n4871 ^ 1'b0 ;
  assign n4874 = n293 & ~n4873 ;
  assign n4875 = ~n4870 & n4874 ;
  assign n4876 = n993 ^ n608 ^ 1'b0 ;
  assign n4877 = n3356 & ~n4876 ;
  assign n4878 = n4877 ^ n820 ^ 1'b0 ;
  assign n4879 = n169 & n300 ;
  assign n4880 = n3523 & ~n4879 ;
  assign n4881 = ~n4878 & n4880 ;
  assign n4882 = n1129 & ~n4881 ;
  assign n4883 = n663 & ~n1053 ;
  assign n4884 = n4883 ^ n601 ^ 1'b0 ;
  assign n4885 = n1760 ^ n1096 ^ n220 ;
  assign n4886 = n2553 & n3636 ;
  assign n4887 = ~n4885 & n4886 ;
  assign n4888 = n4887 ^ n4795 ^ 1'b0 ;
  assign n4889 = n2019 & n4888 ;
  assign n4890 = n1674 | n4433 ;
  assign n4891 = n4890 ^ n2789 ^ n1210 ;
  assign n4892 = ~n2174 & n4235 ;
  assign n4893 = n4891 & n4892 ;
  assign n4894 = n1892 | n4893 ;
  assign n4895 = n4894 ^ n2285 ^ 1'b0 ;
  assign n4896 = n4895 ^ n3674 ^ 1'b0 ;
  assign n4897 = n1499 ^ x35 ^ 1'b0 ;
  assign n4898 = n4897 ^ n1611 ^ n1545 ;
  assign n4899 = n4898 ^ n358 ^ 1'b0 ;
  assign n4900 = ( n1352 & ~n1672 ) | ( n1352 & n2258 ) | ( ~n1672 & n2258 ) ;
  assign n4901 = n4900 ^ n2285 ^ 1'b0 ;
  assign n4902 = n4070 & ~n4584 ;
  assign n4903 = n299 | n794 ;
  assign n4904 = n4903 ^ n721 ^ 1'b0 ;
  assign n4905 = n4904 ^ n4219 ^ 1'b0 ;
  assign n4906 = ( n3831 & n4902 ) | ( n3831 & ~n4905 ) | ( n4902 & ~n4905 ) ;
  assign n4907 = n286 & ~n2002 ;
  assign n4908 = n4907 ^ n265 ^ 1'b0 ;
  assign n4909 = n4908 ^ n4444 ^ n4182 ;
  assign n4910 = n475 | n1906 ;
  assign n4911 = n4910 ^ n1082 ^ 1'b0 ;
  assign n4912 = n4911 ^ n162 ^ 1'b0 ;
  assign n4913 = ~n3798 & n4912 ;
  assign n4914 = ( n901 & ~n1216 ) | ( n901 & n1575 ) | ( ~n1216 & n1575 ) ;
  assign n4915 = ( ~x98 & n415 ) | ( ~x98 & n2237 ) | ( n415 & n2237 ) ;
  assign n4916 = ( n1057 & n4578 ) | ( n1057 & n4915 ) | ( n4578 & n4915 ) ;
  assign n4917 = ( n496 & n1104 ) | ( n496 & n1127 ) | ( n1104 & n1127 ) ;
  assign n4918 = n3038 ^ x79 ^ 1'b0 ;
  assign n4919 = ~n1776 & n4918 ;
  assign n4920 = x91 & ~n2491 ;
  assign n4921 = ~n4919 & n4920 ;
  assign n4922 = n4917 & ~n4921 ;
  assign n4923 = n4922 ^ n4367 ^ 1'b0 ;
  assign n4924 = n746 | n4923 ;
  assign n4925 = n2364 & n3428 ;
  assign n4926 = n2451 ^ n1848 ^ 1'b0 ;
  assign n4927 = n4117 ^ n258 ^ 1'b0 ;
  assign n4928 = ~n909 & n2662 ;
  assign n4929 = ~n2055 & n4928 ;
  assign n4930 = n4927 | n4929 ;
  assign n4931 = n4930 ^ n1546 ^ 1'b0 ;
  assign n4932 = n1593 | n4931 ;
  assign n4933 = n4926 & ~n4932 ;
  assign n4934 = n4394 ^ x43 ^ 1'b0 ;
  assign n4935 = n831 ^ n323 ^ x26 ;
  assign n4936 = n815 & n1744 ;
  assign n4937 = n4936 ^ n808 ^ 1'b0 ;
  assign n4938 = n4935 & n4937 ;
  assign n4939 = ( ~n852 & n1129 ) | ( ~n852 & n3862 ) | ( n1129 & n3862 ) ;
  assign n4940 = n4199 ^ n3854 ^ n485 ;
  assign n4941 = n4940 ^ n1338 ^ n193 ;
  assign n4942 = ( ~n1680 & n3586 ) | ( ~n1680 & n3917 ) | ( n3586 & n3917 ) ;
  assign n4943 = n4942 ^ n4049 ^ 1'b0 ;
  assign n4944 = n1433 | n1834 ;
  assign n4945 = n4944 ^ n2458 ^ 1'b0 ;
  assign n4946 = ~n3539 & n4945 ;
  assign n4947 = ~n578 & n3362 ;
  assign n4948 = ~n4946 & n4947 ;
  assign n4949 = n1720 ^ n1715 ^ 1'b0 ;
  assign n4950 = n2462 & n4949 ;
  assign n4951 = n2562 & n3689 ;
  assign n4952 = n4951 ^ n2415 ^ n285 ;
  assign n4953 = n4359 & n4952 ;
  assign n4954 = ~n4950 & n4953 ;
  assign n4955 = n4593 ^ n827 ^ 1'b0 ;
  assign n4956 = n4081 ^ n312 ^ 1'b0 ;
  assign n4957 = ( n487 & ~n4955 ) | ( n487 & n4956 ) | ( ~n4955 & n4956 ) ;
  assign n4958 = n4957 ^ n4749 ^ n3146 ;
  assign n4959 = ~n755 & n897 ;
  assign n4960 = n4959 ^ n1477 ^ 1'b0 ;
  assign n4961 = n617 & n4960 ;
  assign n4962 = n2203 ^ n471 ^ 1'b0 ;
  assign n4963 = n2148 & n4962 ;
  assign n4964 = ~n3076 & n4963 ;
  assign n4965 = x105 & ~n4483 ;
  assign n4966 = n4965 ^ n3803 ^ 1'b0 ;
  assign n4967 = ( n537 & n3127 ) | ( n537 & ~n4328 ) | ( n3127 & ~n4328 ) ;
  assign n4968 = n3763 ^ n2591 ^ 1'b0 ;
  assign n4969 = ~n2163 & n4968 ;
  assign n4970 = ~n746 & n1216 ;
  assign n4971 = n4000 & n4970 ;
  assign n4972 = n4969 & n4971 ;
  assign n4973 = n4972 ^ n1394 ^ 1'b0 ;
  assign n4974 = n4147 ^ n3921 ^ 1'b0 ;
  assign n4975 = ~n4973 & n4974 ;
  assign n4976 = n4106 ^ n2451 ^ 1'b0 ;
  assign n4977 = n3534 | n4976 ;
  assign n4978 = n4059 & ~n4977 ;
  assign n4979 = n4144 ^ n1152 ^ 1'b0 ;
  assign n4980 = x12 & ~n4178 ;
  assign n4981 = ~n4313 & n4980 ;
  assign n4982 = n2873 ^ n2044 ^ n1575 ;
  assign n4983 = ~n4981 & n4982 ;
  assign n4984 = n4511 ^ n879 ^ 1'b0 ;
  assign n4985 = n4485 & ~n4984 ;
  assign n4986 = n3792 & n4985 ;
  assign n4987 = n4403 ^ x36 ^ 1'b0 ;
  assign n4988 = ~n4184 & n4987 ;
  assign n4989 = ~x64 & n3568 ;
  assign n4990 = n2081 ^ n1382 ^ 1'b0 ;
  assign n4991 = n2418 & n4990 ;
  assign n4992 = ~n601 & n4991 ;
  assign n4993 = n4332 & n4992 ;
  assign n4994 = n4660 ^ n3355 ^ n2615 ;
  assign n4995 = x106 ^ x43 ^ 1'b0 ;
  assign n4996 = ( n261 & n2228 ) | ( n261 & ~n4995 ) | ( n2228 & ~n4995 ) ;
  assign n4997 = n209 & ~n4996 ;
  assign n4998 = n622 ^ n222 ^ 1'b0 ;
  assign n4999 = ~n2971 & n4998 ;
  assign n5000 = x122 & n251 ;
  assign n5001 = n2290 ^ n2072 ^ x40 ;
  assign n5002 = n5000 | n5001 ;
  assign n5003 = ~n1430 & n4449 ;
  assign n5004 = n2137 & ~n4583 ;
  assign n5005 = n5004 ^ n1696 ^ 1'b0 ;
  assign n5006 = n3642 ^ x35 ^ 1'b0 ;
  assign n5007 = n5006 ^ n4654 ^ 1'b0 ;
  assign n5008 = n5007 ^ n355 ^ 1'b0 ;
  assign n5009 = ( x31 & n5005 ) | ( x31 & n5008 ) | ( n5005 & n5008 ) ;
  assign n5010 = n5009 ^ n1529 ^ 1'b0 ;
  assign n5011 = n5010 ^ n726 ^ 1'b0 ;
  assign n5012 = n2188 ^ n1440 ^ 1'b0 ;
  assign n5016 = n1642 ^ n383 ^ 1'b0 ;
  assign n5013 = n740 & ~n1908 ;
  assign n5014 = ( n2795 & n3871 ) | ( n2795 & n5013 ) | ( n3871 & n5013 ) ;
  assign n5015 = n2939 & n5014 ;
  assign n5017 = n5016 ^ n5015 ^ 1'b0 ;
  assign n5018 = ( n1513 & n4218 ) | ( n1513 & n5017 ) | ( n4218 & n5017 ) ;
  assign n5020 = n1797 ^ x58 ^ 1'b0 ;
  assign n5021 = n5020 ^ n2744 ^ 1'b0 ;
  assign n5019 = n1240 | n2800 ;
  assign n5022 = n5021 ^ n5019 ^ 1'b0 ;
  assign n5023 = n3981 ^ n2150 ^ 1'b0 ;
  assign n5024 = n2837 | n5023 ;
  assign n5025 = n4841 & ~n5024 ;
  assign n5026 = ~n1855 & n5025 ;
  assign n5029 = n190 | n4456 ;
  assign n5030 = n5029 ^ n2315 ^ 1'b0 ;
  assign n5031 = n485 & n5030 ;
  assign n5028 = n1855 & n3326 ;
  assign n5032 = n5031 ^ n5028 ^ 1'b0 ;
  assign n5033 = n3951 & ~n5032 ;
  assign n5034 = n252 & ~n2860 ;
  assign n5035 = n5034 ^ n1713 ^ n334 ;
  assign n5036 = n5033 & n5035 ;
  assign n5027 = n1408 ^ n447 ^ 1'b0 ;
  assign n5037 = n5036 ^ n5027 ^ 1'b0 ;
  assign n5038 = n1731 ^ n536 ^ 1'b0 ;
  assign n5039 = n4137 ^ n2628 ^ 1'b0 ;
  assign n5040 = n1035 & ~n5039 ;
  assign n5041 = n4061 ^ n1812 ^ 1'b0 ;
  assign n5042 = n504 | n1014 ;
  assign n5043 = n5042 ^ n2831 ^ 1'b0 ;
  assign n5044 = n5043 ^ n1086 ^ 1'b0 ;
  assign n5045 = n3472 ^ n1800 ^ 1'b0 ;
  assign n5046 = n465 & n1534 ;
  assign n5047 = n1478 | n5046 ;
  assign n5048 = n1588 | n5047 ;
  assign n5049 = n1927 & ~n3533 ;
  assign n5050 = ( ~n631 & n2931 ) | ( ~n631 & n5049 ) | ( n2931 & n5049 ) ;
  assign n5051 = n5050 ^ n402 ^ 1'b0 ;
  assign n5052 = n831 | n3357 ;
  assign n5053 = n3878 & ~n5052 ;
  assign n5054 = ( n3447 & n3830 ) | ( n3447 & ~n4994 ) | ( n3830 & ~n4994 ) ;
  assign n5055 = n1227 & n3017 ;
  assign n5056 = ~n1268 & n5055 ;
  assign n5057 = n424 & n2962 ;
  assign n5058 = n1451 ^ n1089 ^ 1'b0 ;
  assign n5059 = n4263 | n4571 ;
  assign n5060 = ( n5031 & n5058 ) | ( n5031 & n5059 ) | ( n5058 & n5059 ) ;
  assign n5061 = ( n2905 & n5050 ) | ( n2905 & n5060 ) | ( n5050 & n5060 ) ;
  assign n5062 = n3123 | n4220 ;
  assign n5063 = n4429 | n5062 ;
  assign n5064 = ~n3339 & n5063 ;
  assign n5065 = n5064 ^ n4859 ^ 1'b0 ;
  assign n5066 = n3026 ^ x39 ^ 1'b0 ;
  assign n5067 = n2788 | n3262 ;
  assign n5068 = n3050 | n5067 ;
  assign n5069 = n3026 ^ n1993 ^ 1'b0 ;
  assign n5070 = n730 & ~n5069 ;
  assign n5074 = x46 & n2363 ;
  assign n5075 = ( n1626 & n2407 ) | ( n1626 & ~n5074 ) | ( n2407 & ~n5074 ) ;
  assign n5072 = n2039 & n3651 ;
  assign n5071 = ~n2894 & n3445 ;
  assign n5073 = n5072 ^ n5071 ^ 1'b0 ;
  assign n5076 = n5075 ^ n5073 ^ n4318 ;
  assign n5077 = n3978 ^ n3358 ^ n1345 ;
  assign n5078 = ( ~n1045 & n1435 ) | ( ~n1045 & n3291 ) | ( n1435 & n3291 ) ;
  assign n5079 = n4007 ^ n1760 ^ 1'b0 ;
  assign n5080 = n5079 ^ n146 ^ 1'b0 ;
  assign n5081 = ( n5077 & n5078 ) | ( n5077 & ~n5080 ) | ( n5078 & ~n5080 ) ;
  assign n5082 = n746 | n1817 ;
  assign n5083 = n5082 ^ n2133 ^ 1'b0 ;
  assign n5084 = n1996 ^ n349 ^ 1'b0 ;
  assign n5085 = ~n5083 & n5084 ;
  assign n5086 = ~n1496 & n5085 ;
  assign n5087 = n5086 ^ n4919 ^ 1'b0 ;
  assign n5088 = n152 & ~n3005 ;
  assign n5089 = ( n3778 & n4314 ) | ( n3778 & n5088 ) | ( n4314 & n5088 ) ;
  assign n5090 = n3939 ^ n2444 ^ n1057 ;
  assign n5103 = ( n293 & n740 ) | ( n293 & n1654 ) | ( n740 & n1654 ) ;
  assign n5101 = ~n412 & n3045 ;
  assign n5102 = n5101 ^ n4533 ^ 1'b0 ;
  assign n5095 = n1587 | n3482 ;
  assign n5096 = n1383 & ~n5095 ;
  assign n5097 = n1696 & ~n5096 ;
  assign n5098 = ~n2316 & n5097 ;
  assign n5093 = n2567 ^ n2409 ^ 1'b0 ;
  assign n5094 = ( n2054 & n4003 ) | ( n2054 & ~n5093 ) | ( n4003 & ~n5093 ) ;
  assign n5099 = n5098 ^ n5094 ^ n857 ;
  assign n5092 = n1585 & n4032 ;
  assign n5091 = ~n4043 & n4217 ;
  assign n5100 = n5099 ^ n5092 ^ n5091 ;
  assign n5104 = n5103 ^ n5102 ^ n5100 ;
  assign n5105 = n630 | n4249 ;
  assign n5106 = n1205 & ~n5105 ;
  assign n5107 = n3697 & n5106 ;
  assign n5108 = ~n2155 & n5107 ;
  assign n5109 = n2842 | n4927 ;
  assign n5110 = n5109 ^ x82 ^ 1'b0 ;
  assign n5111 = ( n718 & n1861 ) | ( n718 & ~n5110 ) | ( n1861 & ~n5110 ) ;
  assign n5112 = ( ~x56 & n1903 ) | ( ~x56 & n5111 ) | ( n1903 & n5111 ) ;
  assign n5113 = n4615 ^ n3945 ^ 1'b0 ;
  assign n5114 = n1518 ^ x98 ^ 1'b0 ;
  assign n5115 = n4717 & ~n5114 ;
  assign n5116 = n5115 ^ n4284 ^ 1'b0 ;
  assign n5119 = n2624 ^ n644 ^ 1'b0 ;
  assign n5120 = n4393 | n5119 ;
  assign n5121 = n5120 ^ n3485 ^ 1'b0 ;
  assign n5117 = n3791 ^ n3679 ^ n1522 ;
  assign n5118 = ( ~n1046 & n1622 ) | ( ~n1046 & n5117 ) | ( n1622 & n5117 ) ;
  assign n5122 = n5121 ^ n5118 ^ 1'b0 ;
  assign n5123 = n2226 & ~n5122 ;
  assign n5124 = ~n2903 & n5123 ;
  assign n5125 = n5124 ^ n4828 ^ 1'b0 ;
  assign n5128 = n2835 ^ n2243 ^ 1'b0 ;
  assign n5127 = x97 & ~n2233 ;
  assign n5129 = n5128 ^ n5127 ^ 1'b0 ;
  assign n5130 = ~n4336 & n5129 ;
  assign n5126 = ( n1640 & n3136 ) | ( n1640 & ~n4404 ) | ( n3136 & ~n4404 ) ;
  assign n5131 = n5130 ^ n5126 ^ n4710 ;
  assign n5132 = n3311 & ~n3917 ;
  assign n5133 = n847 | n5132 ;
  assign n5134 = n5133 ^ n3037 ^ 1'b0 ;
  assign n5137 = n2990 ^ n1894 ^ x74 ;
  assign n5138 = n5137 ^ n4675 ^ n1712 ;
  assign n5139 = n2285 ^ n2221 ^ n1634 ;
  assign n5140 = n1324 | n5139 ;
  assign n5141 = n5140 ^ n2731 ^ 1'b0 ;
  assign n5142 = n5141 ^ n261 ^ 1'b0 ;
  assign n5143 = n5138 | n5142 ;
  assign n5135 = n893 & ~n4826 ;
  assign n5136 = n2933 | n5135 ;
  assign n5144 = n5143 ^ n5136 ^ 1'b0 ;
  assign n5145 = n2322 & n5144 ;
  assign n5151 = n2056 & n3006 ;
  assign n5147 = ( n768 & n1485 ) | ( n768 & ~n1593 ) | ( n1485 & ~n1593 ) ;
  assign n5148 = n3330 & n5147 ;
  assign n5149 = n4203 & n5148 ;
  assign n5150 = n1731 & ~n5149 ;
  assign n5152 = n5151 ^ n5150 ^ 1'b0 ;
  assign n5146 = n1305 & n3628 ;
  assign n5153 = n5152 ^ n5146 ^ 1'b0 ;
  assign n5154 = n5153 ^ n637 ^ n533 ;
  assign n5155 = ( ~n946 & n2530 ) | ( ~n946 & n4619 ) | ( n2530 & n4619 ) ;
  assign n5156 = x82 & ~n5155 ;
  assign n5157 = n4085 ^ n331 ^ 1'b0 ;
  assign n5158 = n4978 & n5157 ;
  assign n5159 = n2304 ^ n1810 ^ 1'b0 ;
  assign n5160 = n5159 ^ n158 ^ 1'b0 ;
  assign n5161 = ~n571 & n4581 ;
  assign n5162 = n1675 ^ n1461 ^ 1'b0 ;
  assign n5163 = n340 | n3837 ;
  assign n5164 = n3477 & n5163 ;
  assign n5165 = n5162 | n5164 ;
  assign n5166 = n2493 & ~n3975 ;
  assign n5167 = n5166 ^ n4952 ^ n1198 ;
  assign n5169 = ~n1672 & n4462 ;
  assign n5168 = ( n145 & n310 ) | ( n145 & n925 ) | ( n310 & n925 ) ;
  assign n5170 = n5169 ^ n5168 ^ n5149 ;
  assign n5171 = n1020 ^ n177 ^ x79 ;
  assign n5172 = n3118 & n5171 ;
  assign n5175 = ~n579 & n1256 ;
  assign n5173 = n3364 | n4152 ;
  assign n5174 = n5074 | n5173 ;
  assign n5176 = n5175 ^ n5174 ^ 1'b0 ;
  assign n5177 = ( ~n2624 & n4854 ) | ( ~n2624 & n4973 ) | ( n4854 & n4973 ) ;
  assign n5178 = n3545 & n5177 ;
  assign n5179 = n2115 ^ n1906 ^ 1'b0 ;
  assign n5180 = n807 | n5179 ;
  assign n5181 = ( n938 & n1617 ) | ( n938 & ~n2515 ) | ( n1617 & ~n2515 ) ;
  assign n5187 = ( n1179 & n2906 ) | ( n1179 & n3651 ) | ( n2906 & n3651 ) ;
  assign n5182 = n2124 & ~n2413 ;
  assign n5183 = ~n825 & n5182 ;
  assign n5184 = n1929 & ~n5183 ;
  assign n5185 = ~n1931 & n5184 ;
  assign n5186 = ( ~n843 & n4922 ) | ( ~n843 & n5185 ) | ( n4922 & n5185 ) ;
  assign n5188 = n5187 ^ n5186 ^ 1'b0 ;
  assign n5189 = n5181 & ~n5188 ;
  assign n5190 = ~n186 & n3813 ;
  assign n5191 = ~n3278 & n5190 ;
  assign n5192 = n5189 | n5191 ;
  assign n5193 = n201 | n383 ;
  assign n5194 = n746 & ~n5193 ;
  assign n5195 = ~n1947 & n5194 ;
  assign n5196 = ~n620 & n5195 ;
  assign n5197 = ( n193 & ~n1214 ) | ( n193 & n1485 ) | ( ~n1214 & n1485 ) ;
  assign n5198 = n4029 & n5197 ;
  assign n5199 = n1260 & ~n4745 ;
  assign n5200 = n951 & n1897 ;
  assign n5201 = n5200 ^ n2029 ^ 1'b0 ;
  assign n5202 = n3016 & n5201 ;
  assign n5207 = n4234 ^ n3372 ^ x16 ;
  assign n5204 = n1725 & n2828 ;
  assign n5205 = n165 & n5204 ;
  assign n5203 = n2942 | n3482 ;
  assign n5206 = n5205 ^ n5203 ^ 1'b0 ;
  assign n5208 = n5207 ^ n5206 ^ n4191 ;
  assign n5209 = n4099 ^ n3689 ^ 1'b0 ;
  assign n5210 = n1218 & n5209 ;
  assign n5211 = n1205 & ~n1815 ;
  assign n5212 = n5211 ^ n2521 ^ 1'b0 ;
  assign n5213 = ( n1605 & ~n4267 ) | ( n1605 & n5212 ) | ( ~n4267 & n5212 ) ;
  assign n5216 = x1 | n489 ;
  assign n5217 = n5216 ^ n2867 ^ 1'b0 ;
  assign n5218 = n445 & ~n3734 ;
  assign n5219 = ~n5217 & n5218 ;
  assign n5220 = n309 & n1082 ;
  assign n5221 = n5220 ^ n654 ^ 1'b0 ;
  assign n5222 = n5221 ^ n129 ^ 1'b0 ;
  assign n5223 = ~n5219 & n5222 ;
  assign n5214 = n161 | n281 ;
  assign n5215 = n1854 & ~n5214 ;
  assign n5224 = n5223 ^ n5215 ^ 1'b0 ;
  assign n5225 = n3349 ^ n1939 ^ 1'b0 ;
  assign n5226 = n2328 ^ n1393 ^ 1'b0 ;
  assign n5227 = ( n870 & n2617 ) | ( n870 & n5226 ) | ( n2617 & n5226 ) ;
  assign n5230 = n749 | n778 ;
  assign n5228 = n362 & n1528 ;
  assign n5229 = ( n210 & n3961 ) | ( n210 & ~n5228 ) | ( n3961 & ~n5228 ) ;
  assign n5231 = n5230 ^ n5229 ^ n4397 ;
  assign n5232 = n3638 ^ n2262 ^ 1'b0 ;
  assign n5233 = n3186 | n5232 ;
  assign n5234 = n1672 & ~n2535 ;
  assign n5235 = n3323 ^ n256 ^ 1'b0 ;
  assign n5236 = n2127 & ~n4532 ;
  assign n5237 = n2337 ^ n693 ^ 1'b0 ;
  assign n5238 = n347 & n1415 ;
  assign n5239 = n5238 ^ n238 ^ 1'b0 ;
  assign n5240 = n3099 | n4238 ;
  assign n5241 = n5239 | n5240 ;
  assign n5242 = n5241 ^ n4249 ^ n143 ;
  assign n5243 = n4497 ^ n758 ^ n383 ;
  assign n5244 = n646 | n668 ;
  assign n5245 = n3221 ^ n2361 ^ 1'b0 ;
  assign n5246 = ( n4646 & n5244 ) | ( n4646 & ~n5245 ) | ( n5244 & ~n5245 ) ;
  assign n5250 = n5163 ^ n2316 ^ 1'b0 ;
  assign n5251 = n3866 | n5250 ;
  assign n5252 = n5251 ^ n709 ^ 1'b0 ;
  assign n5253 = n882 & ~n3143 ;
  assign n5254 = n3143 & n5253 ;
  assign n5255 = n5252 & n5254 ;
  assign n5247 = n2664 & n2783 ;
  assign n5248 = ~n4956 & n5247 ;
  assign n5249 = n4956 & n5248 ;
  assign n5256 = n5255 ^ n5249 ^ n487 ;
  assign n5261 = ~n1418 & n3600 ;
  assign n5262 = n1665 & n5261 ;
  assign n5263 = n5262 ^ n3019 ^ n1539 ;
  assign n5257 = ( n2395 & n4069 ) | ( n2395 & n5074 ) | ( n4069 & n5074 ) ;
  assign n5258 = n5257 ^ n4329 ^ 1'b0 ;
  assign n5259 = n2246 ^ n2212 ^ n802 ;
  assign n5260 = ( n4408 & n5258 ) | ( n4408 & n5259 ) | ( n5258 & n5259 ) ;
  assign n5264 = n5263 ^ n5260 ^ 1'b0 ;
  assign n5265 = x93 & ~n4110 ;
  assign n5266 = n956 & n3237 ;
  assign n5267 = n5266 ^ n3284 ^ 1'b0 ;
  assign n5268 = ~n2288 & n5267 ;
  assign n5269 = n5265 | n5268 ;
  assign n5270 = ~n211 & n5269 ;
  assign n5271 = n716 & ~n5113 ;
  assign n5272 = n5271 ^ n710 ^ 1'b0 ;
  assign n5273 = n2177 ^ n627 ^ 1'b0 ;
  assign n5274 = ~n494 & n5273 ;
  assign n5275 = n2923 ^ n1140 ^ 1'b0 ;
  assign n5276 = ~n726 & n5275 ;
  assign n5277 = n5276 ^ n2845 ^ 1'b0 ;
  assign n5278 = n2726 & ~n5277 ;
  assign n5279 = n5274 & ~n5278 ;
  assign n5280 = ~n3522 & n4275 ;
  assign n5281 = n4257 & n5280 ;
  assign n5282 = n2662 ^ n510 ^ 1'b0 ;
  assign n5283 = n1477 & ~n5282 ;
  assign n5284 = n2750 ^ n1130 ^ n608 ;
  assign n5285 = n4158 & n5284 ;
  assign n5286 = ( n1651 & n3311 ) | ( n1651 & ~n3416 ) | ( n3311 & ~n3416 ) ;
  assign n5287 = n4113 ^ n1887 ^ 1'b0 ;
  assign n5288 = n3477 & ~n3926 ;
  assign n5289 = n5288 ^ n827 ^ 1'b0 ;
  assign n5290 = n1980 ^ n1692 ^ 1'b0 ;
  assign n5291 = n2912 & n5290 ;
  assign n5292 = n4779 | n5291 ;
  assign n5293 = n5289 | n5292 ;
  assign n5294 = n3189 ^ n1159 ^ 1'b0 ;
  assign n5296 = n1617 ^ x48 ^ 1'b0 ;
  assign n5297 = ~n847 & n5296 ;
  assign n5298 = n2836 & n5297 ;
  assign n5299 = n5298 ^ n4826 ^ 1'b0 ;
  assign n5295 = n3576 ^ n1794 ^ 1'b0 ;
  assign n5300 = n5299 ^ n5295 ^ n951 ;
  assign n5301 = n419 ^ n269 ^ 1'b0 ;
  assign n5302 = n264 | n5301 ;
  assign n5303 = n5302 ^ n4795 ^ 1'b0 ;
  assign n5304 = n979 | n2949 ;
  assign n5305 = n1373 & ~n5304 ;
  assign n5306 = n1537 & n2177 ;
  assign n5307 = ~n1667 & n3935 ;
  assign n5308 = ~n5306 & n5307 ;
  assign n5310 = n2322 ^ n1642 ^ n1375 ;
  assign n5311 = n2641 ^ n142 ^ 1'b0 ;
  assign n5312 = n5310 | n5311 ;
  assign n5309 = n2478 | n3504 ;
  assign n5313 = n5312 ^ n5309 ^ 1'b0 ;
  assign n5314 = n3074 ^ n1096 ^ 1'b0 ;
  assign n5315 = n207 & ~n3701 ;
  assign n5316 = ~n1177 & n2809 ;
  assign n5317 = x38 & n859 ;
  assign n5318 = ( n155 & n2276 ) | ( n155 & n4416 ) | ( n2276 & n4416 ) ;
  assign n5319 = n5317 & n5318 ;
  assign n5320 = n3406 & n5319 ;
  assign n5321 = n3329 | n3353 ;
  assign n5322 = x104 | n5321 ;
  assign n5323 = n5322 ^ n2843 ^ 1'b0 ;
  assign n5324 = n809 & ~n4223 ;
  assign n5325 = ~n1435 & n5324 ;
  assign n5326 = n2624 | n5325 ;
  assign n5327 = n5326 ^ n5119 ^ 1'b0 ;
  assign n5328 = n2915 ^ n1678 ^ 1'b0 ;
  assign n5329 = n3186 ^ n768 ^ 1'b0 ;
  assign n5330 = n4905 & n5051 ;
  assign n5331 = n5330 ^ n330 ^ 1'b0 ;
  assign n5332 = n2809 ^ n242 ^ 1'b0 ;
  assign n5333 = n3697 ^ n3423 ^ n3343 ;
  assign n5334 = n260 | n452 ;
  assign n5335 = n1595 | n5334 ;
  assign n5336 = n3121 ^ n300 ^ 1'b0 ;
  assign n5337 = n5335 & ~n5336 ;
  assign n5338 = n2874 ^ n1051 ^ 1'b0 ;
  assign n5339 = n5338 ^ x13 ^ 1'b0 ;
  assign n5340 = n5337 & n5339 ;
  assign n5341 = ( n945 & n1335 ) | ( n945 & ~n2622 ) | ( n1335 & ~n2622 ) ;
  assign n5342 = n4824 ^ n4281 ^ 1'b0 ;
  assign n5343 = n484 | n5342 ;
  assign n5344 = n5343 ^ n741 ^ 1'b0 ;
  assign n5345 = n3790 | n5344 ;
  assign n5346 = n5341 | n5345 ;
  assign n5347 = n5340 | n5346 ;
  assign n5351 = n2641 ^ n1285 ^ 1'b0 ;
  assign n5348 = n1719 ^ n165 ^ 1'b0 ;
  assign n5349 = ( n420 & n4027 ) | ( n420 & n5348 ) | ( n4027 & n5348 ) ;
  assign n5350 = n3484 & n5349 ;
  assign n5352 = n5351 ^ n5350 ^ 1'b0 ;
  assign n5353 = ~n1106 & n5352 ;
  assign n5354 = ~n2206 & n5353 ;
  assign n5355 = n3624 ^ n1010 ^ x68 ;
  assign n5356 = n1651 & ~n5355 ;
  assign n5357 = ( x109 & n2906 ) | ( x109 & n5356 ) | ( n2906 & n5356 ) ;
  assign n5358 = n5357 ^ n865 ^ 1'b0 ;
  assign n5359 = n2650 & ~n4000 ;
  assign n5360 = ~n5358 & n5359 ;
  assign n5363 = n2932 ^ n654 ^ 1'b0 ;
  assign n5361 = x127 & n2976 ;
  assign n5362 = n438 | n5361 ;
  assign n5364 = n5363 ^ n5362 ^ 1'b0 ;
  assign n5365 = n948 | n5364 ;
  assign n5366 = n3554 & ~n5365 ;
  assign n5367 = n716 & ~n1190 ;
  assign n5368 = x13 & ~n2785 ;
  assign n5369 = ~n5367 & n5368 ;
  assign n5370 = n4578 & n5369 ;
  assign n5371 = n1910 ^ n1336 ^ 1'b0 ;
  assign n5372 = x98 & n5371 ;
  assign n5373 = n1266 & ~n2014 ;
  assign n5374 = n5373 ^ n3684 ^ 1'b0 ;
  assign n5375 = n422 & ~n925 ;
  assign n5376 = ~n5374 & n5375 ;
  assign n5377 = n5376 ^ n4424 ^ 1'b0 ;
  assign n5378 = n1897 | n5377 ;
  assign n5379 = n1995 ^ n748 ^ x89 ;
  assign n5380 = ( n1214 & n1448 ) | ( n1214 & ~n5379 ) | ( n1448 & ~n5379 ) ;
  assign n5381 = n2004 & n5380 ;
  assign n5382 = n3363 & n5381 ;
  assign n5383 = n5382 ^ n1366 ^ 1'b0 ;
  assign n5384 = n541 & n5383 ;
  assign n5385 = ( n247 & ~n252 ) | ( n247 & n494 ) | ( ~n252 & n494 ) ;
  assign n5386 = n1177 & ~n5385 ;
  assign n5387 = n361 & n5386 ;
  assign n5388 = n284 | n1819 ;
  assign n5389 = n5388 ^ n606 ^ 1'b0 ;
  assign n5390 = ( n1034 & n1394 ) | ( n1034 & n2619 ) | ( n1394 & n2619 ) ;
  assign n5391 = n5390 ^ n1805 ^ 1'b0 ;
  assign n5392 = ~n5214 & n5391 ;
  assign n5393 = ( ~n4175 & n5389 ) | ( ~n4175 & n5392 ) | ( n5389 & n5392 ) ;
  assign n5394 = n1556 & n1949 ;
  assign n5395 = n3159 & ~n3298 ;
  assign n5396 = ( ~n965 & n1354 ) | ( ~n965 & n1460 ) | ( n1354 & n1460 ) ;
  assign n5397 = ( ~n133 & n335 ) | ( ~n133 & n5396 ) | ( n335 & n5396 ) ;
  assign n5398 = ~n2974 & n5397 ;
  assign n5399 = ~n5395 & n5398 ;
  assign n5400 = n2278 ^ n298 ^ 1'b0 ;
  assign n5401 = n5400 ^ n3108 ^ 1'b0 ;
  assign n5402 = n5401 ^ n1800 ^ 1'b0 ;
  assign n5403 = n2613 | n5402 ;
  assign n5404 = n2750 & n5170 ;
  assign n5405 = n3689 & ~n5139 ;
  assign n5406 = n5405 ^ n5013 ^ 1'b0 ;
  assign n5410 = n1098 ^ n571 ^ n463 ;
  assign n5411 = n5032 | n5410 ;
  assign n5412 = n5411 ^ n4215 ^ 1'b0 ;
  assign n5407 = n2423 ^ n1251 ^ 1'b0 ;
  assign n5408 = n2334 ^ n1607 ^ 1'b0 ;
  assign n5409 = ~n5407 & n5408 ;
  assign n5413 = n5412 ^ n5409 ^ n5066 ;
  assign n5414 = n5413 ^ n256 ^ 1'b0 ;
  assign n5416 = n551 | n723 ;
  assign n5417 = n5416 ^ n4737 ^ n4527 ;
  assign n5415 = n848 & ~n980 ;
  assign n5418 = n5417 ^ n5415 ^ 1'b0 ;
  assign n5419 = n5418 ^ n4443 ^ n664 ;
  assign n5420 = n1770 & ~n2801 ;
  assign n5421 = ~n5017 & n5420 ;
  assign n5422 = ( n2884 & ~n5366 ) | ( n2884 & n5421 ) | ( ~n5366 & n5421 ) ;
  assign n5423 = ( ~n1156 & n2195 ) | ( ~n1156 & n4003 ) | ( n2195 & n4003 ) ;
  assign n5425 = ( n2253 & n2293 ) | ( n2253 & ~n3900 ) | ( n2293 & ~n3900 ) ;
  assign n5424 = ~n2763 & n4567 ;
  assign n5426 = n5425 ^ n5424 ^ 1'b0 ;
  assign n5427 = n3312 ^ n3111 ^ 1'b0 ;
  assign n5428 = n3149 & n5427 ;
  assign n5429 = n1108 | n4312 ;
  assign n5430 = n5428 | n5429 ;
  assign n5431 = ( n1166 & n4012 ) | ( n1166 & n5430 ) | ( n4012 & n5430 ) ;
  assign n5432 = ( n2286 & ~n3009 ) | ( n2286 & n3505 ) | ( ~n3009 & n3505 ) ;
  assign n5433 = n5432 ^ n4109 ^ 1'b0 ;
  assign n5434 = n4001 | n5433 ;
  assign n5435 = n5431 & ~n5434 ;
  assign n5436 = n5435 ^ n5317 ^ 1'b0 ;
  assign n5437 = n2752 ^ n1728 ^ 1'b0 ;
  assign n5438 = n1481 | n5437 ;
  assign n5439 = n5438 ^ n4802 ^ 1'b0 ;
  assign n5440 = n4857 ^ n4095 ^ n1894 ;
  assign n5441 = n4398 & ~n5440 ;
  assign n5442 = ~n4055 & n5441 ;
  assign n5443 = n4748 | n4997 ;
  assign n5444 = x80 & ~n771 ;
  assign n5445 = n5444 ^ n2723 ^ 1'b0 ;
  assign n5446 = n3637 & n5445 ;
  assign n5447 = ~n531 & n5446 ;
  assign n5448 = ( n456 & ~n5001 ) | ( n456 & n5447 ) | ( ~n5001 & n5447 ) ;
  assign n5449 = ( n323 & n379 ) | ( n323 & ~n2264 ) | ( n379 & ~n2264 ) ;
  assign n5450 = n2870 ^ n1607 ^ 1'b0 ;
  assign n5451 = ~n5449 & n5450 ;
  assign n5452 = n1434 | n5111 ;
  assign n5453 = n5451 | n5452 ;
  assign n5454 = n878 & ~n3898 ;
  assign n5455 = ~n223 & n5454 ;
  assign n5456 = n5455 ^ n2641 ^ 1'b0 ;
  assign n5457 = n5432 | n5456 ;
  assign n5458 = n3440 | n3722 ;
  assign n5459 = ( n967 & n1576 ) | ( n967 & ~n4840 ) | ( n1576 & ~n4840 ) ;
  assign n5461 = ( n530 & ~n787 ) | ( n530 & n3072 ) | ( ~n787 & n3072 ) ;
  assign n5460 = ( n4261 & n4697 ) | ( n4261 & n4856 ) | ( n4697 & n4856 ) ;
  assign n5462 = n5461 ^ n5460 ^ n3384 ;
  assign n5463 = n2242 ^ n1797 ^ 1'b0 ;
  assign n5464 = n1478 ^ n748 ^ 1'b0 ;
  assign n5465 = ~n2563 & n5464 ;
  assign n5466 = n1715 ^ n145 ^ 1'b0 ;
  assign n5467 = n5465 & ~n5466 ;
  assign n5468 = n5467 ^ n4665 ^ 1'b0 ;
  assign n5469 = n5463 & n5468 ;
  assign n5470 = n4969 & ~n4983 ;
  assign n5471 = ~n5469 & n5470 ;
  assign n5472 = n1355 & ~n1692 ;
  assign n5473 = n995 & n5472 ;
  assign n5474 = n3887 ^ n3278 ^ 1'b0 ;
  assign n5475 = n5473 | n5474 ;
  assign n5476 = n2964 ^ n1764 ^ 1'b0 ;
  assign n5477 = n3009 & n5476 ;
  assign n5478 = ( ~n1795 & n3957 ) | ( ~n1795 & n5477 ) | ( n3957 & n5477 ) ;
  assign n5479 = n740 ^ n290 ^ 1'b0 ;
  assign n5480 = ~n1351 & n3335 ;
  assign n5481 = n1214 | n5480 ;
  assign n5482 = n5479 & ~n5481 ;
  assign n5485 = n663 ^ x40 ^ 1'b0 ;
  assign n5486 = n716 & n5485 ;
  assign n5483 = n1389 & n1691 ;
  assign n5484 = n5483 ^ n1874 ^ n1290 ;
  assign n5487 = n5486 ^ n5484 ^ 1'b0 ;
  assign n5488 = ~n2109 & n4013 ;
  assign n5490 = ( ~n139 & n790 ) | ( ~n139 & n1972 ) | ( n790 & n1972 ) ;
  assign n5491 = n5490 ^ n1291 ^ 1'b0 ;
  assign n5492 = n739 & n5491 ;
  assign n5489 = n526 & n3022 ;
  assign n5493 = n5492 ^ n5489 ^ 1'b0 ;
  assign n5494 = n2082 ^ n1874 ^ n330 ;
  assign n5495 = ( n152 & ~n692 ) | ( n152 & n784 ) | ( ~n692 & n784 ) ;
  assign n5496 = n1512 ^ n1368 ^ 1'b0 ;
  assign n5497 = n1678 & n5496 ;
  assign n5498 = ~n5495 & n5497 ;
  assign n5499 = n5498 ^ n1463 ^ 1'b0 ;
  assign n5500 = ( ~n260 & n2739 ) | ( ~n260 & n5499 ) | ( n2739 & n5499 ) ;
  assign n5501 = ( n4868 & n5494 ) | ( n4868 & n5500 ) | ( n5494 & n5500 ) ;
  assign n5502 = ( n1152 & n1455 ) | ( n1152 & ~n2363 ) | ( n1455 & ~n2363 ) ;
  assign n5503 = n5494 & ~n5502 ;
  assign n5504 = n5503 ^ n5276 ^ 1'b0 ;
  assign n5505 = n2653 & ~n3410 ;
  assign n5506 = n4795 & n5505 ;
  assign n5507 = n3965 ^ n2377 ^ 1'b0 ;
  assign n5508 = n1840 | n5507 ;
  assign n5509 = ~n751 & n5221 ;
  assign n5510 = n5509 ^ x66 ^ 1'b0 ;
  assign n5511 = n2377 & ~n5510 ;
  assign n5512 = n5511 ^ n247 ^ 1'b0 ;
  assign n5513 = ( n3989 & ~n5508 ) | ( n3989 & n5512 ) | ( ~n5508 & n5512 ) ;
  assign n5514 = n4292 | n5119 ;
  assign n5515 = n4393 ^ n2737 ^ 1'b0 ;
  assign n5516 = n3043 & n3241 ;
  assign n5517 = n5516 ^ n1924 ^ 1'b0 ;
  assign n5518 = ~n3150 & n5517 ;
  assign n5519 = n5515 & n5518 ;
  assign n5520 = n3261 ^ n1709 ^ n1292 ;
  assign n5521 = n644 & n2576 ;
  assign n5522 = n3587 & n5521 ;
  assign n5523 = n1135 ^ n891 ^ 1'b0 ;
  assign n5525 = ( n2021 & n4900 ) | ( n2021 & ~n5497 ) | ( n4900 & ~n5497 ) ;
  assign n5526 = ~n1008 & n5525 ;
  assign n5524 = n4403 & ~n5106 ;
  assign n5527 = n5526 ^ n5524 ^ 1'b0 ;
  assign n5528 = ( n1999 & ~n5523 ) | ( n1999 & n5527 ) | ( ~n5523 & n5527 ) ;
  assign n5529 = n3905 & ~n5528 ;
  assign n5530 = n5529 ^ n5160 ^ 1'b0 ;
  assign n5531 = n1475 ^ x4 ^ 1'b0 ;
  assign n5532 = n5531 ^ n3792 ^ n2055 ;
  assign n5533 = ( n644 & n1690 ) | ( n644 & ~n4211 ) | ( n1690 & ~n4211 ) ;
  assign n5534 = n2985 ^ n2498 ^ 1'b0 ;
  assign n5535 = n932 | n5534 ;
  assign n5536 = n5535 ^ n5137 ^ n2058 ;
  assign n5537 = n2021 ^ n1164 ^ 1'b0 ;
  assign n5538 = n5537 ^ n312 ^ 1'b0 ;
  assign n5539 = n303 | n3565 ;
  assign n5540 = n5183 ^ n3586 ^ n3553 ;
  assign n5541 = x70 & n5502 ;
  assign n5542 = n5473 & n5541 ;
  assign n5543 = n5123 & n5542 ;
  assign n5544 = ~n2450 & n4959 ;
  assign n5545 = n2278 ^ n890 ^ x72 ;
  assign n5546 = n3102 ^ n2401 ^ n714 ;
  assign n5547 = n1250 | n5438 ;
  assign n5548 = n5547 ^ n1304 ^ 1'b0 ;
  assign n5549 = n5546 & n5548 ;
  assign n5550 = ~n5545 & n5549 ;
  assign n5551 = n4887 ^ n4384 ^ n2034 ;
  assign n5552 = ~n5111 & n5551 ;
  assign n5553 = n4307 & n4960 ;
  assign n5554 = n2906 & n5553 ;
  assign n5555 = ~n2987 & n3254 ;
  assign n5556 = n1501 & n5555 ;
  assign n5557 = n5554 & n5556 ;
  assign n5558 = n1949 & n2078 ;
  assign n5559 = n3368 ^ n1173 ^ n406 ;
  assign n5560 = n4374 ^ n1955 ^ 1'b0 ;
  assign n5561 = ~n5559 & n5560 ;
  assign n5565 = n4779 ^ n744 ^ 1'b0 ;
  assign n5562 = n965 & n1318 ;
  assign n5563 = ~n5242 & n5562 ;
  assign n5564 = n933 & ~n5563 ;
  assign n5566 = n5565 ^ n5564 ^ 1'b0 ;
  assign n5567 = n4115 ^ n1986 ^ n1610 ;
  assign n5568 = n2546 ^ n749 ^ n646 ;
  assign n5569 = n5568 ^ n172 ^ n140 ;
  assign n5570 = ( n3102 & n5567 ) | ( n3102 & ~n5569 ) | ( n5567 & ~n5569 ) ;
  assign n5572 = n2769 ^ n1933 ^ n1327 ;
  assign n5571 = n1649 ^ n876 ^ 1'b0 ;
  assign n5573 = n5572 ^ n5571 ^ n4492 ;
  assign n5574 = ( n3600 & ~n3658 ) | ( n3600 & n5573 ) | ( ~n3658 & n5573 ) ;
  assign n5575 = ( n904 & ~n4362 ) | ( n904 & n5111 ) | ( ~n4362 & n5111 ) ;
  assign n5576 = ( n316 & n4326 ) | ( n316 & ~n5555 ) | ( n4326 & ~n5555 ) ;
  assign n5577 = n1498 | n2173 ;
  assign n5578 = ~n3323 & n5577 ;
  assign n5579 = n731 ^ x80 ^ 1'b0 ;
  assign n5580 = n5312 | n5579 ;
  assign n5581 = ( n2157 & ~n2586 ) | ( n2157 & n3001 ) | ( ~n2586 & n3001 ) ;
  assign n5582 = ~n1234 & n5581 ;
  assign n5583 = n1890 ^ n1860 ^ 1'b0 ;
  assign n5584 = x26 & n5583 ;
  assign n5585 = n5584 ^ x115 ^ 1'b0 ;
  assign n5586 = n4813 ^ n730 ^ 1'b0 ;
  assign n5587 = n3814 | n5075 ;
  assign n5588 = n2730 | n2868 ;
  assign n5589 = n5259 ^ n4760 ^ 1'b0 ;
  assign n5590 = n2217 | n2877 ;
  assign n5591 = n3663 & ~n5590 ;
  assign n5592 = n2520 ^ n1023 ^ 1'b0 ;
  assign n5593 = ~n285 & n5592 ;
  assign n5594 = ~n2530 & n4269 ;
  assign n5595 = ~x36 & n5594 ;
  assign n5596 = n5595 ^ n5380 ^ 1'b0 ;
  assign n5597 = ( n3911 & ~n5593 ) | ( n3911 & n5596 ) | ( ~n5593 & n5596 ) ;
  assign n5598 = n3928 ^ n608 ^ x41 ;
  assign n5599 = n2504 | n4014 ;
  assign n5600 = n504 | n1046 ;
  assign n5601 = n815 | n5600 ;
  assign n5604 = x98 | n3376 ;
  assign n5605 = n458 & ~n5604 ;
  assign n5606 = n4203 ^ n1754 ^ 1'b0 ;
  assign n5607 = ~n1154 & n5606 ;
  assign n5608 = ~n2459 & n5607 ;
  assign n5609 = n5605 & n5608 ;
  assign n5602 = n2481 ^ n1581 ^ n197 ;
  assign n5603 = ( n804 & n1997 ) | ( n804 & n5602 ) | ( n1997 & n5602 ) ;
  assign n5610 = n5609 ^ n5603 ^ n1203 ;
  assign n5611 = ( n5317 & n5601 ) | ( n5317 & ~n5610 ) | ( n5601 & ~n5610 ) ;
  assign n5612 = n3989 ^ n471 ^ 1'b0 ;
  assign n5613 = n3978 ^ n1216 ^ n216 ;
  assign n5614 = n5613 ^ n384 ^ n378 ;
  assign n5615 = n5614 ^ n2635 ^ x90 ;
  assign n5616 = n3023 & ~n4712 ;
  assign n5617 = n3063 ^ n2873 ^ n357 ;
  assign n5618 = n5616 & ~n5617 ;
  assign n5619 = ~x77 & n5618 ;
  assign n5620 = n2056 ^ n1806 ^ 1'b0 ;
  assign n5621 = n2934 ^ n332 ^ 1'b0 ;
  assign n5622 = n1153 | n5473 ;
  assign n5623 = n5622 ^ x2 ^ 1'b0 ;
  assign n5624 = n3117 & ~n5244 ;
  assign n5625 = n5624 ^ n3584 ^ 1'b0 ;
  assign n5626 = n5625 ^ n3329 ^ 1'b0 ;
  assign n5627 = n5623 & n5626 ;
  assign n5628 = n3794 ^ n2355 ^ n1550 ;
  assign n5629 = ~n509 & n5628 ;
  assign n5630 = ~n1836 & n5629 ;
  assign n5631 = n3723 | n5630 ;
  assign n5632 = n5360 & n5460 ;
  assign n5633 = ~n308 & n2813 ;
  assign n5634 = n5633 ^ n356 ^ 1'b0 ;
  assign n5635 = n2371 ^ n1049 ^ 1'b0 ;
  assign n5636 = n5635 ^ n3805 ^ 1'b0 ;
  assign n5637 = ~n5634 & n5636 ;
  assign n5638 = x87 & n1518 ;
  assign n5639 = ~n553 & n5638 ;
  assign n5640 = n3862 & ~n5639 ;
  assign n5641 = ( n3824 & n5114 ) | ( n3824 & ~n5640 ) | ( n5114 & ~n5640 ) ;
  assign n5642 = n1112 & n3190 ;
  assign n5648 = n3271 ^ n3037 ^ n1196 ;
  assign n5643 = n542 ^ n389 ^ 1'b0 ;
  assign n5644 = n2785 | n5643 ;
  assign n5645 = n5644 ^ n2371 ^ 1'b0 ;
  assign n5646 = ~n1107 & n5645 ;
  assign n5647 = ~n4867 & n5646 ;
  assign n5649 = n5648 ^ n5647 ^ 1'b0 ;
  assign n5650 = n2178 ^ n2120 ^ 1'b0 ;
  assign n5651 = n2025 | n2475 ;
  assign n5652 = n5651 ^ n378 ^ 1'b0 ;
  assign n5653 = n4549 ^ n2506 ^ n1205 ;
  assign n5654 = n5653 ^ n4855 ^ n2951 ;
  assign n5655 = n4523 ^ n1752 ^ 1'b0 ;
  assign n5656 = n2246 | n3576 ;
  assign n5657 = n1577 & ~n5656 ;
  assign n5658 = n1461 | n5657 ;
  assign n5659 = ~n3117 & n5658 ;
  assign n5660 = n4710 ^ n2972 ^ 1'b0 ;
  assign n5661 = n243 | n5399 ;
  assign n5662 = n2100 ^ x11 ^ 1'b0 ;
  assign n5663 = n1207 & n1515 ;
  assign n5664 = ( ~n846 & n2435 ) | ( ~n846 & n2708 ) | ( n2435 & n2708 ) ;
  assign n5665 = n4031 | n5664 ;
  assign n5666 = n5665 ^ n3430 ^ 1'b0 ;
  assign n5672 = n3425 ^ n1374 ^ 1'b0 ;
  assign n5673 = n813 & n5672 ;
  assign n5674 = n1444 & ~n1577 ;
  assign n5675 = ~n5673 & n5674 ;
  assign n5669 = ~n1123 & n2156 ;
  assign n5670 = n5669 ^ n2690 ^ 1'b0 ;
  assign n5671 = n2068 & n5670 ;
  assign n5676 = n5675 ^ n5671 ^ 1'b0 ;
  assign n5667 = n4975 ^ n4111 ^ n2731 ;
  assign n5668 = ~n2962 & n5667 ;
  assign n5677 = n5676 ^ n5668 ^ 1'b0 ;
  assign n5678 = n684 ^ n634 ^ 1'b0 ;
  assign n5679 = n1978 ^ n1539 ^ 1'b0 ;
  assign n5680 = n251 & n5679 ;
  assign n5681 = n5680 ^ n1089 ^ 1'b0 ;
  assign n5682 = n4996 | n5681 ;
  assign n5683 = n5678 & ~n5682 ;
  assign n5684 = n1379 & n4216 ;
  assign n5685 = ~n2763 & n5219 ;
  assign n5686 = n2792 ^ n2009 ^ 1'b0 ;
  assign n5687 = n5686 ^ n2034 ^ 1'b0 ;
  assign n5688 = n3335 & ~n5687 ;
  assign n5689 = ~n3597 & n5688 ;
  assign n5690 = ( n1317 & n3476 ) | ( n1317 & ~n5601 ) | ( n3476 & ~n5601 ) ;
  assign n5691 = n810 | n4835 ;
  assign n5692 = n1282 ^ n761 ^ 1'b0 ;
  assign n5693 = ~n227 & n4681 ;
  assign n5694 = ~x111 & n5693 ;
  assign n5696 = ( n1523 & ~n3429 ) | ( n1523 & n3751 ) | ( ~n3429 & n3751 ) ;
  assign n5697 = ( x115 & ~n3418 ) | ( x115 & n5696 ) | ( ~n3418 & n5696 ) ;
  assign n5695 = ~n3174 & n4332 ;
  assign n5698 = n5697 ^ n5695 ^ n2347 ;
  assign n5699 = n5698 ^ n5694 ^ 1'b0 ;
  assign n5700 = ~n3514 & n5699 ;
  assign n5701 = ( x97 & n418 ) | ( x97 & ~n4664 ) | ( n418 & ~n4664 ) ;
  assign n5702 = n5701 ^ n1327 ^ 1'b0 ;
  assign n5703 = n2113 ^ n1205 ^ 1'b0 ;
  assign n5704 = n1473 & n5703 ;
  assign n5705 = n1985 & n5704 ;
  assign n5706 = n5705 ^ n2824 ^ n2695 ;
  assign n5712 = n1262 & ~n2272 ;
  assign n5713 = ~n1262 & n5712 ;
  assign n5707 = ~n841 & n4293 ;
  assign n5708 = n841 & n5707 ;
  assign n5709 = n1192 & ~n1536 ;
  assign n5710 = ~n1192 & n5709 ;
  assign n5711 = n5708 | n5710 ;
  assign n5714 = n5713 ^ n5711 ^ 1'b0 ;
  assign n5715 = n4443 & n4844 ;
  assign n5716 = ( n1714 & ~n1882 ) | ( n1714 & n5715 ) | ( ~n1882 & n5715 ) ;
  assign n5717 = n1320 & ~n2565 ;
  assign n5718 = n5717 ^ n639 ^ 1'b0 ;
  assign n5719 = ~n4142 & n5718 ;
  assign n5720 = n1260 & n5719 ;
  assign n5721 = n5720 ^ n614 ^ 1'b0 ;
  assign n5724 = n2974 | n3244 ;
  assign n5725 = n1037 | n5724 ;
  assign n5722 = n2581 ^ n1049 ^ 1'b0 ;
  assign n5723 = n1645 & n5722 ;
  assign n5726 = n5725 ^ n5723 ^ 1'b0 ;
  assign n5727 = n522 & n2237 ;
  assign n5728 = n1406 & n5727 ;
  assign n5732 = n2306 ^ n292 ^ 1'b0 ;
  assign n5733 = ~n1392 & n5732 ;
  assign n5734 = ~n2654 & n5733 ;
  assign n5729 = n523 & ~n2568 ;
  assign n5730 = ~n2532 & n5729 ;
  assign n5731 = n5730 ^ n4856 ^ n1473 ;
  assign n5735 = n5734 ^ n5731 ^ n1860 ;
  assign n5736 = n3121 ^ n2824 ^ n2504 ;
  assign n5737 = ~n5563 & n5736 ;
  assign n5738 = n1633 & ~n5128 ;
  assign n5739 = ~n154 & n1904 ;
  assign n5740 = x6 & ~n5739 ;
  assign n5741 = n5740 ^ n2181 ^ 1'b0 ;
  assign n5742 = n1636 & ~n2183 ;
  assign n5743 = ~n223 & n5284 ;
  assign n5744 = n4561 ^ n2770 ^ 1'b0 ;
  assign n5745 = n5743 & n5744 ;
  assign n5746 = n763 & n3117 ;
  assign n5747 = n1322 & n3965 ;
  assign n5748 = n2054 & n2709 ;
  assign n5749 = n1254 & ~n5748 ;
  assign n5750 = n2272 & n5749 ;
  assign n5751 = n4313 ^ n3111 ^ 1'b0 ;
  assign n5752 = n5147 & n5751 ;
  assign n5753 = n5752 ^ n2323 ^ n625 ;
  assign n5754 = n548 & n1177 ;
  assign n5755 = ~n4028 & n5754 ;
  assign n5756 = n5755 ^ n4230 ^ n925 ;
  assign n5757 = n3657 ^ n2715 ^ 1'b0 ;
  assign n5758 = ~n5687 & n5757 ;
  assign n5760 = n3524 ^ n1983 ^ 1'b0 ;
  assign n5761 = ~n3455 & n5760 ;
  assign n5762 = ~n1984 & n5761 ;
  assign n5759 = n374 & n1709 ;
  assign n5763 = n5762 ^ n5759 ^ 1'b0 ;
  assign n5764 = n2056 | n5763 ;
  assign n5765 = n5764 ^ n5761 ^ 1'b0 ;
  assign n5766 = n1488 & ~n5510 ;
  assign n5767 = ~n1493 & n5766 ;
  assign n5768 = n1327 & ~n5767 ;
  assign n5769 = n5515 & n5768 ;
  assign n5771 = n3894 ^ n1738 ^ n1680 ;
  assign n5770 = n4221 ^ n4109 ^ n2222 ;
  assign n5772 = n5771 ^ n5770 ^ n5354 ;
  assign n5773 = x75 & ~n2986 ;
  assign n5774 = ( n3180 & n3224 ) | ( n3180 & n5773 ) | ( n3224 & n5773 ) ;
  assign n5775 = ~n238 & n5774 ;
  assign n5776 = n5594 ^ n416 ^ 1'b0 ;
  assign n5777 = n4357 ^ n4066 ^ n4061 ;
  assign n5778 = n2641 ^ n1017 ^ 1'b0 ;
  assign n5779 = x115 & n5778 ;
  assign n5780 = n5779 ^ n3695 ^ 1'b0 ;
  assign n5781 = n5780 ^ n3574 ^ n2519 ;
  assign n5782 = n2034 ^ n201 ^ 1'b0 ;
  assign n5783 = ( n1952 & n2939 ) | ( n1952 & ~n5782 ) | ( n2939 & ~n5782 ) ;
  assign n5784 = n1153 & ~n3965 ;
  assign n5785 = n5783 & n5784 ;
  assign n5786 = x37 | n1320 ;
  assign n5787 = x44 & n1515 ;
  assign n5788 = n5786 & n5787 ;
  assign n5789 = n5788 ^ n1089 ^ 1'b0 ;
  assign n5790 = ~n3320 & n5789 ;
  assign n5791 = ~n3391 & n5790 ;
  assign n5792 = ( n1903 & n2798 ) | ( n1903 & ~n5586 ) | ( n2798 & ~n5586 ) ;
  assign n5793 = n1236 & n4983 ;
  assign n5794 = ( n1101 & ~n5792 ) | ( n1101 & n5793 ) | ( ~n5792 & n5793 ) ;
  assign n5795 = x47 & n1033 ;
  assign n5796 = n131 & n5795 ;
  assign n5797 = n1156 & n2019 ;
  assign n5798 = n5796 & n5797 ;
  assign n5799 = n5798 ^ n681 ^ 1'b0 ;
  assign n5800 = ~x49 & n5799 ;
  assign n5801 = n2559 & ~n4853 ;
  assign n5802 = n935 ^ n381 ^ 1'b0 ;
  assign n5803 = n1084 & n5802 ;
  assign n5804 = n5803 ^ n1779 ^ 1'b0 ;
  assign n5805 = n2712 ^ n480 ^ 1'b0 ;
  assign n5806 = n3015 & ~n5805 ;
  assign n5807 = n5806 ^ n4505 ^ n1460 ;
  assign n5808 = ( n589 & n5785 ) | ( n589 & n5807 ) | ( n5785 & n5807 ) ;
  assign n5809 = n2297 & ~n4746 ;
  assign n5810 = ( n1165 & ~n2344 ) | ( n1165 & n2460 ) | ( ~n2344 & n2460 ) ;
  assign n5811 = ( n1141 & ~n2668 ) | ( n1141 & n3499 ) | ( ~n2668 & n3499 ) ;
  assign n5812 = n5811 ^ n5252 ^ 1'b0 ;
  assign n5813 = n4991 & ~n5812 ;
  assign n5814 = n1062 ^ n501 ^ 1'b0 ;
  assign n5815 = n1230 & n5814 ;
  assign n5816 = n1503 ^ n715 ^ 1'b0 ;
  assign n5817 = n3017 & ~n5816 ;
  assign n5818 = n5817 ^ n3027 ^ 1'b0 ;
  assign n5819 = ~n1186 & n3816 ;
  assign n5820 = n1881 | n3886 ;
  assign n5821 = n4445 | n5820 ;
  assign n5822 = n2540 ^ n1610 ^ n160 ;
  assign n5823 = n3724 | n5822 ;
  assign n5824 = n3844 | n5823 ;
  assign n5825 = n5824 ^ n2242 ^ 1'b0 ;
  assign n5826 = n4179 | n5825 ;
  assign n5827 = ( n1209 & ~n3757 ) | ( n1209 & n5176 ) | ( ~n3757 & n5176 ) ;
  assign n5828 = n891 | n1470 ;
  assign n5829 = ~n579 & n5828 ;
  assign n5831 = n5317 ^ n1900 ^ n250 ;
  assign n5830 = ~n1160 & n2437 ;
  assign n5832 = n5831 ^ n5830 ^ 1'b0 ;
  assign n5833 = n5832 ^ n5132 ^ 1'b0 ;
  assign n5834 = ~n3559 & n5833 ;
  assign n5835 = n2238 ^ x27 ^ 1'b0 ;
  assign n5836 = n5742 & n5835 ;
  assign n5837 = n2361 ^ n2061 ^ n1129 ;
  assign n5838 = n2206 | n3650 ;
  assign n5839 = n3172 & ~n5582 ;
  assign n5840 = ( n281 & n1424 ) | ( n281 & ~n3134 ) | ( n1424 & ~n3134 ) ;
  assign n5841 = ( n157 & n2884 ) | ( n157 & n5840 ) | ( n2884 & n5840 ) ;
  assign n5842 = n5841 ^ n607 ^ 1'b0 ;
  assign n5843 = n1648 & n5842 ;
  assign n5844 = n4578 & n5843 ;
  assign n5854 = n600 & n2018 ;
  assign n5855 = n5854 ^ n3037 ^ n1506 ;
  assign n5856 = n1238 | n5029 ;
  assign n5857 = n5855 & ~n5856 ;
  assign n5847 = ~n993 & n1784 ;
  assign n5848 = n1625 ^ n172 ^ 1'b0 ;
  assign n5849 = ~n480 & n5848 ;
  assign n5850 = ( x59 & ~n3181 ) | ( x59 & n5849 ) | ( ~n3181 & n5849 ) ;
  assign n5851 = n5850 ^ n3669 ^ 1'b0 ;
  assign n5852 = ( n3323 & n5847 ) | ( n3323 & ~n5851 ) | ( n5847 & ~n5851 ) ;
  assign n5853 = n2454 | n5852 ;
  assign n5845 = n3092 ^ n2844 ^ n274 ;
  assign n5846 = ( n2547 & ~n3178 ) | ( n2547 & n5845 ) | ( ~n3178 & n5845 ) ;
  assign n5858 = n5857 ^ n5853 ^ n5846 ;
  assign n5859 = n4125 ^ n3989 ^ 1'b0 ;
  assign n5860 = n1475 ^ n406 ^ 1'b0 ;
  assign n5861 = n5860 ^ n3298 ^ 1'b0 ;
  assign n5862 = n402 ^ x25 ^ 1'b0 ;
  assign n5863 = n5862 ^ n2554 ^ n245 ;
  assign n5865 = n5278 ^ n155 ^ 1'b0 ;
  assign n5864 = n5284 ^ n4834 ^ 1'b0 ;
  assign n5866 = n5865 ^ n5864 ^ 1'b0 ;
  assign n5867 = ~n5863 & n5866 ;
  assign n5868 = n1567 ^ n225 ^ 1'b0 ;
  assign n5869 = n2149 | n5868 ;
  assign n5870 = n5869 ^ n1507 ^ 1'b0 ;
  assign n5871 = n5870 ^ n5421 ^ n2496 ;
  assign n5872 = n210 & ~n2416 ;
  assign n5873 = n2772 ^ n1929 ^ 1'b0 ;
  assign n5874 = n1734 & ~n5873 ;
  assign n5875 = n1273 & n5874 ;
  assign n5876 = n5875 ^ n4382 ^ 1'b0 ;
  assign n5877 = n5770 | n5876 ;
  assign n5878 = n5877 ^ n1082 ^ 1'b0 ;
  assign n5879 = n3400 | n4078 ;
  assign n5880 = n846 & n5879 ;
  assign n5881 = n3931 ^ n276 ^ 1'b0 ;
  assign n5882 = n4113 & n4590 ;
  assign n5883 = ~x113 & n1988 ;
  assign n5884 = ( n909 & n1656 ) | ( n909 & n5883 ) | ( n1656 & n5883 ) ;
  assign n5885 = n2193 & n3375 ;
  assign n5886 = n2767 | n3388 ;
  assign n5887 = n240 & ~n5886 ;
  assign n5888 = n5887 ^ n1436 ^ n1435 ;
  assign n5889 = n820 | n2349 ;
  assign n5890 = n5889 ^ n1946 ^ 1'b0 ;
  assign n5891 = n1200 ^ n1023 ^ 1'b0 ;
  assign n5892 = n1501 & n5891 ;
  assign n5893 = ~n867 & n5892 ;
  assign n5894 = n2873 | n4742 ;
  assign n5895 = n5894 ^ n5657 ^ n2589 ;
  assign n5896 = n1433 & ~n5854 ;
  assign n5897 = n5896 ^ n5826 ^ 1'b0 ;
  assign n5898 = n3009 ^ n2332 ^ 1'b0 ;
  assign n5899 = n2282 & n5898 ;
  assign n5902 = ( x76 & n1905 ) | ( x76 & n4431 ) | ( n1905 & n4431 ) ;
  assign n5903 = n4793 & ~n5902 ;
  assign n5904 = n5903 ^ n470 ^ 1'b0 ;
  assign n5900 = n427 | n1090 ;
  assign n5901 = n5900 ^ n3587 ^ 1'b0 ;
  assign n5905 = n5904 ^ n5901 ^ 1'b0 ;
  assign n5906 = n5899 & n5905 ;
  assign n5907 = n2959 ^ n1519 ^ n270 ;
  assign n5908 = n2625 & n5907 ;
  assign n5909 = ~n5906 & n5908 ;
  assign n5910 = ( ~x106 & n3399 ) | ( ~x106 & n4169 ) | ( n3399 & n4169 ) ;
  assign n5911 = ( n3494 & n3930 ) | ( n3494 & n5910 ) | ( n3930 & n5910 ) ;
  assign n5912 = ~n4292 & n5911 ;
  assign n5913 = n572 | n1335 ;
  assign n5914 = n3971 & ~n5913 ;
  assign n5915 = x107 & n2842 ;
  assign n5916 = n1983 & n5915 ;
  assign n5917 = n3326 ^ n664 ^ 1'b0 ;
  assign n5918 = x17 & ~n5917 ;
  assign n5919 = ~n2063 & n2952 ;
  assign n5920 = n5919 ^ n3767 ^ 1'b0 ;
  assign n5921 = n4211 ^ n1165 ^ 1'b0 ;
  assign n5922 = n1820 & n2500 ;
  assign n5923 = n5922 ^ n3609 ^ 1'b0 ;
  assign n5924 = ~n5921 & n5923 ;
  assign n5925 = ~n3859 & n5924 ;
  assign n5926 = n5925 ^ n3260 ^ 1'b0 ;
  assign n5927 = ~n163 & n2884 ;
  assign n5928 = n5927 ^ n4179 ^ 1'b0 ;
  assign n5929 = n1505 | n1512 ;
  assign n5930 = n5929 ^ n747 ^ 1'b0 ;
  assign n5931 = n3130 ^ n2934 ^ 1'b0 ;
  assign n5934 = n2072 ^ n367 ^ x98 ;
  assign n5932 = n447 & n4055 ;
  assign n5933 = n5932 ^ n3009 ^ 1'b0 ;
  assign n5935 = n5934 ^ n5933 ^ 1'b0 ;
  assign n5936 = n2090 | n3214 ;
  assign n5937 = n5935 | n5936 ;
  assign n5939 = n242 ^ x66 ^ 1'b0 ;
  assign n5940 = ~n760 & n5939 ;
  assign n5941 = n5940 ^ n557 ^ 1'b0 ;
  assign n5942 = n309 & ~n5941 ;
  assign n5943 = ( n946 & ~n2596 ) | ( n946 & n5942 ) | ( ~n2596 & n5942 ) ;
  assign n5938 = n2641 ^ n1505 ^ n576 ;
  assign n5944 = n5943 ^ n5938 ^ x86 ;
  assign n5945 = n358 & ~n5542 ;
  assign n5946 = n571 & ~n2645 ;
  assign n5947 = n5945 & n5946 ;
  assign n5948 = n5392 ^ n3788 ^ 1'b0 ;
  assign n5951 = ( ~n584 & n2546 ) | ( ~n584 & n5238 ) | ( n2546 & n5238 ) ;
  assign n5952 = n5951 ^ n3364 ^ 1'b0 ;
  assign n5953 = n5952 ^ n4675 ^ n713 ;
  assign n5949 = n4375 ^ x53 ^ 1'b0 ;
  assign n5950 = n4490 | n5949 ;
  assign n5954 = n5953 ^ n5950 ^ n963 ;
  assign n5955 = n1485 & n2012 ;
  assign n5956 = ( n2792 & ~n5425 ) | ( n2792 & n5874 ) | ( ~n5425 & n5874 ) ;
  assign n5957 = n5956 ^ n3796 ^ 1'b0 ;
  assign n5958 = n5955 | n5957 ;
  assign n5959 = ( n353 & ~n1481 ) | ( n353 & n2924 ) | ( ~n1481 & n2924 ) ;
  assign n5960 = n5824 ^ n307 ^ 1'b0 ;
  assign n5961 = n5960 ^ n5244 ^ 1'b0 ;
  assign n5962 = n4878 ^ n4144 ^ n3046 ;
  assign n5963 = n3883 | n5962 ;
  assign n5964 = n5914 | n5963 ;
  assign n5965 = n5964 ^ n361 ^ 1'b0 ;
  assign n5966 = n3766 & n5499 ;
  assign n5967 = x0 & n3090 ;
  assign n5968 = n968 & n1793 ;
  assign n5969 = n5968 ^ n1738 ^ n1326 ;
  assign n5970 = n5967 & n5969 ;
  assign n5971 = n718 & ~n755 ;
  assign n5972 = n5971 ^ n1276 ^ 1'b0 ;
  assign n5973 = ( n362 & n5970 ) | ( n362 & n5972 ) | ( n5970 & n5972 ) ;
  assign n5974 = n5973 ^ n3609 ^ 1'b0 ;
  assign n5975 = n954 | n2770 ;
  assign n5980 = n1184 & ~n2930 ;
  assign n5976 = n413 & n2270 ;
  assign n5977 = ~n3218 & n5976 ;
  assign n5978 = n2528 & ~n5977 ;
  assign n5979 = ~n2471 & n5978 ;
  assign n5981 = n5980 ^ n5979 ^ 1'b0 ;
  assign n5982 = n5975 & ~n5981 ;
  assign n5983 = n1221 & n5982 ;
  assign n5984 = n5983 ^ n1284 ^ 1'b0 ;
  assign n5985 = n463 & ~n1761 ;
  assign n5986 = ~n5940 & n5985 ;
  assign n5987 = n1014 & ~n2965 ;
  assign n5988 = ( n2328 & n3771 ) | ( n2328 & ~n5987 ) | ( n3771 & ~n5987 ) ;
  assign n5989 = n2708 ^ n1433 ^ 1'b0 ;
  assign n5990 = n2040 & n5989 ;
  assign n5991 = n1216 | n3676 ;
  assign n5992 = n5990 | n5991 ;
  assign n5993 = ( n2956 & n3211 ) | ( n2956 & n4016 ) | ( n3211 & n4016 ) ;
  assign n5994 = ( n4519 & ~n5680 ) | ( n4519 & n5993 ) | ( ~n5680 & n5993 ) ;
  assign n5995 = ( n3969 & n4908 ) | ( n3969 & ~n5994 ) | ( n4908 & ~n5994 ) ;
  assign n5998 = n2813 ^ n511 ^ 1'b0 ;
  assign n5999 = ~n827 & n5998 ;
  assign n5996 = n2511 ^ n1527 ^ 1'b0 ;
  assign n5997 = n2534 & ~n5996 ;
  assign n6000 = n5999 ^ n5997 ^ 1'b0 ;
  assign n6001 = ~n2530 & n6000 ;
  assign n6008 = n4073 & ~n4538 ;
  assign n6009 = n6008 ^ n2452 ^ 1'b0 ;
  assign n6010 = ( x85 & ~n4434 ) | ( x85 & n6009 ) | ( ~n4434 & n6009 ) ;
  assign n6011 = ~n2406 & n4382 ;
  assign n6012 = ~n6010 & n6011 ;
  assign n6013 = n6012 ^ n4226 ^ 1'b0 ;
  assign n6002 = n1064 ^ n380 ^ 1'b0 ;
  assign n6003 = n5259 & n6002 ;
  assign n6004 = n5325 ^ n3463 ^ 1'b0 ;
  assign n6005 = n6004 ^ n5094 ^ n2631 ;
  assign n6006 = n6005 ^ n4070 ^ 1'b0 ;
  assign n6007 = n6003 & ~n6006 ;
  assign n6014 = n6013 ^ n6007 ^ n3618 ;
  assign n6015 = n5888 ^ n3459 ^ n2744 ;
  assign n6016 = x107 & ~n588 ;
  assign n6017 = n6016 ^ n2382 ^ 1'b0 ;
  assign n6018 = n4770 & n6017 ;
  assign n6019 = n2737 & n6018 ;
  assign n6020 = n654 | n2890 ;
  assign n6021 = n6020 ^ n2979 ^ 1'b0 ;
  assign n6022 = n1272 & n1914 ;
  assign n6023 = ( n1915 & n4172 ) | ( n1915 & ~n6022 ) | ( n4172 & ~n6022 ) ;
  assign n6024 = n4031 ^ n2538 ^ 1'b0 ;
  assign n6025 = n5018 ^ n3143 ^ 1'b0 ;
  assign n6026 = n6025 ^ n5662 ^ n1621 ;
  assign n6027 = n424 & n1460 ;
  assign n6028 = n6027 ^ n918 ^ 1'b0 ;
  assign n6029 = ( n4592 & ~n4856 ) | ( n4592 & n6028 ) | ( ~n4856 & n6028 ) ;
  assign n6030 = n6029 ^ n4126 ^ n1515 ;
  assign n6031 = n456 | n603 ;
  assign n6032 = x106 | n6031 ;
  assign n6033 = n1015 & ~n1150 ;
  assign n6034 = ~n6032 & n6033 ;
  assign n6035 = n6034 ^ n4346 ^ n2187 ;
  assign n6036 = ( n2193 & n4264 ) | ( n2193 & n4900 ) | ( n4264 & n4900 ) ;
  assign n6037 = ( n181 & ~n3090 ) | ( n181 & n6036 ) | ( ~n3090 & n6036 ) ;
  assign n6038 = n6037 ^ n2100 ^ n178 ;
  assign n6039 = n5821 ^ n1851 ^ 1'b0 ;
  assign n6040 = n4422 ^ n3245 ^ 1'b0 ;
  assign n6041 = n5425 ^ n1064 ^ n646 ;
  assign n6042 = ( n2787 & ~n4418 ) | ( n2787 & n6041 ) | ( ~n4418 & n6041 ) ;
  assign n6043 = n4805 ^ n3561 ^ n2554 ;
  assign n6044 = n6043 ^ n5794 ^ 1'b0 ;
  assign n6045 = n3307 ^ n1433 ^ 1'b0 ;
  assign n6046 = n256 & ~n6045 ;
  assign n6047 = n4748 & n6046 ;
  assign n6048 = n4359 ^ n3162 ^ n2875 ;
  assign n6049 = n3969 & ~n6048 ;
  assign n6050 = n3252 ^ n1950 ^ 1'b0 ;
  assign n6051 = n4962 ^ n3019 ^ 1'b0 ;
  assign n6052 = n992 & ~n5535 ;
  assign n6053 = ( n1493 & ~n1678 ) | ( n1493 & n3347 ) | ( ~n1678 & n3347 ) ;
  assign n6054 = n827 | n3864 ;
  assign n6055 = n6053 & ~n6054 ;
  assign n6056 = ( n1297 & n5402 ) | ( n1297 & n6055 ) | ( n5402 & n6055 ) ;
  assign n6057 = ~n169 & n1355 ;
  assign n6058 = n3379 | n6057 ;
  assign n6059 = n6058 ^ n2719 ^ 1'b0 ;
  assign n6060 = n1678 | n6059 ;
  assign n6061 = n6060 ^ n3711 ^ 1'b0 ;
  assign n6062 = n3406 | n4523 ;
  assign n6063 = n3519 & ~n6062 ;
  assign n6064 = n990 ^ x118 ^ 1'b0 ;
  assign n6065 = n3255 & n5125 ;
  assign n6066 = ~n6064 & n6065 ;
  assign n6067 = n2483 & n4876 ;
  assign n6068 = ( ~n260 & n4719 ) | ( ~n260 & n6067 ) | ( n4719 & n6067 ) ;
  assign n6069 = ~n1475 & n3824 ;
  assign n6070 = n6069 ^ n548 ^ 1'b0 ;
  assign n6071 = n5583 ^ n887 ^ 1'b0 ;
  assign n6072 = ~n1086 & n6071 ;
  assign n6073 = ( n3255 & n4746 ) | ( n3255 & ~n6072 ) | ( n4746 & ~n6072 ) ;
  assign n6076 = ( n2349 & n3698 ) | ( n2349 & n4265 ) | ( n3698 & n4265 ) ;
  assign n6074 = n811 & ~n3572 ;
  assign n6075 = n6074 ^ n3887 ^ 1'b0 ;
  assign n6077 = n6076 ^ n6075 ^ n2664 ;
  assign n6078 = n2897 & ~n6077 ;
  assign n6079 = ~n6073 & n6078 ;
  assign n6080 = n6079 ^ n3054 ^ 1'b0 ;
  assign n6081 = n6070 & ~n6080 ;
  assign n6082 = n6081 ^ n5021 ^ 1'b0 ;
  assign n6083 = n1929 & n6082 ;
  assign n6084 = n4951 ^ n2393 ^ n1876 ;
  assign n6085 = n712 | n6084 ;
  assign n6086 = n1799 ^ x30 ^ 1'b0 ;
  assign n6087 = n2508 & n6086 ;
  assign n6088 = n6087 ^ n2640 ^ n1686 ;
  assign n6089 = n6088 ^ n3043 ^ 1'b0 ;
  assign n6090 = n1268 & ~n6089 ;
  assign n6091 = n1456 | n5206 ;
  assign n6092 = n3104 | n6091 ;
  assign n6093 = ~n3471 & n6092 ;
  assign n6094 = ~n1528 & n6093 ;
  assign n6095 = n6094 ^ n4006 ^ 1'b0 ;
  assign n6096 = n423 | n6095 ;
  assign n6098 = n3016 ^ n1054 ^ n267 ;
  assign n6099 = n207 & ~n6098 ;
  assign n6100 = n6099 ^ n6058 ^ 1'b0 ;
  assign n6097 = n3989 | n5537 ;
  assign n6101 = n6100 ^ n6097 ^ 1'b0 ;
  assign n6102 = n1067 & n4308 ;
  assign n6103 = ~n1800 & n6102 ;
  assign n6104 = n6103 ^ n4617 ^ 1'b0 ;
  assign n6105 = ( n3059 & n6101 ) | ( n3059 & ~n6104 ) | ( n6101 & ~n6104 ) ;
  assign n6106 = n2817 ^ x41 ^ 1'b0 ;
  assign n6107 = n2948 ^ n1431 ^ 1'b0 ;
  assign n6108 = ~n6106 & n6107 ;
  assign n6109 = n4498 ^ x97 ^ 1'b0 ;
  assign n6110 = n6108 & ~n6109 ;
  assign n6111 = n4332 & ~n4388 ;
  assign n6120 = n1368 ^ n779 ^ 1'b0 ;
  assign n6121 = n620 & n6120 ;
  assign n6122 = n6121 ^ n2145 ^ 1'b0 ;
  assign n6123 = n3681 & ~n6122 ;
  assign n6112 = n4567 ^ n829 ^ 1'b0 ;
  assign n6115 = ( n543 & ~n1935 ) | ( n543 & n2831 ) | ( ~n1935 & n2831 ) ;
  assign n6116 = n309 & n4143 ;
  assign n6117 = ~n6115 & n6116 ;
  assign n6113 = n5151 ^ n847 ^ 1'b0 ;
  assign n6114 = n2661 & ~n6113 ;
  assign n6118 = n6117 ^ n6114 ^ n2915 ;
  assign n6119 = ~n6112 & n6118 ;
  assign n6124 = n6123 ^ n6119 ^ 1'b0 ;
  assign n6126 = ( n694 & n741 ) | ( n694 & n1990 ) | ( n741 & n1990 ) ;
  assign n6125 = n1370 & n2927 ;
  assign n6127 = n6126 ^ n6125 ^ n4667 ;
  assign n6128 = n6127 ^ n3643 ^ 1'b0 ;
  assign n6129 = n1867 ^ n187 ^ 1'b0 ;
  assign n6130 = ( n3669 & n6128 ) | ( n3669 & n6129 ) | ( n6128 & n6129 ) ;
  assign n6131 = n1104 & n5050 ;
  assign n6132 = n6131 ^ n3988 ^ 1'b0 ;
  assign n6133 = n4758 ^ n3015 ^ x102 ;
  assign n6134 = n3829 & ~n5403 ;
  assign n6135 = n234 ^ n142 ^ 1'b0 ;
  assign n6136 = n6135 ^ n2738 ^ n836 ;
  assign n6137 = n6136 ^ n4397 ^ n474 ;
  assign n6138 = n6137 ^ n1565 ^ 1'b0 ;
  assign n6139 = n5221 ^ n2589 ^ 1'b0 ;
  assign n6140 = n4184 ^ n3756 ^ n2856 ;
  assign n6141 = ~n701 & n6140 ;
  assign n6142 = ~n6139 & n6141 ;
  assign n6143 = n6121 & ~n6142 ;
  assign n6144 = n6143 ^ n843 ^ 1'b0 ;
  assign n6145 = n6138 | n6144 ;
  assign n6146 = n580 & ~n5725 ;
  assign n6147 = ( n2269 & ~n4107 ) | ( n2269 & n6146 ) | ( ~n4107 & n6146 ) ;
  assign n6148 = n563 | n3291 ;
  assign n6149 = ( n2748 & ~n3686 ) | ( n2748 & n6148 ) | ( ~n3686 & n6148 ) ;
  assign n6150 = n6149 ^ n4071 ^ n3850 ;
  assign n6151 = n962 & ~n2120 ;
  assign n6152 = n6151 ^ n4451 ^ 1'b0 ;
  assign n6153 = n1376 & ~n4387 ;
  assign n6154 = n6153 ^ n4207 ^ 1'b0 ;
  assign n6155 = n3026 & n3581 ;
  assign n6156 = n6155 ^ n4364 ^ 1'b0 ;
  assign n6157 = n6156 ^ n1850 ^ 1'b0 ;
  assign n6158 = n677 | n1054 ;
  assign n6159 = n6158 ^ x93 ^ 1'b0 ;
  assign n6160 = ( n935 & ~n6157 ) | ( n935 & n6159 ) | ( ~n6157 & n6159 ) ;
  assign n6161 = n3293 & ~n5963 ;
  assign n6162 = n2524 & ~n4758 ;
  assign n6163 = ~n1190 & n6162 ;
  assign n6164 = ~n4507 & n6163 ;
  assign n6165 = ( n168 & n3908 ) | ( n168 & ~n6164 ) | ( n3908 & ~n6164 ) ;
  assign n6166 = ~x73 & n438 ;
  assign n6167 = n6166 ^ n196 ^ 1'b0 ;
  assign n6168 = ( n1126 & n1691 ) | ( n1126 & ~n4929 ) | ( n1691 & ~n4929 ) ;
  assign n6169 = n4935 | n6168 ;
  assign n6170 = n933 & n6169 ;
  assign n6171 = ~n2111 & n2933 ;
  assign n6172 = ( n2499 & n5482 ) | ( n2499 & n6171 ) | ( n5482 & n6171 ) ;
  assign n6173 = n6158 ^ n3413 ^ 1'b0 ;
  assign n6179 = ( n1003 & n2355 ) | ( n1003 & n2988 ) | ( n2355 & n2988 ) ;
  assign n6177 = ~x37 & n5739 ;
  assign n6174 = n2893 ^ n1394 ^ n1381 ;
  assign n6175 = n6076 ^ n1454 ^ 1'b0 ;
  assign n6176 = ~n6174 & n6175 ;
  assign n6178 = n6177 ^ n6176 ^ n5852 ;
  assign n6180 = n6179 ^ n6178 ^ 1'b0 ;
  assign n6181 = n1283 ^ n696 ^ 1'b0 ;
  assign n6182 = n6181 ^ n3921 ^ 1'b0 ;
  assign n6183 = n4112 ^ n804 ^ 1'b0 ;
  assign n6184 = n2134 ^ n603 ^ 1'b0 ;
  assign n6185 = x83 & n6184 ;
  assign n6186 = n6185 ^ n1317 ^ 1'b0 ;
  assign n6187 = ~n378 & n2542 ;
  assign n6188 = n2031 & ~n6187 ;
  assign n6189 = ~n917 & n6188 ;
  assign n6190 = ( n238 & ~n2044 ) | ( n238 & n2615 ) | ( ~n2044 & n2615 ) ;
  assign n6191 = n6190 ^ n4436 ^ n579 ;
  assign n6194 = n265 & n2575 ;
  assign n6195 = n6194 ^ n1921 ^ 1'b0 ;
  assign n6196 = n1594 & ~n6195 ;
  assign n6192 = n3967 ^ n2761 ^ n1502 ;
  assign n6193 = n6192 ^ n5059 ^ 1'b0 ;
  assign n6197 = n6196 ^ n6193 ^ n1124 ;
  assign n6198 = n3169 ^ n1487 ^ 1'b0 ;
  assign n6199 = n4927 | n6198 ;
  assign n6200 = n2985 & n6199 ;
  assign n6201 = n5526 ^ n531 ^ 1'b0 ;
  assign n6202 = n6201 ^ n5446 ^ 1'b0 ;
  assign n6203 = ~n3169 & n6202 ;
  assign n6204 = x31 & n6121 ;
  assign n6205 = n6204 ^ n3915 ^ 1'b0 ;
  assign n6206 = ( n2705 & n3716 ) | ( n2705 & n6205 ) | ( n3716 & n6205 ) ;
  assign n6207 = n351 | n6206 ;
  assign n6208 = n2248 ^ n1392 ^ x15 ;
  assign n6209 = ( n949 & n2575 ) | ( n949 & n6208 ) | ( n2575 & n6208 ) ;
  assign n6210 = ~n993 & n6209 ;
  assign n6211 = ~n5860 & n6210 ;
  assign n6218 = n2886 ^ n1647 ^ 1'b0 ;
  assign n6219 = n995 | n6218 ;
  assign n6220 = n6219 ^ x59 ^ 1'b0 ;
  assign n6213 = n1856 & ~n2285 ;
  assign n6214 = n6213 ^ n1776 ^ 1'b0 ;
  assign n6215 = ~n1585 & n6214 ;
  assign n6216 = n6215 ^ n3817 ^ 1'b0 ;
  assign n6212 = n725 | n1871 ;
  assign n6217 = n6216 ^ n6212 ^ 1'b0 ;
  assign n6221 = n6220 ^ n6217 ^ n3771 ;
  assign n6222 = ( n3202 & n6211 ) | ( n3202 & ~n6221 ) | ( n6211 & ~n6221 ) ;
  assign n6227 = n2851 ^ n1332 ^ 1'b0 ;
  assign n6228 = n6227 ^ n5680 ^ 1'b0 ;
  assign n6224 = n1915 ^ n209 ^ 1'b0 ;
  assign n6225 = x100 & n6224 ;
  assign n6223 = n397 & ~n1577 ;
  assign n6226 = n6225 ^ n6223 ^ n2115 ;
  assign n6229 = n6228 ^ n6226 ^ n1227 ;
  assign n6230 = n6229 ^ n4689 ^ n1712 ;
  assign n6233 = n1481 ^ n422 ^ 1'b0 ;
  assign n6234 = n6233 ^ n850 ^ n433 ;
  assign n6231 = n3177 ^ n2454 ^ 1'b0 ;
  assign n6232 = n4543 | n6231 ;
  assign n6235 = n6234 ^ n6232 ^ n2624 ;
  assign n6236 = n2063 ^ x54 ^ 1'b0 ;
  assign n6243 = n2791 ^ n546 ^ n240 ;
  assign n6237 = ( n613 & n2315 ) | ( n613 & ~n2512 ) | ( n2315 & ~n2512 ) ;
  assign n6238 = n712 ^ n207 ^ 1'b0 ;
  assign n6239 = ~n3556 & n6238 ;
  assign n6240 = n6239 ^ n1025 ^ n482 ;
  assign n6241 = n2053 & ~n6240 ;
  assign n6242 = n6237 & n6241 ;
  assign n6244 = n6243 ^ n6242 ^ 1'b0 ;
  assign n6245 = n5899 & n6244 ;
  assign n6248 = n1760 ^ n1120 ^ 1'b0 ;
  assign n6249 = ~n995 & n6248 ;
  assign n6246 = n3408 ^ n729 ^ 1'b0 ;
  assign n6247 = n634 & n6246 ;
  assign n6250 = n6249 ^ n6247 ^ n3399 ;
  assign n6253 = ~n1667 & n2408 ;
  assign n6254 = n6253 ^ n3734 ^ 1'b0 ;
  assign n6251 = ~n1673 & n2809 ;
  assign n6252 = n6251 ^ n3314 ^ 1'b0 ;
  assign n6255 = n6254 ^ n6252 ^ n374 ;
  assign n6257 = n811 & n4331 ;
  assign n6258 = n3674 & n6257 ;
  assign n6259 = x8 & ~n1729 ;
  assign n6260 = n6258 & n6259 ;
  assign n6261 = n6260 ^ n4382 ^ 1'b0 ;
  assign n6256 = n3620 & n5770 ;
  assign n6262 = n6261 ^ n6256 ^ 1'b0 ;
  assign n6263 = n1841 | n2180 ;
  assign n6264 = n6263 ^ n327 ^ 1'b0 ;
  assign n6265 = n2586 ^ n2211 ^ n1955 ;
  assign n6266 = n5000 & n5074 ;
  assign n6267 = ~n6265 & n6266 ;
  assign n6273 = n3445 ^ x106 ^ 1'b0 ;
  assign n6274 = n3194 & n6273 ;
  assign n6270 = ~n624 & n1132 ;
  assign n6271 = n6270 ^ n1000 ^ 1'b0 ;
  assign n6268 = n1669 ^ n782 ^ n778 ;
  assign n6269 = n6268 ^ n3088 ^ x83 ;
  assign n6272 = n6271 ^ n6269 ^ 1'b0 ;
  assign n6275 = n6274 ^ n6272 ^ 1'b0 ;
  assign n6276 = n5191 ^ n1937 ^ 1'b0 ;
  assign n6277 = ~n2484 & n5151 ;
  assign n6278 = ~n522 & n6277 ;
  assign n6279 = n1470 ^ n422 ^ 1'b0 ;
  assign n6280 = ~n6278 & n6279 ;
  assign n6281 = n1440 & ~n6280 ;
  assign n6282 = ( ~n1049 & n3894 ) | ( ~n1049 & n6281 ) | ( n3894 & n6281 ) ;
  assign n6283 = n960 & n2587 ;
  assign n6284 = n1615 & ~n6283 ;
  assign n6294 = n2787 ^ n1057 ^ n189 ;
  assign n6292 = n2928 & ~n4734 ;
  assign n6293 = ~n3278 & n6292 ;
  assign n6295 = n6294 ^ n6293 ^ 1'b0 ;
  assign n6291 = n389 & n2267 ;
  assign n6296 = n6295 ^ n6291 ^ 1'b0 ;
  assign n6297 = ( n935 & ~n2068 ) | ( n935 & n6296 ) | ( ~n2068 & n6296 ) ;
  assign n6285 = ( n269 & n767 ) | ( n269 & n918 ) | ( n767 & n918 ) ;
  assign n6286 = n6285 ^ n2445 ^ 1'b0 ;
  assign n6287 = ~n2275 & n6286 ;
  assign n6288 = n6287 ^ n6127 ^ 1'b0 ;
  assign n6289 = n343 & ~n4995 ;
  assign n6290 = ( ~n5801 & n6288 ) | ( ~n5801 & n6289 ) | ( n6288 & n6289 ) ;
  assign n6298 = n6297 ^ n6290 ^ 1'b0 ;
  assign n6299 = ( n798 & n1033 ) | ( n798 & ~n2995 ) | ( n1033 & ~n2995 ) ;
  assign n6300 = n6299 ^ n5335 ^ 1'b0 ;
  assign n6301 = n4234 & n6300 ;
  assign n6302 = n3092 ^ n347 ^ 1'b0 ;
  assign n6303 = ~n817 & n6302 ;
  assign n6304 = n6303 ^ n207 ^ 1'b0 ;
  assign n6305 = n6301 & ~n6304 ;
  assign n6306 = n1649 ^ n1181 ^ 1'b0 ;
  assign n6307 = n706 & ~n1238 ;
  assign n6308 = n2905 & n6307 ;
  assign n6309 = n6308 ^ x2 ^ 1'b0 ;
  assign n6310 = n4945 ^ n995 ^ x80 ;
  assign n6311 = x103 & n2602 ;
  assign n6312 = n6311 ^ n1567 ^ 1'b0 ;
  assign n6313 = n6312 ^ n5982 ^ 1'b0 ;
  assign n6314 = n4561 ^ n528 ^ 1'b0 ;
  assign n6315 = n3238 & ~n6314 ;
  assign n6316 = ( n3020 & n4275 ) | ( n3020 & ~n6315 ) | ( n4275 & ~n6315 ) ;
  assign n6317 = n1231 ^ n1125 ^ n286 ;
  assign n6318 = ( ~n5345 & n6316 ) | ( ~n5345 & n6317 ) | ( n6316 & n6317 ) ;
  assign n6319 = n5259 ^ n929 ^ 1'b0 ;
  assign n6320 = n6319 ^ n3957 ^ n3802 ;
  assign n6321 = n2584 ^ n2074 ^ 1'b0 ;
  assign n6322 = n739 & n6321 ;
  assign n6324 = ( n1928 & ~n3365 ) | ( n1928 & n5759 ) | ( ~n3365 & n5759 ) ;
  assign n6323 = ~n138 & n3238 ;
  assign n6325 = n6324 ^ n6323 ^ 1'b0 ;
  assign n6326 = n6325 ^ n1823 ^ 1'b0 ;
  assign n6331 = n184 & n1218 ;
  assign n6332 = ~n4574 & n6331 ;
  assign n6333 = n6332 ^ n3027 ^ 1'b0 ;
  assign n6334 = n4900 ^ n4275 ^ 1'b0 ;
  assign n6335 = ~n6333 & n6334 ;
  assign n6327 = n4202 ^ n4180 ^ 1'b0 ;
  assign n6328 = n2452 | n6327 ;
  assign n6329 = n2783 | n6328 ;
  assign n6330 = ~n1264 & n6329 ;
  assign n6336 = n6335 ^ n6330 ^ 1'b0 ;
  assign n6337 = n3631 ^ n3410 ^ 1'b0 ;
  assign n6338 = n1126 | n3453 ;
  assign n6339 = n2288 & ~n6338 ;
  assign n6340 = n6339 ^ n1312 ^ 1'b0 ;
  assign n6341 = n6340 ^ n2209 ^ 1'b0 ;
  assign n6342 = n901 & n3999 ;
  assign n6343 = n4542 ^ n4273 ^ 1'b0 ;
  assign n6344 = n2148 & ~n6343 ;
  assign n6345 = n1209 & n3506 ;
  assign n6346 = n5873 ^ n2957 ^ n2647 ;
  assign n6347 = n6345 & ~n6346 ;
  assign n6348 = ( n2109 & n6344 ) | ( n2109 & n6347 ) | ( n6344 & n6347 ) ;
  assign n6349 = ( x15 & n719 ) | ( x15 & n1335 ) | ( n719 & n1335 ) ;
  assign n6350 = n2945 ^ n773 ^ 1'b0 ;
  assign n6351 = ~n6349 & n6350 ;
  assign n6352 = ~n216 & n2898 ;
  assign n6353 = ~n768 & n6352 ;
  assign n6354 = n4061 | n6353 ;
  assign n6355 = ~n6077 & n6354 ;
  assign n6356 = n4494 ^ n4173 ^ 1'b0 ;
  assign n6357 = n6356 ^ n4858 ^ 1'b0 ;
  assign n6358 = n1600 ^ n1493 ^ n489 ;
  assign n6359 = n6163 ^ n4935 ^ 1'b0 ;
  assign n6360 = ~n6358 & n6359 ;
  assign n6361 = n2472 ^ n1538 ^ 1'b0 ;
  assign n6362 = n753 & ~n2638 ;
  assign n6363 = n6362 ^ n2184 ^ 1'b0 ;
  assign n6364 = n6363 ^ n4977 ^ 1'b0 ;
  assign n6365 = ~n6361 & n6364 ;
  assign n6366 = n6365 ^ x100 ^ 1'b0 ;
  assign n6367 = n5235 ^ n2535 ^ n796 ;
  assign n6368 = n1162 & ~n4562 ;
  assign n6369 = n6368 ^ n2069 ^ 1'b0 ;
  assign n6370 = n236 | n6369 ;
  assign n6371 = n6367 & ~n6370 ;
  assign n6372 = n1312 & n6371 ;
  assign n6373 = n3968 ^ n858 ^ 1'b0 ;
  assign n6374 = n4512 ^ n3404 ^ 1'b0 ;
  assign n6375 = n5980 ^ n1907 ^ 1'b0 ;
  assign n6376 = n1274 & n6375 ;
  assign n6377 = n6376 ^ n3953 ^ 1'b0 ;
  assign n6378 = ~n1640 & n6377 ;
  assign n6382 = n2772 ^ n274 ^ 1'b0 ;
  assign n6381 = ( n307 & ~n992 ) | ( n307 & n1127 ) | ( ~n992 & n1127 ) ;
  assign n6379 = n5454 ^ n4114 ^ 1'b0 ;
  assign n6380 = n1082 & n6379 ;
  assign n6383 = n6382 ^ n6381 ^ n6380 ;
  assign n6384 = n3022 & ~n6112 ;
  assign n6385 = ~n670 & n6384 ;
  assign n6386 = n2207 & ~n6385 ;
  assign n6387 = ~n4290 & n6386 ;
  assign n6388 = n2824 ^ n216 ^ 1'b0 ;
  assign n6389 = n4981 ^ n4180 ^ 1'b0 ;
  assign n6390 = n6388 & ~n6389 ;
  assign n6391 = n4119 & n6390 ;
  assign n6392 = ~n5037 & n6391 ;
  assign n6393 = n3517 & ~n5089 ;
  assign n6394 = ( n494 & n797 ) | ( n494 & n1262 ) | ( n797 & n1262 ) ;
  assign n6395 = n2665 | n6394 ;
  assign n6396 = n3121 ^ n3077 ^ n1218 ;
  assign n6397 = n6396 ^ n2209 ^ n1914 ;
  assign n6398 = n6397 ^ n5577 ^ n2416 ;
  assign n6399 = n4355 ^ n1787 ^ 1'b0 ;
  assign n6400 = n1923 | n6399 ;
  assign n6401 = n5642 ^ n3335 ^ n2063 ;
  assign n6402 = ( ~n3448 & n4856 ) | ( ~n3448 & n5266 ) | ( n4856 & n5266 ) ;
  assign n6403 = n3327 ^ n3173 ^ 1'b0 ;
  assign n6404 = n6402 & n6403 ;
  assign n6406 = n3508 ^ n2370 ^ 1'b0 ;
  assign n6407 = ~n211 & n6406 ;
  assign n6408 = ( n2041 & ~n3342 ) | ( n2041 & n6407 ) | ( ~n3342 & n6407 ) ;
  assign n6409 = n6408 ^ n4209 ^ 1'b0 ;
  assign n6405 = n5337 & ~n5508 ;
  assign n6410 = n6409 ^ n6405 ^ 1'b0 ;
  assign n6419 = n6036 ^ n353 ^ 1'b0 ;
  assign n6417 = n763 ^ n652 ^ 1'b0 ;
  assign n6418 = n3716 & ~n6417 ;
  assign n6420 = n6419 ^ n6418 ^ 1'b0 ;
  assign n6421 = ( ~n1488 & n5106 ) | ( ~n1488 & n6420 ) | ( n5106 & n6420 ) ;
  assign n6415 = n4521 ^ n934 ^ n847 ;
  assign n6416 = n2606 & n6415 ;
  assign n6422 = n6421 ^ n6416 ^ 1'b0 ;
  assign n6411 = n1699 & ~n5000 ;
  assign n6412 = n1722 & ~n5306 ;
  assign n6413 = n6412 ^ n3969 ^ n908 ;
  assign n6414 = n6411 | n6413 ;
  assign n6423 = n6422 ^ n6414 ^ 1'b0 ;
  assign n6424 = ( ~n1424 & n1434 ) | ( ~n1424 & n3624 ) | ( n1434 & n3624 ) ;
  assign n6425 = n5407 ^ n4387 ^ n626 ;
  assign n6426 = n1881 | n6425 ;
  assign n6427 = n6424 | n6426 ;
  assign n6428 = n4598 & n5929 ;
  assign n6429 = n649 & ~n2084 ;
  assign n6430 = n6429 ^ n2252 ^ n622 ;
  assign n6431 = n2307 | n3792 ;
  assign n6432 = n4318 & n6431 ;
  assign n6433 = n6432 ^ n3420 ^ n1858 ;
  assign n6434 = n3737 ^ n3173 ^ 1'b0 ;
  assign n6435 = ~n6433 & n6434 ;
  assign n6436 = ( n278 & n778 ) | ( n278 & ~n4614 ) | ( n778 & ~n4614 ) ;
  assign n6437 = n4915 ^ n4657 ^ 1'b0 ;
  assign n6438 = ( ~n1615 & n3030 ) | ( ~n1615 & n6022 ) | ( n3030 & n6022 ) ;
  assign n6440 = ~n1373 & n2688 ;
  assign n6439 = n1186 & n1448 ;
  assign n6441 = n6440 ^ n6439 ^ 1'b0 ;
  assign n6442 = n6438 & ~n6441 ;
  assign n6443 = ~n2937 & n3109 ;
  assign n6444 = ~n3860 & n6443 ;
  assign n6445 = n6442 | n6444 ;
  assign n6446 = ( ~n4259 & n5418 ) | ( ~n4259 & n5945 ) | ( n5418 & n5945 ) ;
  assign n6447 = n3980 ^ n1234 ^ 1'b0 ;
  assign n6448 = n180 & ~n6447 ;
  assign n6449 = n6448 ^ n1194 ^ 1'b0 ;
  assign n6450 = n5928 ^ n5804 ^ 1'b0 ;
  assign n6451 = ~n6268 & n6450 ;
  assign n6452 = n5519 & n6087 ;
  assign n6453 = n2968 ^ n2399 ^ n859 ;
  assign n6454 = n5174 ^ n379 ^ 1'b0 ;
  assign n6455 = n2499 | n6454 ;
  assign n6456 = n6453 & ~n6455 ;
  assign n6457 = n4802 ^ n4501 ^ n1472 ;
  assign n6458 = n4885 ^ n4444 ^ n3045 ;
  assign n6459 = n6457 & ~n6458 ;
  assign n6460 = n223 | n5572 ;
  assign n6461 = n152 & n2265 ;
  assign n6462 = n3108 ^ n493 ^ 1'b0 ;
  assign n6463 = n6462 ^ n2791 ^ 1'b0 ;
  assign n6464 = n2416 & ~n6463 ;
  assign n6465 = n6464 ^ n3417 ^ 1'b0 ;
  assign n6466 = n6163 | n6465 ;
  assign n6467 = n6466 ^ n4351 ^ 1'b0 ;
  assign n6470 = ~n219 & n2868 ;
  assign n6471 = n932 & n6470 ;
  assign n6469 = x63 & ~n2960 ;
  assign n6472 = n6471 ^ n6469 ^ 1'b0 ;
  assign n6468 = n2435 & ~n4527 ;
  assign n6473 = n6472 ^ n6468 ^ 1'b0 ;
  assign n6474 = n4507 ^ n897 ^ 1'b0 ;
  assign n6475 = n6473 & ~n6474 ;
  assign n6476 = n6475 ^ n1643 ^ 1'b0 ;
  assign n6477 = n1656 & n2626 ;
  assign n6478 = ~n4498 & n6477 ;
  assign n6479 = ~n6476 & n6478 ;
  assign n6480 = n3821 ^ n2874 ^ 1'b0 ;
  assign n6481 = n3121 ^ x51 ^ 1'b0 ;
  assign n6482 = ~n1741 & n3718 ;
  assign n6483 = n6482 ^ n1200 ^ 1'b0 ;
  assign n6484 = n613 | n1679 ;
  assign n6485 = ( n4367 & n6483 ) | ( n4367 & ~n6484 ) | ( n6483 & ~n6484 ) ;
  assign n6486 = ( n316 & ~n2971 ) | ( n316 & n5581 ) | ( ~n2971 & n5581 ) ;
  assign n6487 = n2471 & ~n6486 ;
  assign n6488 = n4741 & n6487 ;
  assign n6489 = n1150 | n2971 ;
  assign n6490 = n770 & n4376 ;
  assign n6491 = n6490 ^ n2567 ^ 1'b0 ;
  assign n6492 = ~x121 & n3550 ;
  assign n6493 = n617 | n1682 ;
  assign n6494 = ( n1420 & n1911 ) | ( n1420 & n5038 ) | ( n1911 & n5038 ) ;
  assign n6495 = n2002 ^ n398 ^ 1'b0 ;
  assign n6496 = n1576 & n6495 ;
  assign n6497 = n3824 & ~n6496 ;
  assign n6498 = n2264 | n6497 ;
  assign n6499 = n1907 & ~n3108 ;
  assign n6500 = n2555 & n6499 ;
  assign n6501 = n1625 & ~n6500 ;
  assign n6502 = n6501 ^ n932 ^ 1'b0 ;
  assign n6503 = n6498 & ~n6502 ;
  assign n6504 = n5657 ^ n4286 ^ 1'b0 ;
  assign n6505 = n1527 | n6504 ;
  assign n6506 = n1190 | n6505 ;
  assign n6512 = ( ~n965 & n2280 ) | ( ~n965 & n2965 ) | ( n2280 & n2965 ) ;
  assign n6507 = n4853 ^ n4431 ^ n533 ;
  assign n6508 = ( n1272 & n1403 ) | ( n1272 & ~n6507 ) | ( n1403 & ~n6507 ) ;
  assign n6509 = n1404 & ~n6508 ;
  assign n6510 = n6509 ^ n4015 ^ 1'b0 ;
  assign n6511 = n4172 & n6510 ;
  assign n6513 = n6512 ^ n6511 ^ n148 ;
  assign n6514 = n1943 & n5589 ;
  assign n6515 = n6514 ^ n3416 ^ 1'b0 ;
  assign n6516 = n4814 ^ n2252 ^ 1'b0 ;
  assign n6517 = n6460 & ~n6516 ;
  assign n6518 = n6491 ^ n5845 ^ 1'b0 ;
  assign n6519 = ~n3096 & n6518 ;
  assign n6520 = n1826 & ~n6076 ;
  assign n6521 = n4413 ^ n654 ^ 1'b0 ;
  assign n6522 = ~n2730 & n3515 ;
  assign n6524 = ( ~n2411 & n2470 ) | ( ~n2411 & n5445 ) | ( n2470 & n5445 ) ;
  assign n6523 = ( n843 & n1913 ) | ( n843 & ~n2074 ) | ( n1913 & ~n2074 ) ;
  assign n6525 = n6524 ^ n6523 ^ n3391 ;
  assign n6526 = n6525 ^ n4130 ^ 1'b0 ;
  assign n6527 = n6522 & ~n6526 ;
  assign n6530 = n3423 ^ n2333 ^ 1'b0 ;
  assign n6528 = n2089 & n3005 ;
  assign n6529 = n6528 ^ n6424 ^ 1'b0 ;
  assign n6531 = n6530 ^ n6529 ^ n5089 ;
  assign n6532 = n2957 ^ n2654 ^ 1'b0 ;
  assign n6533 = n1260 | n6532 ;
  assign n6534 = x127 & ~n6533 ;
  assign n6535 = n6534 ^ n971 ^ 1'b0 ;
  assign n6536 = x74 & n6329 ;
  assign n6537 = n4029 ^ n2570 ^ 1'b0 ;
  assign n6538 = n6537 ^ n302 ^ 1'b0 ;
  assign n6539 = n1020 & ~n2698 ;
  assign n6540 = n3765 & n6539 ;
  assign n6541 = n603 & n6540 ;
  assign n6542 = ~x106 & n1507 ;
  assign n6543 = ~n4027 & n6542 ;
  assign n6544 = n578 & n3058 ;
  assign n6545 = n5559 ^ n377 ^ 1'b0 ;
  assign n6546 = n3015 & ~n6545 ;
  assign n6547 = n4675 & n6546 ;
  assign n6548 = n1921 & n6547 ;
  assign n6549 = n2051 & n6548 ;
  assign n6550 = ( n876 & ~n6544 ) | ( n876 & n6549 ) | ( ~n6544 & n6549 ) ;
  assign n6551 = n641 ^ x96 ^ 1'b0 ;
  assign n6552 = n6551 ^ n3438 ^ 1'b0 ;
  assign n6553 = n4617 ^ n684 ^ 1'b0 ;
  assign n6554 = n1728 ^ n286 ^ 1'b0 ;
  assign n6555 = n4119 & n6554 ;
  assign n6556 = n2688 ^ n554 ^ 1'b0 ;
  assign n6557 = n6555 & ~n6556 ;
  assign n6559 = ~n370 & n2312 ;
  assign n6560 = n6559 ^ n153 ^ 1'b0 ;
  assign n6558 = ( n360 & n1415 ) | ( n360 & n2589 ) | ( n1415 & n2589 ) ;
  assign n6561 = n6560 ^ n6558 ^ 1'b0 ;
  assign n6562 = n5655 & n6561 ;
  assign n6563 = n908 & n6562 ;
  assign n6564 = n6563 ^ n3049 ^ 1'b0 ;
  assign n6565 = ~n1233 & n2192 ;
  assign n6566 = n6565 ^ n3122 ^ 1'b0 ;
  assign n6567 = n2182 & n6566 ;
  assign n6568 = n4130 & n6567 ;
  assign n6569 = ~n3332 & n3771 ;
  assign n6570 = n5784 & n6569 ;
  assign n6571 = n6570 ^ n2113 ^ n2016 ;
  assign n6572 = n3452 ^ n2714 ^ 1'b0 ;
  assign n6573 = n6572 ^ n6242 ^ 1'b0 ;
  assign n6574 = ~n540 & n3228 ;
  assign n6575 = ~n4420 & n6574 ;
  assign n6576 = n5314 & n6575 ;
  assign n6577 = n3157 & n6376 ;
  assign n6578 = ~n2418 & n6577 ;
  assign n6583 = ( ~n992 & n2493 ) | ( ~n992 & n4533 ) | ( n2493 & n4533 ) ;
  assign n6584 = n2034 ^ n1254 ^ 1'b0 ;
  assign n6585 = n6583 & n6584 ;
  assign n6586 = n6585 ^ n3521 ^ n1523 ;
  assign n6581 = n1732 ^ n419 ^ 1'b0 ;
  assign n6582 = ~n3651 & n6581 ;
  assign n6587 = n6586 ^ n6582 ^ n2905 ;
  assign n6579 = n4879 ^ n3769 ^ n1141 ;
  assign n6580 = ( ~x86 & n797 ) | ( ~x86 & n6579 ) | ( n797 & n6579 ) ;
  assign n6588 = n6587 ^ n6580 ^ 1'b0 ;
  assign n6589 = n3017 & n6588 ;
  assign n6590 = n4141 ^ n2923 ^ n196 ;
  assign n6591 = ~n761 & n1098 ;
  assign n6592 = n3472 ^ n3113 ^ 1'b0 ;
  assign n6593 = n6591 & ~n6592 ;
  assign n6594 = n6471 ^ n4063 ^ 1'b0 ;
  assign n6595 = n6593 & n6594 ;
  assign n6596 = ~n6590 & n6595 ;
  assign n6597 = n517 & ~n2406 ;
  assign n6598 = ~n2153 & n6597 ;
  assign n6599 = n710 & ~n4641 ;
  assign n6600 = n6599 ^ n2431 ^ 1'b0 ;
  assign n6601 = ( n1152 & n4155 ) | ( n1152 & n6600 ) | ( n4155 & n6600 ) ;
  assign n6602 = n2113 & n6601 ;
  assign n6603 = n3180 & n6602 ;
  assign n6604 = n3574 & ~n6603 ;
  assign n6605 = n1130 & n6604 ;
  assign n6606 = n3830 & ~n6605 ;
  assign n6607 = ~x31 & n6606 ;
  assign n6608 = n6598 | n6607 ;
  assign n6609 = n6608 ^ n4444 ^ 1'b0 ;
  assign n6610 = n3919 | n6221 ;
  assign n6611 = n3785 ^ n3090 ^ 1'b0 ;
  assign n6612 = n6609 ^ n5291 ^ 1'b0 ;
  assign n6620 = ( n340 & ~n5007 ) | ( n340 & n6301 ) | ( ~n5007 & n6301 ) ;
  assign n6615 = ~n429 & n5975 ;
  assign n6616 = ~n2372 & n6615 ;
  assign n6614 = n3037 ^ n203 ^ x97 ;
  assign n6617 = n6616 ^ n6614 ^ n2781 ;
  assign n6618 = n6617 ^ n2167 ^ 1'b0 ;
  assign n6619 = n2942 | n6618 ;
  assign n6613 = ~n2041 & n2275 ;
  assign n6621 = n6620 ^ n6619 ^ n6613 ;
  assign n6622 = n6319 | n6621 ;
  assign n6623 = n6622 ^ n2200 ^ 1'b0 ;
  assign n6624 = n223 | n6354 ;
  assign n6625 = n281 & ~n6624 ;
  assign n6626 = n5131 ^ n3104 ^ 1'b0 ;
  assign n6627 = ~n6625 & n6626 ;
  assign n6628 = n3277 ^ n2377 ^ n288 ;
  assign n6629 = n6168 ^ n5335 ^ n3068 ;
  assign n6630 = ( n3914 & ~n6628 ) | ( n3914 & n6629 ) | ( ~n6628 & n6629 ) ;
  assign n6631 = n3298 | n6630 ;
  assign n6632 = ( n1412 & n1516 ) | ( n1412 & ~n6631 ) | ( n1516 & ~n6631 ) ;
  assign n6633 = ~n3163 & n4142 ;
  assign n6634 = n4380 & ~n6633 ;
  assign n6635 = n5394 ^ n4072 ^ 1'b0 ;
  assign n6636 = n3735 ^ n3023 ^ n1379 ;
  assign n6637 = n5697 ^ n716 ^ 1'b0 ;
  assign n6638 = n6636 | n6637 ;
  assign n6639 = n3767 & n4637 ;
  assign n6640 = ~n1390 & n6639 ;
  assign n6641 = ( n2122 & n6420 ) | ( n2122 & n6640 ) | ( n6420 & n6640 ) ;
  assign n6642 = n251 & n2496 ;
  assign n6643 = n6642 ^ n5864 ^ 1'b0 ;
  assign n6644 = n1542 | n4933 ;
  assign n6645 = n6644 ^ x118 ^ 1'b0 ;
  assign n6646 = n4387 ^ n1725 ^ n1457 ;
  assign n6647 = ( ~n1035 & n1473 ) | ( ~n1035 & n6646 ) | ( n1473 & n6646 ) ;
  assign n6648 = n3529 ^ n344 ^ 1'b0 ;
  assign n6649 = n2127 & ~n3373 ;
  assign n6650 = n6648 | n6649 ;
  assign n6651 = n6647 & ~n6650 ;
  assign n6652 = ~n1184 & n5059 ;
  assign n6653 = n6652 ^ n5168 ^ n4806 ;
  assign n6654 = n6653 ^ n1199 ^ 1'b0 ;
  assign n6655 = n3781 ^ n3714 ^ 1'b0 ;
  assign n6656 = n2536 | n6655 ;
  assign n6658 = n566 & ~n1307 ;
  assign n6659 = ~n3628 & n6658 ;
  assign n6657 = n4029 & ~n4086 ;
  assign n6660 = n6659 ^ n6657 ^ 1'b0 ;
  assign n6661 = ~n561 & n1340 ;
  assign n6662 = n4837 & ~n5863 ;
  assign n6663 = n6662 ^ n370 ^ 1'b0 ;
  assign n6664 = ( n514 & n6661 ) | ( n514 & n6663 ) | ( n6661 & n6663 ) ;
  assign n6665 = n1199 | n4096 ;
  assign n6666 = n6665 ^ n614 ^ 1'b0 ;
  assign n6667 = n540 | n6666 ;
  assign n6668 = n434 & n2976 ;
  assign n6669 = n4876 ^ n3997 ^ 1'b0 ;
  assign n6670 = n6668 | n6669 ;
  assign n6671 = ( n411 & n1282 ) | ( n411 & n4256 ) | ( n1282 & n4256 ) ;
  assign n6672 = n6671 ^ n3836 ^ 1'b0 ;
  assign n6673 = n391 ^ n152 ^ 1'b0 ;
  assign n6674 = n809 & n2738 ;
  assign n6675 = n6674 ^ n480 ^ 1'b0 ;
  assign n6676 = n3549 ^ n1442 ^ n269 ;
  assign n6677 = n1874 & n4591 ;
  assign n6678 = n6676 | n6677 ;
  assign n6679 = n6675 | n6678 ;
  assign n6680 = ( x123 & ~n6673 ) | ( x123 & n6679 ) | ( ~n6673 & n6679 ) ;
  assign n6681 = n892 & ~n2479 ;
  assign n6683 = ~n4163 & n4475 ;
  assign n6684 = n6683 ^ n3005 ^ 1'b0 ;
  assign n6682 = n5786 | n6313 ;
  assign n6685 = n6684 ^ n6682 ^ 1'b0 ;
  assign n6686 = n3828 ^ n1209 ^ 1'b0 ;
  assign n6687 = n1362 & n4636 ;
  assign n6688 = n2751 ^ n1984 ^ n1388 ;
  assign n6689 = n6688 ^ n5746 ^ 1'b0 ;
  assign n6690 = n6687 & n6689 ;
  assign n6691 = ( ~n1469 & n1502 ) | ( ~n1469 & n1710 ) | ( n1502 & n1710 ) ;
  assign n6692 = n2651 & ~n6037 ;
  assign n6693 = ~n2397 & n6692 ;
  assign n6694 = n4219 & n4772 ;
  assign n6695 = n6694 ^ n2122 ^ 1'b0 ;
  assign n6696 = ( n5687 & ~n6646 ) | ( n5687 & n6695 ) | ( ~n6646 & n6695 ) ;
  assign n6697 = ( ~n2126 & n5673 ) | ( ~n2126 & n6696 ) | ( n5673 & n6696 ) ;
  assign n6698 = ~n1933 & n3440 ;
  assign n6699 = ~n2774 & n6072 ;
  assign n6700 = ( n2893 & ~n3926 ) | ( n2893 & n4437 ) | ( ~n3926 & n4437 ) ;
  assign n6701 = n2501 & ~n6700 ;
  assign n6702 = n4564 ^ n3263 ^ 1'b0 ;
  assign n6703 = ( n3477 & n4029 ) | ( n3477 & ~n6702 ) | ( n4029 & ~n6702 ) ;
  assign n6704 = n1036 & n3693 ;
  assign n6705 = ~n511 & n6704 ;
  assign n6706 = ~n2285 & n5942 ;
  assign n6707 = ~n6476 & n6706 ;
  assign n6708 = n6707 ^ n3178 ^ 1'b0 ;
  assign n6709 = ~n6705 & n6708 ;
  assign n6710 = ~n6354 & n6591 ;
  assign n6711 = ( ~n4029 & n5581 ) | ( ~n4029 & n6710 ) | ( n5581 & n6710 ) ;
  assign n6712 = n5045 ^ n2927 ^ n1110 ;
  assign n6714 = ( n836 & n975 ) | ( n836 & n2355 ) | ( n975 & n2355 ) ;
  assign n6713 = ( ~n418 & n4096 ) | ( ~n418 & n5723 ) | ( n4096 & n5723 ) ;
  assign n6715 = n6714 ^ n6713 ^ n5988 ;
  assign n6716 = n4413 ^ n3113 ^ 1'b0 ;
  assign n6720 = n1487 ^ n1037 ^ x113 ;
  assign n6721 = n2448 ^ x49 ^ 1'b0 ;
  assign n6722 = n6720 & ~n6721 ;
  assign n6717 = ~n709 & n1569 ;
  assign n6718 = ( n1078 & n1427 ) | ( n1078 & n6717 ) | ( n1427 & n6717 ) ;
  assign n6719 = ~n5279 & n6718 ;
  assign n6723 = n6722 ^ n6719 ^ 1'b0 ;
  assign n6724 = ( n852 & ~n2617 ) | ( n852 & n4295 ) | ( ~n2617 & n4295 ) ;
  assign n6725 = ( n2034 & ~n2245 ) | ( n2034 & n6724 ) | ( ~n2245 & n6724 ) ;
  assign n6726 = n5726 ^ n5683 ^ n2796 ;
  assign n6727 = n502 & ~n904 ;
  assign n6728 = n1542 & n6727 ;
  assign n6729 = n2217 | n6728 ;
  assign n6730 = n6729 ^ n2862 ^ x113 ;
  assign n6731 = n6730 ^ n1972 ^ 1'b0 ;
  assign n6732 = n6731 ^ n2218 ^ 1'b0 ;
  assign n6733 = n808 & n2947 ;
  assign n6735 = n2818 | n3975 ;
  assign n6736 = n742 | n6735 ;
  assign n6737 = ( n1677 & ~n2044 ) | ( n1677 & n6736 ) | ( ~n2044 & n6736 ) ;
  assign n6738 = ~n5357 & n6737 ;
  assign n6739 = n6738 ^ n809 ^ 1'b0 ;
  assign n6740 = ~n1317 & n6739 ;
  assign n6734 = n1669 & ~n3383 ;
  assign n6741 = n6740 ^ n6734 ^ 1'b0 ;
  assign n6742 = n4016 ^ n1015 ^ 1'b0 ;
  assign n6743 = ~n6659 & n6742 ;
  assign n6745 = ~n551 & n1031 ;
  assign n6746 = n6745 ^ n760 ^ 1'b0 ;
  assign n6744 = n412 ^ n374 ^ 1'b0 ;
  assign n6747 = n6746 ^ n6744 ^ n4012 ;
  assign n6748 = n6747 ^ n2359 ^ 1'b0 ;
  assign n6749 = n6743 & n6748 ;
  assign n6750 = ~n1113 & n1756 ;
  assign n6751 = ( n3674 & ~n4489 ) | ( n3674 & n6750 ) | ( ~n4489 & n6750 ) ;
  assign n6752 = n5701 ^ n2948 ^ 1'b0 ;
  assign n6753 = n1340 & n5737 ;
  assign n6754 = n3952 & n4359 ;
  assign n6757 = x106 & ~n1064 ;
  assign n6758 = n6757 ^ x13 ^ 1'b0 ;
  assign n6755 = n5351 | n6744 ;
  assign n6756 = n6755 ^ x90 ^ 1'b0 ;
  assign n6759 = n6758 ^ n6756 ^ 1'b0 ;
  assign n6760 = n146 | n6759 ;
  assign n6761 = n6280 ^ n4908 ^ n3667 ;
  assign n6762 = n3179 & ~n6761 ;
  assign n6763 = ~n4104 & n6762 ;
  assign n6764 = n6763 ^ n214 ^ 1'b0 ;
  assign n6765 = n3507 & n4180 ;
  assign n6766 = ~n2111 & n6765 ;
  assign n6767 = n6720 ^ n1422 ^ 1'b0 ;
  assign n6768 = ( n4442 & n4593 ) | ( n4442 & ~n6767 ) | ( n4593 & ~n6767 ) ;
  assign n6769 = ( ~n872 & n1425 ) | ( ~n872 & n2581 ) | ( n1425 & n2581 ) ;
  assign n6770 = n5703 ^ n2926 ^ 1'b0 ;
  assign n6771 = n6770 ^ n3751 ^ 1'b0 ;
  assign n6774 = n298 ^ n193 ^ 1'b0 ;
  assign n6772 = n6429 ^ n3372 ^ 1'b0 ;
  assign n6773 = n4170 & n6772 ;
  assign n6775 = n6774 ^ n6773 ^ 1'b0 ;
  assign n6776 = ( n6763 & n6771 ) | ( n6763 & n6775 ) | ( n6771 & n6775 ) ;
  assign n6777 = n1682 | n3613 ;
  assign n6778 = n2813 | n6777 ;
  assign n6779 = n1675 & ~n6778 ;
  assign n6780 = n2586 & ~n6779 ;
  assign n6781 = n6780 ^ n4361 ^ 1'b0 ;
  assign n6782 = ( n648 & n3508 ) | ( n648 & n6781 ) | ( n3508 & n6781 ) ;
  assign n6783 = n5814 ^ n2843 ^ n1881 ;
  assign n6784 = n6783 ^ n1777 ^ 1'b0 ;
  assign n6785 = n1858 & n3817 ;
  assign n6786 = n6785 ^ n2571 ^ 1'b0 ;
  assign n6787 = n4558 & ~n6786 ;
  assign n6788 = n627 & n3493 ;
  assign n6789 = n1898 | n6788 ;
  assign n6790 = n1304 & n2907 ;
  assign n6791 = n6790 ^ n6698 ^ 1'b0 ;
  assign n6792 = n3560 ^ n1811 ^ 1'b0 ;
  assign n6793 = n4425 ^ n1748 ^ 1'b0 ;
  assign n6796 = ~n2291 & n4469 ;
  assign n6797 = ~n4069 & n6796 ;
  assign n6798 = n4462 & n6797 ;
  assign n6794 = n1904 ^ n201 ^ 1'b0 ;
  assign n6795 = n5512 | n6794 ;
  assign n6799 = n6798 ^ n6795 ^ 1'b0 ;
  assign n6800 = n3215 & ~n6513 ;
  assign n6801 = n5652 ^ n1868 ^ n1634 ;
  assign n6802 = ~n646 & n2493 ;
  assign n6803 = n6802 ^ n265 ^ 1'b0 ;
  assign n6804 = n4473 ^ n2090 ^ 1'b0 ;
  assign n6805 = n6803 | n6804 ;
  assign n6806 = n6805 ^ n536 ^ 1'b0 ;
  assign n6810 = n6533 ^ n2134 ^ 1'b0 ;
  assign n6807 = ~n1040 & n3550 ;
  assign n6808 = n4895 & n6807 ;
  assign n6809 = ( x7 & n6720 ) | ( x7 & n6808 ) | ( n6720 & n6808 ) ;
  assign n6811 = n6810 ^ n6809 ^ n2285 ;
  assign n6812 = n1256 | n5879 ;
  assign n6813 = n1969 ^ n665 ^ 1'b0 ;
  assign n6814 = n5652 ^ n3868 ^ 1'b0 ;
  assign n6815 = n4413 & n6235 ;
  assign n6816 = n2695 & n6815 ;
  assign n6817 = n836 | n1118 ;
  assign n6818 = n6817 ^ n927 ^ 1'b0 ;
  assign n6819 = ( ~n614 & n2086 ) | ( ~n614 & n4585 ) | ( n2086 & n4585 ) ;
  assign n6820 = ( n2388 & n6818 ) | ( n2388 & n6819 ) | ( n6818 & n6819 ) ;
  assign n6825 = n1203 & ~n1782 ;
  assign n6826 = ( ~n2260 & n2988 ) | ( ~n2260 & n6825 ) | ( n2988 & n6825 ) ;
  assign n6827 = n6826 ^ n1739 ^ 1'b0 ;
  assign n6828 = n1511 | n6827 ;
  assign n6821 = n2333 ^ x26 ^ 1'b0 ;
  assign n6822 = ( x29 & ~n496 ) | ( x29 & n6821 ) | ( ~n496 & n6821 ) ;
  assign n6823 = n2149 | n6822 ;
  assign n6824 = n6823 ^ n511 ^ 1'b0 ;
  assign n6829 = n6828 ^ n6824 ^ 1'b0 ;
  assign n6830 = ( ~n2085 & n2120 ) | ( ~n2085 & n5756 ) | ( n2120 & n5756 ) ;
  assign n6831 = n160 & n1854 ;
  assign n6832 = n6831 ^ n1544 ^ 1'b0 ;
  assign n6833 = n5425 | n6832 ;
  assign n6834 = n1612 & n6833 ;
  assign n6838 = n1689 & ~n2879 ;
  assign n6835 = n5490 ^ n3160 ^ 1'b0 ;
  assign n6836 = n4130 | n6835 ;
  assign n6837 = n6836 ^ n3583 ^ 1'b0 ;
  assign n6839 = n6838 ^ n6837 ^ 1'b0 ;
  assign n6840 = n6834 & ~n6839 ;
  assign n6841 = n883 | n2844 ;
  assign n6842 = ~n2245 & n6841 ;
  assign n6843 = n1362 & n6842 ;
  assign n6844 = n5999 ^ n4803 ^ 1'b0 ;
  assign n6845 = n6844 ^ n4110 ^ 1'b0 ;
  assign n6846 = n3214 ^ n968 ^ 1'b0 ;
  assign n6847 = ~n1086 & n4746 ;
  assign n6848 = n4057 & n6847 ;
  assign n6849 = n2653 & n4295 ;
  assign n6850 = n6849 ^ n740 ^ 1'b0 ;
  assign n6851 = n3794 & ~n6850 ;
  assign n6854 = n2064 & n3744 ;
  assign n6855 = ( n236 & n2599 ) | ( n236 & n6854 ) | ( n2599 & n6854 ) ;
  assign n6856 = n6855 ^ n3257 ^ 1'b0 ;
  assign n6857 = n5337 & ~n6856 ;
  assign n6852 = ( n4524 & n4748 ) | ( n4524 & ~n5265 ) | ( n4748 & ~n5265 ) ;
  assign n6853 = n6852 ^ n4409 ^ n2241 ;
  assign n6858 = n6857 ^ n6853 ^ 1'b0 ;
  assign n6859 = ( n4783 & n5068 ) | ( n4783 & n6858 ) | ( n5068 & n6858 ) ;
  assign n6861 = n917 | n2933 ;
  assign n6862 = n3625 ^ n1324 ^ n915 ;
  assign n6863 = n6862 ^ n3254 ^ 1'b0 ;
  assign n6864 = n6861 & n6863 ;
  assign n6860 = ( n1318 & ~n2650 ) | ( n1318 & n4793 ) | ( ~n2650 & n4793 ) ;
  assign n6865 = n6864 ^ n6860 ^ n3060 ;
  assign n6866 = n3964 ^ n2717 ^ 1'b0 ;
  assign n6867 = n2719 | n6866 ;
  assign n6868 = n4821 & n6867 ;
  assign n6869 = ( n893 & ~n4124 ) | ( n893 & n5036 ) | ( ~n4124 & n5036 ) ;
  assign n6870 = n6869 ^ n2125 ^ 1'b0 ;
  assign n6875 = n1785 & ~n4685 ;
  assign n6871 = n3821 ^ n1475 ^ 1'b0 ;
  assign n6872 = n1132 & n6871 ;
  assign n6873 = n6872 ^ n1057 ^ 1'b0 ;
  assign n6874 = ~n3954 & n6873 ;
  assign n6876 = n6875 ^ n6874 ^ n6254 ;
  assign n6879 = n510 | n2617 ;
  assign n6880 = n6879 ^ n525 ^ 1'b0 ;
  assign n6877 = n573 & n935 ;
  assign n6878 = n1313 & ~n6877 ;
  assign n6881 = n6880 ^ n6878 ^ n5238 ;
  assign n6882 = n1331 ^ n721 ^ 1'b0 ;
  assign n6883 = ( x1 & ~n6087 ) | ( x1 & n6524 ) | ( ~n6087 & n6524 ) ;
  assign n6884 = n3961 ^ n3805 ^ 1'b0 ;
  assign n6885 = n6209 & n6884 ;
  assign n6886 = n3212 & ~n6885 ;
  assign n6887 = n6886 ^ n1386 ^ 1'b0 ;
  assign n6888 = ~n6883 & n6887 ;
  assign n6889 = ( n155 & n1805 ) | ( n155 & ~n3949 ) | ( n1805 & ~n3949 ) ;
  assign n6890 = ~n2291 & n5798 ;
  assign n6891 = ( ~n4456 & n6889 ) | ( ~n4456 & n6890 ) | ( n6889 & n6890 ) ;
  assign n6892 = n2332 & ~n3126 ;
  assign n6893 = n6892 ^ n2657 ^ 1'b0 ;
  assign n6894 = ~n5299 & n5851 ;
  assign n6895 = n3505 & ~n6264 ;
  assign n6896 = n2913 & n6895 ;
  assign n6897 = ( n4673 & n6651 ) | ( n4673 & n6896 ) | ( n6651 & n6896 ) ;
  assign n6905 = n1120 | n1905 ;
  assign n6898 = x90 & n447 ;
  assign n6899 = n2264 & n6898 ;
  assign n6900 = n2778 ^ x52 ^ 1'b0 ;
  assign n6901 = n6899 | n6900 ;
  assign n6902 = n6901 ^ n4397 ^ 1'b0 ;
  assign n6903 = n2393 | n6902 ;
  assign n6904 = n5497 & ~n6903 ;
  assign n6906 = n6905 ^ n6904 ^ 1'b0 ;
  assign n6907 = n4437 | n4717 ;
  assign n6908 = n6907 ^ n3537 ^ n2961 ;
  assign n6909 = n6651 & ~n6908 ;
  assign n6910 = n975 & n6043 ;
  assign n6911 = n3335 & n6910 ;
  assign n6912 = n6911 ^ n2086 ^ 1'b0 ;
  assign n6913 = n3586 | n6912 ;
  assign n6914 = ( n145 & n1483 ) | ( n145 & ~n2917 ) | ( n1483 & ~n2917 ) ;
  assign n6915 = ( n2772 & n3214 ) | ( n2772 & n6914 ) | ( n3214 & n6914 ) ;
  assign n6916 = n236 & n6915 ;
  assign n6917 = ( n542 & n1463 ) | ( n542 & ~n6551 ) | ( n1463 & ~n6551 ) ;
  assign n6918 = n2597 ^ n145 ^ 1'b0 ;
  assign n6919 = n2819 ^ n322 ^ 1'b0 ;
  assign n6920 = n568 & n6919 ;
  assign n6921 = ~x17 & n2471 ;
  assign n6922 = n4133 ^ n316 ^ 1'b0 ;
  assign n6923 = n4059 & ~n5073 ;
  assign n6924 = n6923 ^ n6269 ^ 1'b0 ;
  assign n6925 = n6922 & n6924 ;
  assign n6933 = ~n1478 & n4756 ;
  assign n6926 = ( n399 & n4092 ) | ( n399 & ~n4316 ) | ( n4092 & ~n4316 ) ;
  assign n6927 = ~n945 & n3093 ;
  assign n6928 = n1958 & n6927 ;
  assign n6929 = n770 | n6928 ;
  assign n6930 = n6929 ^ n5117 ^ n2595 ;
  assign n6931 = ~n6926 & n6930 ;
  assign n6932 = n6931 ^ n1767 ^ 1'b0 ;
  assign n6934 = n6933 ^ n6932 ^ n6106 ;
  assign n6935 = ( n2797 & n3129 ) | ( n2797 & ~n4814 ) | ( n3129 & ~n4814 ) ;
  assign n6936 = n2962 ^ n285 ^ 1'b0 ;
  assign n6937 = n6936 ^ n2995 ^ n684 ;
  assign n6938 = ( n4452 & ~n6779 ) | ( n4452 & n6937 ) | ( ~n6779 & n6937 ) ;
  assign n6939 = ( ~n4202 & n5475 ) | ( ~n4202 & n5821 ) | ( n5475 & n5821 ) ;
  assign n6943 = ~n1659 & n2910 ;
  assign n6944 = n6943 ^ n379 ^ 1'b0 ;
  assign n6941 = n1066 & ~n2580 ;
  assign n6942 = ~n234 & n6941 ;
  assign n6940 = x1 & n5610 ;
  assign n6945 = n6944 ^ n6942 ^ n6940 ;
  assign n6946 = n2862 ^ n614 ^ 1'b0 ;
  assign n6947 = ~n449 & n6946 ;
  assign n6948 = n6947 ^ n606 ^ 1'b0 ;
  assign n6949 = n1528 | n6948 ;
  assign n6950 = n5329 ^ n1224 ^ 1'b0 ;
  assign n6951 = n1758 | n6950 ;
  assign n6952 = n6951 ^ n800 ^ 1'b0 ;
  assign n6953 = ( ~n3244 & n3416 ) | ( ~n3244 & n3471 ) | ( n3416 & n3471 ) ;
  assign n6954 = n5910 ^ n1402 ^ 1'b0 ;
  assign n6955 = ~n6953 & n6954 ;
  assign n6956 = n6955 ^ n5289 ^ 1'b0 ;
  assign n6957 = n3323 ^ x29 ^ 1'b0 ;
  assign n6958 = n6956 | n6957 ;
  assign n6959 = n4216 & n6822 ;
  assign n6960 = ~n6217 & n6959 ;
  assign n6961 = n606 & ~n692 ;
  assign n6962 = n6961 ^ n4639 ^ 1'b0 ;
  assign n6965 = n178 & ~n1969 ;
  assign n6963 = n2328 ^ n1216 ^ 1'b0 ;
  assign n6964 = n1715 & ~n6963 ;
  assign n6966 = n6965 ^ n6964 ^ n5665 ;
  assign n6967 = n6962 & n6966 ;
  assign n6968 = n6633 ^ n5003 ^ 1'b0 ;
  assign n6969 = n3232 ^ n1565 ^ 1'b0 ;
  assign n6970 = n6969 ^ n1023 ^ 1'b0 ;
  assign n6971 = x20 & n6970 ;
  assign n6972 = ( ~n2934 & n4593 ) | ( ~n2934 & n6971 ) | ( n4593 & n6971 ) ;
  assign n6973 = n6916 ^ n6112 ^ 1'b0 ;
  assign n6974 = n4935 ^ n2233 ^ n154 ;
  assign n6975 = n3659 & n6974 ;
  assign n6976 = n6975 ^ n3020 ^ 1'b0 ;
  assign n6980 = n677 | n1202 ;
  assign n6979 = n675 & n1100 ;
  assign n6981 = n6980 ^ n6979 ^ 1'b0 ;
  assign n6977 = n5050 ^ n2668 ^ 1'b0 ;
  assign n6978 = ( x10 & n2733 ) | ( x10 & n6977 ) | ( n2733 & n6977 ) ;
  assign n6982 = n6981 ^ n6978 ^ n3942 ;
  assign n6983 = n684 ^ n164 ^ 1'b0 ;
  assign n6984 = n6983 ^ n4113 ^ n2931 ;
  assign n6985 = n2859 & ~n4708 ;
  assign n6986 = n1311 ^ x77 ^ 1'b0 ;
  assign n6987 = n6986 ^ n2328 ^ 1'b0 ;
  assign n6988 = n6985 & n6987 ;
  assign n6989 = n227 & ~n2971 ;
  assign n6990 = n5870 ^ n4779 ^ 1'b0 ;
  assign n6991 = n6989 | n6990 ;
  assign n6992 = ( n477 & n3914 ) | ( n477 & n6991 ) | ( n3914 & n6991 ) ;
  assign n6993 = n6992 ^ n3842 ^ 1'b0 ;
  assign n6995 = n4066 ^ x48 ^ 1'b0 ;
  assign n6996 = n4571 | n6995 ;
  assign n6997 = n6996 ^ n3701 ^ 1'b0 ;
  assign n6994 = n420 & n1561 ;
  assign n6998 = n6997 ^ n6994 ^ 1'b0 ;
  assign n6999 = n3373 & ~n6998 ;
  assign n7000 = ~n509 & n5463 ;
  assign n7001 = n7000 ^ n1921 ^ 1'b0 ;
  assign n7002 = n4193 | n7001 ;
  assign n7003 = n4084 & ~n4538 ;
  assign n7004 = n6285 ^ n1783 ^ 1'b0 ;
  assign n7005 = n5868 ^ n3490 ^ 1'b0 ;
  assign n7006 = n3341 & n4975 ;
  assign n7007 = ( ~n7004 & n7005 ) | ( ~n7004 & n7006 ) | ( n7005 & n7006 ) ;
  assign n7008 = n2769 & ~n7007 ;
  assign n7009 = n7003 | n7008 ;
  assign n7010 = ~n993 & n4146 ;
  assign n7011 = n7010 ^ n5586 ^ n4404 ;
  assign n7012 = n7011 ^ n6305 ^ 1'b0 ;
  assign n7013 = n6921 & ~n7012 ;
  assign n7014 = ~n1677 & n1892 ;
  assign n7015 = x6 & n7014 ;
  assign n7016 = n7015 ^ n3337 ^ 1'b0 ;
  assign n7017 = n3348 | n7016 ;
  assign n7018 = n685 & ~n3191 ;
  assign n7019 = n4590 ^ n4293 ^ 1'b0 ;
  assign n7020 = n1116 & n3609 ;
  assign n7022 = ( n2221 & n2841 ) | ( n2221 & n5847 ) | ( n2841 & n5847 ) ;
  assign n7021 = n6796 | n6884 ;
  assign n7023 = n7022 ^ n7021 ^ n5477 ;
  assign n7024 = n7020 & ~n7023 ;
  assign n7025 = n6447 & n7024 ;
  assign n7026 = n223 & n644 ;
  assign n7027 = n7026 ^ n4847 ^ 1'b0 ;
  assign n7028 = n4385 | n7027 ;
  assign n7029 = n7028 ^ n744 ^ 1'b0 ;
  assign n7030 = n2118 ^ n2026 ^ 1'b0 ;
  assign n7031 = n7030 ^ n478 ^ n404 ;
  assign n7032 = n6281 ^ n1881 ^ 1'b0 ;
  assign n7033 = n7032 ^ n1280 ^ n356 ;
  assign n7034 = n4538 ^ n1576 ^ n1442 ;
  assign n7035 = n1700 | n5331 ;
  assign n7036 = ( n613 & n7034 ) | ( n613 & ~n7035 ) | ( n7034 & ~n7035 ) ;
  assign n7037 = n832 | n6729 ;
  assign n7038 = n7037 ^ n3291 ^ 1'b0 ;
  assign n7039 = n7038 ^ n3218 ^ 1'b0 ;
  assign n7040 = n7036 | n7039 ;
  assign n7041 = ~n2902 & n5490 ;
  assign n7042 = ~n6736 & n7041 ;
  assign n7043 = n7042 ^ n3974 ^ 1'b0 ;
  assign n7044 = n6960 ^ n809 ^ 1'b0 ;
  assign n7045 = n3878 | n7044 ;
  assign n7046 = ~n3643 & n4857 ;
  assign n7047 = n1929 & n7046 ;
  assign n7048 = n3111 & ~n4844 ;
  assign n7049 = ~n250 & n7048 ;
  assign n7050 = n624 | n7049 ;
  assign n7051 = n7050 ^ n2062 ^ 1'b0 ;
  assign n7052 = n292 | n7051 ;
  assign n7053 = n723 | n2697 ;
  assign n7054 = n7053 ^ n3883 ^ n167 ;
  assign n7055 = n7054 ^ n3682 ^ 1'b0 ;
  assign n7056 = n4419 ^ n1348 ^ n962 ;
  assign n7057 = n523 & n969 ;
  assign n7058 = n7056 & n7057 ;
  assign n7059 = n3866 ^ n1682 ^ n1199 ;
  assign n7060 = n2218 & ~n7059 ;
  assign n7061 = ~n5329 & n7060 ;
  assign n7062 = n7061 ^ n5475 ^ 1'b0 ;
  assign n7063 = n4208 ^ n353 ^ 1'b0 ;
  assign n7064 = n7063 ^ n6135 ^ n1629 ;
  assign n7065 = ( n1078 & ~n4456 ) | ( n1078 & n7064 ) | ( ~n4456 & n7064 ) ;
  assign n7066 = ~n323 & n7065 ;
  assign n7067 = n585 & ~n1767 ;
  assign n7077 = ( x36 & ~n954 ) | ( x36 & n985 ) | ( ~n954 & n985 ) ;
  assign n7078 = n606 & ~n1447 ;
  assign n7079 = n1252 & n7078 ;
  assign n7080 = n4533 | n7079 ;
  assign n7081 = n1006 & ~n7080 ;
  assign n7082 = ( n555 & n6433 ) | ( n555 & ~n7081 ) | ( n6433 & ~n7081 ) ;
  assign n7083 = ( n1728 & n7077 ) | ( n1728 & ~n7082 ) | ( n7077 & ~n7082 ) ;
  assign n7072 = n5317 ^ n380 ^ 1'b0 ;
  assign n7073 = n2947 & ~n7072 ;
  assign n7074 = n2273 & ~n3537 ;
  assign n7075 = ~n7073 & n7074 ;
  assign n7069 = x93 ^ x32 ^ 1'b0 ;
  assign n7070 = n3418 & n7069 ;
  assign n7071 = n7070 ^ n2527 ^ 1'b0 ;
  assign n7076 = n7075 ^ n7071 ^ n699 ;
  assign n7068 = ~n1537 & n3403 ;
  assign n7084 = n7083 ^ n7076 ^ n7068 ;
  assign n7085 = n6810 ^ n4024 ^ 1'b0 ;
  assign n7086 = ~n1260 & n2471 ;
  assign n7087 = ~n866 & n7086 ;
  assign n7088 = ( n920 & ~n6198 ) | ( n920 & n7087 ) | ( ~n6198 & n7087 ) ;
  assign n7090 = n2788 ^ n1400 ^ 1'b0 ;
  assign n7091 = n2820 & ~n7090 ;
  assign n7089 = n1981 & n6288 ;
  assign n7092 = n7091 ^ n7089 ^ 1'b0 ;
  assign n7093 = n6949 | n7092 ;
  assign n7097 = n2041 | n2782 ;
  assign n7098 = ( n880 & n3706 ) | ( n880 & n7097 ) | ( n3706 & n7097 ) ;
  assign n7094 = n3166 ^ n3072 ^ 1'b0 ;
  assign n7095 = n4155 & n7094 ;
  assign n7096 = ~n5888 & n7095 ;
  assign n7099 = n7098 ^ n7096 ^ 1'b0 ;
  assign n7100 = ~n4160 & n5642 ;
  assign n7101 = ( ~n3790 & n5681 ) | ( ~n3790 & n7100 ) | ( n5681 & n7100 ) ;
  assign n7102 = n4170 & ~n4318 ;
  assign n7103 = n1687 & n7102 ;
  assign n7104 = n7103 ^ n923 ^ n238 ;
  assign n7105 = n7104 ^ n1304 ^ 1'b0 ;
  assign n7112 = x66 & n4607 ;
  assign n7113 = n4788 & n7112 ;
  assign n7106 = n1253 | n1766 ;
  assign n7107 = n7106 ^ n1789 ^ 1'b0 ;
  assign n7108 = n4180 ^ n1685 ^ 1'b0 ;
  assign n7109 = ~n2841 & n7108 ;
  assign n7110 = ~n6579 & n7109 ;
  assign n7111 = n7107 & ~n7110 ;
  assign n7114 = n7113 ^ n7111 ^ 1'b0 ;
  assign n7121 = n4913 & n5265 ;
  assign n7116 = ( n582 & n1639 ) | ( n582 & ~n3242 ) | ( n1639 & ~n3242 ) ;
  assign n7117 = n4452 & ~n7116 ;
  assign n7118 = n6295 & n7117 ;
  assign n7119 = ~n918 & n7118 ;
  assign n7120 = n4660 & ~n7119 ;
  assign n7122 = n7121 ^ n7120 ^ 1'b0 ;
  assign n7115 = n445 & ~n4434 ;
  assign n7123 = n7122 ^ n7115 ^ 1'b0 ;
  assign n7124 = n5058 ^ n1769 ^ 1'b0 ;
  assign n7125 = ( n4126 & n4646 ) | ( n4126 & ~n7124 ) | ( n4646 & ~n7124 ) ;
  assign n7126 = ~n4852 & n6332 ;
  assign n7127 = ~n7125 & n7126 ;
  assign n7128 = n6960 & n7127 ;
  assign n7129 = n1040 | n3760 ;
  assign n7130 = n7129 ^ n529 ^ 1'b0 ;
  assign n7131 = n816 & n7130 ;
  assign n7132 = x107 & ~n1940 ;
  assign n7133 = n7132 ^ n3287 ^ 1'b0 ;
  assign n7134 = ~n1080 & n1485 ;
  assign n7135 = n7133 & n7134 ;
  assign n7136 = n1408 | n7135 ;
  assign n7137 = n1310 & ~n7136 ;
  assign n7138 = n5728 | n7137 ;
  assign n7139 = n7138 ^ n3150 ^ 1'b0 ;
  assign n7141 = ( x66 & n3407 ) | ( x66 & n4712 ) | ( n3407 & n4712 ) ;
  assign n7140 = n4430 | n6309 ;
  assign n7142 = n7141 ^ n7140 ^ 1'b0 ;
  assign n7143 = ~n2393 & n7142 ;
  assign n7144 = n1692 & ~n6465 ;
  assign n7145 = n6106 | n7144 ;
  assign n7146 = n7145 ^ n5072 ^ 1'b0 ;
  assign n7147 = n4059 ^ n3871 ^ n3011 ;
  assign n7148 = ( n3816 & n5358 ) | ( n3816 & n7147 ) | ( n5358 & n7147 ) ;
  assign n7149 = n1643 | n4462 ;
  assign n7150 = n7149 ^ n1329 ^ 1'b0 ;
  assign n7151 = n3449 | n4795 ;
  assign n7152 = n3298 | n7151 ;
  assign n7153 = ( n1167 & n6333 ) | ( n1167 & n7152 ) | ( n6333 & n7152 ) ;
  assign n7154 = n2411 ^ n1369 ^ 1'b0 ;
  assign n7155 = n7153 & n7154 ;
  assign n7156 = ~n261 & n7155 ;
  assign n7157 = n1931 & ~n3517 ;
  assign n7158 = n7157 ^ n6098 ^ 1'b0 ;
  assign n7159 = n2430 & ~n5824 ;
  assign n7160 = ~n2528 & n7159 ;
  assign n7161 = n887 & ~n7160 ;
  assign n7162 = n2478 & n7161 ;
  assign n7163 = n4724 ^ n1314 ^ 1'b0 ;
  assign n7164 = ~n7162 & n7163 ;
  assign n7165 = n3063 & ~n4982 ;
  assign n7166 = ~n7164 & n7165 ;
  assign n7167 = n1960 | n7166 ;
  assign n7168 = n7167 ^ n4432 ^ 1'b0 ;
  assign n7169 = n1360 | n1419 ;
  assign n7170 = n7169 ^ n3753 ^ n3421 ;
  assign n7171 = n7170 ^ n4041 ^ n264 ;
  assign n7172 = n4841 ^ n4088 ^ 1'b0 ;
  assign n7173 = n7172 ^ n6573 ^ 1'b0 ;
  assign n7174 = n6632 ^ n4240 ^ n412 ;
  assign n7175 = n6247 ^ n3524 ^ 1'b0 ;
  assign n7176 = ~n5343 & n5400 ;
  assign n7177 = n2215 | n7176 ;
  assign n7178 = ~n1673 & n2984 ;
  assign n7179 = ~n697 & n7178 ;
  assign n7180 = n7179 ^ n2801 ^ 1'b0 ;
  assign n7181 = n3433 ^ x84 ^ 1'b0 ;
  assign n7182 = n2637 | n7181 ;
  assign n7183 = ( n4323 & ~n5678 ) | ( n4323 & n7182 ) | ( ~n5678 & n7182 ) ;
  assign n7184 = ( n169 & n1785 ) | ( n169 & ~n6029 ) | ( n1785 & ~n6029 ) ;
  assign n7185 = n193 | n2619 ;
  assign n7186 = n5569 | n7185 ;
  assign n7187 = ~n3676 & n5767 ;
  assign n7188 = n4801 ^ n2972 ^ 1'b0 ;
  assign n7189 = ~n2719 & n7188 ;
  assign n7190 = n7189 ^ n5345 ^ 1'b0 ;
  assign n7191 = n7187 | n7190 ;
  assign n7192 = n6699 ^ n2023 ^ n1160 ;
  assign n7193 = n212 & ~n960 ;
  assign n7196 = ~n1763 & n3375 ;
  assign n7195 = n5258 & n6176 ;
  assign n7197 = n7196 ^ n7195 ^ 1'b0 ;
  assign n7194 = n5040 | n5827 ;
  assign n7198 = n7197 ^ n7194 ^ 1'b0 ;
  assign n7199 = n1923 | n7198 ;
  assign n7203 = n5455 ^ n3453 ^ 1'b0 ;
  assign n7200 = ( n855 & n1148 ) | ( n855 & ~n2988 ) | ( n1148 & ~n2988 ) ;
  assign n7201 = n1903 & ~n5740 ;
  assign n7202 = n7200 & ~n7201 ;
  assign n7204 = n7203 ^ n7202 ^ 1'b0 ;
  assign n7205 = n2688 & ~n7170 ;
  assign n7206 = n7205 ^ n6515 ^ 1'b0 ;
  assign n7207 = n6730 ^ n2026 ^ 1'b0 ;
  assign n7208 = x123 & ~n7207 ;
  assign n7209 = n490 & n7208 ;
  assign n7210 = ~n1713 & n7209 ;
  assign n7211 = n1605 & n6653 ;
  assign n7212 = n3537 ^ n672 ^ 1'b0 ;
  assign n7213 = n5183 ^ n2083 ^ 1'b0 ;
  assign n7214 = n773 & ~n3779 ;
  assign n7216 = ( n1491 & n1674 ) | ( n1491 & n4499 ) | ( n1674 & n4499 ) ;
  assign n7215 = n1483 & n3059 ;
  assign n7217 = n7216 ^ n7215 ^ 1'b0 ;
  assign n7218 = n5792 & n6198 ;
  assign n7219 = ~n1058 & n7218 ;
  assign n7220 = n7219 ^ n1362 ^ 1'b0 ;
  assign n7221 = n6073 & n7220 ;
  assign n7222 = n6778 & n7221 ;
  assign n7223 = n3691 & n7222 ;
  assign n7224 = n7223 ^ n3851 ^ n3625 ;
  assign n7225 = n180 | n3814 ;
  assign n7226 = n2796 ^ n2105 ^ 1'b0 ;
  assign n7227 = n7226 ^ n3242 ^ n1089 ;
  assign n7228 = n4517 & n5543 ;
  assign n7229 = ~n2650 & n7228 ;
  assign n7230 = n7227 & ~n7229 ;
  assign n7231 = n7230 ^ n836 ^ 1'b0 ;
  assign n7232 = n2651 ^ n1664 ^ 1'b0 ;
  assign n7233 = n7232 ^ n2195 ^ x1 ;
  assign n7234 = n7233 ^ n1496 ^ 1'b0 ;
  assign n7235 = n7234 ^ n540 ^ 1'b0 ;
  assign n7246 = n4521 ^ n494 ^ 1'b0 ;
  assign n7242 = n285 | n701 ;
  assign n7243 = n398 & ~n7242 ;
  assign n7238 = n3670 ^ n578 ^ n307 ;
  assign n7239 = n1806 | n3657 ;
  assign n7240 = n7238 & ~n7239 ;
  assign n7241 = ( n1145 & n4413 ) | ( n1145 & n7240 ) | ( n4413 & n7240 ) ;
  assign n7236 = n2549 ^ n1992 ^ n210 ;
  assign n7237 = ~n2044 & n7236 ;
  assign n7244 = n7243 ^ n7241 ^ n7237 ;
  assign n7245 = n7244 ^ n3903 ^ 1'b0 ;
  assign n7247 = n7246 ^ n7245 ^ n5924 ;
  assign n7248 = n5370 ^ n561 ^ n270 ;
  assign n7249 = n2658 & n7248 ;
  assign n7250 = n1201 & n6252 ;
  assign n7251 = n7250 ^ n4083 ^ 1'b0 ;
  assign n7254 = n4142 ^ n307 ^ 1'b0 ;
  assign n7255 = ( ~n986 & n3613 ) | ( ~n986 & n7254 ) | ( n3613 & n7254 ) ;
  assign n7252 = n422 & ~n1008 ;
  assign n7253 = ~n5982 & n7252 ;
  assign n7256 = n7255 ^ n7253 ^ x119 ;
  assign n7257 = n4286 & n7256 ;
  assign n7258 = ( n551 & n1164 ) | ( n551 & ~n3787 ) | ( n1164 & ~n3787 ) ;
  assign n7259 = n670 & ~n7258 ;
  assign n7260 = n7257 & n7259 ;
  assign n7261 = n6166 ^ n6106 ^ n138 ;
  assign n7262 = n1307 | n5916 ;
  assign n7263 = n6885 & ~n7262 ;
  assign n7264 = n1079 | n1887 ;
  assign n7265 = n7264 ^ n1649 ^ 1'b0 ;
  assign n7266 = n7265 ^ n1394 ^ n443 ;
  assign n7267 = x58 & n5304 ;
  assign n7268 = n6746 & n7267 ;
  assign n7269 = n3160 & ~n7268 ;
  assign n7270 = n7269 ^ n1373 ^ 1'b0 ;
  assign n7271 = ~n2756 & n7270 ;
  assign n7272 = ~n7266 & n7271 ;
  assign n7273 = n1014 & n2744 ;
  assign n7274 = ( ~n5863 & n6833 ) | ( ~n5863 & n7273 ) | ( n6833 & n7273 ) ;
  assign n7276 = n4855 ^ n1971 ^ 1'b0 ;
  assign n7277 = n7276 ^ n2625 ^ n1706 ;
  assign n7275 = ~n2077 & n5072 ;
  assign n7278 = n7277 ^ n7275 ^ 1'b0 ;
  assign n7279 = n7278 ^ n1840 ^ 1'b0 ;
  assign n7280 = n6365 & ~n7279 ;
  assign n7281 = ( n1573 & n5051 ) | ( n1573 & ~n7280 ) | ( n5051 & ~n7280 ) ;
  assign n7282 = n5907 & ~n7281 ;
  assign n7283 = n7282 ^ n5299 ^ 1'b0 ;
  assign n7290 = n1825 | n6881 ;
  assign n7291 = n285 | n7290 ;
  assign n7292 = n3118 | n5276 ;
  assign n7293 = n1269 & ~n2839 ;
  assign n7294 = ( n2459 & ~n4269 ) | ( n2459 & n7293 ) | ( ~n4269 & n7293 ) ;
  assign n7295 = n2355 | n2982 ;
  assign n7296 = n3158 & ~n7295 ;
  assign n7297 = n616 & n7296 ;
  assign n7298 = ( n2121 & n7294 ) | ( n2121 & n7297 ) | ( n7294 & n7297 ) ;
  assign n7299 = n7292 & n7298 ;
  assign n7300 = ~n7291 & n7299 ;
  assign n7284 = ( x108 & n393 ) | ( x108 & ~n535 ) | ( n393 & ~n535 ) ;
  assign n7285 = ~n322 & n7284 ;
  assign n7286 = n7285 ^ n965 ^ 1'b0 ;
  assign n7287 = n4978 & ~n7286 ;
  assign n7288 = n3391 & ~n7287 ;
  assign n7289 = ~n6752 & n7288 ;
  assign n7301 = n7300 ^ n7289 ^ 1'b0 ;
  assign n7302 = n2841 ^ n2158 ^ 1'b0 ;
  assign n7303 = n5781 & n7302 ;
  assign n7306 = ( n846 & ~n1895 ) | ( n846 & n7116 ) | ( ~n1895 & n7116 ) ;
  assign n7304 = n4182 & ~n6036 ;
  assign n7305 = n5919 | n7304 ;
  assign n7307 = n7306 ^ n7305 ^ 1'b0 ;
  assign n7308 = n5929 ^ n3232 ^ n1347 ;
  assign n7309 = ~n6258 & n7308 ;
  assign n7310 = ~n6329 & n7309 ;
  assign n7311 = n3912 & n5685 ;
  assign n7312 = n358 & ~n6408 ;
  assign n7313 = ~n732 & n7312 ;
  assign n7314 = ~n173 & n3589 ;
  assign n7315 = n839 | n1214 ;
  assign n7316 = n1591 & ~n7315 ;
  assign n7317 = ( ~n900 & n4767 ) | ( ~n900 & n7316 ) | ( n4767 & n7316 ) ;
  assign n7318 = n3222 ^ n310 ^ 1'b0 ;
  assign n7319 = ( n555 & n7317 ) | ( n555 & ~n7318 ) | ( n7317 & ~n7318 ) ;
  assign n7320 = n7319 ^ n2670 ^ 1'b0 ;
  assign n7321 = n571 & n7320 ;
  assign n7322 = n1552 | n4926 ;
  assign n7323 = n7322 ^ n5904 ^ 1'b0 ;
  assign n7324 = n4397 ^ n4069 ^ 1'b0 ;
  assign n7325 = n7324 ^ n3356 ^ 1'b0 ;
  assign n7326 = n4269 | n7325 ;
  assign n7327 = ( n719 & ~n4556 ) | ( n719 & n7326 ) | ( ~n4556 & n7326 ) ;
  assign n7328 = n7327 ^ n6034 ^ 1'b0 ;
  assign n7329 = n4003 ^ n3383 ^ 1'b0 ;
  assign n7331 = n2267 ^ n1905 ^ n882 ;
  assign n7332 = n7331 ^ n4717 ^ 1'b0 ;
  assign n7330 = n3655 & n5192 ;
  assign n7333 = n7332 ^ n7330 ^ 1'b0 ;
  assign n7334 = n4451 & ~n7333 ;
  assign n7335 = n4904 ^ n4224 ^ 1'b0 ;
  assign n7336 = n796 & n7335 ;
  assign n7337 = n7336 ^ n4099 ^ 1'b0 ;
  assign n7338 = ( x3 & n2469 ) | ( x3 & n7337 ) | ( n2469 & n7337 ) ;
  assign n7339 = n6986 ^ n4737 ^ x40 ;
  assign n7340 = ~n7221 & n7339 ;
  assign n7341 = ( n259 & n382 ) | ( n259 & n4152 ) | ( n382 & n4152 ) ;
  assign n7342 = n1051 ^ n737 ^ 1'b0 ;
  assign n7343 = n2422 ^ n252 ^ x127 ;
  assign n7344 = ( n2219 & ~n2415 ) | ( n2219 & n4542 ) | ( ~n2415 & n4542 ) ;
  assign n7345 = ~n2847 & n6348 ;
  assign n7346 = n7345 ^ n1376 ^ 1'b0 ;
  assign n7347 = n2759 | n4973 ;
  assign n7348 = n4110 | n7347 ;
  assign n7349 = n7348 ^ x67 ^ 1'b0 ;
  assign n7350 = n1348 | n7342 ;
  assign n7351 = n2278 & n4535 ;
  assign n7353 = n3521 ^ n1936 ^ 1'b0 ;
  assign n7354 = n463 & ~n7353 ;
  assign n7355 = n7354 ^ n6718 ^ x92 ;
  assign n7352 = n945 | n3178 ;
  assign n7356 = n7355 ^ n7352 ^ 1'b0 ;
  assign n7357 = n4179 | n7356 ;
  assign n7358 = n3595 & ~n7357 ;
  assign n7359 = n7358 ^ n6714 ^ 1'b0 ;
  assign n7360 = n5555 ^ n5174 ^ 1'b0 ;
  assign n7361 = n6661 ^ n2229 ^ 1'b0 ;
  assign n7362 = n4037 & ~n4484 ;
  assign n7363 = ~n7361 & n7362 ;
  assign n7364 = n258 & n1112 ;
  assign n7365 = ~n1150 & n7364 ;
  assign n7366 = n7363 & n7365 ;
  assign n7367 = n6828 ^ n1343 ^ 1'b0 ;
  assign n7368 = n7367 ^ n1921 ^ n1726 ;
  assign n7369 = ( n374 & n2895 ) | ( n374 & n3298 ) | ( n2895 & n3298 ) ;
  assign n7370 = n5967 ^ n2219 ^ n1777 ;
  assign n7371 = n7369 & n7370 ;
  assign n7372 = n7371 ^ n4958 ^ 1'b0 ;
  assign n7373 = n1211 ^ n901 ^ 1'b0 ;
  assign n7374 = ( n1348 & n6166 ) | ( n1348 & n7373 ) | ( n6166 & n7373 ) ;
  assign n7375 = n1923 & ~n7374 ;
  assign n7376 = n325 | n7375 ;
  assign n7377 = n4091 ^ n1108 ^ 1'b0 ;
  assign n7378 = n5242 & n7377 ;
  assign n7379 = ~n5588 & n7378 ;
  assign n7384 = x43 & n2443 ;
  assign n7385 = ~n314 & n7384 ;
  assign n7380 = n1055 | n7358 ;
  assign n7381 = n7380 ^ n1882 ^ 1'b0 ;
  assign n7382 = n7381 ^ n5502 ^ 1'b0 ;
  assign n7383 = n4713 | n7382 ;
  assign n7386 = n7385 ^ n7383 ^ 1'b0 ;
  assign n7387 = ~n5046 & n7386 ;
  assign n7388 = n1398 & ~n4314 ;
  assign n7389 = n804 & n7388 ;
  assign n7393 = ( n1079 & ~n1918 ) | ( n1079 & n3874 ) | ( ~n1918 & n3874 ) ;
  assign n7394 = n3581 ^ n2069 ^ 1'b0 ;
  assign n7395 = n7393 & ~n7394 ;
  assign n7390 = ~n5079 & n5594 ;
  assign n7391 = n7390 ^ n6640 ^ 1'b0 ;
  assign n7392 = ~n6281 & n7391 ;
  assign n7396 = n7395 ^ n7392 ^ 1'b0 ;
  assign n7397 = n5597 ^ n3395 ^ 1'b0 ;
  assign n7400 = n2648 ^ n458 ^ 1'b0 ;
  assign n7398 = n1157 & n5128 ;
  assign n7399 = n3082 & n7398 ;
  assign n7401 = n7400 ^ n7399 ^ 1'b0 ;
  assign n7402 = n7401 ^ n1591 ^ 1'b0 ;
  assign n7403 = n319 | n7101 ;
  assign n7404 = n7403 ^ n5857 ^ n3821 ;
  assign n7405 = ( ~n1923 & n2553 ) | ( ~n1923 & n4385 ) | ( n2553 & n4385 ) ;
  assign n7406 = ( n2761 & n4610 ) | ( n2761 & n7405 ) | ( n4610 & n7405 ) ;
  assign n7407 = n3262 | n7054 ;
  assign n7408 = n7407 ^ n365 ^ n180 ;
  assign n7409 = n1414 & ~n7360 ;
  assign n7410 = n1598 ^ n654 ^ 1'b0 ;
  assign n7411 = n6620 ^ n5872 ^ n536 ;
  assign n7412 = ( n161 & n1988 ) | ( n161 & ~n7411 ) | ( n1988 & ~n7411 ) ;
  assign n7416 = ~n1764 & n4609 ;
  assign n7417 = ~n775 & n7416 ;
  assign n7418 = n5000 ^ n4431 ^ n1148 ;
  assign n7419 = ~n7417 & n7418 ;
  assign n7420 = n7419 ^ n708 ^ 1'b0 ;
  assign n7413 = ( ~n4493 & n4706 ) | ( ~n4493 & n5139 ) | ( n4706 & n5139 ) ;
  assign n7414 = n3584 & n7413 ;
  assign n7415 = n4601 & n7414 ;
  assign n7421 = n7420 ^ n7415 ^ 1'b0 ;
  assign n7422 = n5134 ^ n5056 ^ n2517 ;
  assign n7423 = n1065 & ~n7422 ;
  assign n7424 = ~n7421 & n7423 ;
  assign n7425 = n1794 & ~n4855 ;
  assign n7429 = n3116 & ~n5832 ;
  assign n7430 = ~n3933 & n7429 ;
  assign n7426 = n620 | n4233 ;
  assign n7427 = n3772 & ~n7426 ;
  assign n7428 = n7427 ^ n4178 ^ 1'b0 ;
  assign n7431 = n7430 ^ n7428 ^ n5936 ;
  assign n7432 = n591 ^ n422 ^ 1'b0 ;
  assign n7433 = ( n5380 & n5399 ) | ( n5380 & n7432 ) | ( n5399 & n7432 ) ;
  assign n7434 = n7431 | n7433 ;
  assign n7446 = n1856 & ~n5559 ;
  assign n7447 = n7446 ^ n2450 ^ 1'b0 ;
  assign n7448 = n1008 | n7447 ;
  assign n7435 = n6411 ^ n6127 ^ x112 ;
  assign n7436 = n618 | n7435 ;
  assign n7437 = n2395 | n7436 ;
  assign n7438 = n7437 ^ n563 ^ n339 ;
  assign n7439 = x83 & n1933 ;
  assign n7441 = n2374 | n6379 ;
  assign n7442 = n7441 ^ n3664 ^ 1'b0 ;
  assign n7440 = n173 & ~n1483 ;
  assign n7443 = n7442 ^ n7440 ^ 1'b0 ;
  assign n7444 = n7439 & ~n7443 ;
  assign n7445 = n7438 & n7444 ;
  assign n7449 = n7448 ^ n7445 ^ 1'b0 ;
  assign n7450 = n2039 & n7449 ;
  assign n7451 = n7450 ^ n3860 ^ 1'b0 ;
  assign n7452 = ~n5291 & n5573 ;
  assign n7453 = ~n614 & n7452 ;
  assign n7454 = n1502 & ~n1561 ;
  assign n7455 = n7454 ^ n630 ^ 1'b0 ;
  assign n7456 = ~n1622 & n7455 ;
  assign n7457 = n7456 ^ n6149 ^ 1'b0 ;
  assign n7458 = n4603 & n4952 ;
  assign n7459 = n7458 ^ n775 ^ 1'b0 ;
  assign n7460 = n3586 | n7459 ;
  assign n7461 = n432 & n2685 ;
  assign n7462 = n7461 ^ n684 ^ 1'b0 ;
  assign n7463 = ( n356 & n4312 ) | ( n356 & ~n7462 ) | ( n4312 & ~n7462 ) ;
  assign n7464 = n4600 ^ n2179 ^ 1'b0 ;
  assign n7469 = ( x73 & n2759 ) | ( x73 & n6803 ) | ( n2759 & n6803 ) ;
  assign n7470 = n7469 ^ n1338 ^ 1'b0 ;
  assign n7465 = n5199 ^ n2781 ^ 1'b0 ;
  assign n7466 = n3822 | n7465 ;
  assign n7467 = n4768 & n6971 ;
  assign n7468 = n7466 & n7467 ;
  assign n7471 = n7470 ^ n7468 ^ 1'b0 ;
  assign n7472 = n2179 ^ n138 ^ 1'b0 ;
  assign n7473 = n471 & ~n7472 ;
  assign n7474 = ( n477 & n482 ) | ( n477 & n1129 ) | ( n482 & n1129 ) ;
  assign n7475 = n6796 ^ n4472 ^ n730 ;
  assign n7476 = ~n624 & n7475 ;
  assign n7477 = n1747 & n7476 ;
  assign n7478 = n7474 | n7477 ;
  assign n7479 = n7478 ^ n2575 ^ 1'b0 ;
  assign n7482 = n2454 ^ n436 ^ 1'b0 ;
  assign n7480 = n4675 & n6072 ;
  assign n7481 = n477 & n7480 ;
  assign n7483 = n7482 ^ n7481 ^ 1'b0 ;
  assign n7484 = n7479 & ~n7483 ;
  assign n7485 = n1071 & n6284 ;
  assign n7486 = ( x112 & n2012 ) | ( x112 & ~n2751 ) | ( n2012 & ~n2751 ) ;
  assign n7487 = ( n410 & n1731 ) | ( n410 & ~n2335 ) | ( n1731 & ~n2335 ) ;
  assign n7488 = n2510 ^ n1116 ^ n412 ;
  assign n7489 = ( n7486 & ~n7487 ) | ( n7486 & n7488 ) | ( ~n7487 & n7488 ) ;
  assign n7490 = ( ~n4033 & n4220 ) | ( ~n4033 & n6746 ) | ( n4220 & n6746 ) ;
  assign n7491 = n3434 ^ n1441 ^ n828 ;
  assign n7492 = n4182 & ~n7491 ;
  assign n7493 = n7490 & n7492 ;
  assign n7494 = ~n808 & n4776 ;
  assign n7495 = ( n616 & ~n771 ) | ( n616 & n982 ) | ( ~n771 & n982 ) ;
  assign n7496 = ~n3329 & n7495 ;
  assign n7497 = n4128 & n7496 ;
  assign n7498 = n238 | n7497 ;
  assign n7499 = n7498 ^ n4596 ^ 1'b0 ;
  assign n7503 = n351 | n7079 ;
  assign n7504 = n7503 ^ x113 ^ 1'b0 ;
  assign n7505 = n2917 ^ n2857 ^ 1'b0 ;
  assign n7506 = ( n2069 & n2582 ) | ( n2069 & ~n7505 ) | ( n2582 & ~n7505 ) ;
  assign n7507 = n7506 ^ n1560 ^ x23 ;
  assign n7508 = n307 | n1317 ;
  assign n7509 = n2070 & n7508 ;
  assign n7510 = n7509 ^ n4180 ^ 1'b0 ;
  assign n7511 = ( ~n5295 & n7507 ) | ( ~n5295 & n7510 ) | ( n7507 & n7510 ) ;
  assign n7512 = ( ~n1956 & n7504 ) | ( ~n1956 & n7511 ) | ( n7504 & n7511 ) ;
  assign n7500 = n644 & ~n6659 ;
  assign n7501 = n7500 ^ n848 ^ 1'b0 ;
  assign n7502 = n7501 ^ n1448 ^ 1'b0 ;
  assign n7513 = n7512 ^ n7502 ^ 1'b0 ;
  assign n7514 = n7226 ^ n6959 ^ n820 ;
  assign n7515 = n139 & n7514 ;
  assign n7516 = ~n2184 & n7515 ;
  assign n7517 = n3176 | n7516 ;
  assign n7518 = n3693 ^ n243 ^ 1'b0 ;
  assign n7519 = n4362 ^ n3749 ^ 1'b0 ;
  assign n7520 = n585 & n7519 ;
  assign n7521 = n2927 & n4354 ;
  assign n7522 = ~n7520 & n7521 ;
  assign n7523 = n7518 & ~n7522 ;
  assign n7524 = n7523 ^ x18 ^ 1'b0 ;
  assign n7525 = n335 & ~n3856 ;
  assign n7526 = n3552 & n7525 ;
  assign n7527 = n7526 ^ n6729 ^ n3651 ;
  assign n7528 = n7527 ^ n4075 ^ 1'b0 ;
  assign n7529 = n1065 & n3341 ;
  assign n7530 = n1327 & n7529 ;
  assign n7531 = n7530 ^ n2890 ^ 1'b0 ;
  assign n7532 = ~x97 & n7531 ;
  assign n7533 = ~n465 & n928 ;
  assign n7534 = n7533 ^ n497 ^ 1'b0 ;
  assign n7535 = n7534 ^ n2828 ^ 1'b0 ;
  assign n7536 = n7278 & n7535 ;
  assign n7537 = n1622 & n7536 ;
  assign n7538 = n3560 & ~n7537 ;
  assign n7539 = n307 & ~n3319 ;
  assign n7540 = ~n2094 & n7539 ;
  assign n7541 = n5111 & ~n7540 ;
  assign n7552 = ( ~n436 & n1929 ) | ( ~n436 & n2498 ) | ( n1929 & n2498 ) ;
  assign n7551 = ( x78 & n2682 ) | ( x78 & ~n3461 ) | ( n2682 & ~n3461 ) ;
  assign n7548 = n7207 ^ n4356 ^ n866 ;
  assign n7547 = ~n2390 & n3615 ;
  assign n7549 = n7548 ^ n7547 ^ 1'b0 ;
  assign n7545 = n3853 & ~n3986 ;
  assign n7542 = n6034 ^ n1856 ^ 1'b0 ;
  assign n7543 = n2870 | n7542 ;
  assign n7544 = n5818 & ~n7543 ;
  assign n7546 = n7545 ^ n7544 ^ 1'b0 ;
  assign n7550 = n7549 ^ n7546 ^ n5192 ;
  assign n7553 = n7552 ^ n7551 ^ n7550 ;
  assign n7556 = n732 & ~n5162 ;
  assign n7557 = n7556 ^ n2183 ^ 1'b0 ;
  assign n7554 = n1501 & ~n1589 ;
  assign n7555 = n2363 & n7554 ;
  assign n7558 = n7557 ^ n7555 ^ 1'b0 ;
  assign n7559 = ~n3972 & n4402 ;
  assign n7560 = n7559 ^ n677 ^ 1'b0 ;
  assign n7561 = n7560 ^ n1586 ^ 1'b0 ;
  assign n7562 = n7561 ^ n5858 ^ 1'b0 ;
  assign n7563 = n415 | n781 ;
  assign n7564 = n4024 & n7563 ;
  assign n7565 = ( n3981 & n6652 ) | ( n3981 & n7564 ) | ( n6652 & n7564 ) ;
  assign n7566 = n4384 & n7565 ;
  assign n7567 = n3943 & ~n6550 ;
  assign n7570 = n1292 ^ n1261 ^ 1'b0 ;
  assign n7571 = ( ~n2502 & n4505 ) | ( ~n2502 & n7570 ) | ( n4505 & n7570 ) ;
  assign n7568 = n6087 ^ n2660 ^ n1247 ;
  assign n7569 = n175 & n7568 ;
  assign n7572 = n7571 ^ n7569 ^ 1'b0 ;
  assign n7573 = ( n1179 & n6363 ) | ( n1179 & n6865 ) | ( n6363 & n6865 ) ;
  assign n7574 = n7054 ^ n6845 ^ 1'b0 ;
  assign n7575 = n3212 | n4851 ;
  assign n7576 = n1894 & ~n6714 ;
  assign n7577 = n7576 ^ n3798 ^ 1'b0 ;
  assign n7578 = ( n5305 & ~n6475 ) | ( n5305 & n7577 ) | ( ~n6475 & n7577 ) ;
  assign n7579 = n1470 & ~n2746 ;
  assign n7580 = ~n5822 & n7579 ;
  assign n7585 = n2738 & ~n3396 ;
  assign n7586 = n7585 ^ n6986 ^ 1'b0 ;
  assign n7584 = n1273 & n6376 ;
  assign n7587 = n7586 ^ n7584 ^ 1'b0 ;
  assign n7581 = n578 ^ x87 ^ 1'b0 ;
  assign n7582 = ~n2919 & n7581 ;
  assign n7583 = n7582 ^ n6903 ^ 1'b0 ;
  assign n7588 = n7587 ^ n7583 ^ 1'b0 ;
  assign n7589 = ~n3730 & n7588 ;
  assign n7590 = ( n908 & ~n1706 ) | ( n908 & n4787 ) | ( ~n1706 & n4787 ) ;
  assign n7591 = n7590 ^ n3822 ^ 1'b0 ;
  assign n7592 = x5 & ~n7591 ;
  assign n7593 = n7592 ^ n2552 ^ 1'b0 ;
  assign n7594 = n5106 | n6168 ;
  assign n7595 = ( n2062 & n7593 ) | ( n2062 & n7594 ) | ( n7593 & n7594 ) ;
  assign n7596 = n292 | n6885 ;
  assign n7597 = n2740 & n4609 ;
  assign n7598 = n2540 & n7597 ;
  assign n7599 = n2483 & ~n7598 ;
  assign n7600 = n7599 ^ n1162 ^ 1'b0 ;
  assign n7601 = n1470 | n7600 ;
  assign n7602 = n5335 | n7601 ;
  assign n7603 = ~n2976 & n5163 ;
  assign n7604 = ~n7545 & n7603 ;
  assign n7605 = ~n138 & n5490 ;
  assign n7606 = n7605 ^ n4062 ^ n2051 ;
  assign n7607 = ( n523 & n2016 ) | ( n523 & ~n7606 ) | ( n2016 & ~n7606 ) ;
  assign n7611 = n5262 ^ n1259 ^ 1'b0 ;
  assign n7612 = n3674 | n7611 ;
  assign n7609 = n459 & ~n2833 ;
  assign n7610 = n7609 ^ n1381 ^ 1'b0 ;
  assign n7613 = n7612 ^ n7610 ^ n5510 ;
  assign n7608 = n4885 & ~n5410 ;
  assign n7614 = n7613 ^ n7608 ^ 1'b0 ;
  assign n7615 = n7614 ^ n4995 ^ 1'b0 ;
  assign n7616 = n3686 & n7615 ;
  assign n7617 = ( n1076 & n5376 ) | ( n1076 & n6115 ) | ( n5376 & n6115 ) ;
  assign n7618 = n2040 & ~n3408 ;
  assign n7619 = n1058 & n7618 ;
  assign n7620 = ~n7617 & n7619 ;
  assign n7621 = n2290 ^ n2002 ^ 1'b0 ;
  assign n7622 = n1802 & ~n7621 ;
  assign n7626 = n2706 ^ n248 ^ 1'b0 ;
  assign n7627 = n207 & n7626 ;
  assign n7623 = n788 & n2647 ;
  assign n7624 = n7623 ^ n2597 ^ 1'b0 ;
  assign n7625 = ~n5942 & n7624 ;
  assign n7628 = n7627 ^ n7625 ^ 1'b0 ;
  assign n7629 = n4480 | n7628 ;
  assign n7630 = n4308 ^ n3099 ^ 1'b0 ;
  assign n7631 = n3237 & ~n7630 ;
  assign n7632 = n7631 ^ n2258 ^ 1'b0 ;
  assign n7634 = n2514 ^ n2467 ^ 1'b0 ;
  assign n7635 = n7634 ^ n2365 ^ 1'b0 ;
  assign n7633 = n1942 | n5473 ;
  assign n7636 = n7635 ^ n7633 ^ 1'b0 ;
  assign n7639 = n3971 ^ x41 ^ 1'b0 ;
  assign n7640 = n1996 & ~n7639 ;
  assign n7637 = x8 & n1067 ;
  assign n7638 = ~n5230 & n7637 ;
  assign n7641 = n7640 ^ n7638 ^ n5988 ;
  assign n7642 = n4300 ^ x126 ^ 1'b0 ;
  assign n7643 = n1892 ^ n944 ^ n646 ;
  assign n7644 = n5555 & ~n7643 ;
  assign n7645 = n3856 ^ n163 ^ 1'b0 ;
  assign n7646 = n7645 ^ n7240 ^ x70 ;
  assign n7647 = n2182 & n5948 ;
  assign n7648 = n7647 ^ n7537 ^ 1'b0 ;
  assign n7649 = n1972 ^ n331 ^ 1'b0 ;
  assign n7650 = ( n4756 & n5244 ) | ( n4756 & ~n7649 ) | ( n5244 & ~n7649 ) ;
  assign n7651 = n7650 ^ n6223 ^ 1'b0 ;
  assign n7652 = ~n5382 & n7651 ;
  assign n7653 = n4660 & n5349 ;
  assign n7654 = ~n1386 & n7653 ;
  assign n7655 = ( ~n1137 & n3314 ) | ( ~n1137 & n7525 ) | ( n3314 & n7525 ) ;
  assign n7656 = ( ~n3789 & n4431 ) | ( ~n3789 & n4437 ) | ( n4431 & n4437 ) ;
  assign n7657 = ( ~n1168 & n2846 ) | ( ~n1168 & n7656 ) | ( n2846 & n7656 ) ;
  assign n7658 = n7657 ^ n1882 ^ 1'b0 ;
  assign n7659 = n2014 | n7658 ;
  assign n7660 = n1365 & ~n2161 ;
  assign n7661 = n756 & n7660 ;
  assign n7662 = n7661 ^ n2884 ^ 1'b0 ;
  assign n7663 = n7662 ^ n6833 ^ 1'b0 ;
  assign n7664 = n551 | n6149 ;
  assign n7665 = x8 | n7664 ;
  assign n7666 = n3371 & n3707 ;
  assign n7667 = n3447 & n7666 ;
  assign n7668 = n4753 & ~n7667 ;
  assign n7669 = ( x103 & ~n2032 ) | ( x103 & n2999 ) | ( ~n2032 & n2999 ) ;
  assign n7670 = ( x9 & n829 ) | ( x9 & ~n1723 ) | ( n829 & ~n1723 ) ;
  assign n7671 = n2976 & n7670 ;
  assign n7672 = n6868 ^ n3538 ^ 1'b0 ;
  assign n7673 = n4739 ^ n2570 ^ 1'b0 ;
  assign n7674 = ~n2329 & n7673 ;
  assign n7675 = n1589 & n7495 ;
  assign n7676 = n6339 ^ n484 ^ 1'b0 ;
  assign n7677 = n6163 ^ n1639 ^ 1'b0 ;
  assign n7678 = n7676 & n7677 ;
  assign n7679 = ( ~n4561 & n6816 ) | ( ~n4561 & n7678 ) | ( n6816 & n7678 ) ;
  assign n7680 = n3378 | n5602 ;
  assign n7681 = n3349 | n7680 ;
  assign n7682 = n3933 & ~n7681 ;
  assign n7683 = n2108 | n3410 ;
  assign n7684 = n5041 | n6596 ;
  assign n7685 = n7683 | n7684 ;
  assign n7686 = ( ~n1485 & n4430 ) | ( ~n1485 & n5355 ) | ( n4430 & n5355 ) ;
  assign n7687 = n4521 | n6304 ;
  assign n7692 = n4581 ^ n2237 ^ n1511 ;
  assign n7688 = ~n2355 & n3423 ;
  assign n7689 = n7688 ^ n977 ^ 1'b0 ;
  assign n7690 = n3628 & ~n7689 ;
  assign n7691 = n7690 ^ n1921 ^ 1'b0 ;
  assign n7693 = n7692 ^ n7691 ^ 1'b0 ;
  assign n7694 = n1794 & ~n7693 ;
  assign n7695 = n1788 ^ n1248 ^ 1'b0 ;
  assign n7696 = ( n1402 & n2772 ) | ( n1402 & n7695 ) | ( n2772 & n7695 ) ;
  assign n7697 = n3830 ^ n970 ^ 1'b0 ;
  assign n7699 = ( n3879 & n4106 ) | ( n3879 & ~n5163 ) | ( n4106 & ~n5163 ) ;
  assign n7700 = n5258 & ~n7699 ;
  assign n7701 = n7700 ^ n2383 ^ 1'b0 ;
  assign n7702 = n7701 ^ n7216 ^ 1'b0 ;
  assign n7698 = n737 & ~n2228 ;
  assign n7703 = n7702 ^ n7698 ^ 1'b0 ;
  assign n7704 = n5328 ^ n4601 ^ n2956 ;
  assign n7705 = ~n4652 & n7704 ;
  assign n7706 = n7705 ^ n1282 ^ 1'b0 ;
  assign n7707 = n7706 ^ n6861 ^ 1'b0 ;
  assign n7708 = ( n2204 & n2375 ) | ( n2204 & ~n6852 ) | ( n2375 & ~n6852 ) ;
  assign n7709 = ( ~n1946 & n2318 ) | ( ~n1946 & n6659 ) | ( n2318 & n6659 ) ;
  assign n7710 = n2597 ^ n2100 ^ 1'b0 ;
  assign n7711 = n1073 | n7710 ;
  assign n7712 = n344 | n7711 ;
  assign n7713 = n7709 & ~n7712 ;
  assign n7714 = n2353 ^ x91 ^ 1'b0 ;
  assign n7715 = x42 & ~n7714 ;
  assign n7716 = n950 ^ n354 ^ 1'b0 ;
  assign n7717 = n7716 ^ n3364 ^ 1'b0 ;
  assign n7718 = n7715 | n7717 ;
  assign n7719 = n7718 ^ n3398 ^ 1'b0 ;
  assign n7721 = ~n2952 & n4495 ;
  assign n7722 = ~n1388 & n7721 ;
  assign n7723 = ~n2895 & n7722 ;
  assign n7720 = n1515 & n1823 ;
  assign n7724 = n7723 ^ n7720 ^ 1'b0 ;
  assign n7725 = ( n1129 & n3009 ) | ( n1129 & ~n3563 ) | ( n3009 & ~n3563 ) ;
  assign n7726 = n7725 ^ n888 ^ 1'b0 ;
  assign n7727 = n4927 | n7726 ;
  assign n7728 = n4679 & ~n7040 ;
  assign n7729 = n2903 & n7728 ;
  assign n7730 = n6668 ^ n4797 ^ 1'b0 ;
  assign n7732 = n4870 & ~n5783 ;
  assign n7733 = n7732 ^ n1215 ^ 1'b0 ;
  assign n7731 = n131 & ~n2371 ;
  assign n7734 = n7733 ^ n7731 ^ 1'b0 ;
  assign n7735 = ( n727 & n1418 ) | ( n727 & n3100 ) | ( n1418 & n3100 ) ;
  assign n7736 = n411 | n7735 ;
  assign n7739 = ( n2183 & n3624 ) | ( n2183 & ~n3629 ) | ( n3624 & ~n3629 ) ;
  assign n7737 = x108 | n2668 ;
  assign n7738 = n7737 ^ n1084 ^ n593 ;
  assign n7740 = n7739 ^ n7738 ^ n7475 ;
  assign n7741 = n7658 ^ n5167 ^ 1'b0 ;
  assign n7742 = ( ~x50 & n4710 ) | ( ~x50 & n6200 ) | ( n4710 & n6200 ) ;
  assign n7743 = n1750 & n3289 ;
  assign n7744 = n7743 ^ n6994 ^ 1'b0 ;
  assign n7745 = n7744 ^ n5347 ^ n2021 ;
  assign n7746 = x30 & ~n3878 ;
  assign n7747 = ~n3111 & n7746 ;
  assign n7748 = n7697 & n7747 ;
  assign n7753 = n3507 & n5438 ;
  assign n7751 = n1106 | n1455 ;
  assign n7752 = n7751 ^ n1049 ^ 1'b0 ;
  assign n7749 = n205 & n2014 ;
  assign n7750 = ( n2221 & n2965 ) | ( n2221 & n7749 ) | ( n2965 & n7749 ) ;
  assign n7754 = n7753 ^ n7752 ^ n7750 ;
  assign n7755 = ~n5883 & n6752 ;
  assign n7756 = n7755 ^ n4069 ^ 1'b0 ;
  assign n7757 = n7756 ^ n3594 ^ 1'b0 ;
  assign n7758 = ~n4015 & n7757 ;
  assign n7759 = n4519 & n5102 ;
  assign n7760 = n1552 & n7759 ;
  assign n7761 = n7760 ^ n2200 ^ 1'b0 ;
  assign n7762 = n7758 & ~n7761 ;
  assign n7763 = n136 | n5752 ;
  assign n7764 = n7763 ^ n7512 ^ 1'b0 ;
  assign n7765 = ~n3694 & n7764 ;
  assign n7766 = n4632 ^ n4401 ^ n2527 ;
  assign n7767 = n7766 ^ n4440 ^ 1'b0 ;
  assign n7768 = n1508 & n5421 ;
  assign n7769 = n6092 ^ n3221 ^ n2145 ;
  assign n7770 = ~n911 & n3436 ;
  assign n7771 = n7770 ^ n6303 ^ 1'b0 ;
  assign n7772 = ~n3364 & n7771 ;
  assign n7773 = ~n7769 & n7772 ;
  assign n7774 = ~n6258 & n7773 ;
  assign n7775 = ( n2144 & n2349 ) | ( n2144 & n3426 ) | ( n2349 & n3426 ) ;
  assign n7776 = ~n4312 & n7775 ;
  assign n7777 = n7776 ^ n7377 ^ 1'b0 ;
  assign n7778 = n5881 ^ n4099 ^ n3925 ;
  assign n7788 = n7715 ^ n2391 ^ 1'b0 ;
  assign n7789 = ( ~n461 & n3342 ) | ( ~n461 & n7788 ) | ( n3342 & n7788 ) ;
  assign n7790 = ( n5535 & ~n6798 ) | ( n5535 & n7789 ) | ( ~n6798 & n7789 ) ;
  assign n7779 = n4554 ^ n3250 ^ 1'b0 ;
  assign n7780 = ~n2530 & n7779 ;
  assign n7781 = n1902 & n5605 ;
  assign n7782 = n7780 & n7781 ;
  assign n7783 = n2755 | n2971 ;
  assign n7784 = n7783 ^ n3747 ^ 1'b0 ;
  assign n7785 = ( n3681 & n6045 ) | ( n3681 & ~n7784 ) | ( n6045 & ~n7784 ) ;
  assign n7786 = n7785 ^ n7543 ^ 1'b0 ;
  assign n7787 = n7782 & n7786 ;
  assign n7791 = n7790 ^ n7787 ^ n4461 ;
  assign n7794 = n157 & ~n6125 ;
  assign n7792 = n4871 ^ n320 ^ 1'b0 ;
  assign n7793 = n7733 & n7792 ;
  assign n7795 = n7794 ^ n7793 ^ n3864 ;
  assign n7796 = x82 & ~x112 ;
  assign n7797 = ~n2763 & n3503 ;
  assign n7798 = n7796 & n7797 ;
  assign n7799 = n7485 ^ n378 ^ 1'b0 ;
  assign n7800 = n2606 & n7799 ;
  assign n7801 = n2705 & n7598 ;
  assign n7802 = n3038 & ~n6131 ;
  assign n7803 = n7801 & n7802 ;
  assign n7804 = ( n3718 & n5205 ) | ( n3718 & n7803 ) | ( n5205 & n7803 ) ;
  assign n7805 = ~n398 & n6496 ;
  assign n7806 = n3034 ^ n1905 ^ 1'b0 ;
  assign n7807 = n3796 & ~n7806 ;
  assign n7808 = ( n3102 & n3371 ) | ( n3102 & ~n7807 ) | ( n3371 & ~n7807 ) ;
  assign n7809 = n3391 & ~n6783 ;
  assign n7810 = n7809 ^ x65 ^ 1'b0 ;
  assign n7811 = ~n351 & n7810 ;
  assign n7812 = n5565 & n7614 ;
  assign n7813 = n7812 ^ n7295 ^ 1'b0 ;
  assign n7814 = n697 ^ x30 ^ 1'b0 ;
  assign n7815 = ( ~n5390 & n5615 ) | ( ~n5390 & n7814 ) | ( n5615 & n7814 ) ;
  assign n7816 = n5599 & ~n6724 ;
  assign n7817 = n206 & ~n4667 ;
  assign n7818 = n7817 ^ n411 ^ 1'b0 ;
  assign n7823 = n6810 ^ n6169 ^ n2254 ;
  assign n7819 = n334 & n1311 ;
  assign n7820 = ~n2772 & n7819 ;
  assign n7821 = ( n2900 & n4397 ) | ( n2900 & n7820 ) | ( n4397 & n7820 ) ;
  assign n7822 = n7821 ^ n1622 ^ 1'b0 ;
  assign n7824 = n7823 ^ n7822 ^ 1'b0 ;
  assign n7825 = n4858 & n5102 ;
  assign n7826 = n7825 ^ n7277 ^ 1'b0 ;
  assign n7827 = ~n386 & n1655 ;
  assign n7828 = ~n2796 & n7827 ;
  assign n7829 = n5345 | n7828 ;
  assign n7830 = n7826 & n7829 ;
  assign n7831 = ~n5994 & n7830 ;
  assign n7832 = n7373 ^ n6529 ^ 1'b0 ;
  assign n7833 = n4821 ^ n4044 ^ 1'b0 ;
  assign n7836 = n1441 & ~n4826 ;
  assign n7837 = n2002 & n7836 ;
  assign n7834 = n737 & n2358 ;
  assign n7835 = n7834 ^ n7207 ^ x78 ;
  assign n7838 = n7837 ^ n7835 ^ 1'b0 ;
  assign n7839 = n2062 | n6500 ;
  assign n7840 = n389 & ~n7839 ;
  assign n7841 = n4792 & n7840 ;
  assign n7842 = ~n1867 & n6408 ;
  assign n7843 = n5416 ^ n4533 ^ 1'b0 ;
  assign n7844 = n4214 & ~n7843 ;
  assign n7845 = n2018 ^ n886 ^ 1'b0 ;
  assign n7846 = n7844 & ~n7845 ;
  assign n7847 = x43 & ~n1342 ;
  assign n7848 = n7847 ^ n3501 ^ 1'b0 ;
  assign n7849 = n6245 ^ n6111 ^ 1'b0 ;
  assign n7850 = n7848 & ~n7849 ;
  assign n7851 = x111 & n1538 ;
  assign n7852 = n893 & n7851 ;
  assign n7853 = n4785 & ~n5619 ;
  assign n7854 = n7853 ^ n6600 ^ 1'b0 ;
  assign n7855 = n7854 ^ n3128 ^ 1'b0 ;
  assign n7856 = n7852 | n7855 ;
  assign n7857 = n2774 & ~n5484 ;
  assign n7858 = n7857 ^ n7681 ^ 1'b0 ;
  assign n7859 = ( ~n3676 & n4443 ) | ( ~n3676 & n7858 ) | ( n4443 & n7858 ) ;
  assign n7860 = n6394 | n7859 ;
  assign n7861 = n2083 | n4605 ;
  assign n7862 = n990 | n3122 ;
  assign n7863 = n1719 & ~n7862 ;
  assign n7864 = n7863 ^ n2740 ^ 1'b0 ;
  assign n7865 = n1438 & ~n7864 ;
  assign n7866 = n2026 & n7865 ;
  assign n7867 = n7854 & n7866 ;
  assign n7868 = n2719 ^ n635 ^ 1'b0 ;
  assign n7869 = n3310 & ~n7868 ;
  assign n7870 = n4346 ^ n3864 ^ 1'b0 ;
  assign n7871 = ~n2371 & n4761 ;
  assign n7872 = ~n7243 & n7871 ;
  assign n7873 = n7872 ^ n7428 ^ 1'b0 ;
  assign n7874 = n6730 ^ n5266 ^ n1706 ;
  assign n7876 = n1970 | n4160 ;
  assign n7877 = n3503 | n7876 ;
  assign n7875 = n1489 & ~n6649 ;
  assign n7878 = n7877 ^ n7875 ^ 1'b0 ;
  assign n7879 = n5078 ^ n4797 ^ 1'b0 ;
  assign n7880 = n1404 | n7879 ;
  assign n7881 = n7880 ^ n1150 ^ 1'b0 ;
  assign n7882 = ~n4645 & n7881 ;
  assign n7883 = ~n7878 & n7882 ;
  assign n7884 = n2228 & n7883 ;
  assign n7885 = n5740 ^ n4110 ^ 1'b0 ;
  assign n7886 = ~n300 & n7885 ;
  assign n7887 = n6986 & n7207 ;
  assign n7891 = n1633 & n5036 ;
  assign n7892 = n7891 ^ n4665 ^ 1'b0 ;
  assign n7893 = n2421 ^ n1104 ^ 1'b0 ;
  assign n7894 = ~n847 & n7893 ;
  assign n7895 = n4326 & n7894 ;
  assign n7896 = n4761 & n7895 ;
  assign n7897 = ~n7892 & n7896 ;
  assign n7888 = n1913 & ~n4580 ;
  assign n7889 = n422 & ~n7888 ;
  assign n7890 = ~n5660 & n7889 ;
  assign n7898 = n7897 ^ n7890 ^ n3421 ;
  assign n7899 = n7894 ^ n7474 ^ 1'b0 ;
  assign n7900 = n5559 | n7899 ;
  assign n7901 = n885 | n7900 ;
  assign n7902 = n7649 & ~n7901 ;
  assign n7903 = n4263 | n7902 ;
  assign n7904 = n7903 ^ n1116 ^ 1'b0 ;
  assign n7906 = n5262 ^ n4321 ^ n569 ;
  assign n7905 = ~n4908 & n5789 ;
  assign n7907 = n7906 ^ n7905 ^ 1'b0 ;
  assign n7908 = n7904 & n7907 ;
  assign n7909 = ~n1170 & n5653 ;
  assign n7910 = n7909 ^ n314 ^ 1'b0 ;
  assign n7911 = n2181 | n2791 ;
  assign n7912 = ~n7910 & n7911 ;
  assign n7913 = n2771 | n4422 ;
  assign n7914 = n7913 ^ n5823 ^ 1'b0 ;
  assign n7915 = n4733 ^ n4032 ^ 1'b0 ;
  assign n7916 = n927 | n7814 ;
  assign n7917 = n5276 & ~n7916 ;
  assign n7918 = n7801 ^ n2252 ^ n1135 ;
  assign n7919 = n7918 ^ n3286 ^ 1'b0 ;
  assign n7922 = n3265 ^ n154 ^ 1'b0 ;
  assign n7923 = n809 & n7922 ;
  assign n7920 = ( n1280 & ~n3917 ) | ( n1280 & n4029 ) | ( ~n3917 & n4029 ) ;
  assign n7921 = n1684 | n7920 ;
  assign n7924 = n7923 ^ n7921 ^ 1'b0 ;
  assign n7925 = n1615 ^ n652 ^ 1'b0 ;
  assign n7926 = n7925 ^ n4347 ^ 1'b0 ;
  assign n7927 = n7924 & n7926 ;
  assign n7928 = n971 & ~n3830 ;
  assign n7929 = ( n293 & ~n934 ) | ( n293 & n7928 ) | ( ~n934 & n7928 ) ;
  assign n7930 = ~n749 & n7929 ;
  assign n7931 = n1287 | n5198 ;
  assign n7932 = n560 & ~n2772 ;
  assign n7933 = n7932 ^ n3852 ^ 1'b0 ;
  assign n7934 = n1682 | n7933 ;
  assign n7935 = n2974 & ~n7934 ;
  assign n7936 = ~n1067 & n4242 ;
  assign n7937 = n7936 ^ n6264 ^ n5864 ;
  assign n7938 = ( n231 & n1552 ) | ( n231 & n4856 ) | ( n1552 & n4856 ) ;
  assign n7939 = n5522 & ~n6603 ;
  assign n7940 = n7938 | n7939 ;
  assign n7941 = n5399 & ~n7940 ;
  assign n7942 = n7941 ^ n2930 ^ 1'b0 ;
  assign n7943 = n7869 | n7942 ;
  assign n7944 = n986 | n1545 ;
  assign n7945 = n7944 ^ n3597 ^ 1'b0 ;
  assign n7946 = n2496 & n7945 ;
  assign n7947 = ~n3279 & n7946 ;
  assign n7948 = n3871 | n5873 ;
  assign n7949 = n7948 ^ n3732 ^ 1'b0 ;
  assign n7950 = n3511 & ~n7949 ;
  assign n7951 = ( ~n140 & n3363 ) | ( ~n140 & n3688 ) | ( n3363 & n3688 ) ;
  assign n7952 = n3009 & ~n7951 ;
  assign n7953 = ( n686 & ~n2201 ) | ( n686 & n3324 ) | ( ~n2201 & n3324 ) ;
  assign n7954 = n7952 & n7953 ;
  assign n7955 = n6300 ^ n3822 ^ n1826 ;
  assign n7956 = ( ~n418 & n3211 ) | ( ~n418 & n5939 ) | ( n3211 & n5939 ) ;
  assign n7957 = n7956 ^ n2304 ^ x29 ;
  assign n7960 = n3267 ^ n1186 ^ 1'b0 ;
  assign n7961 = n4416 & ~n7960 ;
  assign n7962 = n7961 ^ n5841 ^ 1'b0 ;
  assign n7958 = n1637 ^ n133 ^ 1'b0 ;
  assign n7959 = n761 | n7958 ;
  assign n7963 = n7962 ^ n7959 ^ 1'b0 ;
  assign n7964 = ( n986 & n1947 ) | ( n986 & ~n6605 ) | ( n1947 & ~n6605 ) ;
  assign n7965 = n2939 ^ n1250 ^ 1'b0 ;
  assign n7966 = ( ~n925 & n6143 ) | ( ~n925 & n7965 ) | ( n6143 & n7965 ) ;
  assign n7967 = n7964 & n7966 ;
  assign n7968 = n7967 ^ n6669 ^ 1'b0 ;
  assign n7969 = n5587 | n7237 ;
  assign n7970 = n1353 & ~n7969 ;
  assign n7971 = n1234 | n2612 ;
  assign n7973 = n5317 ^ n1104 ^ n182 ;
  assign n7974 = ( n885 & n1752 ) | ( n885 & ~n7973 ) | ( n1752 & ~n7973 ) ;
  assign n7972 = n1708 | n1914 ;
  assign n7975 = n7974 ^ n7972 ^ 1'b0 ;
  assign n7976 = ( n1581 & ~n2203 ) | ( n1581 & n5822 ) | ( ~n2203 & n5822 ) ;
  assign n7977 = ( ~n445 & n2580 ) | ( ~n445 & n7976 ) | ( n2580 & n7976 ) ;
  assign n7978 = n7977 ^ n3239 ^ 1'b0 ;
  assign n7979 = n7978 ^ n4342 ^ 1'b0 ;
  assign n7980 = ~n2371 & n6503 ;
  assign n7981 = n7980 ^ n6576 ^ 1'b0 ;
  assign n7982 = n3106 ^ n2488 ^ 1'b0 ;
  assign n7983 = n2660 | n7982 ;
  assign n7984 = n7983 ^ n4340 ^ 1'b0 ;
  assign n7985 = ~n1873 & n2712 ;
  assign n7986 = n7985 ^ n7809 ^ n4927 ;
  assign n7987 = ~n3696 & n7952 ;
  assign n7988 = n459 & n3920 ;
  assign n7989 = n4631 & n7988 ;
  assign n7990 = n4221 | n7989 ;
  assign n7995 = ( n846 & n2855 ) | ( n846 & ~n4824 ) | ( n2855 & ~n4824 ) ;
  assign n7996 = n3679 ^ n3375 ^ 1'b0 ;
  assign n7997 = ( n4688 & ~n7995 ) | ( n4688 & n7996 ) | ( ~n7995 & n7996 ) ;
  assign n7991 = n1244 & n3240 ;
  assign n7992 = ~n7370 & n7991 ;
  assign n7993 = n2074 | n7992 ;
  assign n7994 = n692 & ~n7993 ;
  assign n7998 = n7997 ^ n7994 ^ n1721 ;
  assign n7999 = ~n3005 & n7998 ;
  assign n8000 = n5780 | n7182 ;
  assign n8001 = n8000 ^ n2817 ^ 1'b0 ;
  assign n8002 = ( n1506 & n2188 ) | ( n1506 & ~n4144 ) | ( n2188 & ~n4144 ) ;
  assign n8003 = n1971 & ~n8002 ;
  assign n8004 = n8003 ^ n1710 ^ 1'b0 ;
  assign n8005 = n8004 ^ n5331 ^ 1'b0 ;
  assign n8006 = n3583 & n6663 ;
  assign n8007 = n3965 ^ n2349 ^ n1768 ;
  assign n8008 = n5531 ^ n1501 ^ 1'b0 ;
  assign n8009 = n8007 & ~n8008 ;
  assign n8010 = n8009 ^ n7917 ^ n480 ;
  assign n8011 = n6452 & n7785 ;
  assign n8012 = n5598 & n8011 ;
  assign n8013 = n2590 | n3187 ;
  assign n8014 = n8013 ^ n6849 ^ 1'b0 ;
  assign n8015 = n5643 ^ n2245 ^ 1'b0 ;
  assign n8016 = n2771 | n8015 ;
  assign n8017 = n1419 | n2931 ;
  assign n8018 = n4735 ^ n1696 ^ n1368 ;
  assign n8019 = ( n8016 & n8017 ) | ( n8016 & ~n8018 ) | ( n8017 & ~n8018 ) ;
  assign n8020 = ~n2678 & n3434 ;
  assign n8021 = n804 | n2499 ;
  assign n8022 = n8021 ^ n4895 ^ 1'b0 ;
  assign n8023 = n8022 ^ n4401 ^ 1'b0 ;
  assign n8024 = n3654 ^ n2139 ^ 1'b0 ;
  assign n8026 = n1034 | n1159 ;
  assign n8027 = n768 | n8026 ;
  assign n8025 = ~n2741 & n5671 ;
  assign n8028 = n8027 ^ n8025 ^ 1'b0 ;
  assign n8029 = ~n1305 & n3513 ;
  assign n8030 = n8028 & ~n8029 ;
  assign n8031 = n4634 ^ n1157 ^ 1'b0 ;
  assign n8032 = ( n6749 & ~n7110 ) | ( n6749 & n8031 ) | ( ~n7110 & n8031 ) ;
  assign n8033 = n7560 ^ n4795 ^ n936 ;
  assign n8034 = n1894 & ~n2854 ;
  assign n8035 = n3671 & n8034 ;
  assign n8036 = ( n3651 & n8033 ) | ( n3651 & n8035 ) | ( n8033 & n8035 ) ;
  assign n8037 = n8036 ^ n5305 ^ 1'b0 ;
  assign n8038 = ~n1854 & n8037 ;
  assign n8039 = n4124 | n8038 ;
  assign n8040 = n3794 ^ n1159 ^ 1'b0 ;
  assign n8041 = ( n617 & n1846 ) | ( n617 & n8040 ) | ( n1846 & n8040 ) ;
  assign n8042 = n7227 ^ n5001 ^ 1'b0 ;
  assign n8043 = n7462 | n8042 ;
  assign n8044 = n565 & ~n1686 ;
  assign n8045 = n8044 ^ n5096 ^ 1'b0 ;
  assign n8046 = n3865 ^ n1680 ^ 1'b0 ;
  assign n8047 = n3334 & n8046 ;
  assign n8048 = n354 & n8047 ;
  assign n8049 = ~n4588 & n8048 ;
  assign n8050 = n4891 ^ n1090 ^ 1'b0 ;
  assign n8051 = n6401 ^ n5164 ^ 1'b0 ;
  assign n8052 = ~n4425 & n8051 ;
  assign n8053 = n8052 ^ n5928 ^ 1'b0 ;
  assign n8054 = n8017 & n8053 ;
  assign n8055 = n1694 & ~n4564 ;
  assign n8056 = n8055 ^ n4885 ^ 1'b0 ;
  assign n8057 = n2051 | n8056 ;
  assign n8058 = n5851 | n8057 ;
  assign n8059 = n1386 & n2709 ;
  assign n8060 = ( n4733 & n5348 ) | ( n4733 & ~n8059 ) | ( n5348 & ~n8059 ) ;
  assign n8061 = ( n3095 & n5745 ) | ( n3095 & ~n8060 ) | ( n5745 & ~n8060 ) ;
  assign n8062 = n7924 ^ n6378 ^ 1'b0 ;
  assign n8064 = n1584 ^ n822 ^ 1'b0 ;
  assign n8065 = n8064 ^ n7982 ^ 1'b0 ;
  assign n8063 = n6379 ^ n1112 ^ 1'b0 ;
  assign n8066 = n8065 ^ n8063 ^ n4472 ;
  assign n8067 = ( n3896 & n5091 ) | ( n3896 & ~n7238 ) | ( n5091 & ~n7238 ) ;
  assign n8068 = ~n1898 & n8067 ;
  assign n8069 = n8068 ^ n2118 ^ 1'b0 ;
  assign n8070 = n1556 & ~n6746 ;
  assign n8071 = n1561 & n8070 ;
  assign n8072 = n8071 ^ n5734 ^ 1'b0 ;
  assign n8073 = n8069 & ~n8072 ;
  assign n8075 = n3402 ^ x96 ^ 1'b0 ;
  assign n8074 = n1700 & ~n3060 ;
  assign n8076 = n8075 ^ n8074 ^ 1'b0 ;
  assign n8077 = ~n2758 & n5966 ;
  assign n8078 = n8077 ^ n4227 ^ 1'b0 ;
  assign n8079 = n8078 ^ n4580 ^ 1'b0 ;
  assign n8080 = n6914 ^ n5092 ^ 1'b0 ;
  assign n8081 = ~n1739 & n8080 ;
  assign n8082 = n1643 ^ n1029 ^ n916 ;
  assign n8083 = ~n1582 & n8082 ;
  assign n8084 = n8083 ^ n2140 ^ 1'b0 ;
  assign n8085 = n5315 ^ n5141 ^ 1'b0 ;
  assign n8086 = n374 | n8085 ;
  assign n8087 = n2044 & ~n8086 ;
  assign n8088 = ~n8084 & n8087 ;
  assign n8089 = ~n979 & n6486 ;
  assign n8090 = ( ~n1371 & n5033 ) | ( ~n1371 & n8089 ) | ( n5033 & n8089 ) ;
  assign n8091 = n429 & n8090 ;
  assign n8092 = ~n3688 & n8091 ;
  assign n8094 = n2609 ^ n1850 ^ 1'b0 ;
  assign n8095 = ~n2233 & n8094 ;
  assign n8093 = n3814 ^ n1539 ^ n608 ;
  assign n8096 = n8095 ^ n8093 ^ n3024 ;
  assign n8097 = n2156 ^ n1259 ^ 1'b0 ;
  assign n8098 = n8097 ^ n484 ^ 1'b0 ;
  assign n8099 = n1992 | n8098 ;
  assign n8100 = n8099 ^ n739 ^ 1'b0 ;
  assign n8101 = ~n3245 & n8100 ;
  assign n8102 = ( n3466 & n4033 ) | ( n3466 & ~n7598 ) | ( n4033 & ~n7598 ) ;
  assign n8103 = n8102 ^ n954 ^ 1'b0 ;
  assign n8104 = n8101 & n8103 ;
  assign n8105 = n8104 ^ n1075 ^ 1'b0 ;
  assign n8106 = ~n2224 & n8105 ;
  assign n8107 = n2283 & n5017 ;
  assign n8108 = n8107 ^ n4095 ^ 1'b0 ;
  assign n8109 = n8108 ^ n688 ^ 1'b0 ;
  assign n8110 = ~n1577 & n8109 ;
  assign n8111 = n3429 | n4184 ;
  assign n8112 = n4281 | n4798 ;
  assign n8113 = x122 & n8112 ;
  assign n8114 = n5643 ^ n327 ^ 1'b0 ;
  assign n8115 = n8114 ^ n5306 ^ 1'b0 ;
  assign n8116 = ~n2904 & n8115 ;
  assign n8117 = n8116 ^ n3916 ^ n1706 ;
  assign n8118 = n168 & ~n7356 ;
  assign n8119 = ( n2715 & ~n8117 ) | ( n2715 & n8118 ) | ( ~n8117 & n8118 ) ;
  assign n8120 = n3130 & n8119 ;
  assign n8121 = n2962 & ~n3836 ;
  assign n8122 = ( n1262 & n1803 ) | ( n1262 & ~n8121 ) | ( n1803 & ~n8121 ) ;
  assign n8135 = n6064 ^ n824 ^ 1'b0 ;
  assign n8128 = n2487 ^ n2353 ^ 1'b0 ;
  assign n8129 = n3691 | n8128 ;
  assign n8130 = ~n1582 & n2854 ;
  assign n8131 = n4331 & ~n8130 ;
  assign n8132 = ~n3271 & n8131 ;
  assign n8133 = ~n5572 & n8132 ;
  assign n8134 = n8129 | n8133 ;
  assign n8136 = n8135 ^ n8134 ^ 1'b0 ;
  assign n8126 = n1582 | n7135 ;
  assign n8123 = ( n1230 & n3423 ) | ( n1230 & n3817 ) | ( n3423 & n3817 ) ;
  assign n8124 = ~n2929 & n8123 ;
  assign n8125 = n2976 & n8124 ;
  assign n8127 = n8126 ^ n8125 ^ n334 ;
  assign n8137 = n8136 ^ n8127 ^ 1'b0 ;
  assign n8138 = n1552 & n3813 ;
  assign n8139 = ~n1495 & n3533 ;
  assign n8140 = n7400 | n8139 ;
  assign n8141 = n2879 ^ n654 ^ 1'b0 ;
  assign n8142 = n8140 | n8141 ;
  assign n8143 = n599 | n1594 ;
  assign n8144 = n3809 ^ n1483 ^ n755 ;
  assign n8145 = ( n434 & n6684 ) | ( n434 & n8144 ) | ( n6684 & n8144 ) ;
  assign n8146 = n8145 ^ n1022 ^ 1'b0 ;
  assign n8147 = n4376 ^ n2312 ^ n214 ;
  assign n8148 = n5951 & n6228 ;
  assign n8149 = n8148 ^ n1874 ^ 1'b0 ;
  assign n8150 = ( n2014 & n3741 ) | ( n2014 & n5214 ) | ( n3741 & n5214 ) ;
  assign n8151 = ( n1785 & n2272 ) | ( n1785 & n2657 ) | ( n2272 & n2657 ) ;
  assign n8152 = n1986 & ~n8151 ;
  assign n8153 = n8152 ^ n2819 ^ 1'b0 ;
  assign n8154 = ( n4037 & ~n4096 ) | ( n4037 & n8153 ) | ( ~n4096 & n8153 ) ;
  assign n8155 = n644 & ~n3561 ;
  assign n8156 = n8155 ^ n1617 ^ 1'b0 ;
  assign n8157 = n6040 & n8156 ;
  assign n8162 = n3625 ^ n3245 ^ 1'b0 ;
  assign n8163 = n4294 & ~n8162 ;
  assign n8158 = n8114 ^ n855 ^ 1'b0 ;
  assign n8159 = n885 | n1593 ;
  assign n8160 = ( n140 & n2598 ) | ( n140 & n8159 ) | ( n2598 & n8159 ) ;
  assign n8161 = ( n915 & ~n8158 ) | ( n915 & n8160 ) | ( ~n8158 & n8160 ) ;
  assign n8164 = n8163 ^ n8161 ^ n7785 ;
  assign n8165 = n5355 ^ x69 ^ 1'b0 ;
  assign n8166 = n8165 ^ n6527 ^ n6437 ;
  assign n8167 = n8164 | n8166 ;
  assign n8170 = ~n3591 & n4824 ;
  assign n8171 = n1238 | n1428 ;
  assign n8172 = n8170 & ~n8171 ;
  assign n8168 = ~n4554 & n5207 ;
  assign n8169 = n8168 ^ n2527 ^ 1'b0 ;
  assign n8173 = n8172 ^ n8169 ^ 1'b0 ;
  assign n8174 = n7520 ^ n138 ^ x15 ;
  assign n8175 = n8174 ^ n6686 ^ 1'b0 ;
  assign n8176 = ~n1704 & n8175 ;
  assign n8177 = n800 ^ x43 ^ 1'b0 ;
  assign n8178 = n819 & ~n8177 ;
  assign n8179 = n719 | n1990 ;
  assign n8180 = n608 | n8179 ;
  assign n8181 = n8180 ^ n138 ^ 1'b0 ;
  assign n8182 = n8181 ^ n7005 ^ 1'b0 ;
  assign n8183 = n3525 ^ n2965 ^ n1160 ;
  assign n8184 = ( n1542 & ~n1602 ) | ( n1542 & n3749 ) | ( ~n1602 & n3749 ) ;
  assign n8185 = ( n2449 & ~n4580 ) | ( n2449 & n7570 ) | ( ~n4580 & n7570 ) ;
  assign n8186 = n8185 ^ n7817 ^ 1'b0 ;
  assign n8187 = n8186 ^ n2902 ^ n1170 ;
  assign n8188 = n370 & n7260 ;
  assign n8189 = n1565 ^ n1251 ^ 1'b0 ;
  assign n8190 = n4563 | n8189 ;
  assign n8191 = n4445 & ~n7525 ;
  assign n8192 = n2690 & n8191 ;
  assign n8193 = n8192 ^ n5403 ^ x23 ;
  assign n8194 = n3656 ^ n1621 ^ n397 ;
  assign n8195 = n3926 | n8194 ;
  assign n8196 = n1365 | n8195 ;
  assign n8197 = n8193 & ~n8196 ;
  assign n8199 = n6803 ^ n2451 ^ 1'b0 ;
  assign n8200 = n8199 ^ n1666 ^ 1'b0 ;
  assign n8198 = ( n1865 & ~n3735 ) | ( n1865 & n6301 ) | ( ~n3735 & n6301 ) ;
  assign n8201 = n8200 ^ n8198 ^ 1'b0 ;
  assign n8202 = n8201 ^ n6267 ^ n2315 ;
  assign n8204 = n950 & ~n1179 ;
  assign n8203 = n746 & ~n3792 ;
  assign n8205 = n8204 ^ n8203 ^ 1'b0 ;
  assign n8206 = n1666 & ~n8205 ;
  assign n8207 = n7821 & n8206 ;
  assign n8212 = n1696 ^ n158 ^ 1'b0 ;
  assign n8213 = ( ~n530 & n7477 ) | ( ~n530 & n8212 ) | ( n7477 & n8212 ) ;
  assign n8208 = n434 | n1523 ;
  assign n8209 = x17 | n8208 ;
  assign n8210 = n8209 ^ n2377 ^ 1'b0 ;
  assign n8211 = n7038 | n8210 ;
  assign n8214 = n8213 ^ n8211 ^ 1'b0 ;
  assign n8215 = n252 & n882 ;
  assign n8216 = ~n3160 & n8215 ;
  assign n8217 = ( ~n838 & n3933 ) | ( ~n838 & n8216 ) | ( n3933 & n8216 ) ;
  assign n8218 = ( n143 & ~n6691 ) | ( n143 & n8217 ) | ( ~n6691 & n8217 ) ;
  assign n8219 = ( n1190 & n5072 ) | ( n1190 & n8218 ) | ( n5072 & n8218 ) ;
  assign n8220 = n4180 ^ n1324 ^ 1'b0 ;
  assign n8221 = n194 & n8220 ;
  assign n8222 = n1832 & n8058 ;
  assign n8223 = n1020 & ~n3255 ;
  assign n8224 = ~n2425 & n8223 ;
  assign n8225 = ~n3391 & n8224 ;
  assign n8226 = n7865 ^ n3158 ^ 1'b0 ;
  assign n8227 = n8226 ^ n3599 ^ 1'b0 ;
  assign n8229 = n6758 ^ n2056 ^ 1'b0 ;
  assign n8228 = n765 & ~n2469 ;
  assign n8230 = n8229 ^ n8228 ^ 1'b0 ;
  assign n8231 = ( n970 & n2242 ) | ( n970 & ~n8230 ) | ( n2242 & ~n8230 ) ;
  assign n8232 = ~n2637 & n8231 ;
  assign n8233 = n8232 ^ n5878 ^ n4597 ;
  assign n8234 = ( n1973 & n4926 ) | ( n1973 & ~n5480 ) | ( n4926 & ~n5480 ) ;
  assign n8235 = n1544 ^ n982 ^ 1'b0 ;
  assign n8236 = n711 | n8235 ;
  assign n8237 = ( n456 & n2787 ) | ( n456 & n8236 ) | ( n2787 & n8236 ) ;
  assign n8238 = n173 | n4181 ;
  assign n8239 = n8237 & ~n8238 ;
  assign n8240 = ( ~x60 & n2086 ) | ( ~x60 & n2726 ) | ( n2086 & n2726 ) ;
  assign n8241 = n3103 ^ n909 ^ 1'b0 ;
  assign n8242 = n6550 & n8241 ;
  assign n8243 = n8240 & n8242 ;
  assign n8244 = n5670 ^ n3766 ^ 1'b0 ;
  assign n8245 = n1049 & n8244 ;
  assign n8246 = n3149 ^ n1626 ^ 1'b0 ;
  assign n8247 = n7077 ^ n1937 ^ 1'b0 ;
  assign n8248 = ~n3854 & n8247 ;
  assign n8249 = n3173 ^ n1249 ^ 1'b0 ;
  assign n8250 = n627 | n8249 ;
  assign n8251 = n1431 & n3523 ;
  assign n8252 = n8251 ^ n2060 ^ 1'b0 ;
  assign n8255 = n900 ^ n565 ^ 1'b0 ;
  assign n8254 = ( n313 & n2965 ) | ( n313 & ~n6139 ) | ( n2965 & ~n6139 ) ;
  assign n8256 = n8255 ^ n8254 ^ n3540 ;
  assign n8257 = n8256 ^ n5202 ^ n1743 ;
  assign n8253 = n1932 | n5123 ;
  assign n8258 = n8257 ^ n8253 ^ n5517 ;
  assign n8259 = n5768 ^ n256 ^ 1'b0 ;
  assign n8260 = ~n8258 & n8259 ;
  assign n8261 = n5943 ^ n4758 ^ n2654 ;
  assign n8262 = ( n1207 & n2335 ) | ( n1207 & n2999 ) | ( n2335 & n2999 ) ;
  assign n8263 = n3123 ^ n846 ^ 1'b0 ;
  assign n8264 = n8263 ^ n5851 ^ 1'b0 ;
  assign n8265 = n299 | n8264 ;
  assign n8266 = n6179 & n6944 ;
  assign n8267 = n7433 & n8266 ;
  assign n8268 = ( n5241 & n6271 ) | ( n5241 & n8267 ) | ( n6271 & n8267 ) ;
  assign n8269 = n2977 | n5748 ;
  assign n8270 = n595 & ~n8269 ;
  assign n8271 = n8270 ^ n5036 ^ n727 ;
  assign n8272 = n3506 ^ n3236 ^ x103 ;
  assign n8273 = ( n3955 & n7807 ) | ( n3955 & n8272 ) | ( n7807 & n8272 ) ;
  assign n8274 = n8273 ^ n4473 ^ n2388 ;
  assign n8275 = n1626 | n8274 ;
  assign n8276 = n4945 | n8275 ;
  assign n8277 = ~n462 & n6264 ;
  assign n8278 = n8277 ^ n7580 ^ 1'b0 ;
  assign n8279 = n834 & n8278 ;
  assign n8280 = ~n2337 & n8279 ;
  assign n8281 = n8280 ^ n2298 ^ n1252 ;
  assign n8282 = n3827 | n4909 ;
  assign n8283 = ( n804 & n1210 ) | ( n804 & n1728 ) | ( n1210 & n1728 ) ;
  assign n8284 = n7448 ^ n2387 ^ 1'b0 ;
  assign n8285 = n2957 | n8284 ;
  assign n8286 = n8283 & n8285 ;
  assign n8287 = n7455 ^ n3961 ^ 1'b0 ;
  assign n8288 = ~n2827 & n4717 ;
  assign n8289 = n4451 & ~n4552 ;
  assign n8290 = n8289 ^ n1690 ^ 1'b0 ;
  assign n8291 = n8232 | n8290 ;
  assign n8292 = n173 & ~n8291 ;
  assign n8293 = n5230 & ~n7490 ;
  assign n8294 = n911 & n8293 ;
  assign n8295 = n8294 ^ n2715 ^ 1'b0 ;
  assign n8296 = n5031 ^ n4216 ^ n529 ;
  assign n8297 = n7284 ^ n667 ^ 1'b0 ;
  assign n8298 = n1927 | n8297 ;
  assign n8299 = n3483 & ~n8114 ;
  assign n8300 = n8298 & ~n8299 ;
  assign n8301 = n4955 ^ n4546 ^ 1'b0 ;
  assign n8302 = n578 & ~n8301 ;
  assign n8303 = ~n164 & n4521 ;
  assign n8304 = n8302 & n8303 ;
  assign n8305 = n5907 ^ n2719 ^ 1'b0 ;
  assign n8306 = n3890 | n7814 ;
  assign n8307 = n7534 ^ n4256 ^ n2740 ;
  assign n8308 = n4450 ^ n1842 ^ 1'b0 ;
  assign n8309 = n4376 ^ n4088 ^ 1'b0 ;
  assign n8310 = n1598 & ~n8309 ;
  assign n8311 = n8310 ^ n1964 ^ 1'b0 ;
  assign n8312 = n8311 ^ n347 ^ n272 ;
  assign n8313 = n2081 ^ n1272 ^ n445 ;
  assign n8314 = n4057 | n8313 ;
  assign n8315 = n7769 ^ n1433 ^ 1'b0 ;
  assign n8316 = ~n2930 & n8315 ;
  assign n8317 = x49 | n2252 ;
  assign n8318 = n8317 ^ n3734 ^ 1'b0 ;
  assign n8319 = n1845 | n8318 ;
  assign n8320 = n8319 ^ n4148 ^ 1'b0 ;
  assign n8321 = ~n4571 & n8320 ;
  assign n8322 = ~n6754 & n8321 ;
  assign n8323 = n1708 & n8322 ;
  assign n8324 = n2574 | n2580 ;
  assign n8325 = n1020 | n8324 ;
  assign n8326 = n1593 ^ n937 ^ 1'b0 ;
  assign n8327 = x112 & ~n8326 ;
  assign n8328 = x81 & ~n8327 ;
  assign n8329 = n2338 | n8328 ;
  assign n8330 = n8329 ^ n3430 ^ 1'b0 ;
  assign n8331 = ( ~n7612 & n8325 ) | ( ~n7612 & n8330 ) | ( n8325 & n8330 ) ;
  assign n8332 = n2500 & n4805 ;
  assign n8333 = n7557 & ~n8332 ;
  assign n8334 = n8333 ^ n4993 ^ 1'b0 ;
  assign n8335 = ( n3726 & n3822 ) | ( n3726 & n6252 ) | ( n3822 & n6252 ) ;
  assign n8336 = ~n2467 & n8335 ;
  assign n8337 = ~n8334 & n8336 ;
  assign n8338 = n8337 ^ n4114 ^ 1'b0 ;
  assign n8339 = n6299 ^ n5944 ^ 1'b0 ;
  assign n8340 = n1288 & ~n8339 ;
  assign n8341 = n1199 & ~n3875 ;
  assign n8344 = ~n3822 & n5151 ;
  assign n8345 = n8344 ^ n1358 ^ 1'b0 ;
  assign n8346 = ~n1423 & n8345 ;
  assign n8347 = n5134 | n8346 ;
  assign n8342 = ( n442 & n1373 ) | ( n442 & n6219 ) | ( n1373 & n6219 ) ;
  assign n8343 = n4941 | n8342 ;
  assign n8348 = n8347 ^ n8343 ^ n4860 ;
  assign n8352 = ~n2985 & n3632 ;
  assign n8353 = ~n3999 & n8352 ;
  assign n8349 = n131 | n3566 ;
  assign n8350 = n4000 & ~n8349 ;
  assign n8351 = n8350 ^ n2880 ^ 1'b0 ;
  assign n8354 = n8353 ^ n8351 ^ 1'b0 ;
  assign n8355 = ~n8348 & n8354 ;
  assign n8356 = n2596 ^ n1244 ^ 1'b0 ;
  assign n8357 = n5792 & ~n8356 ;
  assign n8358 = n8357 ^ n4749 ^ n511 ;
  assign n8359 = n4057 ^ n3522 ^ 1'b0 ;
  assign n8360 = n150 | n7725 ;
  assign n8361 = n8360 ^ n6928 ^ 1'b0 ;
  assign n8362 = n2447 ^ n197 ^ 1'b0 ;
  assign n8363 = n8361 | n8362 ;
  assign n8364 = n2219 & ~n8363 ;
  assign n8365 = ~n256 & n8364 ;
  assign n8366 = n5416 ^ n560 ^ 1'b0 ;
  assign n8367 = n8366 ^ n3237 ^ n3030 ;
  assign n8368 = ~n3640 & n8367 ;
  assign n8373 = n6361 ^ n3859 ^ n768 ;
  assign n8374 = ~n3472 & n8373 ;
  assign n8369 = ~n654 & n2382 ;
  assign n8370 = n5901 & ~n8369 ;
  assign n8371 = n7513 & ~n8370 ;
  assign n8372 = ~n6894 & n8371 ;
  assign n8375 = n8374 ^ n8372 ^ x97 ;
  assign n8376 = n2409 | n4592 ;
  assign n8377 = ~n2770 & n4307 ;
  assign n8378 = ~n8376 & n8377 ;
  assign n8379 = n449 | n3864 ;
  assign n8380 = n8379 ^ n1167 ^ 1'b0 ;
  assign n8381 = ~n2741 & n8380 ;
  assign n8382 = n8381 ^ n1368 ^ 1'b0 ;
  assign n8383 = ~n6614 & n8382 ;
  assign n8384 = ~n8378 & n8383 ;
  assign n8385 = n2120 & n8384 ;
  assign n8386 = ( n3656 & ~n5920 ) | ( n3656 & n6225 ) | ( ~n5920 & n6225 ) ;
  assign n8387 = ( n1300 & n1797 ) | ( n1300 & ~n8386 ) | ( n1797 & ~n8386 ) ;
  assign n8388 = n302 & n5185 ;
  assign n8389 = n3281 ^ n2597 ^ 1'b0 ;
  assign n8390 = ~n8388 & n8389 ;
  assign n8391 = n1379 ^ n522 ^ 1'b0 ;
  assign n8392 = n6299 & ~n8391 ;
  assign n8393 = ~n2133 & n8392 ;
  assign n8394 = n8393 ^ n1254 ^ 1'b0 ;
  assign n8395 = ~n1508 & n4865 ;
  assign n8396 = n8395 ^ n8353 ^ n4167 ;
  assign n8397 = ( ~n1981 & n7064 ) | ( ~n1981 & n7317 ) | ( n7064 & n7317 ) ;
  assign n8398 = n8397 ^ x98 ^ 1'b0 ;
  assign n8399 = n874 & n8398 ;
  assign n8400 = n5950 & n8399 ;
  assign n8401 = n3600 & n6946 ;
  assign n8402 = n8401 ^ n6132 ^ 1'b0 ;
  assign n8403 = n2915 | n6284 ;
  assign n8404 = ( n5213 & n6104 ) | ( n5213 & ~n8403 ) | ( n6104 & ~n8403 ) ;
  assign n8405 = n8380 ^ n3632 ^ 1'b0 ;
  assign n8406 = ~n384 & n8405 ;
  assign n8407 = n1649 ^ n909 ^ 1'b0 ;
  assign n8408 = n8406 & ~n8407 ;
  assign n8409 = n1781 | n7716 ;
  assign n8410 = n7932 ^ n4161 ^ x98 ;
  assign n8411 = n8410 ^ n4484 ^ n245 ;
  assign n8412 = n8411 ^ n7407 ^ 1'b0 ;
  assign n8413 = ( ~n210 & n2423 ) | ( ~n210 & n2698 ) | ( n2423 & n2698 ) ;
  assign n8414 = n4191 | n8413 ;
  assign n8415 = n7788 ^ n3863 ^ 1'b0 ;
  assign n8417 = n4717 ^ n1950 ^ 1'b0 ;
  assign n8416 = n1331 & ~n4749 ;
  assign n8418 = n8417 ^ n8416 ^ 1'b0 ;
  assign n8419 = n1890 ^ n504 ^ 1'b0 ;
  assign n8420 = n6494 & ~n8419 ;
  assign n8421 = ~n7455 & n8420 ;
  assign n8422 = n8421 ^ n1491 ^ 1'b0 ;
  assign n8423 = n6245 & ~n8422 ;
  assign n8424 = ~n8418 & n8423 ;
  assign n8425 = n3446 & n4488 ;
  assign n8426 = n7703 ^ n4231 ^ 1'b0 ;
  assign n8427 = n6158 & n7398 ;
  assign n8428 = n3349 & n3659 ;
  assign n8429 = n8428 ^ n4997 ^ 1'b0 ;
  assign n8430 = ( n2172 & ~n8424 ) | ( n2172 & n8429 ) | ( ~n8424 & n8429 ) ;
  assign n8431 = ( ~n2903 & n3751 ) | ( ~n2903 & n8236 ) | ( n3751 & n8236 ) ;
  assign n8432 = n2763 & n4358 ;
  assign n8433 = ( n2078 & n2206 ) | ( n2078 & ~n5390 ) | ( n2206 & ~n5390 ) ;
  assign n8434 = ( ~n5546 & n5572 ) | ( ~n5546 & n8433 ) | ( n5572 & n8433 ) ;
  assign n8435 = ~n3763 & n8434 ;
  assign n8436 = n6444 & n8435 ;
  assign n8437 = n1386 ^ n927 ^ n813 ;
  assign n8438 = n8437 ^ n2361 ^ 1'b0 ;
  assign n8439 = n1505 & n8438 ;
  assign n8440 = n1739 ^ n521 ^ n491 ;
  assign n8441 = n1890 ^ n1442 ^ 1'b0 ;
  assign n8442 = n8440 | n8441 ;
  assign n8443 = ~n5523 & n8042 ;
  assign n8447 = n2120 & n2397 ;
  assign n8444 = n5241 ^ n1595 ^ 1'b0 ;
  assign n8445 = n8444 ^ n594 ^ 1'b0 ;
  assign n8446 = ( n654 & n2192 ) | ( n654 & ~n8445 ) | ( n2192 & ~n8445 ) ;
  assign n8448 = n8447 ^ n8446 ^ 1'b0 ;
  assign n8449 = n4290 & n5111 ;
  assign n8450 = ( n3583 & n4103 ) | ( n3583 & ~n8449 ) | ( n4103 & ~n8449 ) ;
  assign n8451 = n1608 & ~n8450 ;
  assign n8452 = n325 & n8451 ;
  assign n8453 = n1639 ^ n1575 ^ 1'b0 ;
  assign n8454 = ~n1199 & n8432 ;
  assign n8455 = ~n3189 & n8454 ;
  assign n8456 = ~n2549 & n3621 ;
  assign n8457 = ( ~n2968 & n6960 ) | ( ~n2968 & n8456 ) | ( n6960 & n8456 ) ;
  assign n8458 = n593 | n4027 ;
  assign n8459 = n2452 | n5559 ;
  assign n8460 = n8459 ^ n5078 ^ 1'b0 ;
  assign n8461 = ( n3964 & n4581 ) | ( n3964 & n8460 ) | ( n4581 & n8460 ) ;
  assign n8462 = n8458 & n8461 ;
  assign n8463 = ~n1167 & n8462 ;
  assign n8467 = n1959 ^ n1003 ^ n249 ;
  assign n8465 = n4095 ^ n1470 ^ 1'b0 ;
  assign n8466 = ~n3327 & n8465 ;
  assign n8468 = n8467 ^ n8466 ^ 1'b0 ;
  assign n8464 = n836 & n2884 ;
  assign n8469 = n8468 ^ n8464 ^ n4043 ;
  assign n8472 = n7784 ^ n1200 ^ 1'b0 ;
  assign n8470 = n3488 ^ n3169 ^ 1'b0 ;
  assign n8471 = ~n5088 & n8470 ;
  assign n8473 = n8472 ^ n8471 ^ 1'b0 ;
  assign n8474 = n5020 ^ n1644 ^ n568 ;
  assign n8475 = ( ~n892 & n5250 ) | ( ~n892 & n8474 ) | ( n5250 & n8474 ) ;
  assign n8476 = n8475 ^ n3483 ^ n245 ;
  assign n8477 = ~n2986 & n7346 ;
  assign n8478 = n3961 ^ n2008 ^ 1'b0 ;
  assign n8479 = n8478 ^ n6525 ^ n1890 ;
  assign n8481 = ~n2491 & n5669 ;
  assign n8482 = n8481 ^ x55 ^ 1'b0 ;
  assign n8483 = ~n8125 & n8482 ;
  assign n8480 = n1796 & n1960 ;
  assign n8484 = n8483 ^ n8480 ^ 1'b0 ;
  assign n8485 = n303 | n6295 ;
  assign n8486 = n7820 ^ n949 ^ n790 ;
  assign n8487 = n8486 ^ n768 ^ 1'b0 ;
  assign n8488 = n8487 ^ n3745 ^ 1'b0 ;
  assign n8489 = ( n3874 & ~n5921 ) | ( n3874 & n6117 ) | ( ~n5921 & n6117 ) ;
  assign n8490 = ~n526 & n8489 ;
  assign n8491 = n1330 ^ x87 ^ 1'b0 ;
  assign n8492 = n8491 ^ n4734 ^ n2056 ;
  assign n8493 = ( n1654 & n8490 ) | ( n1654 & n8492 ) | ( n8490 & n8492 ) ;
  assign n8494 = n8493 ^ n2853 ^ 1'b0 ;
  assign n8495 = n3513 ^ x13 ^ 1'b0 ;
  assign n8496 = ~n2999 & n8495 ;
  assign n8497 = n8496 ^ n4261 ^ n1498 ;
  assign n8498 = n2364 | n4617 ;
  assign n8499 = n6036 & ~n8498 ;
  assign n8500 = n8499 ^ n6258 ^ 1'b0 ;
  assign n8501 = ( ~n4158 & n8486 ) | ( ~n4158 & n8500 ) | ( n8486 & n8500 ) ;
  assign n8502 = ( n2304 & n2582 ) | ( n2304 & ~n4608 ) | ( n2582 & ~n4608 ) ;
  assign n8506 = n4035 ^ n340 ^ 1'b0 ;
  assign n8507 = n1754 | n8506 ;
  assign n8505 = ~n1653 & n2342 ;
  assign n8508 = n8507 ^ n8505 ^ 1'b0 ;
  assign n8509 = x18 & n2416 ;
  assign n8510 = n8509 ^ n1283 ^ 1'b0 ;
  assign n8511 = n8510 ^ n6152 ^ n600 ;
  assign n8512 = x126 & ~n8511 ;
  assign n8513 = ~n8508 & n8512 ;
  assign n8503 = n2248 ^ n1793 ^ n383 ;
  assign n8504 = ( n4879 & n5198 ) | ( n4879 & ~n8503 ) | ( n5198 & ~n8503 ) ;
  assign n8514 = n8513 ^ n8504 ^ 1'b0 ;
  assign n8515 = n8502 & ~n8514 ;
  assign n8518 = ~n820 & n7769 ;
  assign n8519 = ~n5822 & n8518 ;
  assign n8516 = n8468 ^ n3270 ^ 1'b0 ;
  assign n8517 = n6793 & ~n8516 ;
  assign n8520 = n8519 ^ n8517 ^ 1'b0 ;
  assign n8521 = n3615 | n6341 ;
  assign n8523 = n4959 ^ n758 ^ n270 ;
  assign n8524 = ( n3880 & ~n3949 ) | ( n3880 & n8523 ) | ( ~n3949 & n8523 ) ;
  assign n8522 = n3257 | n5057 ;
  assign n8525 = n8524 ^ n8522 ^ n7695 ;
  assign n8526 = n7189 & ~n7286 ;
  assign n8527 = ~n358 & n1521 ;
  assign n8528 = n2948 ^ n2342 ^ 1'b0 ;
  assign n8529 = n8528 ^ n5916 ^ 1'b0 ;
  assign n8530 = n600 | n6788 ;
  assign n8531 = n8529 & ~n8530 ;
  assign n8538 = n2438 ^ n813 ^ 1'b0 ;
  assign n8532 = n2371 ^ n914 ^ 1'b0 ;
  assign n8533 = n8532 ^ n5854 ^ 1'b0 ;
  assign n8534 = n1171 & ~n3345 ;
  assign n8535 = n8534 ^ n4243 ^ 1'b0 ;
  assign n8536 = ( n3941 & n4094 ) | ( n3941 & ~n8535 ) | ( n4094 & ~n8535 ) ;
  assign n8537 = n8533 & ~n8536 ;
  assign n8539 = n8538 ^ n8537 ^ 1'b0 ;
  assign n8540 = n8539 ^ n6012 ^ 1'b0 ;
  assign n8541 = n6477 & ~n8540 ;
  assign n8542 = n4704 | n5049 ;
  assign n8543 = n8542 ^ x37 ^ 1'b0 ;
  assign n8544 = n3894 & ~n7552 ;
  assign n8545 = n8544 ^ n2536 ^ 1'b0 ;
  assign n8546 = n2416 & n8545 ;
  assign n8547 = ( n7312 & n8543 ) | ( n7312 & n8546 ) | ( n8543 & n8546 ) ;
  assign n8548 = n399 & n2761 ;
  assign n8549 = ~n1160 & n8548 ;
  assign n8550 = n1216 & n8549 ;
  assign n8551 = n8550 ^ n8410 ^ n4055 ;
  assign n8552 = n3316 ^ n193 ^ 1'b0 ;
  assign n8553 = n8552 ^ n6012 ^ n1210 ;
  assign n8554 = n4215 | n8553 ;
  assign n8555 = n8554 ^ n8295 ^ 1'b0 ;
  assign n8556 = n4584 | n5963 ;
  assign n8557 = n6057 ^ n4567 ^ n3013 ;
  assign n8558 = ~n423 & n8557 ;
  assign n8559 = n6730 | n8558 ;
  assign n8560 = n8559 ^ n5938 ^ 1'b0 ;
  assign n8561 = n5822 ^ n1400 ^ 1'b0 ;
  assign n8562 = n6242 | n8561 ;
  assign n8563 = n4033 | n4083 ;
  assign n8564 = n8563 ^ n2850 ^ 1'b0 ;
  assign n8565 = ( n557 & ~n8562 ) | ( n557 & n8564 ) | ( ~n8562 & n8564 ) ;
  assign n8566 = n5977 ^ n3951 ^ n1740 ;
  assign n8567 = ~n8565 & n8566 ;
  assign n8568 = ( n667 & n7980 ) | ( n667 & ~n8567 ) | ( n7980 & ~n8567 ) ;
  assign n8569 = n2421 ^ n529 ^ 1'b0 ;
  assign n8570 = ~n219 & n8569 ;
  assign n8571 = ~x31 & n8570 ;
  assign n8572 = n354 & ~n3100 ;
  assign n8573 = n8572 ^ n5959 ^ n1485 ;
  assign n8574 = ( ~n836 & n1133 ) | ( ~n836 & n2882 ) | ( n1133 & n2882 ) ;
  assign n8575 = n8574 ^ n5168 ^ n1659 ;
  assign n8576 = ( ~n1537 & n3753 ) | ( ~n1537 & n7244 ) | ( n3753 & n7244 ) ;
  assign n8577 = ( n8573 & n8575 ) | ( n8573 & n8576 ) | ( n8575 & n8576 ) ;
  assign n8583 = n1093 | n5361 ;
  assign n8584 = n8583 ^ n8229 ^ n3574 ;
  assign n8585 = n5488 | n8584 ;
  assign n8578 = n3709 & n4120 ;
  assign n8579 = ~n374 & n1846 ;
  assign n8580 = n8578 & n8579 ;
  assign n8581 = n3478 & ~n8580 ;
  assign n8582 = n8581 ^ n3661 ^ 1'b0 ;
  assign n8586 = n8585 ^ n8582 ^ n6198 ;
  assign n8587 = ( ~n154 & n1154 ) | ( ~n154 & n2783 ) | ( n1154 & n2783 ) ;
  assign n8588 = ~n2180 & n6562 ;
  assign n8589 = n8588 ^ n7360 ^ 1'b0 ;
  assign n8590 = n5070 ^ n3118 ^ 1'b0 ;
  assign n8591 = ~n6905 & n8590 ;
  assign n8592 = n2300 ^ n950 ^ n477 ;
  assign n8593 = ~n4310 & n8592 ;
  assign n8594 = ~n3163 & n4581 ;
  assign n8595 = ~n4581 & n8594 ;
  assign n8596 = n8595 ^ x38 ^ 1'b0 ;
  assign n8597 = n751 | n8596 ;
  assign n8598 = n1257 | n8597 ;
  assign n8599 = n367 & ~n1209 ;
  assign n8600 = n8599 ^ n4095 ^ 1'b0 ;
  assign n8601 = n1173 & ~n8600 ;
  assign n8602 = n4557 ^ x79 ^ 1'b0 ;
  assign n8603 = n5236 | n8602 ;
  assign n8604 = n4029 & ~n8603 ;
  assign n8605 = n8604 ^ n6169 ^ 1'b0 ;
  assign n8606 = n1512 | n2092 ;
  assign n8607 = n8606 ^ n4221 ^ 1'b0 ;
  assign n8608 = ( n1690 & n7970 ) | ( n1690 & ~n8607 ) | ( n7970 & ~n8607 ) ;
  assign n8609 = n3961 ^ n383 ^ n206 ;
  assign n8610 = n8609 ^ n1305 ^ 1'b0 ;
  assign n8611 = n518 & n8610 ;
  assign n8612 = n1779 | n8611 ;
  assign n8613 = n5902 & n8612 ;
  assign n8614 = n801 | n7298 ;
  assign n8615 = ~n2165 & n2275 ;
  assign n8616 = ( x28 & n1887 ) | ( x28 & ~n2917 ) | ( n1887 & ~n2917 ) ;
  assign n8617 = n8616 ^ n2791 ^ 1'b0 ;
  assign n8618 = n8617 ^ n1083 ^ 1'b0 ;
  assign n8619 = n8236 ^ n4103 ^ 1'b0 ;
  assign n8620 = n3701 & ~n3905 ;
  assign n8621 = ( n1392 & n7804 ) | ( n1392 & n8620 ) | ( n7804 & n8620 ) ;
  assign n8622 = n6718 ^ n1960 ^ 1'b0 ;
  assign n8623 = n4264 | n8622 ;
  assign n8624 = n1928 | n8623 ;
  assign n8625 = n860 & ~n8624 ;
  assign n8629 = ~n362 & n4437 ;
  assign n8630 = n8629 ^ n2538 ^ 1'b0 ;
  assign n8626 = n4532 ^ n3606 ^ n625 ;
  assign n8627 = ( n6758 & ~n8413 ) | ( n6758 & n8626 ) | ( ~n8413 & n8626 ) ;
  assign n8628 = n5323 & n8627 ;
  assign n8631 = n8630 ^ n8628 ^ 1'b0 ;
  assign n8632 = ( n585 & n2597 ) | ( n585 & n7317 ) | ( n2597 & n7317 ) ;
  assign n8633 = n8632 ^ n4118 ^ 1'b0 ;
  assign n8634 = n940 & ~n1162 ;
  assign n8635 = ~n4347 & n6075 ;
  assign n8636 = n5814 & n7122 ;
  assign n8637 = ( ~x22 & n1058 ) | ( ~x22 & n1927 ) | ( n1058 & n1927 ) ;
  assign n8638 = n1979 ^ x97 ^ 1'b0 ;
  assign n8639 = n8637 | n8638 ;
  assign n8640 = x17 & ~n1073 ;
  assign n8641 = n8639 & n8640 ;
  assign n8642 = ~n859 & n3015 ;
  assign n8643 = n8642 ^ n5335 ^ 1'b0 ;
  assign n8644 = n8643 ^ n6821 ^ 1'b0 ;
  assign n8645 = n8644 ^ n6382 ^ n4461 ;
  assign n8646 = n1884 | n2580 ;
  assign n8647 = n8645 & ~n8646 ;
  assign n8648 = ( n3390 & ~n5175 ) | ( n3390 & n8538 ) | ( ~n5175 & n8538 ) ;
  assign n8649 = n3376 & ~n3559 ;
  assign n8650 = n8649 ^ n2740 ^ 1'b0 ;
  assign n8651 = n8648 | n8650 ;
  assign n8652 = n8608 | n8651 ;
  assign n8653 = n5575 ^ n462 ^ 1'b0 ;
  assign n8654 = ( n296 & n5966 ) | ( n296 & ~n8653 ) | ( n5966 & ~n8653 ) ;
  assign n8655 = ~n4387 & n7146 ;
  assign n8656 = ( n4265 & ~n8654 ) | ( n4265 & n8655 ) | ( ~n8654 & n8655 ) ;
  assign n8657 = n5012 | n6521 ;
  assign n8658 = ~n2763 & n6965 ;
  assign n8659 = n3094 ^ n2427 ^ 1'b0 ;
  assign n8660 = n8658 & ~n8659 ;
  assign n8661 = n940 & ~n3453 ;
  assign n8662 = n393 & n8661 ;
  assign n8663 = n8662 ^ n3595 ^ 1'b0 ;
  assign n8666 = n2431 ^ n734 ^ 1'b0 ;
  assign n8667 = n1716 & n8666 ;
  assign n8665 = x25 & n2115 ;
  assign n8668 = n8667 ^ n8665 ^ 1'b0 ;
  assign n8664 = n4398 ^ n3176 ^ 1'b0 ;
  assign n8669 = n8668 ^ n8664 ^ 1'b0 ;
  assign n8670 = n4642 ^ n1435 ^ 1'b0 ;
  assign n8671 = n2286 | n8670 ;
  assign n8672 = ~n1610 & n2779 ;
  assign n8673 = n8671 & n8672 ;
  assign n8674 = n6484 | n8673 ;
  assign n8675 = n8669 & ~n8674 ;
  assign n8676 = n8675 ^ n4576 ^ 1'b0 ;
  assign n8677 = n2264 ^ n708 ^ x124 ;
  assign n8678 = n8193 & ~n8677 ;
  assign n8679 = n6325 & n8678 ;
  assign n8680 = n3508 & ~n7865 ;
  assign n8681 = n6845 ^ n3608 ^ 1'b0 ;
  assign n8682 = ~n8680 & n8681 ;
  assign n8683 = n1993 ^ n1833 ^ 1'b0 ;
  assign n8684 = n3962 & ~n8683 ;
  assign n8685 = n6661 ^ n4991 ^ n1110 ;
  assign n8686 = n2999 | n4663 ;
  assign n8687 = ( ~n1747 & n8685 ) | ( ~n1747 & n8686 ) | ( n8685 & n8686 ) ;
  assign n8688 = n8687 ^ n2137 ^ 1'b0 ;
  assign n8689 = n6651 ^ n4158 ^ n2547 ;
  assign n8690 = x70 & n7197 ;
  assign n8691 = ~n3484 & n8690 ;
  assign n8692 = n3058 ^ n1752 ^ n701 ;
  assign n8693 = n3413 | n8692 ;
  assign n8694 = n8693 ^ n6828 ^ 1'b0 ;
  assign n8695 = n3581 & n8694 ;
  assign n8696 = ~n4163 & n8695 ;
  assign n8697 = n8696 ^ n650 ^ 1'b0 ;
  assign n8699 = n3621 | n6605 ;
  assign n8700 = n7317 | n8699 ;
  assign n8698 = n1489 & n4382 ;
  assign n8701 = n8700 ^ n8698 ^ 1'b0 ;
  assign n8702 = n1114 & n1585 ;
  assign n8703 = n6605 ^ n6381 ^ 1'b0 ;
  assign n8704 = n8702 & ~n8703 ;
  assign n8705 = ( n3063 & n4201 ) | ( n3063 & n6182 ) | ( n4201 & n6182 ) ;
  assign n8717 = n1637 & n2528 ;
  assign n8715 = n1448 & n3482 ;
  assign n8716 = n4840 | n8715 ;
  assign n8718 = n8717 ^ n8716 ^ n5484 ;
  assign n8706 = n6731 ^ n5428 ^ 1'b0 ;
  assign n8707 = n3697 ^ n2929 ^ 1'b0 ;
  assign n8709 = n490 | n608 ;
  assign n8710 = n316 & n8709 ;
  assign n8711 = n8710 ^ n3311 ^ 1'b0 ;
  assign n8708 = n5315 ^ n657 ^ 1'b0 ;
  assign n8712 = n8711 ^ n8708 ^ n345 ;
  assign n8713 = n8707 & n8712 ;
  assign n8714 = n8706 & n8713 ;
  assign n8719 = n8718 ^ n8714 ^ n160 ;
  assign n8720 = n1952 | n2708 ;
  assign n8721 = n8720 ^ n832 ^ 1'b0 ;
  assign n8722 = n8721 ^ n5736 ^ 1'b0 ;
  assign n8726 = n1491 & ~n2028 ;
  assign n8727 = n8726 ^ n5703 ^ 1'b0 ;
  assign n8728 = n8727 ^ n3465 ^ n3390 ;
  assign n8723 = n2666 | n2697 ;
  assign n8724 = n8723 ^ n1855 ^ 1'b0 ;
  assign n8725 = n1502 & n8724 ;
  assign n8729 = n8728 ^ n8725 ^ 1'b0 ;
  assign n8730 = n4664 ^ n3853 ^ n585 ;
  assign n8731 = n7128 ^ n5118 ^ n2979 ;
  assign n8732 = n6712 & n8731 ;
  assign n8734 = x39 & ~n3775 ;
  assign n8735 = n8734 ^ n1880 ^ 1'b0 ;
  assign n8736 = ( n3172 & ~n5951 ) | ( n3172 & n8735 ) | ( ~n5951 & n8735 ) ;
  assign n8733 = ~n6989 & n7894 ;
  assign n8737 = n8736 ^ n8733 ^ 1'b0 ;
  assign n8738 = n8737 ^ x113 ^ 1'b0 ;
  assign n8739 = n8738 ^ n904 ^ 1'b0 ;
  assign n8740 = ~n2176 & n8739 ;
  assign n8741 = n8740 ^ x1 ^ 1'b0 ;
  assign n8742 = n2613 ^ n1096 ^ 1'b0 ;
  assign n8743 = n6878 & n7670 ;
  assign n8744 = n8743 ^ n2391 ^ 1'b0 ;
  assign n8745 = n1972 ^ n1302 ^ 1'b0 ;
  assign n8746 = n1366 | n8745 ;
  assign n8747 = n7393 | n8746 ;
  assign n8748 = n8747 ^ n4126 ^ 1'b0 ;
  assign n8749 = n3076 & ~n8748 ;
  assign n8750 = ~n8744 & n8749 ;
  assign n8751 = n1503 | n5973 ;
  assign n8752 = n7435 ^ n614 ^ 1'b0 ;
  assign n8753 = n5605 | n8752 ;
  assign n8754 = x31 | n8753 ;
  assign n8756 = n269 ^ x17 ^ 1'b0 ;
  assign n8755 = n2440 & ~n6409 ;
  assign n8757 = n8756 ^ n8755 ^ 1'b0 ;
  assign n8758 = n3501 | n5205 ;
  assign n8759 = n5824 & ~n8758 ;
  assign n8760 = n4027 & ~n4598 ;
  assign n8761 = ~n8503 & n8760 ;
  assign n8762 = ( ~n3503 & n6409 ) | ( ~n3503 & n8761 ) | ( n6409 & n8761 ) ;
  assign n8763 = n8762 ^ n270 ^ 1'b0 ;
  assign n8764 = n1497 & ~n8763 ;
  assign n8765 = ~n5804 & n8764 ;
  assign n8766 = n7430 ^ n4229 ^ n2201 ;
  assign n8767 = n4458 ^ n163 ^ x31 ;
  assign n8771 = n968 & n5653 ;
  assign n8772 = n4554 & n8771 ;
  assign n8773 = n8772 ^ n1607 ^ 1'b0 ;
  assign n8768 = n4224 ^ n2179 ^ 1'b0 ;
  assign n8769 = ( ~n2626 & n2702 ) | ( ~n2626 & n8768 ) | ( n2702 & n8768 ) ;
  assign n8770 = n4594 & n8769 ;
  assign n8774 = n8773 ^ n8770 ^ 1'b0 ;
  assign n8775 = ~n4881 & n5879 ;
  assign n8776 = n1054 & n8775 ;
  assign n8777 = n8776 ^ n661 ^ 1'b0 ;
  assign n8778 = n2999 & n3434 ;
  assign n8779 = ~n5936 & n8778 ;
  assign n8780 = n8779 ^ n443 ^ 1'b0 ;
  assign n8781 = n2590 & ~n8780 ;
  assign n8782 = n1445 | n2279 ;
  assign n8783 = n3363 & ~n8782 ;
  assign n8784 = n8783 ^ n8363 ^ n4475 ;
  assign n8785 = ( n4620 & ~n6600 ) | ( n4620 & n7621 ) | ( ~n6600 & n7621 ) ;
  assign n8786 = n8785 ^ n6854 ^ 1'b0 ;
  assign n8787 = n7732 & n8786 ;
  assign n8788 = n3391 & ~n3546 ;
  assign n8789 = ~n1962 & n8788 ;
  assign n8790 = n6756 & n8789 ;
  assign n8791 = n8487 & n8790 ;
  assign n8792 = ~n1900 & n3371 ;
  assign n8793 = n8792 ^ n4185 ^ 1'b0 ;
  assign n8794 = n6903 & n8793 ;
  assign n8795 = ( n1725 & ~n1967 ) | ( n1725 & n2217 ) | ( ~n1967 & n2217 ) ;
  assign n8796 = n7570 & n8795 ;
  assign n8797 = n1507 & ~n8796 ;
  assign n8798 = n8797 ^ n2977 ^ 1'b0 ;
  assign n8799 = ( n2462 & n7938 ) | ( n2462 & ~n8798 ) | ( n7938 & ~n8798 ) ;
  assign n8806 = ~n3670 & n5257 ;
  assign n8807 = ~n2945 & n8806 ;
  assign n8803 = n4150 & ~n4571 ;
  assign n8804 = ~n1425 & n8803 ;
  assign n8805 = n8804 ^ n1617 ^ 1'b0 ;
  assign n8808 = n8807 ^ n8805 ^ n3999 ;
  assign n8809 = n8808 ^ n5530 ^ n4163 ;
  assign n8800 = n533 | n3564 ;
  assign n8801 = n4824 | n8800 ;
  assign n8802 = ~n5045 & n8801 ;
  assign n8810 = n8809 ^ n8802 ^ 1'b0 ;
  assign n8811 = n8810 ^ n6444 ^ n2290 ;
  assign n8812 = n1369 & n1726 ;
  assign n8813 = ( n2698 & n2772 ) | ( n2698 & n3932 ) | ( n2772 & n3932 ) ;
  assign n8814 = ( n8440 & n8812 ) | ( n8440 & n8813 ) | ( n8812 & n8813 ) ;
  assign n8815 = ~n2366 & n2645 ;
  assign n8817 = n925 ^ n613 ^ 1'b0 ;
  assign n8818 = n8817 ^ n5358 ^ 1'b0 ;
  assign n8816 = n250 & n6539 ;
  assign n8819 = n8818 ^ n8816 ^ 1'b0 ;
  assign n8820 = n8819 ^ n7593 ^ 1'b0 ;
  assign n8821 = n1964 & n8820 ;
  assign n8822 = n232 & n936 ;
  assign n8823 = n1290 & n8822 ;
  assign n8824 = ( ~n575 & n2882 ) | ( ~n575 & n8823 ) | ( n2882 & n8823 ) ;
  assign n8825 = ~n2873 & n4437 ;
  assign n8826 = ~n8824 & n8825 ;
  assign n8827 = n1139 | n8826 ;
  assign n8828 = ( n201 & n4252 ) | ( n201 & ~n6587 ) | ( n4252 & ~n6587 ) ;
  assign n8829 = ~n1768 & n2534 ;
  assign n8830 = ( n2174 & ~n6533 ) | ( n2174 & n8829 ) | ( ~n6533 & n8829 ) ;
  assign n8831 = n1722 & n8830 ;
  assign n8832 = n8831 ^ n8768 ^ 1'b0 ;
  assign n8833 = n1420 & n1457 ;
  assign n8834 = n8833 ^ n4552 ^ 1'b0 ;
  assign n8835 = ~n8832 & n8834 ;
  assign n8836 = n6656 ^ n4785 ^ n3263 ;
  assign n8837 = n1594 | n2462 ;
  assign n8838 = n6992 ^ n4372 ^ 1'b0 ;
  assign n8839 = ( n730 & n804 ) | ( n730 & n7255 ) | ( n804 & n7255 ) ;
  assign n8840 = n4527 ^ n1614 ^ n1259 ;
  assign n8841 = n8840 ^ n5377 ^ 1'b0 ;
  assign n8842 = n1721 & n8841 ;
  assign n8843 = n8839 & n8842 ;
  assign n8844 = n8843 ^ n4296 ^ 1'b0 ;
  assign n8845 = n2755 ^ n1588 ^ 1'b0 ;
  assign n8846 = n5639 ^ n2006 ^ 1'b0 ;
  assign n8847 = ( ~n6317 & n8845 ) | ( ~n6317 & n8846 ) | ( n8845 & n8846 ) ;
  assign n8848 = n3009 | n3209 ;
  assign n8849 = ~n849 & n882 ;
  assign n8850 = ~n8848 & n8849 ;
  assign n8854 = ( ~n210 & n2820 ) | ( ~n210 & n4107 ) | ( n2820 & n4107 ) ;
  assign n8852 = n345 | n1781 ;
  assign n8851 = n2106 & ~n7507 ;
  assign n8853 = n8852 ^ n8851 ^ 1'b0 ;
  assign n8855 = n8854 ^ n8853 ^ n7354 ;
  assign n8856 = ( ~n1752 & n2599 ) | ( ~n1752 & n2614 ) | ( n2599 & n2614 ) ;
  assign n8857 = ~n5725 & n8856 ;
  assign n8858 = n2120 | n4959 ;
  assign n8859 = n5010 ^ n349 ^ 1'b0 ;
  assign n8864 = n3270 & ~n7373 ;
  assign n8860 = n3483 | n4917 ;
  assign n8861 = ( x44 & ~n2913 ) | ( x44 & n6079 ) | ( ~n2913 & n6079 ) ;
  assign n8862 = n3926 | n8861 ;
  assign n8863 = n8860 | n8862 ;
  assign n8865 = n8864 ^ n8863 ^ 1'b0 ;
  assign n8868 = ( n4269 & ~n4367 ) | ( n4269 & n4576 ) | ( ~n4367 & n4576 ) ;
  assign n8869 = n8868 ^ n2426 ^ 1'b0 ;
  assign n8866 = ~n1704 & n1869 ;
  assign n8867 = n8866 ^ n1593 ^ 1'b0 ;
  assign n8870 = n8869 ^ n8867 ^ 1'b0 ;
  assign n8871 = n8870 ^ n8288 ^ 1'b0 ;
  assign n8872 = n5155 ^ n4813 ^ 1'b0 ;
  assign n8873 = n6878 ^ n5577 ^ 1'b0 ;
  assign n8874 = ~n862 & n8873 ;
  assign n8875 = ~n383 & n8874 ;
  assign n8876 = x112 & ~n2165 ;
  assign n8877 = n8876 ^ n1485 ^ 1'b0 ;
  assign n8878 = ( n5640 & ~n7221 ) | ( n5640 & n8877 ) | ( ~n7221 & n8877 ) ;
  assign n8879 = n3762 ^ n1988 ^ 1'b0 ;
  assign n8880 = n8644 & n8879 ;
  assign n8881 = n4475 & ~n5815 ;
  assign n8882 = n8881 ^ n7862 ^ 1'b0 ;
  assign n8883 = n2163 ^ n1069 ^ 1'b0 ;
  assign n8884 = n812 | n8883 ;
  assign n8885 = n2268 & ~n8884 ;
  assign n8886 = n3783 & ~n8885 ;
  assign n8887 = ~n8882 & n8886 ;
  assign n8888 = ~n2837 & n2929 ;
  assign n8889 = n152 & n2115 ;
  assign n8890 = ~n444 & n8889 ;
  assign n8891 = n1773 | n8890 ;
  assign n8892 = n1542 & ~n4751 ;
  assign n8893 = n1290 | n8892 ;
  assign n8894 = n8891 & ~n8893 ;
  assign n8895 = n425 | n1046 ;
  assign n8896 = n6930 | n8895 ;
  assign n8897 = n1200 & ~n1369 ;
  assign n8899 = n8728 ^ n4935 ^ 1'b0 ;
  assign n8900 = n172 | n8899 ;
  assign n8898 = ~n2333 & n3207 ;
  assign n8901 = n8900 ^ n8898 ^ 1'b0 ;
  assign n8902 = n8901 ^ n4211 ^ 1'b0 ;
  assign n8903 = n3260 | n8902 ;
  assign n8904 = ( n4757 & n7788 ) | ( n4757 & ~n8903 ) | ( n7788 & ~n8903 ) ;
  assign n8905 = ( ~n5399 & n6946 ) | ( ~n5399 & n8706 ) | ( n6946 & n8706 ) ;
  assign n8907 = n3772 & ~n6395 ;
  assign n8908 = n5844 & n8907 ;
  assign n8906 = n4554 | n5523 ;
  assign n8909 = n8908 ^ n8906 ^ 1'b0 ;
  assign n8910 = n8861 ^ n3695 ^ 1'b0 ;
  assign n8911 = n8909 & n8910 ;
  assign n8912 = n4204 ^ n2151 ^ 1'b0 ;
  assign n8913 = ~n6763 & n8912 ;
  assign n8914 = n2816 ^ n1831 ^ 1'b0 ;
  assign n8915 = n8914 ^ n386 ^ 1'b0 ;
  assign n8916 = n4554 | n8915 ;
  assign n8917 = n8916 ^ n1555 ^ 1'b0 ;
  assign n8918 = n679 & n8917 ;
  assign n8919 = n6402 ^ n1731 ^ 1'b0 ;
  assign n8920 = n2880 ^ n1342 ^ 1'b0 ;
  assign n8921 = n1848 & ~n8920 ;
  assign n8922 = ~n6149 & n6315 ;
  assign n8923 = n4661 | n8922 ;
  assign n8924 = n719 | n4313 ;
  assign n8925 = n8924 ^ n1376 ^ n353 ;
  assign n8926 = n8198 | n8925 ;
  assign n8927 = n2913 ^ n2036 ^ n1660 ;
  assign n8928 = n2498 & n5502 ;
  assign n8929 = n8928 ^ n3907 ^ 1'b0 ;
  assign n8930 = n1822 & ~n8929 ;
  assign n8931 = n6783 & n8930 ;
  assign n8940 = ~n649 & n962 ;
  assign n8941 = ~n5297 & n8940 ;
  assign n8933 = n916 ^ n637 ^ n463 ;
  assign n8934 = n8933 ^ n8065 ^ 1'b0 ;
  assign n8935 = ~n1587 & n8934 ;
  assign n8932 = n768 & ~n6425 ;
  assign n8936 = n8935 ^ n8932 ^ 1'b0 ;
  assign n8937 = n8936 ^ n5003 ^ 1'b0 ;
  assign n8938 = n5931 | n6271 ;
  assign n8939 = n8937 | n8938 ;
  assign n8942 = n8941 ^ n8939 ^ n8038 ;
  assign n8943 = n8942 ^ n5340 ^ 1'b0 ;
  assign n8944 = n8931 | n8943 ;
  assign n8945 = n2472 | n6229 ;
  assign n8946 = n6731 ^ n3299 ^ 1'b0 ;
  assign n8947 = n2493 & n8946 ;
  assign n8948 = n5196 ^ n3493 ^ 1'b0 ;
  assign n8949 = n4586 & n8948 ;
  assign n8950 = n8066 ^ n296 ^ 1'b0 ;
  assign n8951 = n878 & n8950 ;
  assign n8952 = n6183 ^ n4663 ^ n4401 ;
  assign n8953 = n4498 & ~n8952 ;
  assign n8954 = n3009 ^ n485 ^ 1'b0 ;
  assign n8955 = n2269 & n8954 ;
  assign n8956 = x108 & n8955 ;
  assign n8957 = n8956 ^ n3056 ^ 1'b0 ;
  assign n8958 = n4216 ^ n1805 ^ 1'b0 ;
  assign n8959 = n4269 & ~n4738 ;
  assign n8960 = n1110 | n5355 ;
  assign n8961 = n8959 | n8960 ;
  assign n8962 = n4318 ^ n1116 ^ 1'b0 ;
  assign n8963 = n8961 | n8962 ;
  assign n8964 = n6198 ^ n5378 ^ 1'b0 ;
  assign n8965 = ~n2660 & n8964 ;
  assign n8966 = n1114 & ~n2293 ;
  assign n8967 = n1495 & n8966 ;
  assign n8968 = n3180 ^ n2218 ^ 1'b0 ;
  assign n8969 = ~n8967 & n8968 ;
  assign n8970 = ~n5948 & n8969 ;
  assign n8971 = n8970 ^ n8856 ^ 1'b0 ;
  assign n8972 = n8931 | n8971 ;
  assign n8974 = n822 & n1480 ;
  assign n8973 = n6926 | n8761 ;
  assign n8975 = n8974 ^ n8973 ^ 1'b0 ;
  assign n8976 = ~n4281 & n8975 ;
  assign n8977 = n1947 & n4995 ;
  assign n8978 = n8977 ^ n1079 ^ 1'b0 ;
  assign n8979 = n8978 ^ n3616 ^ n2450 ;
  assign n8980 = n1706 ^ n154 ^ 1'b0 ;
  assign n8981 = ( ~n3317 & n7229 ) | ( ~n3317 & n8980 ) | ( n7229 & n8980 ) ;
  assign n8982 = n8981 ^ n7820 ^ n5110 ;
  assign n8983 = n4134 ^ n2125 ^ 1'b0 ;
  assign n8984 = ~n5552 & n8983 ;
  assign n8985 = n8984 ^ n6546 ^ n6496 ;
  assign n8986 = ~n5715 & n7295 ;
  assign n8987 = n8985 & n8986 ;
  assign n8988 = ( ~n502 & n1843 ) | ( ~n502 & n2523 ) | ( n1843 & n2523 ) ;
  assign n8989 = n7428 & ~n8988 ;
  assign n8990 = ~n6070 & n8989 ;
  assign n8991 = n2563 ^ n477 ^ 1'b0 ;
  assign n8992 = n2780 ^ n502 ^ 1'b0 ;
  assign n8993 = ~n8991 & n8992 ;
  assign n8994 = ( n2276 & ~n2686 ) | ( n2276 & n8993 ) | ( ~n2686 & n8993 ) ;
  assign n8995 = n8599 ^ n6243 ^ n4710 ;
  assign n8996 = ( n2173 & n2816 ) | ( n2173 & n8995 ) | ( n2816 & n8995 ) ;
  assign n8997 = n898 | n3806 ;
  assign n8998 = n1485 | n8997 ;
  assign n8999 = n1895 ^ x54 ^ 1'b0 ;
  assign n9000 = n1183 | n8999 ;
  assign n9001 = x39 & n2568 ;
  assign n9002 = n9001 ^ n1034 ^ 1'b0 ;
  assign n9003 = n8860 ^ n1615 ^ 1'b0 ;
  assign n9004 = n1466 & ~n9003 ;
  assign n9005 = n9004 ^ n5942 ^ n4434 ;
  assign n9006 = n9005 ^ n8814 ^ 1'b0 ;
  assign n9007 = n8102 & n9006 ;
  assign n9012 = x68 & ~n1014 ;
  assign n9013 = n9012 ^ n514 ^ 1'b0 ;
  assign n9014 = ( n3395 & n7612 ) | ( n3395 & n9013 ) | ( n7612 & n9013 ) ;
  assign n9015 = ( ~n606 & n4384 ) | ( ~n606 & n5060 ) | ( n4384 & n5060 ) ;
  assign n9016 = ( n2511 & n9014 ) | ( n2511 & ~n9015 ) | ( n9014 & ~n9015 ) ;
  assign n9008 = ( n170 & n3864 ) | ( n170 & n5001 ) | ( n3864 & n5001 ) ;
  assign n9009 = n1674 | n9008 ;
  assign n9010 = n6833 | n9009 ;
  assign n9011 = n4849 & n9010 ;
  assign n9017 = n9016 ^ n9011 ^ 1'b0 ;
  assign n9018 = n7976 ^ n418 ^ 1'b0 ;
  assign n9019 = n6344 ^ n2297 ^ 1'b0 ;
  assign n9021 = ~n4599 & n7098 ;
  assign n9022 = n9021 ^ n4472 ^ n328 ;
  assign n9023 = n9022 ^ n2839 ^ 1'b0 ;
  assign n9024 = n5455 ^ n2053 ^ 1'b0 ;
  assign n9025 = n9023 & n9024 ;
  assign n9020 = n4890 ^ n4042 ^ 1'b0 ;
  assign n9026 = n9025 ^ n9020 ^ 1'b0 ;
  assign n9027 = n5263 ^ n3503 ^ n3393 ;
  assign n9028 = n1354 ^ n867 ^ 1'b0 ;
  assign n9029 = ( n2494 & n5814 ) | ( n2494 & ~n9028 ) | ( n5814 & ~n9028 ) ;
  assign n9030 = n2187 & ~n7981 ;
  assign n9031 = n2338 & n9030 ;
  assign n9033 = ~n705 & n3016 ;
  assign n9032 = n5578 & ~n7243 ;
  assign n9034 = n9033 ^ n9032 ^ 1'b0 ;
  assign n9035 = n5904 ^ n4994 ^ 1'b0 ;
  assign n9036 = n7238 | n9035 ;
  assign n9037 = ~n3257 & n9036 ;
  assign n9038 = n9037 ^ n3864 ^ n971 ;
  assign n9039 = ( n1731 & ~n1935 ) | ( n1731 & n2186 ) | ( ~n1935 & n2186 ) ;
  assign n9040 = ~n3090 & n9039 ;
  assign n9041 = n9038 & n9040 ;
  assign n9042 = ( ~n2915 & n2982 ) | ( ~n2915 & n5967 ) | ( n2982 & n5967 ) ;
  assign n9043 = n2872 & ~n9042 ;
  assign n9044 = n8615 & n9043 ;
  assign n9045 = n1236 & ~n2455 ;
  assign n9046 = n7669 ^ n2021 ^ 1'b0 ;
  assign n9047 = n4688 & n9046 ;
  assign n9048 = n5448 ^ n819 ^ 1'b0 ;
  assign n9049 = ~n4005 & n4443 ;
  assign n9050 = n9049 ^ x13 ^ 1'b0 ;
  assign n9055 = ~n1199 & n2710 ;
  assign n9051 = ~n843 & n1833 ;
  assign n9052 = n9051 ^ n8648 ^ 1'b0 ;
  assign n9053 = n2692 & n9052 ;
  assign n9054 = n9053 ^ n2200 ^ 1'b0 ;
  assign n9056 = n9055 ^ n9054 ^ 1'b0 ;
  assign n9057 = n4697 | n9056 ;
  assign n9058 = n5013 ^ n3848 ^ 1'b0 ;
  assign n9059 = n3957 | n9058 ;
  assign n9060 = ~n260 & n6684 ;
  assign n9061 = n4778 & n7331 ;
  assign n9062 = n9061 ^ n5544 ^ 1'b0 ;
  assign n9063 = n4902 & n9062 ;
  assign n9064 = n2520 & n8690 ;
  assign n9065 = ( ~n4887 & n8250 ) | ( ~n4887 & n9064 ) | ( n8250 & n9064 ) ;
  assign n9066 = ( ~n1586 & n3657 ) | ( ~n1586 & n4256 ) | ( n3657 & n4256 ) ;
  assign n9067 = n648 | n9066 ;
  assign n9068 = n9067 ^ n586 ^ 1'b0 ;
  assign n9069 = n6696 ^ n1102 ^ 1'b0 ;
  assign n9070 = n9068 & ~n9069 ;
  assign n9071 = n9070 ^ n5715 ^ 1'b0 ;
  assign n9072 = n4440 & ~n9071 ;
  assign n9073 = n5554 ^ n3792 ^ 1'b0 ;
  assign n9074 = ~n1927 & n9073 ;
  assign n9075 = n9074 ^ n7998 ^ 1'b0 ;
  assign n9076 = n8746 ^ n2574 ^ 1'b0 ;
  assign n9077 = n568 & n5781 ;
  assign n9078 = n8237 ^ n3063 ^ n3040 ;
  assign n9079 = n4220 ^ n715 ^ 1'b0 ;
  assign n9080 = n3258 | n9079 ;
  assign n9081 = n6527 | n9080 ;
  assign n9082 = n7449 ^ n7123 ^ 1'b0 ;
  assign n9083 = ~n8701 & n9082 ;
  assign n9084 = x78 & ~n2256 ;
  assign n9085 = ~n2066 & n8363 ;
  assign n9086 = n9085 ^ n4770 ^ n4704 ;
  assign n9087 = ( n3886 & n6096 ) | ( n3886 & n9086 ) | ( n6096 & n9086 ) ;
  assign n9088 = n5436 | n7119 ;
  assign n9089 = n8089 | n9088 ;
  assign n9090 = n5876 & n9089 ;
  assign n9091 = ( x13 & n1340 ) | ( x13 & ~n5377 ) | ( n1340 & ~n5377 ) ;
  assign n9092 = ~n865 & n2377 ;
  assign n9093 = n9092 ^ n7828 ^ n1858 ;
  assign n9094 = ( ~n4817 & n6230 ) | ( ~n4817 & n9093 ) | ( n6230 & n9093 ) ;
  assign n9095 = n3448 | n4118 ;
  assign n9096 = n776 | n9095 ;
  assign n9097 = n9096 ^ n1633 ^ n1246 ;
  assign n9103 = n3130 ^ n1893 ^ 1'b0 ;
  assign n9104 = n9073 ^ n2393 ^ 1'b0 ;
  assign n9105 = n9103 | n9104 ;
  assign n9099 = n1326 | n5024 ;
  assign n9100 = n9099 ^ n8519 ^ 1'b0 ;
  assign n9101 = ~n2011 & n9100 ;
  assign n9098 = n266 & n6198 ;
  assign n9102 = n9101 ^ n9098 ^ 1'b0 ;
  assign n9106 = n9105 ^ n9102 ^ n4837 ;
  assign n9107 = n4256 ^ n3597 ^ 1'b0 ;
  assign n9108 = n3203 & ~n9107 ;
  assign n9109 = n9108 ^ n2860 ^ 1'b0 ;
  assign n9110 = n5980 ^ n4065 ^ 1'b0 ;
  assign n9111 = n9110 ^ n8521 ^ n8447 ;
  assign n9114 = n1498 ^ n901 ^ 1'b0 ;
  assign n9112 = ( ~n1974 & n2034 ) | ( ~n1974 & n4826 ) | ( n2034 & n4826 ) ;
  assign n9113 = ( ~n3842 & n5392 ) | ( ~n3842 & n9112 ) | ( n5392 & n9112 ) ;
  assign n9115 = n9114 ^ n9113 ^ 1'b0 ;
  assign n9116 = n8560 & ~n9115 ;
  assign n9117 = n5264 ^ n3507 ^ n1427 ;
  assign n9119 = n5943 ^ n4337 ^ 1'b0 ;
  assign n9120 = n2734 & ~n9119 ;
  assign n9121 = n9120 ^ n1537 ^ 1'b0 ;
  assign n9122 = ( n3905 & n4817 ) | ( n3905 & ~n9121 ) | ( n4817 & ~n9121 ) ;
  assign n9118 = ( ~n1176 & n4753 ) | ( ~n1176 & n5080 ) | ( n4753 & n5080 ) ;
  assign n9123 = n9122 ^ n9118 ^ 1'b0 ;
  assign n9124 = n1272 & n1680 ;
  assign n9125 = n9124 ^ n2734 ^ 1'b0 ;
  assign n9126 = n2851 ^ n2560 ^ n254 ;
  assign n9127 = n1487 & ~n2158 ;
  assign n9128 = n9127 ^ n6149 ^ n3250 ;
  assign n9129 = ~n2898 & n9128 ;
  assign n9130 = n5202 ^ n4952 ^ 1'b0 ;
  assign n9131 = x109 | n3576 ;
  assign n9132 = ( n4955 & n5139 ) | ( n4955 & n9131 ) | ( n5139 & n9131 ) ;
  assign n9134 = n1915 ^ n1741 ^ 1'b0 ;
  assign n9133 = n7490 ^ n878 ^ 1'b0 ;
  assign n9135 = n9134 ^ n9133 ^ n430 ;
  assign n9136 = n9135 ^ n5594 ^ n585 ;
  assign n9137 = ( ~n1715 & n9132 ) | ( ~n1715 & n9136 ) | ( n9132 & n9136 ) ;
  assign n9138 = n7212 & ~n9137 ;
  assign n9139 = n2702 ^ n1448 ^ n809 ;
  assign n9140 = ~n2357 & n9139 ;
  assign n9141 = n9140 ^ n8555 ^ 1'b0 ;
  assign n9142 = n6783 | n9141 ;
  assign n9143 = n2967 | n4935 ;
  assign n9144 = n7894 | n9143 ;
  assign n9145 = n9144 ^ n7455 ^ n3459 ;
  assign n9146 = n9145 ^ n7156 ^ 1'b0 ;
  assign n9147 = ~n3173 & n9146 ;
  assign n9148 = n5500 & n6481 ;
  assign n9149 = ~n9147 & n9148 ;
  assign n9150 = ~n477 & n8856 ;
  assign n9151 = n143 & ~n6654 ;
  assign n9152 = n9151 ^ n7169 ^ n3931 ;
  assign n9153 = ( n4601 & n6835 ) | ( n4601 & ~n9152 ) | ( n6835 & ~n9152 ) ;
  assign n9154 = ( n7301 & n9150 ) | ( n7301 & ~n9153 ) | ( n9150 & ~n9153 ) ;
  assign n9155 = n8255 | n8763 ;
  assign n9157 = n3265 | n4712 ;
  assign n9158 = ~n1358 & n9157 ;
  assign n9156 = n7468 ^ n1800 ^ n880 ;
  assign n9159 = n9158 ^ n9156 ^ n5499 ;
  assign n9160 = n4601 ^ n2609 ^ 1'b0 ;
  assign n9161 = ~n746 & n2614 ;
  assign n9162 = n6462 & n9161 ;
  assign n9163 = n9162 ^ n2688 ^ n520 ;
  assign n9164 = n7377 | n8064 ;
  assign n9165 = n9163 | n9164 ;
  assign n9170 = ~n6525 & n7911 ;
  assign n9167 = n1586 ^ n868 ^ 1'b0 ;
  assign n9166 = n4277 & ~n7038 ;
  assign n9168 = n9167 ^ n9166 ^ 1'b0 ;
  assign n9169 = n9168 ^ n4172 ^ 1'b0 ;
  assign n9171 = n9170 ^ n9169 ^ 1'b0 ;
  assign n9173 = n1610 | n4570 ;
  assign n9172 = n3082 & ~n6132 ;
  assign n9174 = n9173 ^ n9172 ^ 1'b0 ;
  assign n9175 = n1091 & n2421 ;
  assign n9176 = ~n447 & n8724 ;
  assign n9177 = n637 | n9176 ;
  assign n9186 = n6739 ^ n3614 ^ n1262 ;
  assign n9178 = n1186 ^ n843 ^ n649 ;
  assign n9179 = n3865 ^ n3370 ^ 1'b0 ;
  assign n9180 = ~n9178 & n9179 ;
  assign n9181 = n4884 ^ n4472 ^ 1'b0 ;
  assign n9182 = n9180 & ~n9181 ;
  assign n9183 = n9182 ^ n1153 ^ n790 ;
  assign n9184 = ~n5980 & n9183 ;
  assign n9185 = n349 | n9184 ;
  assign n9187 = n9186 ^ n9185 ^ 1'b0 ;
  assign n9188 = ~n6317 & n9187 ;
  assign n9189 = ~n7835 & n9188 ;
  assign n9190 = ~n9177 & n9189 ;
  assign n9191 = n9190 ^ n5355 ^ 1'b0 ;
  assign n9192 = n9175 & n9191 ;
  assign n9193 = ( n7286 & n7916 ) | ( n7286 & n9192 ) | ( n7916 & n9192 ) ;
  assign n9194 = ~n449 & n4123 ;
  assign n9195 = n5056 & n9194 ;
  assign n9196 = ( ~n1420 & n2487 ) | ( ~n1420 & n6477 ) | ( n2487 & n6477 ) ;
  assign n9197 = n6344 ^ n5075 ^ 1'b0 ;
  assign n9198 = n5720 ^ n5317 ^ 1'b0 ;
  assign n9199 = n2489 ^ n1596 ^ 1'b0 ;
  assign n9200 = n9199 ^ n6339 ^ 1'b0 ;
  assign n9201 = n6641 ^ n3239 ^ 1'b0 ;
  assign n9202 = n475 & ~n5139 ;
  assign n9203 = n9202 ^ n7238 ^ 1'b0 ;
  assign n9204 = ( n6571 & n9201 ) | ( n6571 & ~n9203 ) | ( n9201 & ~n9203 ) ;
  assign n9205 = n1495 & n1691 ;
  assign n9206 = n7375 ^ n3430 ^ 1'b0 ;
  assign n9207 = n3969 & ~n9206 ;
  assign n9208 = ~n9205 & n9207 ;
  assign n9209 = n6083 & n8159 ;
  assign n9210 = n2246 ^ n1311 ^ 1'b0 ;
  assign n9211 = n8760 ^ n3330 ^ 1'b0 ;
  assign n9212 = n3248 & ~n9211 ;
  assign n9213 = ~n3731 & n8922 ;
  assign n9214 = ( ~n3652 & n7505 ) | ( ~n3652 & n7820 ) | ( n7505 & n7820 ) ;
  assign n9215 = n9214 ^ n2388 ^ 1'b0 ;
  assign n9216 = n8828 ^ n5272 ^ n4294 ;
  assign n9217 = n3484 ^ n3431 ^ n1370 ;
  assign n9218 = n9216 & n9217 ;
  assign n9219 = n1664 | n4694 ;
  assign n9220 = n5113 & ~n9219 ;
  assign n9221 = ( n1076 & n2618 ) | ( n1076 & ~n8634 ) | ( n2618 & ~n8634 ) ;
  assign n9222 = n9221 ^ n4216 ^ 1'b0 ;
  assign n9223 = ~n2796 & n2893 ;
  assign n9224 = n9013 ^ n4482 ^ 1'b0 ;
  assign n9225 = n882 & ~n9224 ;
  assign n9226 = ( n1678 & ~n5502 ) | ( n1678 & n9225 ) | ( ~n5502 & n9225 ) ;
  assign n9227 = n9223 & n9226 ;
  assign n9229 = n1295 & n3265 ;
  assign n9228 = ( n874 & n1531 ) | ( n874 & n2139 ) | ( n1531 & n2139 ) ;
  assign n9230 = n9229 ^ n9228 ^ 1'b0 ;
  assign n9232 = n891 ^ n515 ^ 1'b0 ;
  assign n9233 = n8877 & n9232 ;
  assign n9231 = n5217 ^ n3834 ^ 1'b0 ;
  assign n9234 = n9233 ^ n9231 ^ 1'b0 ;
  assign n9235 = n3363 ^ x80 ^ 1'b0 ;
  assign n9236 = n189 | n9235 ;
  assign n9237 = n4675 & n9236 ;
  assign n9238 = n9237 ^ n4355 ^ n713 ;
  assign n9239 = n6948 ^ n4621 ^ 1'b0 ;
  assign n9240 = ~n9238 & n9239 ;
  assign n9241 = n658 & n8335 ;
  assign n9242 = n9241 ^ n2066 ^ 1'b0 ;
  assign n9243 = n606 & ~n1579 ;
  assign n9244 = n9243 ^ n2216 ^ 1'b0 ;
  assign n9245 = n1829 & ~n3790 ;
  assign n9246 = n9245 ^ n5502 ^ 1'b0 ;
  assign n9247 = ( n2889 & n9244 ) | ( n2889 & n9246 ) | ( n9244 & n9246 ) ;
  assign n9248 = n152 & ~n284 ;
  assign n9249 = n510 & n9248 ;
  assign n9250 = n2252 ^ n1152 ^ 1'b0 ;
  assign n9251 = n5876 | n9250 ;
  assign n9252 = n2542 & ~n9251 ;
  assign n9253 = n186 | n4792 ;
  assign n9254 = n9253 ^ n7369 ^ 1'b0 ;
  assign n9255 = n4973 ^ n3159 ^ n1015 ;
  assign n9256 = ( n1152 & ~n1617 ) | ( n1152 & n2245 ) | ( ~n1617 & n2245 ) ;
  assign n9257 = n3987 | n9256 ;
  assign n9258 = n2296 & ~n9257 ;
  assign n9259 = ( n4757 & ~n9255 ) | ( n4757 & n9258 ) | ( ~n9255 & n9258 ) ;
  assign n9260 = n5661 ^ n2964 ^ 1'b0 ;
  assign n9261 = n4616 & ~n7075 ;
  assign n9262 = n9261 ^ n289 ^ 1'b0 ;
  assign n9263 = n1175 & n7911 ;
  assign n9264 = n9262 & n9263 ;
  assign n9265 = ~n2858 & n7844 ;
  assign n9266 = n911 & n9265 ;
  assign n9267 = n8086 ^ n7701 ^ x87 ;
  assign n9268 = n4820 ^ n2304 ^ 1'b0 ;
  assign n9269 = n2995 & ~n6258 ;
  assign n9270 = n9269 ^ n9200 ^ 1'b0 ;
  assign n9271 = n3315 ^ n2596 ^ n1626 ;
  assign n9272 = n1843 | n3271 ;
  assign n9273 = n9272 ^ n1027 ^ 1'b0 ;
  assign n9274 = n9273 ^ n1618 ^ 1'b0 ;
  assign n9275 = n9271 & ~n9274 ;
  assign n9276 = n1826 & n9275 ;
  assign n9277 = n9276 ^ n4126 ^ 1'b0 ;
  assign n9278 = n522 & ~n1672 ;
  assign n9279 = n9278 ^ n2551 ^ 1'b0 ;
  assign n9280 = n7621 & ~n9279 ;
  assign n9282 = n1469 | n3898 ;
  assign n9283 = n298 & ~n9282 ;
  assign n9281 = x93 & ~n2619 ;
  assign n9284 = n9283 ^ n9281 ^ 1'b0 ;
  assign n9285 = n7060 ^ n6918 ^ n3104 ;
  assign n9286 = n8099 ^ n6798 ^ n928 ;
  assign n9287 = ~n964 & n4589 ;
  assign n9288 = n8116 & n9287 ;
  assign n9289 = n9288 ^ n2192 ^ 1'b0 ;
  assign n9290 = n773 | n3898 ;
  assign n9291 = n4915 & ~n9290 ;
  assign n9292 = n9291 ^ n2633 ^ n1869 ;
  assign n9293 = n9292 ^ n8773 ^ 1'b0 ;
  assign n9294 = ~n760 & n3789 ;
  assign n9295 = n442 & ~n7160 ;
  assign n9296 = n2083 & n9295 ;
  assign n9297 = n6881 | n9296 ;
  assign n9298 = n9294 & ~n9297 ;
  assign n9299 = n9203 ^ n2361 ^ 1'b0 ;
  assign n9300 = n4521 & n9299 ;
  assign n9310 = ( n781 & ~n2957 ) | ( n781 & n7781 ) | ( ~n2957 & n7781 ) ;
  assign n9301 = n5185 | n7316 ;
  assign n9302 = n1020 | n9301 ;
  assign n9303 = n9302 ^ n3224 ^ n1978 ;
  assign n9304 = n5928 ^ n3174 ^ n2447 ;
  assign n9305 = n509 | n5482 ;
  assign n9306 = n7758 | n9305 ;
  assign n9307 = ~n9304 & n9306 ;
  assign n9308 = n9307 ^ n8486 ^ 1'b0 ;
  assign n9309 = ~n9303 & n9308 ;
  assign n9311 = n9310 ^ n9309 ^ 1'b0 ;
  assign n9312 = n5573 ^ n3483 ^ 1'b0 ;
  assign n9313 = n5612 ^ n4607 ^ n998 ;
  assign n9314 = n3704 ^ n2697 ^ n1480 ;
  assign n9315 = ( n163 & n3352 ) | ( n163 & ~n7006 ) | ( n3352 & ~n7006 ) ;
  assign n9317 = n1512 ^ n967 ^ n304 ;
  assign n9318 = n9317 ^ n2501 ^ 1'b0 ;
  assign n9316 = n6716 ^ n2124 ^ n692 ;
  assign n9319 = n9318 ^ n9316 ^ 1'b0 ;
  assign n9321 = n2032 | n2972 ;
  assign n9322 = n5147 & n9321 ;
  assign n9323 = n1840 & n9322 ;
  assign n9320 = n3410 | n6347 ;
  assign n9324 = n9323 ^ n9320 ^ 1'b0 ;
  assign n9325 = n6262 ^ n4242 ^ n4207 ;
  assign n9326 = n1770 ^ n794 ^ 1'b0 ;
  assign n9327 = n1158 & ~n9326 ;
  assign n9328 = ( ~x41 & n6143 ) | ( ~x41 & n9327 ) | ( n6143 & n9327 ) ;
  assign n9329 = n8543 ^ n2787 ^ n2654 ;
  assign n9330 = n9329 ^ n4614 ^ n1485 ;
  assign n9334 = n2580 ^ n1086 ^ 1'b0 ;
  assign n9335 = ~n7356 & n9334 ;
  assign n9331 = n6605 ^ n5975 ^ 1'b0 ;
  assign n9332 = n3719 | n9331 ;
  assign n9333 = n5008 & ~n9332 ;
  assign n9336 = n9335 ^ n9333 ^ 1'b0 ;
  assign n9337 = n4616 ^ n1653 ^ 1'b0 ;
  assign n9338 = n6810 ^ n4801 ^ 1'b0 ;
  assign n9339 = n2566 & n9338 ;
  assign n9340 = n1368 & n9339 ;
  assign n9341 = n6752 ^ n2382 ^ 1'b0 ;
  assign n9342 = n8179 | n9341 ;
  assign n9343 = n4675 ^ n1397 ^ 1'b0 ;
  assign n9344 = n4530 ^ n209 ^ 1'b0 ;
  assign n9345 = n9343 & n9344 ;
  assign n9346 = n2800 ^ n1799 ^ 1'b0 ;
  assign n9347 = n540 | n9346 ;
  assign n9348 = n8299 ^ n3950 ^ n1715 ;
  assign n9350 = n4724 & ~n5378 ;
  assign n9349 = n4403 & n9058 ;
  assign n9351 = n9350 ^ n9349 ^ 1'b0 ;
  assign n9352 = n2196 & ~n9351 ;
  assign n9353 = n1078 & ~n1575 ;
  assign n9354 = n9353 ^ n4392 ^ 1'b0 ;
  assign n9355 = n2987 & ~n9354 ;
  assign n9356 = n9355 ^ n4349 ^ 1'b0 ;
  assign n9357 = n6125 ^ n4995 ^ 1'b0 ;
  assign n9358 = n9357 ^ x73 ^ 1'b0 ;
  assign n9359 = n9358 ^ n1914 ^ 1'b0 ;
  assign n9360 = n4564 | n8483 ;
  assign n9361 = n9360 ^ n6128 ^ 1'b0 ;
  assign n9362 = n9361 ^ n5360 ^ n4221 ;
  assign n9366 = n3529 | n4264 ;
  assign n9363 = ~n172 & n6365 ;
  assign n9364 = ~n5358 & n9363 ;
  assign n9365 = n6679 & ~n9364 ;
  assign n9367 = n9366 ^ n9365 ^ 1'b0 ;
  assign n9368 = n1689 & n5340 ;
  assign n9369 = n9368 ^ n2326 ^ 1'b0 ;
  assign n9370 = ( ~n2990 & n7375 ) | ( ~n2990 & n9369 ) | ( n7375 & n9369 ) ;
  assign n9371 = n7958 | n9370 ;
  assign n9372 = n6326 ^ n6309 ^ 1'b0 ;
  assign n9373 = n251 & ~n1449 ;
  assign n9374 = n9373 ^ n9342 ^ 1'b0 ;
  assign n9375 = n927 | n6084 ;
  assign n9376 = n4925 & ~n9375 ;
  assign n9377 = ( ~n614 & n2399 ) | ( ~n614 & n9376 ) | ( n2399 & n9376 ) ;
  assign n9378 = n5849 ^ n1776 ^ 1'b0 ;
  assign n9379 = n5453 & ~n9378 ;
  assign n9380 = n9379 ^ n8103 ^ 1'b0 ;
  assign n9381 = n9380 ^ n1794 ^ 1'b0 ;
  assign n9382 = ( n3070 & ~n9110 ) | ( n3070 & n9381 ) | ( ~n9110 & n9381 ) ;
  assign n9385 = n2706 ^ n462 ^ 1'b0 ;
  assign n9383 = n8319 & ~n8817 ;
  assign n9384 = n3563 & ~n9383 ;
  assign n9386 = n9385 ^ n9384 ^ 1'b0 ;
  assign n9387 = n6837 ^ n1485 ^ 1'b0 ;
  assign n9388 = n5961 & ~n9387 ;
  assign n9389 = n2278 & n3686 ;
  assign n9390 = n9389 ^ n2530 ^ 1'b0 ;
  assign n9391 = n9390 ^ n2236 ^ 1'b0 ;
  assign n9392 = n1969 | n9391 ;
  assign n9393 = n1162 & ~n2389 ;
  assign n9394 = n9393 ^ n8113 ^ 1'b0 ;
  assign n9395 = n9392 | n9394 ;
  assign n9396 = n4556 | n5354 ;
  assign n9397 = n9396 ^ n6282 ^ 1'b0 ;
  assign n9398 = n8539 ^ n3059 ^ 1'b0 ;
  assign n9399 = ( n1714 & n3323 ) | ( n1714 & ~n7695 ) | ( n3323 & ~n7695 ) ;
  assign n9400 = n1706 ^ n1375 ^ 1'b0 ;
  assign n9401 = n3012 ^ n1972 ^ n1312 ;
  assign n9402 = ( ~n5873 & n8328 ) | ( ~n5873 & n9401 ) | ( n8328 & n9401 ) ;
  assign n9403 = n2397 & ~n4757 ;
  assign n9404 = n9402 & n9403 ;
  assign n9405 = ~n4853 & n5385 ;
  assign n9411 = ~n692 & n2553 ;
  assign n9412 = ~n1131 & n9411 ;
  assign n9406 = n5128 ^ n5094 ^ n3616 ;
  assign n9407 = n4161 ^ n4045 ^ n1861 ;
  assign n9408 = n9407 ^ n531 ^ 1'b0 ;
  assign n9409 = n9406 & ~n9408 ;
  assign n9410 = ~n4938 & n9409 ;
  assign n9413 = n9412 ^ n9410 ^ 1'b0 ;
  assign n9414 = ~n2761 & n9413 ;
  assign n9415 = n2817 | n3030 ;
  assign n9416 = n9415 ^ n5561 ^ 1'b0 ;
  assign n9417 = n9416 ^ n4862 ^ 1'b0 ;
  assign n9418 = n1360 & n9417 ;
  assign n9419 = n9418 ^ n5356 ^ 1'b0 ;
  assign n9420 = n1851 | n9419 ;
  assign n9421 = ( ~n5372 & n6756 ) | ( ~n5372 & n9420 ) | ( n6756 & n9420 ) ;
  assign n9422 = n9421 ^ n9077 ^ 1'b0 ;
  assign n9423 = n1220 ^ n146 ^ 1'b0 ;
  assign n9424 = n2449 & n9423 ;
  assign n9425 = n9424 ^ n1679 ^ 1'b0 ;
  assign n9426 = n1218 & ~n9425 ;
  assign n9427 = ( ~n3155 & n3384 ) | ( ~n3155 & n7510 ) | ( n3384 & n7510 ) ;
  assign n9428 = n704 | n9427 ;
  assign n9429 = n9428 ^ n143 ^ 1'b0 ;
  assign n9430 = n9429 ^ n9081 ^ 1'b0 ;
  assign n9431 = n9426 & ~n9430 ;
  assign n9432 = ( n2335 & n2425 ) | ( n2335 & n3342 ) | ( n2425 & n3342 ) ;
  assign n9433 = ( ~n607 & n9271 ) | ( ~n607 & n9432 ) | ( n9271 & n9432 ) ;
  assign n9435 = n7266 ^ n1074 ^ 1'b0 ;
  assign n9436 = n9435 ^ n1851 ^ n1498 ;
  assign n9437 = n9436 ^ n8988 ^ n7524 ;
  assign n9434 = n5548 ^ n4139 ^ n2011 ;
  assign n9438 = n9437 ^ n9434 ^ n7097 ;
  assign n9439 = n3140 ^ n2772 ^ n903 ;
  assign n9440 = n1718 & n9439 ;
  assign n9441 = n2909 ^ n1588 ^ n936 ;
  assign n9442 = n3955 ^ n1049 ^ 1'b0 ;
  assign n9443 = n9441 & ~n9442 ;
  assign n9444 = ~n2236 & n3058 ;
  assign n9445 = n9444 ^ n974 ^ 1'b0 ;
  assign n9446 = n6059 | n9445 ;
  assign n9447 = n9446 ^ n3114 ^ 1'b0 ;
  assign n9448 = ~n2127 & n9447 ;
  assign n9449 = n8953 | n9448 ;
  assign n9450 = n6370 ^ n5901 ^ n893 ;
  assign n9451 = ( n3950 & n3968 ) | ( n3950 & n6268 ) | ( n3968 & n6268 ) ;
  assign n9452 = n617 | n9451 ;
  assign n9453 = n1514 & n9452 ;
  assign n9454 = n9453 ^ n4810 ^ 1'b0 ;
  assign n9459 = ~n474 & n6851 ;
  assign n9460 = ~n4864 & n9459 ;
  assign n9455 = n3016 ^ n2460 ^ n1352 ;
  assign n9456 = n9455 ^ n8386 ^ n3063 ;
  assign n9457 = n9456 ^ n5702 ^ 1'b0 ;
  assign n9458 = ~n681 & n9457 ;
  assign n9461 = n9460 ^ n9458 ^ n1280 ;
  assign n9462 = n1582 & n2386 ;
  assign n9463 = n5306 & n9462 ;
  assign n9464 = n9463 ^ n3095 ^ 1'b0 ;
  assign n9465 = n9464 ^ n6462 ^ 1'b0 ;
  assign n9466 = n2869 | n3044 ;
  assign n9467 = n8746 & ~n9466 ;
  assign n9468 = n5320 | n9467 ;
  assign n9469 = n7077 & ~n9468 ;
  assign n9470 = n9465 | n9469 ;
  assign n9471 = n3157 ^ n320 ^ 1'b0 ;
  assign n9472 = n2090 & n9471 ;
  assign n9473 = n7238 | n9472 ;
  assign n9474 = n9473 ^ n7258 ^ 1'b0 ;
  assign n9475 = ( ~n4065 & n4753 ) | ( ~n4065 & n7034 ) | ( n4753 & n7034 ) ;
  assign n9476 = n4158 & ~n9475 ;
  assign n9477 = n9476 ^ n4250 ^ n1577 ;
  assign n9482 = n3406 | n3713 ;
  assign n9479 = ~n440 & n3104 ;
  assign n9480 = n9479 ^ n232 ^ 1'b0 ;
  assign n9481 = n8933 & n9480 ;
  assign n9483 = n9482 ^ n9481 ^ n4104 ;
  assign n9478 = ( ~n2435 & n2930 ) | ( ~n2435 & n4249 ) | ( n2930 & n4249 ) ;
  assign n9484 = n9483 ^ n9478 ^ 1'b0 ;
  assign n9485 = n9477 | n9484 ;
  assign n9487 = ( n5915 & ~n7355 ) | ( n5915 & n9401 ) | ( ~n7355 & n9401 ) ;
  assign n9486 = ( n232 & n6982 ) | ( n232 & n7618 ) | ( n6982 & n7618 ) ;
  assign n9488 = n9487 ^ n9486 ^ n3946 ;
  assign n9489 = n7392 & n9233 ;
  assign n9490 = n8536 & n9489 ;
  assign n9491 = ~n1603 & n2395 ;
  assign n9492 = n9491 ^ n260 ^ 1'b0 ;
  assign n9493 = n2926 ^ n1709 ^ n1374 ;
  assign n9494 = ( n7130 & ~n9492 ) | ( n7130 & n9493 ) | ( ~n9492 & n9493 ) ;
  assign n9495 = n7603 ^ n4102 ^ 1'b0 ;
  assign n9496 = n1545 & n2268 ;
  assign n9497 = ( n9303 & n9495 ) | ( n9303 & n9496 ) | ( n9495 & n9496 ) ;
  assign n9502 = n867 | n1521 ;
  assign n9503 = ( ~n2098 & n4385 ) | ( ~n2098 & n9502 ) | ( n4385 & n9502 ) ;
  assign n9504 = n9503 ^ n654 ^ 1'b0 ;
  assign n9498 = n1988 & ~n2877 ;
  assign n9499 = ~n2527 & n9498 ;
  assign n9500 = n1525 & ~n9499 ;
  assign n9501 = ~n3726 & n9500 ;
  assign n9505 = n9504 ^ n9501 ^ n2054 ;
  assign n9506 = n2215 & n2658 ;
  assign n9507 = n9506 ^ n2679 ^ 1'b0 ;
  assign n9508 = n1868 ^ n485 ^ 1'b0 ;
  assign n9509 = n778 | n9508 ;
  assign n9510 = ( ~n6047 & n8736 ) | ( ~n6047 & n9509 ) | ( n8736 & n9509 ) ;
  assign n9511 = n3465 | n9510 ;
  assign n9512 = n9507 & ~n9511 ;
  assign n9513 = n616 & n4966 ;
  assign n9514 = n2030 | n9513 ;
  assign n9515 = n4686 ^ n4147 ^ 1'b0 ;
  assign n9516 = n3856 & ~n9515 ;
  assign n9517 = ~n6321 & n9516 ;
  assign n9518 = n9517 ^ n3753 ^ 1'b0 ;
  assign n9519 = n9480 ^ n207 ^ 1'b0 ;
  assign n9520 = n2060 & ~n2172 ;
  assign n9521 = n9520 ^ n1207 ^ 1'b0 ;
  assign n9522 = n2021 | n7254 ;
  assign n9523 = ( n6255 & n6654 ) | ( n6255 & n9522 ) | ( n6654 & n9522 ) ;
  assign n9524 = ~n6103 & n7716 ;
  assign n9525 = n3722 | n9524 ;
  assign n9526 = n9525 ^ n3482 ^ 1'b0 ;
  assign n9527 = n9526 ^ n6746 ^ 1'b0 ;
  assign n9528 = n9523 | n9527 ;
  assign n9529 = n6603 ^ n6367 ^ 1'b0 ;
  assign n9530 = n6315 & ~n9529 ;
  assign n9532 = x80 & n6586 ;
  assign n9533 = ( n2504 & n2961 ) | ( n2504 & ~n9532 ) | ( n2961 & ~n9532 ) ;
  assign n9534 = ~n836 & n1506 ;
  assign n9535 = n9533 & n9534 ;
  assign n9531 = n1999 | n6169 ;
  assign n9536 = n9535 ^ n9531 ^ 1'b0 ;
  assign n9537 = n9536 ^ n8615 ^ 1'b0 ;
  assign n9538 = n9530 & n9537 ;
  assign n9539 = n4726 ^ n1629 ^ 1'b0 ;
  assign n9540 = n9539 ^ n3802 ^ 1'b0 ;
  assign n9541 = n8686 ^ n3652 ^ 1'b0 ;
  assign n9542 = n4887 | n9541 ;
  assign n9543 = n1740 ^ n1108 ^ 1'b0 ;
  assign n9544 = n4881 | n9543 ;
  assign n9545 = n9544 ^ n1633 ^ 1'b0 ;
  assign n9546 = n7331 ^ n6628 ^ n1008 ;
  assign n9548 = ( n786 & ~n1190 ) | ( n786 & n5565 ) | ( ~n1190 & n5565 ) ;
  assign n9549 = n6609 ^ n3337 ^ 1'b0 ;
  assign n9550 = n9548 & ~n9549 ;
  assign n9547 = ( n5409 & n6198 ) | ( n5409 & n8929 ) | ( n6198 & n8929 ) ;
  assign n9551 = n9550 ^ n9547 ^ 1'b0 ;
  assign n9552 = ~n9546 & n9551 ;
  assign n9555 = n2923 ^ n2300 ^ 1'b0 ;
  assign n9553 = n3017 ^ n2687 ^ 1'b0 ;
  assign n9554 = n553 | n9553 ;
  assign n9556 = n9555 ^ n9554 ^ 1'b0 ;
  assign n9557 = n7507 ^ n1969 ^ 1'b0 ;
  assign n9558 = n4174 ^ n1272 ^ 1'b0 ;
  assign n9559 = n1304 & ~n1927 ;
  assign n9560 = n509 & n9559 ;
  assign n9561 = n9560 ^ n7938 ^ 1'b0 ;
  assign n9562 = n9558 & n9561 ;
  assign n9563 = n9557 & ~n9562 ;
  assign n9564 = n9563 ^ n3766 ^ 1'b0 ;
  assign n9565 = ( ~n2099 & n3482 ) | ( ~n2099 & n9564 ) | ( n3482 & n9564 ) ;
  assign n9566 = ( n5300 & ~n6437 ) | ( n5300 & n8875 ) | ( ~n6437 & n8875 ) ;
  assign n9568 = n3050 & n6285 ;
  assign n9569 = n4102 & n9568 ;
  assign n9567 = n1220 & n6792 ;
  assign n9570 = n9569 ^ n9567 ^ 1'b0 ;
  assign n9571 = n2759 ^ n1300 ^ n1185 ;
  assign n9572 = n1041 & ~n9571 ;
  assign n9573 = n6527 ^ n4352 ^ n3753 ;
  assign n9574 = n9451 & ~n9573 ;
  assign n9575 = ~n2706 & n9574 ;
  assign n9576 = n9527 & ~n9575 ;
  assign n9577 = ~n1043 & n9576 ;
  assign n9578 = n2250 | n2515 ;
  assign n9579 = n2247 | n9578 ;
  assign n9580 = ~n1651 & n9579 ;
  assign n9581 = n3501 | n9580 ;
  assign n9582 = n3252 & ~n4811 ;
  assign n9583 = ~n487 & n9582 ;
  assign n9584 = n3831 ^ n1878 ^ 1'b0 ;
  assign n9585 = n4148 & n9584 ;
  assign n9586 = ( n1905 & n3834 ) | ( n1905 & ~n5522 ) | ( n3834 & ~n5522 ) ;
  assign n9587 = n3410 & n9586 ;
  assign n9588 = n5369 & n8511 ;
  assign n9589 = ( n344 & n6228 ) | ( n344 & n8796 ) | ( n6228 & n8796 ) ;
  assign n9590 = n9073 ^ n6521 ^ 1'b0 ;
  assign n9591 = n197 & ~n2706 ;
  assign n9592 = n6634 | n9591 ;
  assign n9593 = n5335 | n9592 ;
  assign n9594 = ~n7839 & n9593 ;
  assign n9595 = n7760 & n9594 ;
  assign n9596 = n675 & n9595 ;
  assign n9597 = n442 & ~n1240 ;
  assign n9598 = n9597 ^ n173 ^ 1'b0 ;
  assign n9599 = ~x101 & n9598 ;
  assign n9600 = n9599 ^ n3159 ^ 1'b0 ;
  assign n9601 = n1386 & n6852 ;
  assign n9602 = n1666 & n5845 ;
  assign n9603 = n9601 & n9602 ;
  assign n9605 = ( n1205 & n3140 ) | ( n1205 & n4419 ) | ( n3140 & n4419 ) ;
  assign n9604 = n7928 ^ n3567 ^ x84 ;
  assign n9606 = n9605 ^ n9604 ^ 1'b0 ;
  assign n9607 = n3679 ^ n358 ^ 1'b0 ;
  assign n9608 = n2614 & n6072 ;
  assign n9609 = n9608 ^ n6258 ^ 1'b0 ;
  assign n9610 = n9609 ^ n6045 ^ 1'b0 ;
  assign n9611 = n4806 & n4946 ;
  assign n9612 = n5740 & n9611 ;
  assign n9613 = ~n3189 & n9612 ;
  assign n9614 = n4069 ^ x65 ^ 1'b0 ;
  assign n9615 = n1152 & n5665 ;
  assign n9616 = n9615 ^ n4631 ^ 1'b0 ;
  assign n9617 = n4757 & n9616 ;
  assign n9618 = ( ~n936 & n5131 ) | ( ~n936 & n9617 ) | ( n5131 & n9617 ) ;
  assign n9619 = n4419 ^ n397 ^ 1'b0 ;
  assign n9620 = ( ~n968 & n2806 ) | ( ~n968 & n9619 ) | ( n2806 & n9619 ) ;
  assign n9621 = n1057 & ~n9620 ;
  assign n9622 = n9621 ^ n6794 ^ 1'b0 ;
  assign n9623 = n3218 ^ n308 ^ 1'b0 ;
  assign n9624 = n2009 | n9623 ;
  assign n9625 = n1084 | n9624 ;
  assign n9626 = n2527 ^ n1279 ^ n925 ;
  assign n9627 = n2315 ^ n491 ^ 1'b0 ;
  assign n9628 = n6288 & n9627 ;
  assign n9629 = n2721 & ~n3560 ;
  assign n9630 = ~n9628 & n9629 ;
  assign n9631 = n2984 ^ n2316 ^ 1'b0 ;
  assign n9632 = n971 & n9631 ;
  assign n9633 = ( n2291 & n3436 ) | ( n2291 & ~n9632 ) | ( n3436 & ~n9632 ) ;
  assign n9634 = n9630 | n9633 ;
  assign n9635 = n9409 ^ n8186 ^ 1'b0 ;
  assign n9638 = n3796 ^ n1608 ^ n831 ;
  assign n9636 = n4018 ^ n411 ^ 1'b0 ;
  assign n9637 = n3941 & n9636 ;
  assign n9639 = n9638 ^ n9637 ^ n839 ;
  assign n9640 = n2364 & n7782 ;
  assign n9641 = n6500 ^ n917 ^ 1'b0 ;
  assign n9642 = n8097 ^ n4190 ^ 1'b0 ;
  assign n9643 = n1125 & ~n9642 ;
  assign n9644 = n8856 ^ n727 ^ 1'b0 ;
  assign n9646 = n8473 ^ n903 ^ 1'b0 ;
  assign n9645 = n9072 ^ n4469 ^ n1079 ;
  assign n9647 = n9646 ^ n9645 ^ 1'b0 ;
  assign n9649 = n3630 ^ n2758 ^ n1023 ;
  assign n9650 = ~n4404 & n9649 ;
  assign n9651 = ~n3477 & n9650 ;
  assign n9648 = n1677 & n7166 ;
  assign n9652 = n9651 ^ n9648 ^ 1'b0 ;
  assign n9653 = n4644 | n9652 ;
  assign n9654 = ~n2574 & n3359 ;
  assign n9655 = n9654 ^ n2478 ^ 1'b0 ;
  assign n9656 = n9383 ^ n5937 ^ 1'b0 ;
  assign n9657 = ( ~n6572 & n8390 ) | ( ~n6572 & n9656 ) | ( n8390 & n9656 ) ;
  assign n9658 = n5671 ^ n847 ^ 1'b0 ;
  assign n9659 = ( n853 & n5053 ) | ( n853 & n9658 ) | ( n5053 & n9658 ) ;
  assign n9660 = ( ~n2417 & n3563 ) | ( ~n2417 & n4607 ) | ( n3563 & n4607 ) ;
  assign n9661 = n6010 & ~n8891 ;
  assign n9662 = ~n6143 & n9661 ;
  assign n9663 = n9662 ^ n5260 ^ 1'b0 ;
  assign n9664 = n9660 & ~n9663 ;
  assign n9665 = ( n381 & n3694 ) | ( n381 & n6407 ) | ( n3694 & n6407 ) ;
  assign n9666 = n3294 ^ n3082 ^ 1'b0 ;
  assign n9667 = n9665 | n9666 ;
  assign n9668 = n7170 ^ n2023 ^ 1'b0 ;
  assign n9669 = n3955 ^ n2121 ^ 1'b0 ;
  assign n9670 = ( n7479 & n9668 ) | ( n7479 & ~n9669 ) | ( n9668 & ~n9669 ) ;
  assign n9677 = ~n1920 & n7293 ;
  assign n9678 = n154 & n9677 ;
  assign n9679 = ( ~n2492 & n3726 ) | ( ~n2492 & n9678 ) | ( n3726 & n9678 ) ;
  assign n9680 = n4593 ^ n2976 ^ 1'b0 ;
  assign n9681 = n9680 ^ n4562 ^ 1'b0 ;
  assign n9682 = n9679 | n9681 ;
  assign n9683 = n7702 & ~n9682 ;
  assign n9673 = n1490 & ~n8319 ;
  assign n9674 = ( n8900 & n9668 ) | ( n8900 & n9673 ) | ( n9668 & n9673 ) ;
  assign n9671 = n6256 ^ n2680 ^ 1'b0 ;
  assign n9672 = ~n5417 & n9671 ;
  assign n9675 = n9674 ^ n9672 ^ 1'b0 ;
  assign n9676 = n9675 ^ n4988 ^ 1'b0 ;
  assign n9684 = n9683 ^ n9676 ^ 1'b0 ;
  assign n9685 = n5119 | n9684 ;
  assign n9686 = n1633 & ~n4061 ;
  assign n9687 = n9686 ^ n1201 ^ 1'b0 ;
  assign n9688 = ( ~n290 & n715 ) | ( ~n290 & n4793 ) | ( n715 & n4793 ) ;
  assign n9689 = n4367 | n5159 ;
  assign n9690 = n4724 & n9689 ;
  assign n9691 = ~n9688 & n9690 ;
  assign n9692 = ~n5059 & n5676 ;
  assign n9693 = n8310 ^ n6084 ^ x31 ;
  assign n9694 = ~n614 & n4447 ;
  assign n9695 = n9694 ^ n692 ^ 1'b0 ;
  assign n9696 = ~n1664 & n9447 ;
  assign n9697 = n1729 | n6924 ;
  assign n9698 = n5548 & n9697 ;
  assign n9699 = n9698 ^ n585 ^ 1'b0 ;
  assign n9700 = n5962 ^ n609 ^ 1'b0 ;
  assign n9701 = n9700 ^ n6169 ^ n5715 ;
  assign n9702 = n307 | n2640 ;
  assign n9703 = n143 & ~n4717 ;
  assign n9704 = n9703 ^ n5754 ^ 1'b0 ;
  assign n9705 = n9704 ^ n8523 ^ 1'b0 ;
  assign n9706 = ~n6454 & n9705 ;
  assign n9707 = ~n9702 & n9706 ;
  assign n9708 = n7255 | n9707 ;
  assign n9709 = ( n948 & ~n1418 ) | ( n948 & n2695 ) | ( ~n1418 & n2695 ) ;
  assign n9710 = n897 & ~n9709 ;
  assign n9711 = n3023 ^ n2654 ^ 1'b0 ;
  assign n9712 = n4263 ^ n1760 ^ 1'b0 ;
  assign n9713 = ~n9711 & n9712 ;
  assign n9714 = ~n9710 & n9713 ;
  assign n9715 = n9628 ^ n5552 ^ n5045 ;
  assign n9716 = n9715 ^ n908 ^ 1'b0 ;
  assign n9717 = ~n1810 & n7916 ;
  assign n9718 = n6724 ^ n6230 ^ 1'b0 ;
  assign n9719 = n6600 & ~n9718 ;
  assign n9720 = n4296 ^ n974 ^ 1'b0 ;
  assign n9721 = n1535 & ~n9720 ;
  assign n9722 = ~n2826 & n5018 ;
  assign n9723 = n9722 ^ n6297 ^ 1'b0 ;
  assign n9724 = n2905 ^ n2115 ^ 1'b0 ;
  assign n9725 = n6872 & ~n9724 ;
  assign n9726 = ( n143 & n3575 ) | ( n143 & n9725 ) | ( n3575 & n9725 ) ;
  assign n9727 = ( n893 & n1552 ) | ( n893 & n8004 ) | ( n1552 & n8004 ) ;
  assign n9728 = ( n2191 & n5078 ) | ( n2191 & n5984 ) | ( n5078 & n5984 ) ;
  assign n9729 = n6508 | n9728 ;
  assign n9732 = n8125 ^ n4382 ^ 1'b0 ;
  assign n9730 = n9384 ^ n5847 ^ n1378 ;
  assign n9731 = ( n2406 & ~n5178 ) | ( n2406 & n9730 ) | ( ~n5178 & n9730 ) ;
  assign n9733 = n9732 ^ n9731 ^ 1'b0 ;
  assign n9734 = n3716 ^ n3704 ^ n1695 ;
  assign n9735 = x125 ^ x23 ^ 1'b0 ;
  assign n9736 = ~n4051 & n9735 ;
  assign n9737 = n1037 & n9736 ;
  assign n9738 = ~n1740 & n9737 ;
  assign n9739 = n4016 & n4286 ;
  assign n9740 = n9739 ^ n9452 ^ 1'b0 ;
  assign n9741 = n3905 & n4753 ;
  assign n9742 = ~n1226 & n9741 ;
  assign n9743 = n8823 ^ n4922 ^ n4104 ;
  assign n9744 = n5426 & ~n9743 ;
  assign n9745 = n4708 | n9744 ;
  assign n9746 = ~n2323 & n5650 ;
  assign n9747 = n4121 ^ n3154 ^ n1718 ;
  assign n9748 = ( n881 & n9746 ) | ( n881 & ~n9747 ) | ( n9746 & ~n9747 ) ;
  assign n9749 = ~n182 & n1080 ;
  assign n9750 = n4824 & ~n8631 ;
  assign n9751 = n9750 ^ n4909 ^ 1'b0 ;
  assign n9752 = n8112 ^ n6758 ^ n6648 ;
  assign n9753 = ~n9577 & n9752 ;
  assign n9754 = n1508 & n3856 ;
  assign n9755 = n9754 ^ n5299 ^ 1'b0 ;
  assign n9756 = n8237 & ~n9755 ;
  assign n9758 = n1327 | n2965 ;
  assign n9759 = n9758 ^ n4236 ^ 1'b0 ;
  assign n9757 = n2997 & n3610 ;
  assign n9760 = n9759 ^ n9757 ^ 1'b0 ;
  assign n9761 = n391 | n9760 ;
  assign n9762 = n8040 & ~n9761 ;
  assign n9763 = ( n6497 & n6629 ) | ( n6497 & ~n9762 ) | ( n6629 & ~n9762 ) ;
  assign n9764 = n5399 ^ n1154 ^ n600 ;
  assign n9765 = n9764 ^ n5074 ^ 1'b0 ;
  assign n9766 = ~n8580 & n9765 ;
  assign n9767 = n1887 & n3568 ;
  assign n9768 = ~n2462 & n9767 ;
  assign n9770 = n4012 ^ n2407 ^ n1691 ;
  assign n9769 = n4057 | n6388 ;
  assign n9771 = n9770 ^ n9769 ^ n9447 ;
  assign n9774 = n5121 ^ n4562 ^ 1'b0 ;
  assign n9775 = n8174 & ~n9774 ;
  assign n9772 = ~n3845 & n8376 ;
  assign n9773 = ~n4161 & n9772 ;
  assign n9776 = n9775 ^ n9773 ^ 1'b0 ;
  assign n9777 = n7141 & n9505 ;
  assign n9778 = ~n5500 & n9777 ;
  assign n9779 = n7864 ^ n1918 ^ 1'b0 ;
  assign n9780 = n2040 & n9779 ;
  assign n9781 = n9780 ^ n3058 ^ n1498 ;
  assign n9782 = n576 | n9781 ;
  assign n9783 = n9782 ^ n5013 ^ 1'b0 ;
  assign n9784 = n6273 ^ n5921 ^ 1'b0 ;
  assign n9785 = ( n4967 & n5397 ) | ( n4967 & ~n7087 ) | ( n5397 & ~n7087 ) ;
  assign n9786 = n9784 & n9785 ;
  assign n9788 = ( n1274 & ~n1791 ) | ( n1274 & n2105 ) | ( ~n1791 & n2105 ) ;
  assign n9787 = n8532 ^ n7650 ^ n1444 ;
  assign n9789 = n9788 ^ n9787 ^ 1'b0 ;
  assign n9790 = n4091 & ~n9789 ;
  assign n9791 = n3988 ^ n1110 ^ 1'b0 ;
  assign n9792 = ( n465 & ~n9352 ) | ( n465 & n9791 ) | ( ~n9352 & n9791 ) ;
  assign n9793 = n5732 ^ n1714 ^ n353 ;
  assign n9794 = ( n1867 & n1929 ) | ( n1867 & n2614 ) | ( n1929 & n2614 ) ;
  assign n9795 = n6237 ^ n857 ^ 1'b0 ;
  assign n9796 = n9795 ^ n1218 ^ 1'b0 ;
  assign n9797 = ~n9794 & n9796 ;
  assign n9798 = n9793 & n9797 ;
  assign n9799 = n9792 & n9798 ;
  assign n9800 = ~n1615 & n3964 ;
  assign n9801 = n950 & n9800 ;
  assign n9802 = n9801 ^ n7718 ^ n1665 ;
  assign n9803 = n3198 & ~n9802 ;
  assign n9804 = n1782 ^ n1029 ^ 1'b0 ;
  assign n9805 = n9803 & ~n9804 ;
  assign n9806 = n4029 & ~n7534 ;
  assign n9807 = n6200 ^ n2740 ^ n160 ;
  assign n9808 = ~n1776 & n6198 ;
  assign n9809 = n9808 ^ n2056 ^ 1'b0 ;
  assign n9810 = n9809 ^ n2462 ^ 1'b0 ;
  assign n9811 = n8569 ^ n1249 ^ 1'b0 ;
  assign n9812 = x105 & ~n9811 ;
  assign n9813 = n2580 | n9812 ;
  assign n9820 = n1936 | n3589 ;
  assign n9818 = n794 | n2641 ;
  assign n9819 = n7170 | n9818 ;
  assign n9821 = n9820 ^ n9819 ^ 1'b0 ;
  assign n9822 = n9464 ^ n3140 ^ 1'b0 ;
  assign n9823 = n9821 | n9822 ;
  assign n9814 = n3203 & ~n6325 ;
  assign n9815 = n9814 ^ n3616 ^ 1'b0 ;
  assign n9816 = n7740 & ~n9815 ;
  assign n9817 = ~n8669 & n9816 ;
  assign n9824 = n9823 ^ n9817 ^ 1'b0 ;
  assign n9825 = n7223 ^ n2422 ^ 1'b0 ;
  assign n9826 = n6088 ^ n2183 ^ n225 ;
  assign n9827 = n7063 ^ n4679 ^ n219 ;
  assign n9828 = ( ~n7572 & n9015 ) | ( ~n7572 & n9127 ) | ( n9015 & n9127 ) ;
  assign n9830 = n444 & ~n608 ;
  assign n9831 = n9830 ^ n1744 ^ 1'b0 ;
  assign n9832 = n9831 ^ n3615 ^ 1'b0 ;
  assign n9833 = ~n938 & n9832 ;
  assign n9834 = n4694 ^ n3999 ^ 1'b0 ;
  assign n9835 = n9833 & ~n9834 ;
  assign n9829 = n265 & n1201 ;
  assign n9836 = n9835 ^ n9829 ^ 1'b0 ;
  assign n9837 = n6875 | n8812 ;
  assign n9838 = n7475 ^ n2665 ^ n782 ;
  assign n9839 = n9838 ^ n4710 ^ 1'b0 ;
  assign n9840 = ~n473 & n9839 ;
  assign n9841 = n9840 ^ n438 ^ 1'b0 ;
  assign n9842 = n2999 | n5883 ;
  assign n9843 = n7133 & ~n9842 ;
  assign n9844 = ( n6796 & n9841 ) | ( n6796 & n9843 ) | ( n9841 & n9843 ) ;
  assign n9845 = ( ~x102 & n402 ) | ( ~x102 & n1956 ) | ( n402 & n1956 ) ;
  assign n9846 = ( n5104 & n8253 ) | ( n5104 & n9845 ) | ( n8253 & n9845 ) ;
  assign n9847 = n1136 ^ n778 ^ n694 ;
  assign n9848 = ~n3648 & n9847 ;
  assign n9849 = n6862 & n9848 ;
  assign n9850 = ~n9846 & n9849 ;
  assign n9851 = ( n3446 & n5139 ) | ( n3446 & ~n9850 ) | ( n5139 & ~n9850 ) ;
  assign n9852 = n7873 ^ n3710 ^ 1'b0 ;
  assign n9853 = n7703 ^ n5721 ^ n2860 ;
  assign n9854 = n6515 ^ n2846 ^ n1199 ;
  assign n9855 = ( n3343 & n5681 ) | ( n3343 & ~n7834 ) | ( n5681 & ~n7834 ) ;
  assign n9856 = n9855 ^ n3040 ^ n1125 ;
  assign n9864 = n2026 ^ n1970 ^ n1519 ;
  assign n9865 = n3195 | n9864 ;
  assign n9866 = n9865 ^ n2264 ^ 1'b0 ;
  assign n9867 = n897 & ~n9866 ;
  assign n9868 = n9867 ^ n309 ^ 1'b0 ;
  assign n9859 = n381 ^ x125 ^ 1'b0 ;
  assign n9860 = ( n1045 & n4026 ) | ( n1045 & ~n9859 ) | ( n4026 & ~n9859 ) ;
  assign n9857 = n2200 ^ n337 ^ 1'b0 ;
  assign n9858 = n8991 | n9857 ;
  assign n9861 = n9860 ^ n9858 ^ 1'b0 ;
  assign n9862 = n8884 | n9861 ;
  assign n9863 = n3449 | n9862 ;
  assign n9869 = n9868 ^ n9863 ^ 1'b0 ;
  assign n9870 = ~n885 & n2653 ;
  assign n9871 = n9870 ^ n4252 ^ 1'b0 ;
  assign n9872 = n143 ^ x38 ^ x4 ;
  assign n9873 = ( n920 & n1316 ) | ( n920 & n9872 ) | ( n1316 & n9872 ) ;
  assign n9874 = n9873 ^ n1476 ^ n729 ;
  assign n9875 = n3215 ^ n3001 ^ 1'b0 ;
  assign n9876 = n9875 ^ n7516 ^ n2000 ;
  assign n9877 = n5517 | n6818 ;
  assign n9878 = n9876 | n9877 ;
  assign n9879 = n9878 ^ n631 ^ 1'b0 ;
  assign n9880 = n207 | n3037 ;
  assign n9881 = ( ~n3974 & n5610 ) | ( ~n3974 & n7860 ) | ( n5610 & n7860 ) ;
  assign n9882 = n4206 & n6423 ;
  assign n9883 = ~n9881 & n9882 ;
  assign n9884 = n9883 ^ n1692 ^ 1'b0 ;
  assign n9886 = n2118 & n5990 ;
  assign n9887 = ~n521 & n9886 ;
  assign n9885 = n5074 & ~n7613 ;
  assign n9888 = n9887 ^ n9885 ^ 1'b0 ;
  assign n9889 = n5130 ^ n4498 ^ 1'b0 ;
  assign n9890 = n620 | n9889 ;
  assign n9891 = n9890 ^ n181 ^ 1'b0 ;
  assign n9892 = n8170 ^ n1141 ^ 1'b0 ;
  assign n9893 = n2902 ^ n1999 ^ 1'b0 ;
  assign n9894 = n9892 & n9893 ;
  assign n9895 = n9894 ^ n199 ^ 1'b0 ;
  assign n9896 = n673 & n9493 ;
  assign n9897 = n7713 & ~n8304 ;
  assign n9898 = n9897 ^ n1463 ^ 1'b0 ;
  assign n9899 = n3423 ^ n3166 ^ 1'b0 ;
  assign n9900 = n8487 | n9899 ;
  assign n9901 = n3166 ^ n1488 ^ n709 ;
  assign n9902 = ~n8868 & n9901 ;
  assign n9903 = n5123 ^ n1472 ^ n1139 ;
  assign n9904 = ( n4256 & ~n4876 ) | ( n4256 & n9903 ) | ( ~n4876 & n9903 ) ;
  assign n9905 = n9732 | n9904 ;
  assign n9906 = n9905 ^ n7671 ^ 1'b0 ;
  assign n9907 = n983 & ~n1935 ;
  assign n9908 = ~n2445 & n9907 ;
  assign n9909 = ( n1065 & n1659 ) | ( n1065 & ~n6424 ) | ( n1659 & ~n6424 ) ;
  assign n9913 = ~n2823 & n3816 ;
  assign n9914 = n9913 ^ n2204 ^ 1'b0 ;
  assign n9910 = ~n1911 & n3844 ;
  assign n9911 = n9910 ^ n2507 ^ 1'b0 ;
  assign n9912 = ~n9866 & n9911 ;
  assign n9915 = n9914 ^ n9912 ^ 1'b0 ;
  assign n9916 = n8013 & n9915 ;
  assign n9917 = n4332 | n4704 ;
  assign n9918 = n8562 & ~n9917 ;
  assign n9919 = n3543 ^ n209 ^ 1'b0 ;
  assign n9920 = n9919 ^ n5804 ^ n2905 ;
  assign n9921 = n4473 ^ n4458 ^ n1248 ;
  assign n9922 = n9921 ^ n8845 ^ 1'b0 ;
  assign n9923 = n9922 ^ n3045 ^ n1731 ;
  assign n9924 = n8752 & n9923 ;
  assign n9925 = ~n3207 & n9913 ;
  assign n9926 = n9925 ^ n5904 ^ n853 ;
  assign n9927 = n9926 ^ n5754 ^ 1'b0 ;
  assign n9928 = n2064 & n5873 ;
  assign n9929 = n4003 ^ n3347 ^ 1'b0 ;
  assign n9930 = ~n5118 & n9929 ;
  assign n9931 = ( n1094 & ~n9928 ) | ( n1094 & n9930 ) | ( ~n9928 & n9930 ) ;
  assign n9932 = n9931 ^ n9897 ^ 1'b0 ;
  assign n9933 = n4387 & n8853 ;
  assign n9934 = n4178 | n5566 ;
  assign n9935 = n4687 & ~n9934 ;
  assign n9936 = n9935 ^ n7191 ^ n1388 ;
  assign n9937 = n9821 ^ n3975 ^ 1'b0 ;
  assign n9938 = ~n725 & n9937 ;
  assign n9939 = n580 & ~n7482 ;
  assign n9940 = n6567 ^ n5574 ^ n1299 ;
  assign n9941 = ~n1729 & n9940 ;
  assign n9942 = n8335 & ~n9941 ;
  assign n9946 = n155 & ~n2145 ;
  assign n9943 = n1089 & n8226 ;
  assign n9944 = n1272 ^ n820 ^ 1'b0 ;
  assign n9945 = n9943 | n9944 ;
  assign n9947 = n9946 ^ n9945 ^ n614 ;
  assign n9948 = n7425 ^ n4893 ^ 1'b0 ;
  assign n9949 = n7311 & ~n9948 ;
  assign n9950 = n4498 & ~n9090 ;
  assign n9951 = ~n9949 & n9950 ;
  assign n9954 = x54 & n6048 ;
  assign n9955 = n9954 ^ n4610 ^ 1'b0 ;
  assign n9956 = n3791 ^ n2741 ^ 1'b0 ;
  assign n9957 = ~n9955 & n9956 ;
  assign n9958 = n646 & n9957 ;
  assign n9952 = n7685 ^ n7376 ^ x0 ;
  assign n9953 = n5723 & n9952 ;
  assign n9959 = n9958 ^ n9953 ^ 1'b0 ;
  assign n9960 = n9390 ^ n3157 ^ n2487 ;
  assign n9961 = ( ~n1863 & n5051 ) | ( ~n1863 & n9960 ) | ( n5051 & n9960 ) ;
  assign n9962 = n7758 ^ n7718 ^ 1'b0 ;
  assign n9963 = ~n9961 & n9962 ;
  assign n9964 = n9959 & ~n9963 ;
  assign n9965 = n3796 | n6926 ;
  assign n9966 = n3184 & n6498 ;
  assign n9967 = n6425 & n9966 ;
  assign n9968 = ~n380 & n9967 ;
  assign n9969 = n7189 & ~n8257 ;
  assign n9970 = n3416 ^ n2252 ^ 1'b0 ;
  assign n9971 = ( n3838 & n9969 ) | ( n3838 & n9970 ) | ( n9969 & n9970 ) ;
  assign n9972 = n6100 & n7280 ;
  assign n9973 = n1025 & n9972 ;
  assign n9974 = n4465 | n9973 ;
  assign n9975 = n2891 | n9974 ;
  assign n9976 = n5473 ^ n3926 ^ 1'b0 ;
  assign n9977 = n5730 ^ n3876 ^ 1'b0 ;
  assign n9978 = ~n9976 & n9977 ;
  assign n9979 = n2615 & ~n8024 ;
  assign n9980 = ( n5705 & n6560 ) | ( n5705 & n9979 ) | ( n6560 & n9979 ) ;
  assign n9981 = ~n5780 & n8492 ;
  assign n9982 = ~n8027 & n9981 ;
  assign n9983 = n9982 ^ n7340 ^ 1'b0 ;
  assign n9984 = x55 | n9983 ;
  assign n9985 = n9984 ^ n7219 ^ 1'b0 ;
  assign n9986 = n8089 ^ n2467 ^ n773 ;
  assign n9987 = n3237 & n4673 ;
  assign n9988 = n9987 ^ n2668 ^ 1'b0 ;
  assign n9989 = n5443 ^ n199 ^ 1'b0 ;
  assign n9990 = n6003 & n9989 ;
  assign n9991 = ~n1252 & n4413 ;
  assign n9992 = n9991 ^ n820 ^ 1'b0 ;
  assign n9993 = n2243 | n9992 ;
  assign n9994 = ~n7580 & n9993 ;
  assign n9995 = n2228 & n9994 ;
  assign n9996 = n9995 ^ n1247 ^ 1'b0 ;
  assign n9997 = x116 & ~n2117 ;
  assign n9998 = n9997 ^ n2597 ^ 1'b0 ;
  assign n9999 = ~n3108 & n6264 ;
  assign n10000 = n9999 ^ n5139 ^ 1'b0 ;
  assign n10001 = n3171 ^ x13 ^ 1'b0 ;
  assign n10002 = n8522 | n10001 ;
  assign n10003 = n1598 & n5137 ;
  assign n10004 = n5793 ^ n2804 ^ 1'b0 ;
  assign n10005 = ~n4179 & n10004 ;
  assign n10006 = ( n5395 & n10003 ) | ( n5395 & ~n10005 ) | ( n10003 & ~n10005 ) ;
  assign n10007 = n4501 & n10006 ;
  assign n10008 = n9619 & n10007 ;
  assign n10009 = n10008 ^ n313 ^ 1'b0 ;
  assign n10017 = ( ~n1633 & n5225 ) | ( ~n1633 & n6881 ) | ( n5225 & n6881 ) ;
  assign n10011 = n140 & ~n2624 ;
  assign n10012 = n2488 & n2592 ;
  assign n10013 = n10012 ^ n594 ^ 1'b0 ;
  assign n10014 = n10011 & ~n10013 ;
  assign n10015 = n10014 ^ n7377 ^ x116 ;
  assign n10010 = ~n7565 & n7716 ;
  assign n10016 = n10015 ^ n10010 ^ 1'b0 ;
  assign n10018 = n10017 ^ n10016 ^ n5702 ;
  assign n10019 = n5771 ^ n3717 ^ 1'b0 ;
  assign n10020 = ~n4215 & n10019 ;
  assign n10021 = n10020 ^ n7524 ^ n491 ;
  assign n10022 = n7241 ^ n4914 ^ x103 ;
  assign n10023 = n3964 & n4449 ;
  assign n10024 = n4828 & n10023 ;
  assign n10025 = n10024 ^ n5284 ^ 1'b0 ;
  assign n10026 = ~n10022 & n10025 ;
  assign n10027 = n7439 ^ n4754 ^ 1'b0 ;
  assign n10028 = ~n2888 & n10027 ;
  assign n10029 = ~n1113 & n4654 ;
  assign n10030 = n10029 ^ n4507 ^ 1'b0 ;
  assign n10031 = ( n1039 & n5057 ) | ( n1039 & ~n10030 ) | ( n5057 & ~n10030 ) ;
  assign n10032 = n6368 & ~n10031 ;
  assign n10033 = n10032 ^ n5808 ^ n2233 ;
  assign n10038 = n1065 | n9770 ;
  assign n10039 = ( n1456 & n1546 ) | ( n1456 & n10038 ) | ( n1546 & n10038 ) ;
  assign n10035 = n8067 ^ n3539 ^ 1'b0 ;
  assign n10036 = n2221 & ~n10035 ;
  assign n10037 = n3809 & n10036 ;
  assign n10040 = n10039 ^ n10037 ^ 1'b0 ;
  assign n10041 = ~n9801 & n10040 ;
  assign n10042 = n2086 & n10041 ;
  assign n10043 = n4931 ^ n4527 ^ 1'b0 ;
  assign n10044 = n10042 | n10043 ;
  assign n10034 = n6126 & ~n8216 ;
  assign n10045 = n10044 ^ n10034 ^ 1'b0 ;
  assign n10046 = ( ~n990 & n3343 ) | ( ~n990 & n9601 ) | ( n3343 & n9601 ) ;
  assign n10051 = n1796 & n2604 ;
  assign n10052 = n386 & n10051 ;
  assign n10047 = n7844 ^ n816 ^ 1'b0 ;
  assign n10048 = n3329 & ~n10047 ;
  assign n10049 = n10048 ^ n6928 ^ n2532 ;
  assign n10050 = n10049 ^ n9345 ^ n4135 ;
  assign n10053 = n10052 ^ n10050 ^ 1'b0 ;
  assign n10054 = n10053 ^ n4161 ^ 1'b0 ;
  assign n10055 = ~n694 & n933 ;
  assign n10056 = n10055 ^ n7605 ^ 1'b0 ;
  assign n10057 = n7442 & n8230 ;
  assign n10058 = n10057 ^ n8404 ^ 1'b0 ;
  assign n10059 = n2415 & n10058 ;
  assign n10060 = n2308 & n6855 ;
  assign n10061 = n10060 ^ n1469 ^ 1'b0 ;
  assign n10062 = ~n3615 & n10061 ;
  assign n10063 = n10062 ^ n4765 ^ n2167 ;
  assign n10064 = n730 & n2115 ;
  assign n10065 = n10064 ^ x13 ^ 1'b0 ;
  assign n10066 = n129 & n1507 ;
  assign n10067 = ~n1713 & n10066 ;
  assign n10068 = n10067 ^ n4434 ^ 1'b0 ;
  assign n10069 = n9467 ^ n322 ^ 1'b0 ;
  assign n10070 = n4035 & n4369 ;
  assign n10071 = n10070 ^ n7432 ^ 1'b0 ;
  assign n10072 = n3037 & n8217 ;
  assign n10073 = n10071 & ~n10072 ;
  assign n10074 = ( n3908 & n3986 ) | ( n3908 & n8634 ) | ( n3986 & n8634 ) ;
  assign n10075 = n685 | n9619 ;
  assign n10076 = n10075 ^ n6324 ^ 1'b0 ;
  assign n10077 = n4691 & n10061 ;
  assign n10078 = ~n10076 & n10077 ;
  assign n10079 = ( n848 & n2267 ) | ( n848 & n9028 ) | ( n2267 & n9028 ) ;
  assign n10080 = n2557 | n3398 ;
  assign n10081 = n10079 & ~n10080 ;
  assign n10082 = n2124 & ~n8231 ;
  assign n10083 = n10082 ^ n7318 ^ 1'b0 ;
  assign n10084 = n332 & ~n5412 ;
  assign n10085 = n9510 & n10084 ;
  assign n10086 = n5995 ^ n2192 ^ 1'b0 ;
  assign n10087 = ( n634 & n1316 ) | ( n634 & n5784 ) | ( n1316 & n5784 ) ;
  assign n10088 = ( ~n302 & n8655 ) | ( ~n302 & n10087 ) | ( n8655 & n10087 ) ;
  assign n10089 = n7075 ^ n2844 ^ 1'b0 ;
  assign n10090 = x2 & n10089 ;
  assign n10091 = ( n963 & ~n3865 ) | ( n963 & n4102 ) | ( ~n3865 & n4102 ) ;
  assign n10092 = n10091 ^ n8969 ^ 1'b0 ;
  assign n10093 = n6517 & n7121 ;
  assign n10094 = n2105 ^ n1862 ^ 1'b0 ;
  assign n10095 = n2178 & ~n10094 ;
  assign n10096 = n10095 ^ n1240 ^ 1'b0 ;
  assign n10097 = n1146 & ~n10096 ;
  assign n10098 = n790 & ~n9240 ;
  assign n10099 = x61 | n8885 ;
  assign n10100 = n6854 & ~n9327 ;
  assign n10101 = n7514 ^ n4665 ^ n1613 ;
  assign n10102 = n5134 | n10101 ;
  assign n10103 = n6968 ^ n4054 ^ n1116 ;
  assign n10104 = n3307 & n5930 ;
  assign n10105 = n10104 ^ n9343 ^ 1'b0 ;
  assign n10106 = n2791 ^ n473 ^ 1'b0 ;
  assign n10107 = ~n9467 & n10106 ;
  assign n10108 = n6687 & n10107 ;
  assign n10109 = ~n5901 & n10108 ;
  assign n10110 = n887 & n3015 ;
  assign n10111 = n1731 & n10110 ;
  assign n10112 = n4935 & n10111 ;
  assign n10113 = n356 & ~n10112 ;
  assign n10114 = ~n4316 & n10113 ;
  assign n10115 = n10114 ^ n5467 ^ 1'b0 ;
  assign n10119 = n2804 ^ n2260 ^ 1'b0 ;
  assign n10118 = ~n3316 & n3362 ;
  assign n10116 = n1498 & ~n5425 ;
  assign n10117 = n10116 ^ n6567 ^ n1476 ;
  assign n10120 = n10119 ^ n10118 ^ n10117 ;
  assign n10121 = n1983 ^ n1745 ^ n193 ;
  assign n10122 = n10121 ^ n6349 ^ n2445 ;
  assign n10123 = n9332 ^ n9068 ^ n3258 ;
  assign n10124 = n10123 ^ n3114 ^ 1'b0 ;
  assign n10125 = n1894 & n10124 ;
  assign n10126 = n8196 ^ n514 ^ 1'b0 ;
  assign n10127 = n10125 & ~n10126 ;
  assign n10128 = n7989 & ~n8960 ;
  assign n10133 = n4491 ^ n3751 ^ n2120 ;
  assign n10131 = n5784 ^ n1653 ^ x50 ;
  assign n10132 = n4461 | n10131 ;
  assign n10134 = n10133 ^ n10132 ^ 1'b0 ;
  assign n10135 = n10134 ^ n6190 ^ 1'b0 ;
  assign n10136 = ~n9841 & n10135 ;
  assign n10129 = n5372 | n6632 ;
  assign n10130 = ~n6480 & n10129 ;
  assign n10137 = n10136 ^ n10130 ^ 1'b0 ;
  assign n10138 = n2151 & ~n2520 ;
  assign n10139 = ~x95 & n10138 ;
  assign n10140 = n5654 & ~n10139 ;
  assign n10141 = n7060 & ~n7234 ;
  assign n10142 = n10141 ^ n4273 ^ 1'b0 ;
  assign n10143 = n10142 ^ n1203 ^ n823 ;
  assign n10146 = ~n2801 & n3926 ;
  assign n10144 = n1438 & n4216 ;
  assign n10145 = n2687 & n10144 ;
  assign n10147 = n10146 ^ n10145 ^ n8441 ;
  assign n10148 = n1699 | n7868 ;
  assign n10149 = n10148 ^ n5822 ^ n4326 ;
  assign n10150 = n240 | n2969 ;
  assign n10151 = n308 & ~n10150 ;
  assign n10152 = n10151 ^ n9911 ^ n6112 ;
  assign n10153 = n10152 ^ n4085 ^ 1'b0 ;
  assign n10154 = n1910 ^ n1308 ^ n668 ;
  assign n10155 = ~n4057 & n10154 ;
  assign n10156 = n2816 & n10155 ;
  assign n10157 = n4713 & n10156 ;
  assign n10158 = ( ~n3660 & n4523 ) | ( ~n3660 & n5099 ) | ( n4523 & n5099 ) ;
  assign n10159 = n3482 & n10158 ;
  assign n10160 = n10159 ^ n4916 ^ 1'b0 ;
  assign n10161 = ( n4761 & n10157 ) | ( n4761 & n10160 ) | ( n10157 & n10160 ) ;
  assign n10162 = n6269 ^ n673 ^ 1'b0 ;
  assign n10163 = n5213 & ~n10162 ;
  assign n10164 = n8334 & ~n10163 ;
  assign n10166 = n1312 ^ n350 ^ 1'b0 ;
  assign n10165 = n1573 & n4172 ;
  assign n10167 = n10166 ^ n10165 ^ n5829 ;
  assign n10173 = ( ~n2753 & n8529 ) | ( ~n2753 & n9532 ) | ( n8529 & n9532 ) ;
  assign n10168 = n2986 | n3423 ;
  assign n10169 = n10168 ^ n7618 ^ 1'b0 ;
  assign n10170 = n210 | n1125 ;
  assign n10171 = ( n2761 & ~n10169 ) | ( n2761 & n10170 ) | ( ~n10169 & n10170 ) ;
  assign n10172 = ( ~n3315 & n8181 ) | ( ~n3315 & n10171 ) | ( n8181 & n10171 ) ;
  assign n10174 = n10173 ^ n10172 ^ 1'b0 ;
  assign n10175 = n9762 ^ n8500 ^ 1'b0 ;
  assign n10176 = n2335 | n10175 ;
  assign n10177 = n7406 ^ n7040 ^ 1'b0 ;
  assign n10178 = n5731 & ~n10177 ;
  assign n10179 = ~n3128 & n10178 ;
  assign n10180 = n2560 ^ n2515 ^ 1'b0 ;
  assign n10181 = n6491 & ~n10180 ;
  assign n10182 = n508 | n1918 ;
  assign n10183 = n10182 ^ n1819 ^ 1'b0 ;
  assign n10184 = n2590 | n10053 ;
  assign n10185 = n8350 | n10184 ;
  assign n10186 = n5994 | n10185 ;
  assign n10187 = n6491 ^ x96 ^ 1'b0 ;
  assign n10188 = n1493 & n10187 ;
  assign n10189 = n1425 & ~n4878 ;
  assign n10190 = n6243 & ~n6573 ;
  assign n10191 = ~n10189 & n10190 ;
  assign n10192 = n3111 & n4816 ;
  assign n10193 = ~n8539 & n10192 ;
  assign n10194 = n3090 ^ n2177 ^ 1'b0 ;
  assign n10195 = x51 & ~n10194 ;
  assign n10196 = n1162 | n1459 ;
  assign n10197 = n1162 & ~n10196 ;
  assign n10198 = n10197 ^ n3299 ^ 1'b0 ;
  assign n10199 = n5032 & ~n5073 ;
  assign n10200 = n2625 & ~n10199 ;
  assign n10201 = ~n10198 & n10200 ;
  assign n10202 = ( ~n233 & n1331 ) | ( ~n233 & n5374 ) | ( n1331 & n5374 ) ;
  assign n10203 = n10202 ^ n10072 ^ 1'b0 ;
  assign n10204 = n4487 & n10203 ;
  assign n10205 = ( n4548 & ~n4962 ) | ( n4548 & n7823 ) | ( ~n4962 & n7823 ) ;
  assign n10206 = n10173 ^ n6070 ^ 1'b0 ;
  assign n10207 = n10205 & n10206 ;
  assign n10208 = n2040 ^ n613 ^ 1'b0 ;
  assign n10209 = n3402 | n10208 ;
  assign n10211 = n3999 ^ n1163 ^ x118 ;
  assign n10212 = ( x56 & n1143 ) | ( x56 & n1829 ) | ( n1143 & n1829 ) ;
  assign n10213 = ( n935 & n10211 ) | ( n935 & ~n10212 ) | ( n10211 & ~n10212 ) ;
  assign n10210 = n1659 | n2500 ;
  assign n10214 = n10213 ^ n10210 ^ n431 ;
  assign n10215 = ~n10209 & n10214 ;
  assign n10216 = n1354 & n10215 ;
  assign n10217 = n9775 ^ n3763 ^ n3699 ;
  assign n10218 = n1527 | n2381 ;
  assign n10219 = ~n618 & n6388 ;
  assign n10220 = n10218 & n10219 ;
  assign n10221 = n1368 | n10220 ;
  assign n10222 = n4214 | n10221 ;
  assign n10223 = n1150 & n1642 ;
  assign n10224 = n10223 ^ n5032 ^ 1'b0 ;
  assign n10225 = n10222 & n10224 ;
  assign n10226 = n8941 ^ x107 ^ 1'b0 ;
  assign n10227 = n10225 | n10226 ;
  assign n10228 = n225 | n600 ;
  assign n10229 = n10228 ^ n1084 ^ 1'b0 ;
  assign n10230 = ( ~n6047 & n9306 ) | ( ~n6047 & n9630 ) | ( n9306 & n9630 ) ;
  assign n10231 = n6605 ^ n2597 ^ 1'b0 ;
  assign n10232 = n4352 & n10231 ;
  assign n10233 = n10232 ^ n5703 ^ n3104 ;
  assign n10234 = ~n5593 & n10233 ;
  assign n10235 = n6749 & n8731 ;
  assign n10240 = n825 & ~n3821 ;
  assign n10241 = ( n3953 & n8466 ) | ( n3953 & n10240 ) | ( n8466 & n10240 ) ;
  assign n10236 = ~n693 & n9840 ;
  assign n10237 = n693 & n10236 ;
  assign n10238 = n2107 | n10237 ;
  assign n10239 = n10237 & ~n10238 ;
  assign n10242 = n10241 ^ n10239 ^ 1'b0 ;
  assign n10243 = n1017 & ~n4458 ;
  assign n10244 = ( n8780 & n8798 ) | ( n8780 & ~n10243 ) | ( n8798 & ~n10243 ) ;
  assign n10245 = n2188 | n2968 ;
  assign n10246 = n2188 & ~n10245 ;
  assign n10247 = n10246 ^ n2931 ^ 1'b0 ;
  assign n10248 = n9792 | n10247 ;
  assign n10251 = n714 & ~n8491 ;
  assign n10252 = n8491 & n10251 ;
  assign n10253 = n1913 & n10252 ;
  assign n10249 = n4492 ^ n4418 ^ 1'b0 ;
  assign n10250 = n1760 | n10249 ;
  assign n10254 = n10253 ^ n10250 ^ 1'b0 ;
  assign n10256 = n1960 ^ n618 ^ 1'b0 ;
  assign n10257 = n4169 & n10256 ;
  assign n10258 = n3033 ^ n701 ^ 1'b0 ;
  assign n10259 = n10257 & n10258 ;
  assign n10260 = ( n146 & n5168 ) | ( n146 & n9308 ) | ( n5168 & n9308 ) ;
  assign n10261 = n6452 & ~n10260 ;
  assign n10262 = ~n10259 & n10261 ;
  assign n10255 = n4306 | n7333 ;
  assign n10263 = n10262 ^ n10255 ^ 1'b0 ;
  assign n10264 = n3043 ^ n340 ^ 1'b0 ;
  assign n10265 = n10264 ^ n951 ^ 1'b0 ;
  assign n10267 = n2776 ^ n2554 ^ 1'b0 ;
  assign n10268 = ~n4265 & n10267 ;
  assign n10266 = n7877 ^ n627 ^ 1'b0 ;
  assign n10269 = n10268 ^ n10266 ^ x121 ;
  assign n10270 = n209 | n2211 ;
  assign n10271 = n4955 ^ n1628 ^ n219 ;
  assign n10272 = ~n3317 & n10271 ;
  assign n10273 = n4207 & ~n10272 ;
  assign n10274 = ~n10270 & n10273 ;
  assign n10275 = n10274 ^ n4275 ^ n3363 ;
  assign n10276 = n10275 ^ n8310 ^ 1'b0 ;
  assign n10279 = n3444 ^ n2515 ^ 1'b0 ;
  assign n10280 = n2510 & ~n10279 ;
  assign n10277 = n1748 ^ n1406 ^ 1'b0 ;
  assign n10278 = n3279 & ~n10277 ;
  assign n10281 = n10280 ^ n10278 ^ 1'b0 ;
  assign n10282 = n3357 ^ n855 ^ n657 ;
  assign n10283 = n7363 ^ n5312 ^ 1'b0 ;
  assign n10284 = n1784 & n10283 ;
  assign n10285 = n10284 ^ n3783 ^ 1'b0 ;
  assign n10286 = ~n1034 & n10285 ;
  assign n10287 = ( n8564 & n10282 ) | ( n8564 & n10286 ) | ( n10282 & n10286 ) ;
  assign n10288 = n6034 | n6744 ;
  assign n10289 = n5648 | n6427 ;
  assign n10290 = ( n1029 & n1863 ) | ( n1029 & n5301 ) | ( n1863 & n5301 ) ;
  assign n10291 = n10290 ^ n4835 ^ 1'b0 ;
  assign n10292 = ~n3498 & n10291 ;
  assign n10293 = n10292 ^ n9637 ^ 1'b0 ;
  assign n10294 = ~x64 & n8223 ;
  assign n10295 = ( n432 & n1680 ) | ( n432 & ~n9218 ) | ( n1680 & ~n9218 ) ;
  assign n10296 = n5517 ^ n4397 ^ n533 ;
  assign n10297 = n8106 | n10296 ;
  assign n10298 = n7226 ^ n3345 ^ n1046 ;
  assign n10299 = ~n3719 & n10154 ;
  assign n10300 = n438 & n10299 ;
  assign n10301 = ~n4133 & n6312 ;
  assign n10302 = n10300 & n10301 ;
  assign n10303 = n5703 ^ n4772 ^ n356 ;
  assign n10304 = n1108 ^ n131 ^ 1'b0 ;
  assign n10305 = n10304 ^ n6635 ^ x98 ;
  assign n10306 = n3416 | n10305 ;
  assign n10307 = n10303 & ~n10306 ;
  assign n10309 = n245 ^ x107 ^ 1'b0 ;
  assign n10308 = n1466 ^ x12 ^ 1'b0 ;
  assign n10310 = n10309 ^ n10308 ^ x62 ;
  assign n10311 = ~n2081 & n6226 ;
  assign n10312 = n10311 ^ n4119 ^ 1'b0 ;
  assign n10313 = ( n5665 & ~n8840 ) | ( n5665 & n10312 ) | ( ~n8840 & n10312 ) ;
  assign n10314 = n841 & n5934 ;
  assign n10315 = ~n3819 & n10314 ;
  assign n10316 = n485 & n2743 ;
  assign n10317 = n4593 & n10316 ;
  assign n10318 = n10317 ^ n8848 ^ n2843 ;
  assign n10319 = n1473 & ~n1867 ;
  assign n10320 = n3719 & n10319 ;
  assign n10321 = n5351 ^ n4135 ^ 1'b0 ;
  assign n10322 = ~n10320 & n10321 ;
  assign n10323 = ( ~n8532 & n8776 ) | ( ~n8532 & n10322 ) | ( n8776 & n10322 ) ;
  assign n10324 = n6106 ^ n3778 ^ 1'b0 ;
  assign n10325 = n9025 & ~n10324 ;
  assign n10326 = ~n6781 & n10325 ;
  assign n10327 = n7860 & ~n10326 ;
  assign n10328 = n10323 & n10327 ;
  assign n10329 = n187 & n6585 ;
  assign n10330 = ~n5469 & n10329 ;
  assign n10331 = ( n3771 & ~n10328 ) | ( n3771 & n10330 ) | ( ~n10328 & n10330 ) ;
  assign n10332 = n4942 & n5054 ;
  assign n10333 = n10332 ^ n4716 ^ 1'b0 ;
  assign n10335 = ( n2647 & ~n3232 ) | ( n2647 & n5780 ) | ( ~n3232 & n5780 ) ;
  assign n10334 = n3981 & ~n5400 ;
  assign n10336 = n10335 ^ n10334 ^ 1'b0 ;
  assign n10337 = n10333 & n10336 ;
  assign n10338 = n7130 ^ n4295 ^ 1'b0 ;
  assign n10339 = n8823 ^ n4566 ^ 1'b0 ;
  assign n10341 = n5806 ^ n3921 ^ 1'b0 ;
  assign n10340 = n5689 ^ n2686 ^ n438 ;
  assign n10342 = n10341 ^ n10340 ^ n1756 ;
  assign n10343 = n7725 ^ n2269 ^ n1515 ;
  assign n10344 = n10343 ^ n6552 ^ 1'b0 ;
  assign n10345 = n3863 & n4018 ;
  assign n10346 = n9105 ^ n8078 ^ n4052 ;
  assign n10347 = n8491 ^ n3548 ^ 1'b0 ;
  assign n10348 = n8900 ^ x74 ^ 1'b0 ;
  assign n10349 = n938 & ~n7233 ;
  assign n10350 = n6609 ^ n3355 ^ 1'b0 ;
  assign n10351 = x2 & n10350 ;
  assign n10352 = ( n509 & n5135 ) | ( n509 & ~n5377 ) | ( n5135 & ~n5377 ) ;
  assign n10353 = n10148 & n10352 ;
  assign n10354 = n10353 ^ n4099 ^ 1'b0 ;
  assign n10355 = ~n6401 & n6521 ;
  assign n10356 = n10355 ^ n5973 ^ 1'b0 ;
  assign n10357 = n3088 & n5241 ;
  assign n10358 = n8521 ^ n4921 ^ 1'b0 ;
  assign n10361 = n9042 ^ n6064 ^ 1'b0 ;
  assign n10362 = n7403 & n10361 ;
  assign n10359 = n358 | n4638 ;
  assign n10360 = n10359 ^ n9892 ^ 1'b0 ;
  assign n10363 = n10362 ^ n10360 ^ 1'b0 ;
  assign n10364 = ~n10358 & n10363 ;
  assign n10365 = n1863 & ~n5152 ;
  assign n10366 = n10365 ^ n1725 ^ 1'b0 ;
  assign n10370 = n2597 ^ x36 ^ 1'b0 ;
  assign n10371 = ~n1354 & n1720 ;
  assign n10372 = n10371 ^ n3910 ^ 1'b0 ;
  assign n10373 = n10370 | n10372 ;
  assign n10367 = n4856 & n7140 ;
  assign n10368 = n7363 | n9679 ;
  assign n10369 = n10367 | n10368 ;
  assign n10374 = n10373 ^ n10369 ^ n5555 ;
  assign n10375 = n3002 | n4524 ;
  assign n10376 = ( x116 & n773 ) | ( x116 & n2099 ) | ( n773 & n2099 ) ;
  assign n10377 = n798 & n10376 ;
  assign n10378 = n1093 & n10377 ;
  assign n10379 = n7917 & ~n10378 ;
  assign n10380 = n8445 & n10379 ;
  assign n10381 = x83 & ~n6609 ;
  assign n10382 = ( n5127 & n7011 ) | ( n5127 & n10381 ) | ( n7011 & n10381 ) ;
  assign n10383 = n4275 ^ n1542 ^ 1'b0 ;
  assign n10384 = n10383 ^ n960 ^ 1'b0 ;
  assign n10385 = n6864 ^ n614 ^ 1'b0 ;
  assign n10386 = n6034 | n10385 ;
  assign n10390 = n3127 ^ n298 ^ 1'b0 ;
  assign n10387 = ~n490 & n1783 ;
  assign n10388 = n10387 ^ n6205 ^ n1422 ;
  assign n10389 = n9988 & n10388 ;
  assign n10391 = n10390 ^ n10389 ^ 1'b0 ;
  assign n10393 = n4553 | n7934 ;
  assign n10392 = n5502 & ~n7400 ;
  assign n10394 = n10393 ^ n10392 ^ 1'b0 ;
  assign n10395 = n7311 ^ n6230 ^ 1'b0 ;
  assign n10396 = n497 | n10395 ;
  assign n10397 = n684 & n1631 ;
  assign n10398 = n1611 & n10397 ;
  assign n10399 = n10398 ^ n5341 ^ 1'b0 ;
  assign n10400 = ( n2708 & ~n4837 ) | ( n2708 & n7245 ) | ( ~n4837 & n7245 ) ;
  assign n10401 = n10400 ^ n5658 ^ n572 ;
  assign n10402 = n1979 ^ n1516 ^ 1'b0 ;
  assign n10403 = n1312 | n10402 ;
  assign n10404 = n4862 ^ n920 ^ 1'b0 ;
  assign n10405 = n3121 & n5980 ;
  assign n10406 = ~n1470 & n10405 ;
  assign n10407 = n10406 ^ n6260 ^ 1'b0 ;
  assign n10408 = n7341 & n10407 ;
  assign n10409 = ~n10404 & n10408 ;
  assign n10410 = ( n3950 & n5435 ) | ( n3950 & ~n9914 ) | ( n5435 & ~n9914 ) ;
  assign n10411 = ( n2502 & n5458 ) | ( n2502 & ~n10410 ) | ( n5458 & ~n10410 ) ;
  assign n10412 = ( n6112 & n8535 ) | ( n6112 & ~n10411 ) | ( n8535 & ~n10411 ) ;
  assign n10413 = n6110 ^ n685 ^ 1'b0 ;
  assign n10414 = n6810 & n10413 ;
  assign n10415 = n2029 & n10414 ;
  assign n10416 = ( n4452 & ~n9784 ) | ( n4452 & n10415 ) | ( ~n9784 & n10415 ) ;
  assign n10417 = n5499 & ~n6764 ;
  assign n10418 = n6934 & n10417 ;
  assign n10419 = n10418 ^ n173 ^ 1'b0 ;
  assign n10420 = n2213 & n10419 ;
  assign n10421 = ( n4414 & n5322 ) | ( n4414 & ~n9846 ) | ( n5322 & ~n9846 ) ;
  assign n10422 = n4492 ^ n4261 ^ 1'b0 ;
  assign n10423 = n4193 | n10422 ;
  assign n10424 = n494 & ~n10423 ;
  assign n10425 = n7801 | n10424 ;
  assign n10426 = x14 & ~n1370 ;
  assign n10427 = n10426 ^ n4571 ^ 1'b0 ;
  assign n10428 = ( n3244 & n4159 ) | ( n3244 & ~n10427 ) | ( n4159 & ~n10427 ) ;
  assign n10429 = ( x10 & n4286 ) | ( x10 & ~n4328 ) | ( n4286 & ~n4328 ) ;
  assign n10430 = n1023 | n10429 ;
  assign n10431 = ( n1323 & n6393 ) | ( n1323 & ~n8522 ) | ( n6393 & ~n8522 ) ;
  assign n10432 = ~n3002 & n10431 ;
  assign n10433 = ( n8669 & n10430 ) | ( n8669 & ~n10432 ) | ( n10430 & ~n10432 ) ;
  assign n10434 = n1575 ^ n1521 ^ 1'b0 ;
  assign n10435 = n2363 ^ x86 ^ 1'b0 ;
  assign n10436 = n822 & ~n6772 ;
  assign n10437 = n6412 & n10436 ;
  assign n10438 = ~n10435 & n10437 ;
  assign n10439 = n4216 ^ n4077 ^ 1'b0 ;
  assign n10440 = n10439 ^ n8243 ^ n325 ;
  assign n10441 = ( n932 & n7045 ) | ( n932 & n10440 ) | ( n7045 & n10440 ) ;
  assign n10442 = n2352 | n9503 ;
  assign n10443 = n10142 | n10442 ;
  assign n10444 = n5958 ^ n5768 ^ 1'b0 ;
  assign n10445 = n2102 & ~n2431 ;
  assign n10446 = n822 & n10445 ;
  assign n10447 = n10446 ^ n4358 ^ 1'b0 ;
  assign n10448 = n10444 & ~n10447 ;
  assign n10449 = n3821 & ~n7302 ;
  assign n10450 = n7769 & n10449 ;
  assign n10451 = n10450 ^ n7789 ^ 1'b0 ;
  assign n10454 = ~n3375 & n4440 ;
  assign n10453 = n8033 & ~n8194 ;
  assign n10452 = n2703 & n8799 ;
  assign n10455 = n10454 ^ n10453 ^ n10452 ;
  assign n10456 = n4221 & n9527 ;
  assign n10457 = n9002 ^ n5145 ^ 1'b0 ;
  assign n10458 = n9153 ^ n5011 ^ n2432 ;
  assign n10459 = n7156 ^ n1964 ^ 1'b0 ;
  assign n10460 = n6617 ^ n3701 ^ n2580 ;
  assign n10461 = ~n1252 & n10460 ;
  assign n10462 = n1653 ^ n138 ^ x17 ;
  assign n10463 = n10462 ^ n448 ^ 1'b0 ;
  assign n10464 = n2855 & ~n10463 ;
  assign n10465 = n10398 | n10464 ;
  assign n10466 = n327 & ~n6195 ;
  assign n10467 = n10466 ^ n6724 ^ n3274 ;
  assign n10468 = n3608 & ~n10467 ;
  assign n10469 = n154 | n5011 ;
  assign n10470 = ~n7984 & n10446 ;
  assign n10471 = n7099 ^ n5527 ^ 1'b0 ;
  assign n10472 = n6705 | n10471 ;
  assign n10473 = n8122 | n8413 ;
  assign n10474 = n10473 ^ n5661 ^ 1'b0 ;
  assign n10475 = ~n7526 & n10474 ;
  assign n10476 = n3056 ^ n3030 ^ 1'b0 ;
  assign n10477 = ~n540 & n3813 ;
  assign n10478 = ~n2012 & n10477 ;
  assign n10479 = n10478 ^ n3349 ^ 1'b0 ;
  assign n10480 = n10476 | n10479 ;
  assign n10481 = n9097 ^ n8157 ^ n6609 ;
  assign n10482 = n9099 ^ n3222 ^ n2077 ;
  assign n10483 = n5740 ^ n1227 ^ 1'b0 ;
  assign n10484 = n10483 ^ n6885 ^ n1958 ;
  assign n10485 = ( n4682 & n6853 ) | ( n4682 & n10484 ) | ( n6853 & n10484 ) ;
  assign n10486 = n3953 ^ n1811 ^ 1'b0 ;
  assign n10487 = n10486 ^ n3681 ^ n2491 ;
  assign n10488 = ( x20 & n267 ) | ( x20 & ~n543 ) | ( n267 & ~n543 ) ;
  assign n10489 = ( n4141 & n9409 ) | ( n4141 & ~n10488 ) | ( n9409 & ~n10488 ) ;
  assign n10490 = ~n1809 & n10489 ;
  assign n10491 = n10490 ^ n2581 ^ 1'b0 ;
  assign n10493 = ( n606 & n3260 ) | ( n606 & n4583 ) | ( n3260 & n4583 ) ;
  assign n10494 = n10493 ^ n9495 ^ n1445 ;
  assign n10492 = ( n1622 & ~n3319 ) | ( n1622 & n8694 ) | ( ~n3319 & n8694 ) ;
  assign n10495 = n10494 ^ n10492 ^ n9802 ;
  assign n10496 = n7771 ^ n3390 ^ 1'b0 ;
  assign n10497 = n1167 & ~n2406 ;
  assign n10498 = n6223 ^ n5258 ^ 1'b0 ;
  assign n10503 = n2956 ^ n2549 ^ 1'b0 ;
  assign n10500 = n3868 ^ n3307 ^ n2554 ;
  assign n10501 = n4286 | n10500 ;
  assign n10499 = ( n1588 & n2358 ) | ( n1588 & ~n3341 ) | ( n2358 & ~n3341 ) ;
  assign n10502 = n10501 ^ n10499 ^ 1'b0 ;
  assign n10504 = n10503 ^ n10502 ^ 1'b0 ;
  assign n10505 = ~n6336 & n10504 ;
  assign n10506 = ~n10498 & n10505 ;
  assign n10507 = ( n6225 & ~n10497 ) | ( n6225 & n10506 ) | ( ~n10497 & n10506 ) ;
  assign n10508 = n10507 ^ n1014 ^ 1'b0 ;
  assign n10509 = n7952 & ~n10508 ;
  assign n10510 = n4554 ^ n595 ^ 1'b0 ;
  assign n10511 = n3391 | n10510 ;
  assign n10512 = n1384 & n4458 ;
  assign n10513 = ( n3330 & n8522 ) | ( n3330 & ~n9709 ) | ( n8522 & ~n9709 ) ;
  assign n10514 = n1260 | n3467 ;
  assign n10515 = n10514 ^ n4554 ^ 1'b0 ;
  assign n10516 = n1084 & n8059 ;
  assign n10517 = n10516 ^ n2051 ^ 1'b0 ;
  assign n10518 = n8493 ^ n4051 ^ 1'b0 ;
  assign n10519 = ~n2660 & n9151 ;
  assign n10520 = ( ~n3770 & n6859 ) | ( ~n3770 & n10519 ) | ( n6859 & n10519 ) ;
  assign n10521 = n3337 | n10520 ;
  assign n10522 = ~n841 & n6586 ;
  assign n10523 = n10522 ^ n2693 ^ 1'b0 ;
  assign n10524 = n3699 | n8231 ;
  assign n10525 = n10523 | n10524 ;
  assign n10526 = ( x113 & n177 ) | ( x113 & ~n5096 ) | ( n177 & ~n5096 ) ;
  assign n10527 = n8801 & ~n10526 ;
  assign n10528 = n10525 & ~n10527 ;
  assign n10529 = n1862 & n2323 ;
  assign n10530 = ~n10528 & n10529 ;
  assign n10531 = n9501 ^ n4369 ^ 1'b0 ;
  assign n10541 = n5461 ^ n822 ^ 1'b0 ;
  assign n10542 = n7721 & ~n10541 ;
  assign n10543 = n4670 & n10542 ;
  assign n10540 = n4609 ^ n3491 ^ n3066 ;
  assign n10532 = n1071 | n2324 ;
  assign n10533 = n2931 ^ n665 ^ 1'b0 ;
  assign n10534 = n5058 & ~n10533 ;
  assign n10535 = ~n182 & n10534 ;
  assign n10536 = ~n10532 & n10535 ;
  assign n10537 = ( n2745 & n3127 ) | ( n2745 & ~n8301 ) | ( n3127 & ~n8301 ) ;
  assign n10538 = ~n1430 & n10537 ;
  assign n10539 = n10536 & n10538 ;
  assign n10544 = n10543 ^ n10540 ^ n10539 ;
  assign n10545 = ( n3323 & ~n10531 ) | ( n3323 & n10544 ) | ( ~n10531 & n10544 ) ;
  assign n10546 = n10545 ^ n383 ^ 1'b0 ;
  assign n10549 = n1470 & ~n5369 ;
  assign n10547 = ~n2929 & n9875 ;
  assign n10548 = n10547 ^ n8411 ^ 1'b0 ;
  assign n10550 = n10549 ^ n10548 ^ n368 ;
  assign n10551 = n4525 & ~n6447 ;
  assign n10552 = n10551 ^ n1231 ^ 1'b0 ;
  assign n10557 = n692 | n5510 ;
  assign n10558 = n2081 & ~n10557 ;
  assign n10559 = n10558 ^ n10322 ^ n2662 ;
  assign n10553 = n1294 & n4356 ;
  assign n10554 = n9504 ^ n285 ^ 1'b0 ;
  assign n10555 = n10554 ^ n1649 ^ 1'b0 ;
  assign n10556 = n10553 & n10555 ;
  assign n10560 = n10559 ^ n10556 ^ 1'b0 ;
  assign n10561 = n9845 & n10560 ;
  assign n10562 = ~n3628 & n8830 ;
  assign n10563 = n10562 ^ n6568 ^ 1'b0 ;
  assign n10564 = ~n1307 & n10563 ;
  assign n10565 = n3262 | n6880 ;
  assign n10566 = n10565 ^ n3874 ^ 1'b0 ;
  assign n10567 = n6523 ^ n1744 ^ 1'b0 ;
  assign n10568 = ~n3373 & n3961 ;
  assign n10569 = n10567 & n10568 ;
  assign n10570 = n2932 | n10569 ;
  assign n10571 = n3610 | n10570 ;
  assign n10572 = ( n2231 & n6196 ) | ( n2231 & n7510 ) | ( n6196 & n7510 ) ;
  assign n10573 = n1252 | n6101 ;
  assign n10574 = x113 & ~n4737 ;
  assign n10575 = n10573 & n10574 ;
  assign n10576 = ( n1858 & ~n5138 ) | ( n1858 & n10575 ) | ( ~n5138 & n10575 ) ;
  assign n10577 = n10576 ^ n4193 ^ 1'b0 ;
  assign n10578 = n5515 & ~n10577 ;
  assign n10581 = n6273 ^ n882 ^ 1'b0 ;
  assign n10582 = ~n3467 & n10581 ;
  assign n10583 = ~n5428 & n10582 ;
  assign n10579 = ( n1512 & ~n3704 ) | ( n1512 & n6986 ) | ( ~n3704 & n6986 ) ;
  assign n10580 = ~n4876 & n10579 ;
  assign n10584 = n10583 ^ n10580 ^ 1'b0 ;
  assign n10585 = n8286 ^ n4555 ^ 1'b0 ;
  assign n10586 = n723 & ~n10585 ;
  assign n10587 = n7681 ^ n4229 ^ n1338 ;
  assign n10592 = n2723 | n2818 ;
  assign n10590 = n8458 ^ n2320 ^ 1'b0 ;
  assign n10591 = ~n693 & n10590 ;
  assign n10593 = n10592 ^ n10591 ^ n9736 ;
  assign n10588 = n563 & ~n6114 ;
  assign n10589 = n7935 | n10588 ;
  assign n10594 = n10593 ^ n10589 ^ 1'b0 ;
  assign n10595 = n3009 & n10142 ;
  assign n10596 = ~n7828 & n10595 ;
  assign n10597 = ( n1511 & n3958 ) | ( n1511 & ~n7355 ) | ( n3958 & ~n7355 ) ;
  assign n10598 = n9533 ^ n3218 ^ 1'b0 ;
  assign n10599 = n2962 | n9561 ;
  assign n10600 = n7747 ^ n6722 ^ 1'b0 ;
  assign n10601 = n10599 | n10600 ;
  assign n10602 = n3854 | n3967 ;
  assign n10603 = ( n4490 & ~n5016 ) | ( n4490 & n10602 ) | ( ~n5016 & n10602 ) ;
  assign n10604 = n9580 | n10603 ;
  assign n10605 = n1700 ^ n443 ^ 1'b0 ;
  assign n10606 = n3147 & n10605 ;
  assign n10607 = n10606 ^ n2445 ^ 1'b0 ;
  assign n10608 = ( n972 & n1141 ) | ( n972 & n1960 ) | ( n1141 & n1960 ) ;
  assign n10610 = n2457 ^ n650 ^ 1'b0 ;
  assign n10609 = n4261 ^ n4211 ^ n1628 ;
  assign n10611 = n10610 ^ n10609 ^ n650 ;
  assign n10612 = ( n4217 & n10608 ) | ( n4217 & ~n10611 ) | ( n10608 & ~n10611 ) ;
  assign n10613 = n6560 ^ n5155 ^ 1'b0 ;
  assign n10614 = n10613 ^ n10080 ^ 1'b0 ;
  assign n10615 = ~n3048 & n10614 ;
  assign n10616 = n1316 | n7307 ;
  assign n10617 = n10616 ^ n416 ^ 1'b0 ;
  assign n10622 = n1814 | n9609 ;
  assign n10623 = n10622 ^ n3144 ^ 1'b0 ;
  assign n10618 = ~n210 & n445 ;
  assign n10619 = n7852 ^ n653 ^ 1'b0 ;
  assign n10620 = n10618 | n10619 ;
  assign n10621 = n10620 ^ n4397 ^ n3248 ;
  assign n10624 = n10623 ^ n10621 ^ n9469 ;
  assign n10625 = n4743 ^ n958 ^ 1'b0 ;
  assign n10627 = ~n201 & n1795 ;
  assign n10628 = n10627 ^ n993 ^ 1'b0 ;
  assign n10629 = n3312 & ~n10628 ;
  assign n10626 = ~n2084 & n2643 ;
  assign n10630 = n10629 ^ n10626 ^ n10151 ;
  assign n10631 = ~n10625 & n10630 ;
  assign n10632 = n10380 & n10631 ;
  assign n10633 = ( n692 & ~n3946 ) | ( n692 & n4248 ) | ( ~n3946 & n4248 ) ;
  assign n10634 = n10633 ^ n3599 ^ n1104 ;
  assign n10635 = n5958 ^ n5132 ^ n3202 ;
  assign n10636 = n3522 | n6303 ;
  assign n10637 = ( ~n984 & n4511 ) | ( ~n984 & n10636 ) | ( n4511 & n10636 ) ;
  assign n10638 = n2187 & n3017 ;
  assign n10639 = n10638 ^ n438 ^ 1'b0 ;
  assign n10640 = n10639 ^ n7370 ^ n2320 ;
  assign n10641 = n10640 ^ n5409 ^ n566 ;
  assign n10643 = n528 | n1810 ;
  assign n10642 = ~n210 & n5070 ;
  assign n10644 = n10643 ^ n10642 ^ 1'b0 ;
  assign n10645 = ( n4647 & ~n5113 ) | ( n4647 & n7739 ) | ( ~n5113 & n7739 ) ;
  assign n10646 = n10645 ^ n1207 ^ 1'b0 ;
  assign n10647 = ~n8386 & n10646 ;
  assign n10648 = ( n1436 & n3284 ) | ( n1436 & ~n10647 ) | ( n3284 & ~n10647 ) ;
  assign n10649 = ~n1006 & n3873 ;
  assign n10650 = n4916 | n5049 ;
  assign n10651 = n10649 & ~n10650 ;
  assign n10652 = n1425 & ~n5904 ;
  assign n10653 = ~n4135 & n10652 ;
  assign n10654 = n10611 ^ n4210 ^ 1'b0 ;
  assign n10655 = n5266 | n10654 ;
  assign n10660 = n6237 ^ n3734 ^ n3611 ;
  assign n10656 = n525 & n2897 ;
  assign n10657 = ( n1228 & n1725 ) | ( n1228 & ~n10656 ) | ( n1725 & ~n10656 ) ;
  assign n10658 = n3933 ^ n3587 ^ n3287 ;
  assign n10659 = n10657 & ~n10658 ;
  assign n10661 = n10660 ^ n10659 ^ n2195 ;
  assign n10663 = n8592 ^ n1283 ^ 1'b0 ;
  assign n10662 = n4734 | n10260 ;
  assign n10664 = n10663 ^ n10662 ^ 1'b0 ;
  assign n10665 = n5860 ^ n949 ^ 1'b0 ;
  assign n10666 = n10665 ^ n5012 ^ n729 ;
  assign n10667 = n1477 ^ n1378 ^ n1175 ;
  assign n10668 = ( n7350 & n7822 ) | ( n7350 & ~n10667 ) | ( n7822 & ~n10667 ) ;
  assign n10669 = n10666 | n10668 ;
  assign n10670 = n1373 & n10669 ;
  assign n10671 = n4361 ^ n2315 ^ 1'b0 ;
  assign n10672 = n1112 & n10671 ;
  assign n10673 = n7868 ^ n7557 ^ 1'b0 ;
  assign n10674 = n6131 | n9619 ;
  assign n10675 = n6744 | n10674 ;
  assign n10676 = n10673 & ~n10675 ;
  assign n10677 = n2158 ^ n599 ^ 1'b0 ;
  assign n10678 = n1545 | n10677 ;
  assign n10679 = ( ~n742 & n1829 ) | ( ~n742 & n10678 ) | ( n1829 & n10678 ) ;
  assign n10680 = n4298 ^ n3795 ^ 1'b0 ;
  assign n10681 = n10680 ^ n1075 ^ n1065 ;
  assign n10682 = n4906 | n10272 ;
  assign n10683 = n3611 & ~n10682 ;
  assign n10684 = n4861 | n10683 ;
  assign n10685 = n10684 ^ n7796 ^ 1'b0 ;
  assign n10686 = ~n3827 & n7117 ;
  assign n10687 = ~n6294 & n10686 ;
  assign n10689 = n7771 ^ n2733 ^ n298 ;
  assign n10688 = n8114 ^ n7203 ^ 1'b0 ;
  assign n10690 = n10689 ^ n10688 ^ n3553 ;
  assign n10691 = n9370 ^ n2710 ^ 1'b0 ;
  assign n10692 = n6829 | n10691 ;
  assign n10693 = n10692 ^ n7083 ^ n5328 ;
  assign n10694 = n10693 ^ n10335 ^ 1'b0 ;
  assign n10695 = n7785 ^ n1575 ^ 1'b0 ;
  assign n10696 = n4793 & n10695 ;
  assign n10698 = n8538 ^ n6294 ^ n5382 ;
  assign n10699 = n10698 ^ n3760 ^ 1'b0 ;
  assign n10700 = n10699 ^ n1162 ^ 1'b0 ;
  assign n10697 = n5141 | n7187 ;
  assign n10701 = n10700 ^ n10697 ^ 1'b0 ;
  assign n10702 = n10101 ^ n725 ^ 1'b0 ;
  assign n10703 = n6055 | n10702 ;
  assign n10704 = n3387 & ~n5432 ;
  assign n10714 = n2702 ^ x83 ^ 1'b0 ;
  assign n10715 = n7894 & n10714 ;
  assign n10710 = x28 & ~n631 ;
  assign n10711 = ~n4521 & n10710 ;
  assign n10712 = n9569 | n10711 ;
  assign n10713 = n5070 | n10712 ;
  assign n10706 = ( x19 & n1047 ) | ( x19 & n1733 ) | ( n1047 & n1733 ) ;
  assign n10707 = ~n4114 & n10706 ;
  assign n10708 = n10707 ^ n3425 ^ 1'b0 ;
  assign n10705 = n7949 & ~n8064 ;
  assign n10709 = n10708 ^ n10705 ^ 1'b0 ;
  assign n10716 = n10715 ^ n10713 ^ n10709 ;
  assign n10717 = n2053 & n10716 ;
  assign n10718 = ~n10704 & n10717 ;
  assign n10719 = ~n2296 & n2449 ;
  assign n10720 = n10719 ^ n8507 ^ 1'b0 ;
  assign n10721 = n908 & n2316 ;
  assign n10722 = ~n10720 & n10721 ;
  assign n10723 = n3009 ^ n518 ^ n153 ;
  assign n10724 = n3755 & n10723 ;
  assign n10725 = n7147 | n10724 ;
  assign n10726 = ( ~n5438 & n10526 ) | ( ~n5438 & n10558 ) | ( n10526 & n10558 ) ;
  assign n10727 = ( n3954 & n9710 ) | ( n3954 & ~n10726 ) | ( n9710 & ~n10726 ) ;
  assign n10728 = ~n1073 & n3218 ;
  assign n10729 = ~n6718 & n10728 ;
  assign n10730 = n3300 ^ n155 ^ 1'b0 ;
  assign n10731 = ~n10729 & n10730 ;
  assign n10732 = n6199 & ~n10211 ;
  assign n10733 = n1828 | n10732 ;
  assign n10734 = n10731 | n10733 ;
  assign n10735 = n6424 ^ n2798 ^ 1'b0 ;
  assign n10736 = n10734 & ~n10735 ;
  assign n10737 = ~n5596 & n9628 ;
  assign n10738 = n3693 ^ n1513 ^ 1'b0 ;
  assign n10739 = n8804 | n10738 ;
  assign n10740 = n10737 & ~n10739 ;
  assign n10741 = n1163 & n10740 ;
  assign n10742 = n8105 ^ n3916 ^ n1695 ;
  assign n10744 = n4154 & ~n9509 ;
  assign n10745 = n10744 ^ n193 ^ 1'b0 ;
  assign n10743 = n356 & n1725 ;
  assign n10746 = n10745 ^ n10743 ^ 1'b0 ;
  assign n10747 = ( n4698 & n8049 ) | ( n4698 & n8229 ) | ( n8049 & n8229 ) ;
  assign n10748 = n10747 ^ n8988 ^ 1'b0 ;
  assign n10749 = ~n1940 & n10748 ;
  assign n10750 = ~n2265 & n10749 ;
  assign n10756 = n9919 ^ n1733 ^ n1713 ;
  assign n10757 = ( ~n3932 & n5003 ) | ( ~n3932 & n10756 ) | ( n5003 & n10756 ) ;
  assign n10751 = n4585 ^ n3287 ^ n1386 ;
  assign n10752 = n3763 & n6402 ;
  assign n10753 = n3015 | n10752 ;
  assign n10754 = ~n10751 & n10753 ;
  assign n10755 = ~n1207 & n10754 ;
  assign n10758 = n10757 ^ n10755 ^ 1'b0 ;
  assign n10759 = ~n1266 & n2171 ;
  assign n10760 = n4716 | n4797 ;
  assign n10761 = n2712 & ~n3264 ;
  assign n10762 = n10761 ^ n1512 ^ 1'b0 ;
  assign n10763 = ~n4673 & n9409 ;
  assign n10764 = n10763 ^ n8654 ^ 1'b0 ;
  assign n10765 = ~n7462 & n10764 ;
  assign n10766 = n10765 ^ n4970 ^ 1'b0 ;
  assign n10767 = n10762 & n10766 ;
  assign n10768 = n2086 | n3734 ;
  assign n10769 = n950 | n7960 ;
  assign n10770 = n5423 ^ x10 ^ 1'b0 ;
  assign n10771 = n10769 & n10770 ;
  assign n10772 = n10768 & n10771 ;
  assign n10773 = n1431 | n10772 ;
  assign n10779 = n3109 & ~n7716 ;
  assign n10780 = n10779 ^ n992 ^ 1'b0 ;
  assign n10774 = ~n626 & n2085 ;
  assign n10775 = ( n4091 & n5559 ) | ( n4091 & n6158 ) | ( n5559 & n6158 ) ;
  assign n10776 = n10775 ^ n7827 ^ 1'b0 ;
  assign n10777 = n3574 & n10776 ;
  assign n10778 = n10774 & n10777 ;
  assign n10781 = n10780 ^ n10778 ^ 1'b0 ;
  assign n10782 = ( n5230 & n8425 ) | ( n5230 & n10781 ) | ( n8425 & n10781 ) ;
  assign n10783 = n4356 ^ n3294 ^ n131 ;
  assign n10784 = n7413 | n10783 ;
  assign n10785 = ( ~n2493 & n9862 ) | ( ~n2493 & n10784 ) | ( n9862 & n10784 ) ;
  assign n10788 = n9233 ^ n735 ^ 1'b0 ;
  assign n10789 = n10788 ^ n8709 ^ n8334 ;
  assign n10790 = n10789 ^ n4527 ^ 1'b0 ;
  assign n10786 = n6668 | n8418 ;
  assign n10787 = n1542 | n10786 ;
  assign n10791 = n10790 ^ n10787 ^ 1'b0 ;
  assign n10794 = ( n497 & n3274 ) | ( n497 & n5252 ) | ( n3274 & n5252 ) ;
  assign n10795 = n10794 ^ n4810 ^ 1'b0 ;
  assign n10792 = n597 | n9591 ;
  assign n10793 = n10792 ^ n1802 ^ 1'b0 ;
  assign n10796 = n10795 ^ n10793 ^ n3505 ;
  assign n10797 = n611 | n9943 ;
  assign n10798 = n2960 | n10797 ;
  assign n10799 = n5522 & ~n10798 ;
  assign n10800 = n5617 ^ n1868 ^ 1'b0 ;
  assign n10801 = n10800 ^ n7116 ^ 1'b0 ;
  assign n10802 = n9887 | n10801 ;
  assign n10803 = n3037 | n8780 ;
  assign n10804 = n2432 | n10803 ;
  assign n10805 = n5349 & ~n10804 ;
  assign n10806 = n10805 ^ n5995 ^ n2335 ;
  assign n10807 = n881 | n909 ;
  assign n10808 = ( n1222 & n1992 ) | ( n1222 & n10807 ) | ( n1992 & n10807 ) ;
  assign n10809 = n8082 ^ n6032 ^ n1100 ;
  assign n10810 = n6382 & ~n7796 ;
  assign n10811 = ~n10809 & n10810 ;
  assign n10812 = n267 | n1196 ;
  assign n10813 = n10812 ^ n2466 ^ 1'b0 ;
  assign n10814 = n4404 | n4463 ;
  assign n10815 = n2456 | n10814 ;
  assign n10816 = n10813 & n10815 ;
  assign n10817 = n10816 ^ n6614 ^ 1'b0 ;
  assign n10818 = ( x102 & n2512 ) | ( x102 & ~n9271 ) | ( n2512 & ~n9271 ) ;
  assign n10819 = n243 & ~n10818 ;
  assign n10820 = n10819 ^ n3241 ^ 1'b0 ;
  assign n10821 = x90 & n160 ;
  assign n10822 = n1884 | n2552 ;
  assign n10823 = n7152 & n10822 ;
  assign n10824 = n730 & n6645 ;
  assign n10825 = n1216 | n1795 ;
  assign n10826 = n10824 | n10825 ;
  assign n10827 = n8656 & ~n10826 ;
  assign n10828 = n8145 | n8526 ;
  assign n10829 = n9475 | n10828 ;
  assign n10830 = n10613 ^ n5960 ^ 1'b0 ;
  assign n10831 = x85 & n10830 ;
  assign n10832 = ~n529 & n10831 ;
  assign n10833 = n8021 ^ n7640 ^ 1'b0 ;
  assign n10834 = ( x70 & ~n1998 ) | ( x70 & n8071 ) | ( ~n1998 & n8071 ) ;
  assign n10835 = ~n1107 & n6826 ;
  assign n10836 = n1511 & n10835 ;
  assign n10837 = ( n1165 & n1832 ) | ( n1165 & n10836 ) | ( n1832 & n10836 ) ;
  assign n10838 = n7094 ^ n322 ^ 1'b0 ;
  assign n10839 = n2304 & ~n10838 ;
  assign n10840 = ( n8508 & n10837 ) | ( n8508 & n10839 ) | ( n10837 & n10839 ) ;
  assign n10841 = ( n548 & ~n1101 ) | ( n548 & n1348 ) | ( ~n1101 & n1348 ) ;
  assign n10842 = n10142 & ~n10841 ;
  assign n10843 = ~n10840 & n10842 ;
  assign n10844 = n10834 | n10843 ;
  assign n10845 = n10833 & ~n10844 ;
  assign n10849 = ~n708 & n1791 ;
  assign n10846 = n1184 ^ n832 ^ 1'b0 ;
  assign n10847 = n5952 | n7989 ;
  assign n10848 = ( n3096 & ~n10846 ) | ( n3096 & n10847 ) | ( ~n10846 & n10847 ) ;
  assign n10850 = n10849 ^ n10848 ^ 1'b0 ;
  assign n10851 = ~n2246 & n10850 ;
  assign n10852 = n1552 | n10284 ;
  assign n10853 = n6163 ^ n729 ^ 1'b0 ;
  assign n10854 = n4445 ^ n3090 ^ 1'b0 ;
  assign n10855 = n5451 ^ n2948 ^ n1748 ;
  assign n10856 = ( n441 & ~n10854 ) | ( n441 & n10855 ) | ( ~n10854 & n10855 ) ;
  assign n10857 = n6558 ^ n5376 ^ n3169 ;
  assign n10858 = n10078 | n10857 ;
  assign n10859 = n1722 & ~n6671 ;
  assign n10862 = ( ~n2905 & n4937 ) | ( ~n2905 & n6128 ) | ( n4937 & n6128 ) ;
  assign n10860 = n967 & ~n8763 ;
  assign n10861 = n4370 & n10860 ;
  assign n10863 = n10862 ^ n10861 ^ 1'b0 ;
  assign n10864 = ~n7241 & n9557 ;
  assign n10865 = n587 & n2731 ;
  assign n10866 = n587 & n3731 ;
  assign n10867 = n719 & n10866 ;
  assign n10868 = n10867 ^ n7359 ^ 1'b0 ;
  assign n10869 = n824 | n10868 ;
  assign n10870 = ( ~n10864 & n10865 ) | ( ~n10864 & n10869 ) | ( n10865 & n10869 ) ;
  assign n10871 = n2090 & n7292 ;
  assign n10872 = n5449 ^ n4979 ^ 1'b0 ;
  assign n10873 = ~n2917 & n10872 ;
  assign n10874 = n2345 | n2497 ;
  assign n10875 = n6004 & ~n10874 ;
  assign n10876 = n1706 | n10875 ;
  assign n10877 = n10873 | n10876 ;
  assign n10878 = n5870 & n10877 ;
  assign n10879 = n9260 | n10302 ;
  assign n10880 = n9924 & ~n10879 ;
  assign n10881 = n2076 ^ n1719 ^ n381 ;
  assign n10882 = n3442 & ~n10881 ;
  assign n10888 = ~n1481 & n1677 ;
  assign n10889 = n3942 & n10888 ;
  assign n10890 = n10889 ^ n697 ^ 1'b0 ;
  assign n10883 = n1581 & n2167 ;
  assign n10884 = n10883 ^ n3540 ^ 1'b0 ;
  assign n10885 = ~n6172 & n10884 ;
  assign n10886 = n254 & n10885 ;
  assign n10887 = n10886 ^ n3062 ^ 1'b0 ;
  assign n10891 = n10890 ^ n10887 ^ n7935 ;
  assign n10892 = n2264 & n7225 ;
  assign n10893 = n9533 ^ n2251 ^ n1633 ;
  assign n10894 = n2422 & ~n10139 ;
  assign n10895 = n1888 ^ n1233 ^ 1'b0 ;
  assign n10896 = n9560 | n10895 ;
  assign n10897 = n1515 & ~n6993 ;
  assign n10898 = n10207 ^ n6201 ^ 1'b0 ;
  assign n10899 = n1817 | n9325 ;
  assign n10900 = n9144 | n10899 ;
  assign n10901 = n5448 & n10900 ;
  assign n10902 = n1865 | n1911 ;
  assign n10903 = n10902 ^ n5792 ^ 1'b0 ;
  assign n10904 = n8637 ^ n2731 ^ 1'b0 ;
  assign n10905 = ~n10903 & n10904 ;
  assign n10906 = n10905 ^ n2960 ^ 1'b0 ;
  assign n10907 = n8437 & ~n10906 ;
  assign n10908 = n5228 ^ n2995 ^ x1 ;
  assign n10909 = n5103 | n10908 ;
  assign n10910 = n704 | n4204 ;
  assign n10913 = n256 & ~n2310 ;
  assign n10914 = n10913 ^ n181 ^ 1'b0 ;
  assign n10911 = n1257 & n3423 ;
  assign n10912 = n10911 ^ n3871 ^ 1'b0 ;
  assign n10915 = n10914 ^ n10912 ^ 1'b0 ;
  assign n10916 = n10910 & n10915 ;
  assign n10917 = n954 & n5517 ;
  assign n10918 = n3470 & n10917 ;
  assign n10919 = n10462 ^ n7491 ^ n6283 ;
  assign n10920 = n9203 & ~n10919 ;
  assign n10921 = n10920 ^ n327 ^ 1'b0 ;
  assign n10922 = n8121 ^ n4879 ^ n2202 ;
  assign n10923 = ( n9013 & ~n10503 ) | ( n9013 & n10922 ) | ( ~n10503 & n10922 ) ;
  assign n10924 = n10923 ^ n7023 ^ 1'b0 ;
  assign n10925 = n637 & n4422 ;
  assign n10926 = n7640 ^ n5291 ^ n5214 ;
  assign n10927 = n4365 & ~n6034 ;
  assign n10928 = ~n10926 & n10927 ;
  assign n10929 = n3372 ^ n2182 ^ 1'b0 ;
  assign n10930 = n5050 ^ n5014 ^ 1'b0 ;
  assign n10931 = n10929 | n10930 ;
  assign n10932 = n3392 ^ n905 ^ 1'b0 ;
  assign n10933 = n9913 ^ x6 ^ 1'b0 ;
  assign n10934 = n8801 & n10933 ;
  assign n10935 = ~n5021 & n10934 ;
  assign n10936 = n7605 & ~n10610 ;
  assign n10937 = n10936 ^ n4686 ^ 1'b0 ;
  assign n10938 = ~n9728 & n10937 ;
  assign n10939 = n410 | n1918 ;
  assign n10940 = n10939 ^ n712 ^ 1'b0 ;
  assign n10942 = n1104 ^ n361 ^ 1'b0 ;
  assign n10943 = n4865 & ~n10942 ;
  assign n10941 = n5725 ^ n5382 ^ n4649 ;
  assign n10944 = n10943 ^ n10941 ^ 1'b0 ;
  assign n10945 = ~n9667 & n10944 ;
  assign n10946 = n10777 ^ n1567 ^ 1'b0 ;
  assign n10947 = n4815 ^ n219 ^ 1'b0 ;
  assign n10948 = n10581 ^ n1920 ^ 1'b0 ;
  assign n10949 = n1325 | n10948 ;
  assign n10950 = n10949 ^ n2296 ^ 1'b0 ;
  assign n10951 = n10950 ^ n768 ^ 1'b0 ;
  assign n10952 = n10951 ^ n1567 ^ n1093 ;
  assign n10953 = ~n1748 & n3017 ;
  assign n10954 = n10953 ^ n5327 ^ 1'b0 ;
  assign n10955 = ~n6498 & n8728 ;
  assign n10956 = n9242 & ~n10955 ;
  assign n10957 = n2111 | n6881 ;
  assign n10958 = n10957 ^ n5196 ^ 1'b0 ;
  assign n10959 = ( ~n1331 & n2180 ) | ( ~n1331 & n10958 ) | ( n2180 & n10958 ) ;
  assign n10960 = n9649 ^ n971 ^ 1'b0 ;
  assign n10961 = ~n10959 & n10960 ;
  assign n10962 = ~n4860 & n9178 ;
  assign n10963 = n4793 & ~n8882 ;
  assign n10964 = n6225 & ~n8987 ;
  assign n10965 = n5965 & n10964 ;
  assign n10966 = ( ~n354 & n8176 ) | ( ~n354 & n10965 ) | ( n8176 & n10965 ) ;
  assign n10967 = n6229 & ~n9112 ;
  assign n10968 = n187 & ~n3345 ;
  assign n10969 = n7711 & n10968 ;
  assign n10970 = n252 & ~n10969 ;
  assign n10971 = n10970 ^ n7277 ^ n6861 ;
  assign n10972 = ( n1700 & ~n5925 ) | ( n1700 & n6447 ) | ( ~n5925 & n6447 ) ;
  assign n10973 = n10971 | n10972 ;
  assign n10974 = ( n139 & n1398 ) | ( n139 & n1798 ) | ( n1398 & n1798 ) ;
  assign n10975 = n10974 ^ n8562 ^ n1322 ;
  assign n10976 = ~n9912 & n10975 ;
  assign n10977 = n10976 ^ n5235 ^ 1'b0 ;
  assign n10978 = n3860 ^ n1493 ^ 1'b0 ;
  assign n10979 = n5332 ^ n4083 ^ 1'b0 ;
  assign n10980 = n10978 & ~n10979 ;
  assign n10981 = ( n1244 & n5740 ) | ( n1244 & ~n10980 ) | ( n5740 & ~n10980 ) ;
  assign n10982 = n7557 ^ n6992 ^ n186 ;
  assign n10983 = n4231 & ~n10982 ;
  assign n10984 = n10983 ^ n2004 ^ 1'b0 ;
  assign n10985 = n4070 ^ n4048 ^ 1'b0 ;
  assign n10986 = ( n721 & n1895 ) | ( n721 & n2651 ) | ( n1895 & n2651 ) ;
  assign n10987 = n1722 | n8721 ;
  assign n10988 = ( n3658 & ~n10986 ) | ( n3658 & n10987 ) | ( ~n10986 & n10987 ) ;
  assign n10989 = ~n1563 & n3823 ;
  assign n10990 = ~n436 & n10989 ;
  assign n10991 = ~n5152 & n6928 ;
  assign n10992 = n353 & n3221 ;
  assign n10993 = n10991 & n10992 ;
  assign n10994 = n10993 ^ n10723 ^ 1'b0 ;
  assign n10995 = n10994 ^ n2544 ^ 1'b0 ;
  assign n10997 = x116 & ~n758 ;
  assign n10998 = n10997 ^ n1887 ^ 1'b0 ;
  assign n10996 = ~n2538 & n6527 ;
  assign n10999 = n10998 ^ n10996 ^ 1'b0 ;
  assign n11000 = n10497 ^ n4521 ^ 1'b0 ;
  assign n11001 = n429 & ~n535 ;
  assign n11002 = ( n1279 & ~n9496 ) | ( n1279 & n11001 ) | ( ~n9496 & n11001 ) ;
  assign n11006 = n1718 | n4754 ;
  assign n11007 = n11006 ^ n2930 ^ 1'b0 ;
  assign n11003 = n1567 ^ n892 ^ 1'b0 ;
  assign n11004 = n1629 | n11003 ;
  assign n11005 = n11004 ^ n6924 ^ n1663 ;
  assign n11008 = n11007 ^ n11005 ^ n4995 ;
  assign n11009 = n7105 ^ n6760 ^ 1'b0 ;
  assign n11010 = n11008 & ~n11009 ;
  assign n11011 = n11010 ^ n5128 ^ 1'b0 ;
  assign n11012 = n824 & n11011 ;
  assign n11013 = n3383 | n5061 ;
  assign n11014 = n8960 ^ n2769 ^ 1'b0 ;
  assign n11015 = n1167 & ~n11014 ;
  assign n11016 = ( n6552 & n8158 ) | ( n6552 & n11015 ) | ( n8158 & n11015 ) ;
  assign n11026 = ~n569 & n2496 ;
  assign n11027 = ~n988 & n11026 ;
  assign n11028 = ( ~n3456 & n5610 ) | ( ~n3456 & n11027 ) | ( n5610 & n11027 ) ;
  assign n11019 = n2457 & n7246 ;
  assign n11020 = ~n395 & n11019 ;
  assign n11021 = n11020 ^ n3317 ^ 1'b0 ;
  assign n11018 = n1829 & ~n6969 ;
  assign n11022 = n11021 ^ n11018 ^ 1'b0 ;
  assign n11023 = n1890 | n4411 ;
  assign n11024 = n11022 | n11023 ;
  assign n11025 = ~n5425 & n11024 ;
  assign n11029 = n11028 ^ n11025 ^ 1'b0 ;
  assign n11017 = n620 | n6493 ;
  assign n11030 = n11029 ^ n11017 ^ 1'b0 ;
  assign n11031 = n3413 | n6229 ;
  assign n11032 = n7468 ^ n3724 ^ 1'b0 ;
  assign n11033 = n1299 | n11032 ;
  assign n11034 = n11031 | n11033 ;
  assign n11035 = n4252 ^ n3925 ^ 1'b0 ;
  assign n11036 = x5 & ~n11035 ;
  assign n11037 = ~n4107 & n11036 ;
  assign n11038 = n7366 & ~n11037 ;
  assign n11039 = ~n7939 & n10255 ;
  assign n11040 = n5703 ^ n5180 ^ n4756 ;
  assign n11041 = n131 & n5920 ;
  assign n11042 = n6917 & n11041 ;
  assign n11043 = n11040 & ~n11042 ;
  assign n11044 = ~n11039 & n11043 ;
  assign n11049 = n9772 ^ n3365 ^ n220 ;
  assign n11050 = ( n1825 & n9673 ) | ( n1825 & ~n11049 ) | ( n9673 & ~n11049 ) ;
  assign n11051 = n1283 | n3472 ;
  assign n11052 = ~n4238 & n11051 ;
  assign n11053 = ~n11050 & n11052 ;
  assign n11045 = n2527 ^ n131 ^ 1'b0 ;
  assign n11046 = ( n1722 & n2083 ) | ( n1722 & ~n4473 ) | ( n2083 & ~n4473 ) ;
  assign n11047 = n11046 ^ n7083 ^ 1'b0 ;
  assign n11048 = ( n1390 & ~n11045 ) | ( n1390 & n11047 ) | ( ~n11045 & n11047 ) ;
  assign n11054 = n11053 ^ n11048 ^ n3202 ;
  assign n11057 = ~n1354 & n3076 ;
  assign n11058 = n11057 ^ n4884 ^ 1'b0 ;
  assign n11059 = ~n2868 & n4035 ;
  assign n11060 = n11058 & n11059 ;
  assign n11055 = ( n1200 & ~n4897 ) | ( n1200 & n7992 ) | ( ~n4897 & n7992 ) ;
  assign n11056 = n11055 ^ n415 ^ 1'b0 ;
  assign n11061 = n11060 ^ n11056 ^ 1'b0 ;
  assign n11062 = x13 | n883 ;
  assign n11063 = n6076 ^ n5680 ^ 1'b0 ;
  assign n11064 = n8668 | n9933 ;
  assign n11065 = n11063 | n11064 ;
  assign n11066 = ~n4179 & n9872 ;
  assign n11067 = n11066 ^ n6272 ^ 1'b0 ;
  assign n11068 = n11067 ^ n9710 ^ 1'b0 ;
  assign n11069 = n4211 ^ n4085 ^ n1946 ;
  assign n11070 = n11069 ^ n6600 ^ n3661 ;
  assign n11071 = n9544 | n11070 ;
  assign n11072 = n11071 ^ n5615 ^ 1'b0 ;
  assign n11073 = n2653 ^ n2025 ^ 1'b0 ;
  assign n11074 = n11072 & ~n11073 ;
  assign n11075 = n4169 & ~n11074 ;
  assign n11076 = n2332 & ~n9062 ;
  assign n11077 = n2859 & ~n5681 ;
  assign n11078 = n11077 ^ n2738 ^ 1'b0 ;
  assign n11079 = n11078 ^ n5108 ^ 1'b0 ;
  assign n11081 = n8630 ^ n5973 ^ n467 ;
  assign n11080 = n1157 & ~n4103 ;
  assign n11082 = n11081 ^ n11080 ^ 1'b0 ;
  assign n11083 = n2335 & n11082 ;
  assign n11084 = n11083 ^ x60 ^ 1'b0 ;
  assign n11085 = n5653 & ~n10139 ;
  assign n11086 = n384 & n11085 ;
  assign n11087 = n11086 ^ n7842 ^ 1'b0 ;
  assign n11088 = ~n11084 & n11087 ;
  assign n11089 = ( ~n920 & n3550 ) | ( ~n920 & n5257 ) | ( n3550 & n5257 ) ;
  assign n11090 = n6638 | n11089 ;
  assign n11091 = n8936 ^ n5056 ^ 1'b0 ;
  assign n11092 = n2303 & n11091 ;
  assign n11094 = n1704 | n2986 ;
  assign n11095 = n2715 & ~n11094 ;
  assign n11093 = ~n270 & n746 ;
  assign n11096 = n11095 ^ n11093 ^ 1'b0 ;
  assign n11097 = ( x54 & ~n1772 ) | ( x54 & n7162 ) | ( ~n1772 & n7162 ) ;
  assign n11098 = n11097 ^ n5686 ^ 1'b0 ;
  assign n11099 = n11098 ^ n7268 ^ n158 ;
  assign n11100 = n6283 & n11099 ;
  assign n11101 = ( ~n7193 & n9244 ) | ( ~n7193 & n11100 ) | ( n9244 & n11100 ) ;
  assign n11102 = n2197 & n11101 ;
  assign n11103 = n9014 & n11102 ;
  assign n11104 = n6156 & ~n10376 ;
  assign n11108 = ( n4561 & n5589 ) | ( n4561 & ~n6575 ) | ( n5589 & ~n6575 ) ;
  assign n11109 = n11108 ^ n4724 ^ n395 ;
  assign n11105 = n2397 & ~n10883 ;
  assign n11106 = n6885 & n11105 ;
  assign n11107 = n11106 ^ n3184 ^ 1'b0 ;
  assign n11110 = n11109 ^ n11107 ^ n8037 ;
  assign n11111 = n10602 ^ n172 ^ 1'b0 ;
  assign n11112 = ~n5219 & n11111 ;
  assign n11113 = n4674 ^ x118 ^ 1'b0 ;
  assign n11114 = n6640 | n11113 ;
  assign n11115 = n9623 ^ n1915 ^ n1776 ;
  assign n11116 = ~n5554 & n6915 ;
  assign n11117 = n11116 ^ n3173 ^ 1'b0 ;
  assign n11118 = ~n11115 & n11117 ;
  assign n11119 = n5423 & n11118 ;
  assign n11120 = n6083 & ~n11119 ;
  assign n11121 = n11120 ^ n1763 ^ 1'b0 ;
  assign n11122 = ~n1483 & n10118 ;
  assign n11123 = n11122 ^ n6882 ^ 1'b0 ;
  assign n11124 = n9229 & ~n11123 ;
  assign n11125 = n5665 & ~n10415 ;
  assign n11126 = n1850 | n9630 ;
  assign n11127 = ( n3650 & n8888 ) | ( n3650 & n11126 ) | ( n8888 & n11126 ) ;
  assign n11128 = ~n634 & n9223 ;
  assign n11129 = ~n5935 & n6269 ;
  assign n11130 = n7321 & ~n11129 ;
  assign n11131 = n11130 ^ n3060 ^ 1'b0 ;
  assign n11132 = ( ~n1874 & n4498 ) | ( ~n1874 & n8139 ) | ( n4498 & n8139 ) ;
  assign n11133 = n11132 ^ n3522 ^ 1'b0 ;
  assign n11134 = n9298 | n11133 ;
  assign n11135 = ~n3060 & n3634 ;
  assign n11136 = n11135 ^ x43 ^ 1'b0 ;
  assign n11137 = n11136 ^ n2182 ^ 1'b0 ;
  assign n11138 = n11137 ^ n7551 ^ n2131 ;
  assign n11139 = ( n3254 & n5104 ) | ( n3254 & n7945 ) | ( n5104 & n7945 ) ;
  assign n11140 = ( n2169 & ~n5016 ) | ( n2169 & n6796 ) | ( ~n5016 & n6796 ) ;
  assign n11141 = ( ~n650 & n7020 ) | ( ~n650 & n8645 ) | ( n7020 & n8645 ) ;
  assign n11142 = n6798 ^ n4214 ^ 1'b0 ;
  assign n11148 = n5396 ^ n4437 ^ 1'b0 ;
  assign n11143 = ~n2014 & n3384 ;
  assign n11144 = n11143 ^ n6452 ^ 1'b0 ;
  assign n11145 = n7449 & ~n11144 ;
  assign n11146 = n3172 ^ n2140 ^ 1'b0 ;
  assign n11147 = n11145 & ~n11146 ;
  assign n11149 = n11148 ^ n11147 ^ 1'b0 ;
  assign n11150 = ~n10620 & n11149 ;
  assign n11152 = n9028 ^ n2912 ^ 1'b0 ;
  assign n11153 = n1672 | n11152 ;
  assign n11154 = n11153 ^ n4669 ^ 1'b0 ;
  assign n11155 = ~n5765 & n11154 ;
  assign n11156 = ~n1531 & n3261 ;
  assign n11157 = n1692 & n11156 ;
  assign n11158 = ~n7268 & n11157 ;
  assign n11159 = n11158 ^ n2819 ^ 1'b0 ;
  assign n11160 = n11155 & ~n11159 ;
  assign n11151 = n809 & n8341 ;
  assign n11161 = n11160 ^ n11151 ^ n5354 ;
  assign n11162 = ( n3525 & n10496 ) | ( n3525 & n11161 ) | ( n10496 & n11161 ) ;
  assign n11163 = n6388 ^ x115 ^ 1'b0 ;
  assign n11164 = n11163 ^ n5822 ^ n809 ;
  assign n11165 = n1893 ^ n332 ^ 1'b0 ;
  assign n11166 = n11165 ^ n7125 ^ n4594 ;
  assign n11167 = n4349 ^ n1856 ^ 1'b0 ;
  assign n11168 = n1444 & n11167 ;
  assign n11169 = ~n11166 & n11168 ;
  assign n11170 = n7837 & n11169 ;
  assign n11171 = ( ~n9665 & n11164 ) | ( ~n9665 & n11170 ) | ( n11164 & n11170 ) ;
  assign n11172 = ~n6049 & n9759 ;
  assign n11173 = n4826 & n11172 ;
  assign n11174 = n211 & ~n3722 ;
  assign n11175 = n11045 ^ n3999 ^ 1'b0 ;
  assign n11176 = n4821 & n11175 ;
  assign n11177 = ( n2890 & n8467 ) | ( n2890 & n10268 ) | ( n8467 & n10268 ) ;
  assign n11178 = n11177 ^ n9215 ^ 1'b0 ;
  assign n11179 = n2598 & ~n11178 ;
  assign n11180 = n11179 ^ n4131 ^ 1'b0 ;
  assign n11181 = n11176 & ~n11180 ;
  assign n11182 = ( x125 & n601 ) | ( x125 & ~n8592 ) | ( n601 & ~n8592 ) ;
  assign n11183 = n11182 ^ n5858 ^ 1'b0 ;
  assign n11184 = ( n2992 & n5587 ) | ( n2992 & n8809 ) | ( n5587 & n8809 ) ;
  assign n11185 = ~n475 & n6133 ;
  assign n11186 = n11185 ^ x70 ^ 1'b0 ;
  assign n11187 = ( n1000 & n7604 ) | ( n1000 & n11186 ) | ( n7604 & n11186 ) ;
  assign n11188 = n11187 ^ n8173 ^ 1'b0 ;
  assign n11189 = n3274 & n11188 ;
  assign n11190 = n9847 ^ n4696 ^ n4106 ;
  assign n11191 = n4915 | n11190 ;
  assign n11192 = n11189 | n11191 ;
  assign n11193 = n165 & n6306 ;
  assign n11194 = n6110 & ~n11193 ;
  assign n11195 = n11194 ^ n6072 ^ 1'b0 ;
  assign n11196 = n4209 | n11195 ;
  assign n11197 = n383 | n843 ;
  assign n11198 = n4213 & ~n11197 ;
  assign n11199 = n11198 ^ n10190 ^ n5730 ;
  assign n11200 = ~n1733 & n10188 ;
  assign n11201 = ~n9380 & n11200 ;
  assign n11202 = n6104 ^ n6088 ^ 1'b0 ;
  assign n11204 = n1517 | n3142 ;
  assign n11205 = n11204 ^ n4456 ^ 1'b0 ;
  assign n11206 = n4037 & ~n11205 ;
  assign n11207 = n11206 ^ n10202 ^ n2148 ;
  assign n11203 = n10881 ^ n10040 ^ n882 ;
  assign n11208 = n11207 ^ n11203 ^ n6032 ;
  assign n11209 = n3615 ^ n3103 ^ n236 ;
  assign n11210 = n11209 ^ n6999 ^ n5792 ;
  assign n11211 = n1845 | n8553 ;
  assign n11212 = n3610 & ~n11211 ;
  assign n11213 = ~n8664 & n11212 ;
  assign n11214 = n6946 & ~n8871 ;
  assign n11215 = ~n9797 & n11214 ;
  assign n11216 = n4946 & ~n11215 ;
  assign n11217 = n11216 ^ n949 ^ 1'b0 ;
  assign n11218 = n7650 ^ n2976 ^ 1'b0 ;
  assign n11219 = n6919 ^ n911 ^ 1'b0 ;
  assign n11220 = ~n956 & n7614 ;
  assign n11221 = n11220 ^ n4126 ^ 1'b0 ;
  assign n11222 = ~n4250 & n11221 ;
  assign n11223 = n11219 & n11222 ;
  assign n11224 = n747 | n2566 ;
  assign n11225 = ( n1675 & ~n10028 ) | ( n1675 & n11224 ) | ( ~n10028 & n11224 ) ;
  assign n11226 = n8955 ^ n8724 ^ n4708 ;
  assign n11227 = ( ~n6260 & n7834 ) | ( ~n6260 & n11226 ) | ( n7834 & n11226 ) ;
  assign n11228 = n2760 | n4346 ;
  assign n11229 = n11228 ^ n8004 ^ 1'b0 ;
  assign n11230 = n1274 & ~n11229 ;
  assign n11231 = x10 & ~n3543 ;
  assign n11232 = n11231 ^ n3035 ^ 1'b0 ;
  assign n11233 = n1371 & n3975 ;
  assign n11234 = n4618 ^ n2053 ^ 1'b0 ;
  assign n11235 = n3710 & ~n11234 ;
  assign n11236 = n279 & n11235 ;
  assign n11237 = n11236 ^ n3575 ^ 1'b0 ;
  assign n11238 = n11233 & n11237 ;
  assign n11239 = ~n11232 & n11238 ;
  assign n11240 = n11230 & n11239 ;
  assign n11241 = n6796 ^ n1201 ^ 1'b0 ;
  assign n11242 = n11241 ^ n5417 ^ n1448 ;
  assign n11243 = n1675 & n5894 ;
  assign n11244 = n11242 & n11243 ;
  assign n11245 = n10833 ^ n6068 ^ 1'b0 ;
  assign n11246 = n3299 & ~n11245 ;
  assign n11247 = n319 & n3686 ;
  assign n11249 = n11230 ^ n7437 ^ n4605 ;
  assign n11248 = n5293 & ~n5537 ;
  assign n11250 = n11249 ^ n11248 ^ 1'b0 ;
  assign n11251 = n3420 & n5641 ;
  assign n11252 = n8522 ^ n2200 ^ 1'b0 ;
  assign n11254 = ( x112 & n700 ) | ( x112 & ~n1528 ) | ( n700 & ~n1528 ) ;
  assign n11253 = n7554 ^ n5860 ^ n3689 ;
  assign n11255 = n11254 ^ n11253 ^ 1'b0 ;
  assign n11256 = n3961 & ~n10613 ;
  assign n11257 = n3826 | n4263 ;
  assign n11258 = n11256 | n11257 ;
  assign n11259 = ~n2974 & n4917 ;
  assign n11260 = n5611 & n11259 ;
  assign n11261 = ( ~n5092 & n8263 ) | ( ~n5092 & n11259 ) | ( n8263 & n11259 ) ;
  assign n11262 = n10338 | n11261 ;
  assign n11263 = n7311 | n11262 ;
  assign n11264 = n6123 ^ n2927 ^ n2191 ;
  assign n11265 = n8503 ^ n953 ^ 1'b0 ;
  assign n11266 = n7479 & n11265 ;
  assign n11267 = n11266 ^ n9702 ^ n7174 ;
  assign n11268 = ( ~n885 & n1861 ) | ( ~n885 & n3382 ) | ( n1861 & n3382 ) ;
  assign n11269 = n684 ^ n576 ^ 1'b0 ;
  assign n11270 = ~n4790 & n11269 ;
  assign n11271 = n11270 ^ n5118 ^ 1'b0 ;
  assign n11272 = n9271 ^ n8076 ^ 1'b0 ;
  assign n11273 = n7488 & ~n11272 ;
  assign n11274 = n11273 ^ n2926 ^ 1'b0 ;
  assign n11275 = n7970 ^ n6264 ^ 1'b0 ;
  assign n11276 = n9072 & ~n11275 ;
  assign n11277 = n7856 & n11276 ;
  assign n11278 = ~n1304 & n5870 ;
  assign n11279 = n11278 ^ n4159 ^ 1'b0 ;
  assign n11280 = n11070 & n11279 ;
  assign n11281 = n2087 | n5879 ;
  assign n11282 = ( n1760 & n3778 ) | ( n1760 & n11281 ) | ( n3778 & n11281 ) ;
  assign n11283 = ( ~n231 & n5776 ) | ( ~n231 & n11282 ) | ( n5776 & n11282 ) ;
  assign n11284 = n11283 ^ n9244 ^ n7670 ;
  assign n11285 = n4554 ^ x115 ^ 1'b0 ;
  assign n11286 = n6783 | n11285 ;
  assign n11287 = n6729 ^ n6207 ^ n1065 ;
  assign n11288 = ( n818 & n9911 ) | ( n818 & ~n11287 ) | ( n9911 & ~n11287 ) ;
  assign n11289 = n11288 ^ n2736 ^ 1'b0 ;
  assign n11290 = n1140 ^ x104 ^ 1'b0 ;
  assign n11291 = n2954 & ~n11290 ;
  assign n11292 = ( ~n1527 & n1772 ) | ( ~n1527 & n8129 ) | ( n1772 & n8129 ) ;
  assign n11293 = n5057 & ~n11292 ;
  assign n11294 = n11291 & ~n11293 ;
  assign n11295 = n11294 ^ n5116 ^ 1'b0 ;
  assign n11296 = n1233 ^ n265 ^ 1'b0 ;
  assign n11297 = ( n232 & ~n1386 ) | ( n232 & n11296 ) | ( ~n1386 & n11296 ) ;
  assign n11298 = ( n817 & n11295 ) | ( n817 & ~n11297 ) | ( n11295 & ~n11297 ) ;
  assign n11299 = ~n2808 & n8995 ;
  assign n11303 = n1929 | n7502 ;
  assign n11304 = n4753 & ~n11303 ;
  assign n11305 = n5583 ^ n739 ^ 1'b0 ;
  assign n11306 = ~n11304 & n11305 ;
  assign n11300 = ~n2333 & n3521 ;
  assign n11301 = ~n726 & n11300 ;
  assign n11302 = n2183 & n11301 ;
  assign n11307 = n11306 ^ n11302 ^ n1880 ;
  assign n11308 = n11307 ^ n10507 ^ 1'b0 ;
  assign n11309 = n2549 | n5847 ;
  assign n11310 = n3182 | n11309 ;
  assign n11311 = n6118 ^ n167 ^ 1'b0 ;
  assign n11312 = n8702 & ~n11311 ;
  assign n11313 = ( n8223 & ~n11310 ) | ( n8223 & n11312 ) | ( ~n11310 & n11312 ) ;
  assign n11314 = ( x92 & n6830 ) | ( x92 & ~n7537 ) | ( n6830 & ~n7537 ) ;
  assign n11315 = n129 & ~n6395 ;
  assign n11316 = n5609 ^ n1788 ^ n882 ;
  assign n11317 = ( ~n1248 & n5447 ) | ( ~n1248 & n11316 ) | ( n5447 & n11316 ) ;
  assign n11318 = n6193 | n6275 ;
  assign n11319 = n5798 | n6628 ;
  assign n11320 = n7763 | n11319 ;
  assign n11321 = n5217 ^ n4566 ^ n1589 ;
  assign n11322 = n1162 | n11321 ;
  assign n11323 = n1090 | n11322 ;
  assign n11324 = ~n1586 & n11323 ;
  assign n11325 = n11324 ^ n316 ^ 1'b0 ;
  assign n11326 = n2991 & ~n3199 ;
  assign n11327 = n10264 ^ n6593 ^ 1'b0 ;
  assign n11328 = ~n10732 & n11327 ;
  assign n11329 = n1079 & n11328 ;
  assign n11330 = n11329 ^ n3961 ^ 1'b0 ;
  assign n11331 = n11326 | n11330 ;
  assign n11332 = n6177 | n6885 ;
  assign n11333 = x100 | n11332 ;
  assign n11334 = n11333 ^ n10665 ^ 1'b0 ;
  assign n11335 = n1712 ^ x78 ^ 1'b0 ;
  assign n11336 = ~n6788 & n11335 ;
  assign n11337 = n10965 ^ n2400 ^ n270 ;
  assign n11348 = n3666 ^ n1442 ^ 1'b0 ;
  assign n11349 = ~n6884 & n11348 ;
  assign n11338 = n7625 | n9139 ;
  assign n11339 = n11338 ^ n10987 ^ 1'b0 ;
  assign n11340 = n1205 ^ x125 ^ 1'b0 ;
  assign n11343 = n2253 ^ n1202 ^ n822 ;
  assign n11341 = n3231 ^ n1327 ^ 1'b0 ;
  assign n11342 = n8164 & n11341 ;
  assign n11344 = n11343 ^ n11342 ^ 1'b0 ;
  assign n11345 = n11340 & ~n11344 ;
  assign n11346 = n11345 ^ n6812 ^ 1'b0 ;
  assign n11347 = n11339 & n11346 ;
  assign n11350 = n11349 ^ n11347 ^ n5132 ;
  assign n11351 = n1495 | n10146 ;
  assign n11352 = n11351 ^ n2523 ^ 1'b0 ;
  assign n11353 = n11352 ^ n816 ^ 1'b0 ;
  assign n11354 = n2913 & ~n11353 ;
  assign n11355 = n10142 ^ n4884 ^ 1'b0 ;
  assign n11356 = ~n484 & n11355 ;
  assign n11357 = n11356 ^ n3592 ^ n210 ;
  assign n11358 = n3334 & n11357 ;
  assign n11359 = n4738 ^ n3262 ^ n1621 ;
  assign n11360 = n5804 ^ n2124 ^ 1'b0 ;
  assign n11361 = n11360 ^ n5785 ^ 1'b0 ;
  assign n11362 = n6412 & n11361 ;
  assign n11363 = n11362 ^ n6675 ^ 1'b0 ;
  assign n11364 = n2125 & ~n7897 ;
  assign n11365 = n11364 ^ n9872 ^ 1'b0 ;
  assign n11366 = n11363 | n11365 ;
  assign n11367 = n4826 ^ n4443 ^ 1'b0 ;
  assign n11368 = n6075 & ~n11367 ;
  assign n11369 = n1517 & n5577 ;
  assign n11370 = n11369 ^ n4829 ^ 1'b0 ;
  assign n11371 = n10476 | n11370 ;
  assign n11372 = n11368 | n11371 ;
  assign n11373 = n6472 ^ n1424 ^ 1'b0 ;
  assign n11374 = n6169 ^ n3181 ^ 1'b0 ;
  assign n11375 = ~n1012 & n11374 ;
  assign n11376 = n11375 ^ n7403 ^ 1'b0 ;
  assign n11377 = n8133 | n11376 ;
  assign n11378 = ( n4636 & n7670 ) | ( n4636 & ~n11193 ) | ( n7670 & ~n11193 ) ;
  assign n11379 = n2172 & n4035 ;
  assign n11380 = n2416 & n11379 ;
  assign n11381 = n11380 ^ n4833 ^ 1'b0 ;
  assign n11382 = n9655 ^ n4527 ^ 1'b0 ;
  assign n11383 = x110 & ~n11382 ;
  assign n11384 = ( n3643 & ~n11381 ) | ( n3643 & n11383 ) | ( ~n11381 & n11383 ) ;
  assign n11385 = n11384 ^ n3821 ^ 1'b0 ;
  assign n11386 = n9401 ^ n1876 ^ 1'b0 ;
  assign n11387 = ( n1448 & ~n3211 ) | ( n1448 & n6953 ) | ( ~n3211 & n6953 ) ;
  assign n11388 = ~n11386 & n11387 ;
  assign n11389 = n11388 ^ n5502 ^ 1'b0 ;
  assign n11390 = ( n6150 & n6258 ) | ( n6150 & n11389 ) | ( n6258 & n11389 ) ;
  assign n11391 = ~x49 & n2591 ;
  assign n11393 = n157 | n5581 ;
  assign n11394 = n3139 & ~n11393 ;
  assign n11392 = n4411 ^ n4242 ^ n809 ;
  assign n11395 = n11394 ^ n11392 ^ n322 ;
  assign n11396 = n7667 | n11395 ;
  assign n11397 = n11391 & ~n11396 ;
  assign n11398 = n3211 | n11397 ;
  assign n11399 = n11398 ^ n10640 ^ 1'b0 ;
  assign n11400 = ~n4867 & n9364 ;
  assign n11401 = n6617 & ~n11400 ;
  assign n11402 = n11399 & n11401 ;
  assign n11403 = n2944 ^ n462 ^ 1'b0 ;
  assign n11404 = n4407 ^ n3748 ^ 1'b0 ;
  assign n11405 = n9402 ^ n7726 ^ 1'b0 ;
  assign n11406 = n4649 & ~n11405 ;
  assign n11407 = ~n9742 & n11406 ;
  assign n11408 = n2163 | n3096 ;
  assign n11409 = n1371 | n11408 ;
  assign n11410 = n6731 ^ n6288 ^ n1702 ;
  assign n11411 = ~n11409 & n11410 ;
  assign n11412 = n11411 ^ n381 ^ 1'b0 ;
  assign n11413 = n2717 ^ n1397 ^ 1'b0 ;
  assign n11414 = ~n6038 & n11413 ;
  assign n11415 = ( n10753 & n11412 ) | ( n10753 & n11414 ) | ( n11412 & n11414 ) ;
  assign n11416 = n9501 ^ n4310 ^ 1'b0 ;
  assign n11417 = n3732 & n11416 ;
  assign n11418 = ~n5915 & n10780 ;
  assign n11419 = n11418 ^ n4552 ^ 1'b0 ;
  assign n11420 = x22 & ~n11419 ;
  assign n11421 = n11420 ^ n11261 ^ 1'b0 ;
  assign n11423 = n3418 & n6609 ;
  assign n11424 = n5798 & n11423 ;
  assign n11422 = n6524 ^ n3965 ^ 1'b0 ;
  assign n11425 = n11424 ^ n11422 ^ n2484 ;
  assign n11426 = n6936 & ~n9215 ;
  assign n11427 = n8894 ^ n3441 ^ n2200 ;
  assign n11428 = n365 & ~n10335 ;
  assign n11430 = n2174 | n4176 ;
  assign n11431 = n11430 ^ n9393 ^ 1'b0 ;
  assign n11432 = n154 | n11431 ;
  assign n11433 = n11432 ^ n2335 ^ n643 ;
  assign n11434 = ( ~n6921 & n6938 ) | ( ~n6921 & n11433 ) | ( n6938 & n11433 ) ;
  assign n11429 = n3875 & n6105 ;
  assign n11435 = n11434 ^ n11429 ^ 1'b0 ;
  assign n11436 = n11435 ^ n3634 ^ 1'b0 ;
  assign n11437 = n6177 | n11436 ;
  assign n11438 = n2831 | n11186 ;
  assign n11439 = n11438 ^ n3095 ^ 1'b0 ;
  assign n11440 = n2863 ^ n2849 ^ 1'b0 ;
  assign n11441 = n816 | n7448 ;
  assign n11442 = n11441 ^ n2773 ^ 1'b0 ;
  assign n11443 = ( ~n10376 & n11440 ) | ( ~n10376 & n11442 ) | ( n11440 & n11442 ) ;
  assign n11444 = n5741 | n8515 ;
  assign n11445 = ( n7655 & n11443 ) | ( n7655 & ~n11444 ) | ( n11443 & ~n11444 ) ;
  assign n11451 = n4594 & ~n5692 ;
  assign n11452 = n3299 & n11451 ;
  assign n11449 = ( x86 & n2995 ) | ( x86 & ~n3625 ) | ( n2995 & ~n3625 ) ;
  assign n11447 = ~n2831 & n3370 ;
  assign n11448 = n11447 ^ n2809 ^ 1'b0 ;
  assign n11450 = n11449 ^ n11448 ^ 1'b0 ;
  assign n11446 = n4742 ^ n3628 ^ n3042 ;
  assign n11453 = n11452 ^ n11450 ^ n11446 ;
  assign n11474 = n11310 ^ n1373 ^ 1'b0 ;
  assign n11475 = ~n3820 & n11474 ;
  assign n11457 = n4995 ^ n4328 ^ n846 ;
  assign n11454 = ( ~n922 & n1419 ) | ( ~n922 & n2347 ) | ( n1419 & n2347 ) ;
  assign n11455 = ~n465 & n2207 ;
  assign n11456 = ~n11454 & n11455 ;
  assign n11458 = n11457 ^ n11456 ^ 1'b0 ;
  assign n11459 = n2521 & n3002 ;
  assign n11460 = n882 & n2380 ;
  assign n11461 = n11460 ^ n6129 ^ 1'b0 ;
  assign n11462 = n2167 | n4430 ;
  assign n11463 = n11461 | n11462 ;
  assign n11466 = ~n5098 & n7169 ;
  assign n11467 = n11466 ^ x127 ^ 1'b0 ;
  assign n11464 = n3947 ^ n2715 ^ 1'b0 ;
  assign n11465 = n11464 ^ n713 ^ 1'b0 ;
  assign n11468 = n11467 ^ n11465 ^ n1806 ;
  assign n11469 = n7177 ^ n4966 ^ n2144 ;
  assign n11470 = n11468 & ~n11469 ;
  assign n11471 = ( n11459 & n11463 ) | ( n11459 & ~n11470 ) | ( n11463 & ~n11470 ) ;
  assign n11472 = ~n11458 & n11471 ;
  assign n11473 = n11472 ^ n10559 ^ 1'b0 ;
  assign n11476 = n11475 ^ n11473 ^ x126 ;
  assign n11477 = n5128 ^ n3591 ^ 1'b0 ;
  assign n11478 = ~n1345 & n11477 ;
  assign n11479 = n258 & n3032 ;
  assign n11480 = ~n11478 & n11479 ;
  assign n11481 = n8605 & ~n9173 ;
  assign n11482 = n5351 & n11481 ;
  assign n11483 = ( n7607 & n9431 ) | ( n7607 & ~n11482 ) | ( n9431 & ~n11482 ) ;
  assign n11484 = n2782 ^ n2086 ^ 1'b0 ;
  assign n11485 = ~n9925 & n11484 ;
  assign n11486 = n11485 ^ n10177 ^ n2072 ;
  assign n11487 = ( n443 & n2145 ) | ( n443 & ~n5756 ) | ( n2145 & ~n5756 ) ;
  assign n11488 = n2458 & ~n3174 ;
  assign n11489 = n11488 ^ n10887 ^ 1'b0 ;
  assign n11490 = n11489 ^ n10435 ^ 1'b0 ;
  assign n11491 = ~n6995 & n8101 ;
  assign n11492 = n7206 & n11491 ;
  assign n11493 = n8614 ^ n6230 ^ 1'b0 ;
  assign n11494 = n2578 & n4625 ;
  assign n11497 = n1305 & n2040 ;
  assign n11498 = ~n2924 & n11497 ;
  assign n11496 = n1311 & n4380 ;
  assign n11499 = n11498 ^ n11496 ^ n2507 ;
  assign n11500 = n11499 ^ n6824 ^ 1'b0 ;
  assign n11495 = n7719 & ~n8014 ;
  assign n11501 = n11500 ^ n11495 ^ 1'b0 ;
  assign n11502 = n11494 & n11501 ;
  assign n11503 = n5098 ^ n491 ^ 1'b0 ;
  assign n11504 = n7383 ^ n5278 ^ n3612 ;
  assign n11505 = n11504 ^ n7532 ^ 1'b0 ;
  assign n11506 = ~n2016 & n11505 ;
  assign n11507 = n1967 ^ n832 ^ 1'b0 ;
  assign n11508 = n11507 ^ n1306 ^ 1'b0 ;
  assign n11509 = n6744 ^ n6234 ^ 1'b0 ;
  assign n11510 = n11509 ^ n9429 ^ 1'b0 ;
  assign n11511 = n3856 & n11510 ;
  assign n11512 = n9329 ^ n1577 ^ x11 ;
  assign n11513 = ~n1513 & n7571 ;
  assign n11514 = n3832 & ~n10974 ;
  assign n11515 = n11514 ^ n4803 ^ n2242 ;
  assign n11516 = ~n2149 & n5257 ;
  assign n11517 = n11516 ^ n6427 ^ 1'b0 ;
  assign n11518 = n161 & ~n7900 ;
  assign n11519 = n9064 ^ n7837 ^ n5000 ;
  assign n11520 = n6835 | n10971 ;
  assign n11521 = n11520 ^ n3302 ^ 1'b0 ;
  assign n11522 = n11521 ^ n5244 ^ n1960 ;
  assign n11523 = n6112 ^ n528 ^ 1'b0 ;
  assign n11524 = n796 & ~n11523 ;
  assign n11525 = n2980 & n11524 ;
  assign n11526 = n9113 & ~n11525 ;
  assign n11527 = n9046 ^ n4048 ^ 1'b0 ;
  assign n11528 = n11527 ^ n5318 ^ 1'b0 ;
  assign n11529 = n7695 & ~n11528 ;
  assign n11532 = x106 | n1822 ;
  assign n11533 = n150 | n6959 ;
  assign n11534 = n11532 | n11533 ;
  assign n11530 = n673 ^ x31 ^ 1'b0 ;
  assign n11531 = ~n2409 & n11530 ;
  assign n11535 = n11534 ^ n11531 ^ n8942 ;
  assign n11539 = n8325 ^ n2099 ^ n847 ;
  assign n11537 = n3837 ^ n3758 ^ n2833 ;
  assign n11538 = ( n4819 & n7789 ) | ( n4819 & n11537 ) | ( n7789 & n11537 ) ;
  assign n11536 = ~n3129 & n10398 ;
  assign n11540 = n11539 ^ n11538 ^ n11536 ;
  assign n11541 = ( ~n714 & n4437 ) | ( ~n714 & n7778 ) | ( n4437 & n7778 ) ;
  assign n11542 = n11541 ^ n7473 ^ 1'b0 ;
  assign n11543 = n4102 & ~n10031 ;
  assign n11544 = n11542 & ~n11543 ;
  assign n11545 = n7667 ^ n773 ^ 1'b0 ;
  assign n11546 = n3371 & n5050 ;
  assign n11547 = n3012 & n11546 ;
  assign n11548 = ( n2235 & n7482 ) | ( n2235 & n11547 ) | ( n7482 & n11547 ) ;
  assign n11551 = n6935 ^ n4617 ^ n2452 ;
  assign n11550 = ~n3383 & n4062 ;
  assign n11549 = ~n2019 & n11465 ;
  assign n11552 = n11551 ^ n11550 ^ n11549 ;
  assign n11553 = ~n7021 & n7721 ;
  assign n11554 = n1625 | n8445 ;
  assign n11555 = ~n11553 & n11554 ;
  assign n11556 = n2221 & n2952 ;
  assign n11557 = n11556 ^ n7268 ^ 1'b0 ;
  assign n11558 = ~n6655 & n11557 ;
  assign n11559 = n1536 & n11558 ;
  assign n11560 = n4737 ^ n2262 ^ 1'b0 ;
  assign n11561 = n5845 & ~n11560 ;
  assign n11562 = ~n1042 & n11561 ;
  assign n11563 = n310 & ~n11562 ;
  assign n11564 = n11563 ^ n1918 ^ 1'b0 ;
  assign n11565 = n189 | n4323 ;
  assign n11566 = ( n243 & n4227 ) | ( n243 & ~n11565 ) | ( n4227 & ~n11565 ) ;
  assign n11567 = n11566 ^ n3611 ^ 1'b0 ;
  assign n11568 = n11564 & n11567 ;
  assign n11569 = ~n164 & n4927 ;
  assign n11570 = ~n7964 & n11569 ;
  assign n11571 = n6255 | n11570 ;
  assign n11572 = n5821 ^ n2964 ^ 1'b0 ;
  assign n11573 = ~n9021 & n11572 ;
  assign n11574 = n11573 ^ n2207 ^ 1'b0 ;
  assign n11575 = n6305 ^ n4436 ^ 1'b0 ;
  assign n11576 = n5723 & ~n11575 ;
  assign n11577 = ( ~n3943 & n10918 ) | ( ~n3943 & n11576 ) | ( n10918 & n11576 ) ;
  assign n11578 = n3726 ^ n1091 ^ n514 ;
  assign n11579 = ( ~n2469 & n4847 ) | ( ~n2469 & n9831 ) | ( n4847 & n9831 ) ;
  assign n11580 = n917 & ~n11579 ;
  assign n11581 = n4369 & n6962 ;
  assign n11582 = ~n3128 & n11581 ;
  assign n11583 = n1719 & ~n1828 ;
  assign n11584 = n7612 & n11583 ;
  assign n11585 = n4420 | n11584 ;
  assign n11586 = n5076 ^ n3894 ^ n1636 ;
  assign n11587 = n11586 ^ n7718 ^ n4364 ;
  assign n11588 = n8618 ^ n7189 ^ n5258 ;
  assign n11593 = ( n2145 & n5343 ) | ( n2145 & ~n8985 ) | ( n5343 & ~n8985 ) ;
  assign n11589 = n5114 & ~n7906 ;
  assign n11590 = n790 & ~n7527 ;
  assign n11591 = n11589 & n11590 ;
  assign n11592 = n4805 | n11591 ;
  assign n11594 = n11593 ^ n11592 ^ 1'b0 ;
  assign n11595 = n265 & n3234 ;
  assign n11596 = n9293 ^ n4342 ^ n1911 ;
  assign n11597 = ( n5667 & n11595 ) | ( n5667 & n11596 ) | ( n11595 & n11596 ) ;
  assign n11598 = ~n5479 & n7063 ;
  assign n11599 = ~n4090 & n11598 ;
  assign n11600 = n7920 ^ n718 ^ 1'b0 ;
  assign n11601 = n1438 & ~n11600 ;
  assign n11602 = n3048 | n11601 ;
  assign n11603 = n4405 | n7526 ;
  assign n11605 = ~n1631 & n3450 ;
  assign n11604 = n4797 & ~n5546 ;
  assign n11606 = n11605 ^ n11604 ^ n6376 ;
  assign n11607 = n5593 & ~n8857 ;
  assign n11608 = n2370 & n6720 ;
  assign n11609 = ~n4654 & n11608 ;
  assign n11610 = n10204 & ~n11609 ;
  assign n11611 = n2416 & ~n3971 ;
  assign n11612 = n2285 & n11611 ;
  assign n11613 = n7822 | n8748 ;
  assign n11614 = n7528 ^ n281 ^ 1'b0 ;
  assign n11615 = n10501 | n11614 ;
  assign n11616 = ( n727 & n5017 ) | ( n727 & ~n5338 ) | ( n5017 & ~n5338 ) ;
  assign n11617 = n2894 ^ n554 ^ 1'b0 ;
  assign n11618 = n658 & n11617 ;
  assign n11619 = ~n447 & n11618 ;
  assign n11620 = ( n9844 & n11616 ) | ( n9844 & n11619 ) | ( n11616 & n11619 ) ;
  assign n11621 = n3828 | n5502 ;
  assign n11622 = n6182 & ~n11621 ;
  assign n11623 = n6770 ^ n2954 ^ x55 ;
  assign n11624 = n7718 & ~n11623 ;
  assign n11625 = n11624 ^ n1850 ^ 1'b0 ;
  assign n11626 = n11625 ^ n4087 ^ 1'b0 ;
  assign n11627 = ~n4201 & n11626 ;
  assign n11628 = n5755 | n11627 ;
  assign n11630 = ( n257 & n2374 ) | ( n257 & ~n3257 ) | ( n2374 & ~n3257 ) ;
  assign n11629 = n2444 & n3022 ;
  assign n11631 = n11630 ^ n11629 ^ 1'b0 ;
  assign n11632 = ( n3908 & n5962 ) | ( n3908 & n11631 ) | ( n5962 & n11631 ) ;
  assign n11633 = ( n3408 & n6667 ) | ( n3408 & ~n8997 ) | ( n6667 & ~n8997 ) ;
  assign n11634 = n2408 & ~n4154 ;
  assign n11635 = ~x56 & n10095 ;
  assign n11636 = n6505 ^ n1083 ^ n1022 ;
  assign n11637 = n5586 & n6300 ;
  assign n11638 = n11637 ^ n3154 ^ 1'b0 ;
  assign n11639 = ~n2375 & n11638 ;
  assign n11640 = n7992 | n8066 ;
  assign n11641 = n9557 | n11640 ;
  assign n11642 = ( n1326 & n1895 ) | ( n1326 & ~n6607 ) | ( n1895 & ~n6607 ) ;
  assign n11643 = n1600 ^ x79 ^ 1'b0 ;
  assign n11644 = ~n9985 & n11643 ;
  assign n11646 = n3958 ^ n2253 ^ 1'b0 ;
  assign n11647 = n2105 | n11646 ;
  assign n11645 = n4549 & ~n8184 ;
  assign n11648 = n11647 ^ n11645 ^ 1'b0 ;
  assign n11649 = n3228 & ~n11648 ;
  assign n11650 = n594 & ~n4063 ;
  assign n11651 = n11650 ^ n1841 ^ 1'b0 ;
  assign n11652 = n5201 & ~n11651 ;
  assign n11653 = n6919 ^ n5723 ^ 1'b0 ;
  assign n11654 = ~n2084 & n11653 ;
  assign n11655 = ~n3751 & n11654 ;
  assign n11656 = n1382 | n8414 ;
  assign n11658 = n2708 | n4492 ;
  assign n11657 = n675 & ~n7667 ;
  assign n11659 = n11658 ^ n11657 ^ 1'b0 ;
  assign n11660 = n11659 ^ n8178 ^ 1'b0 ;
  assign n11661 = n9073 & ~n11660 ;
  assign n11662 = n11449 ^ n7053 ^ n2781 ;
  assign n11663 = n3514 ^ x89 ^ 1'b0 ;
  assign n11664 = n3345 | n11448 ;
  assign n11665 = n1725 | n11664 ;
  assign n11666 = ~n7858 & n11665 ;
  assign n11667 = n11352 ^ n6332 ^ 1'b0 ;
  assign n11668 = n11666 & n11667 ;
  assign n11669 = ~n9669 & n11668 ;
  assign n11670 = n10240 ^ n7141 ^ 1'b0 ;
  assign n11671 = x67 & ~n11670 ;
  assign n11672 = x14 & n11671 ;
  assign n11673 = n6394 & n11672 ;
  assign n11674 = n9630 | n11673 ;
  assign n11675 = n8142 & ~n11674 ;
  assign n11676 = ( n660 & n8658 ) | ( n660 & ~n11675 ) | ( n8658 & ~n11675 ) ;
  assign n11677 = ~n9496 & n11676 ;
  assign n11678 = n11677 ^ n1478 ^ 1'b0 ;
  assign n11679 = n1699 & ~n9236 ;
  assign n11680 = n11679 ^ n1715 ^ 1'b0 ;
  assign n11681 = n11678 & n11680 ;
  assign n11683 = n138 & n3431 ;
  assign n11684 = n11683 ^ n250 ^ 1'b0 ;
  assign n11682 = n7079 ^ n6496 ^ n480 ;
  assign n11685 = n11684 ^ n11682 ^ 1'b0 ;
  assign n11686 = n8018 | n11685 ;
  assign n11687 = n1990 | n4316 ;
  assign n11689 = n8241 ^ n5822 ^ 1'b0 ;
  assign n11688 = n6988 ^ n4931 ^ n2267 ;
  assign n11690 = n11689 ^ n11688 ^ 1'b0 ;
  assign n11693 = n1640 ^ n1167 ^ 1'b0 ;
  assign n11694 = n11693 ^ n5912 ^ n5046 ;
  assign n11691 = n2077 & ~n2923 ;
  assign n11692 = n11691 ^ n4558 ^ 1'b0 ;
  assign n11695 = n11694 ^ n11692 ^ n9564 ;
  assign n11696 = ~n1974 & n2940 ;
  assign n11697 = n11695 & n11696 ;
  assign n11698 = x41 & ~n1920 ;
  assign n11699 = n11698 ^ n10112 ^ 1'b0 ;
  assign n11700 = ~n10199 & n11699 ;
  assign n11701 = ~n10898 & n11700 ;
  assign n11702 = n3800 ^ n948 ^ 1'b0 ;
  assign n11703 = n1554 ^ n1420 ^ 1'b0 ;
  assign n11704 = n11703 ^ n11044 ^ 1'b0 ;
  assign n11706 = ~n2974 & n3130 ;
  assign n11707 = n3408 & n11706 ;
  assign n11708 = n2021 & ~n5088 ;
  assign n11709 = n11707 & n11708 ;
  assign n11705 = ~n2224 & n3022 ;
  assign n11710 = n11709 ^ n11705 ^ 1'b0 ;
  assign n11711 = ~n4480 & n11707 ;
  assign n11712 = n9465 & ~n9971 ;
  assign n11713 = ~n1093 & n2372 ;
  assign n11714 = n11713 ^ n8860 ^ 1'b0 ;
  assign n11715 = n1252 & ~n2905 ;
  assign n11716 = ( ~n325 & n1759 ) | ( ~n325 & n11715 ) | ( n1759 & n11715 ) ;
  assign n11719 = ( ~n2448 & n7274 ) | ( ~n2448 & n8017 ) | ( n7274 & n8017 ) ;
  assign n11717 = n3592 & n4901 ;
  assign n11718 = n2364 & n11717 ;
  assign n11720 = n11719 ^ n11718 ^ n11597 ;
  assign n11721 = n274 | n7173 ;
  assign n11722 = ~n8150 & n10313 ;
  assign n11723 = ~x120 & n11722 ;
  assign n11724 = n11721 | n11723 ;
  assign n11725 = n11724 ^ n3722 ^ 1'b0 ;
  assign n11726 = n2571 | n7206 ;
  assign n11727 = n553 | n11726 ;
  assign n11728 = n11727 ^ x124 ^ 1'b0 ;
  assign n11729 = n10769 & n11728 ;
  assign n11730 = n7827 ^ n5643 ^ 1'b0 ;
  assign n11731 = n7023 | n8476 ;
  assign n11733 = n10121 & ~n10540 ;
  assign n11732 = n719 | n6500 ;
  assign n11734 = n11733 ^ n11732 ^ 1'b0 ;
  assign n11735 = ( n11730 & n11731 ) | ( n11730 & n11734 ) | ( n11731 & n11734 ) ;
  assign n11736 = n5873 & n10162 ;
  assign n11737 = n4475 & n11736 ;
  assign n11738 = n11737 ^ n9192 ^ 1'b0 ;
  assign n11739 = x120 & n9755 ;
  assign n11741 = n5461 ^ n2353 ^ 1'b0 ;
  assign n11740 = n8630 ^ n7834 ^ n5130 ;
  assign n11742 = n11741 ^ n11740 ^ n2783 ;
  assign n11744 = n7766 ^ n1499 ^ 1'b0 ;
  assign n11743 = n5161 & ~n7656 ;
  assign n11745 = n11744 ^ n11743 ^ 1'b0 ;
  assign n11746 = n9096 & ~n11745 ;
  assign n11747 = ~n2017 & n9736 ;
  assign n11748 = n11747 ^ n3026 ^ 1'b0 ;
  assign n11749 = n11748 ^ n3758 ^ 1'b0 ;
  assign n11750 = n1528 | n1741 ;
  assign n11751 = n11750 ^ n712 ^ 1'b0 ;
  assign n11752 = n5973 & n11751 ;
  assign n11753 = n384 & n10821 ;
  assign n11754 = ~n1327 & n7200 ;
  assign n11755 = n11754 ^ n704 ^ 1'b0 ;
  assign n11756 = n6150 & n11755 ;
  assign n11757 = n11756 ^ n4772 ^ 1'b0 ;
  assign n11758 = n10136 ^ n5632 ^ 1'b0 ;
  assign n11759 = n542 | n5234 ;
  assign n11760 = n11759 ^ n4170 ^ 1'b0 ;
  assign n11761 = n11760 ^ n1831 ^ 1'b0 ;
  assign n11762 = n11758 | n11761 ;
  assign n11764 = n11027 ^ n5338 ^ n256 ;
  assign n11763 = n1818 & ~n5725 ;
  assign n11765 = n11764 ^ n11763 ^ 1'b0 ;
  assign n11766 = n967 | n11765 ;
  assign n11767 = ( n4399 & n9075 ) | ( n4399 & n11766 ) | ( n9075 & n11766 ) ;
  assign n11768 = x6 & n5850 ;
  assign n11769 = n3048 & n11768 ;
  assign n11770 = n11769 ^ n6072 ^ n3665 ;
  assign n11771 = n11770 ^ n3954 ^ 1'b0 ;
  assign n11772 = n8160 ^ n2344 ^ n888 ;
  assign n11773 = ( ~n918 & n1173 ) | ( ~n918 & n11772 ) | ( n1173 & n11772 ) ;
  assign n11774 = n6726 ^ n4590 ^ 1'b0 ;
  assign n11775 = n3016 & ~n11774 ;
  assign n11776 = n5630 | n9105 ;
  assign n11777 = n11776 ^ n11548 ^ 1'b0 ;
  assign n11778 = n1201 & ~n6361 ;
  assign n11779 = n11778 ^ n9806 ^ 1'b0 ;
  assign n11780 = ~n7992 & n11779 ;
  assign n11781 = n9343 & n11780 ;
  assign n11782 = n3615 ^ n1201 ^ 1'b0 ;
  assign n11783 = n11782 ^ n11301 ^ 1'b0 ;
  assign n11784 = n10886 & n11783 ;
  assign n11785 = n3925 ^ n3650 ^ 1'b0 ;
  assign n11786 = n8785 ^ n3871 ^ n1546 ;
  assign n11787 = n1092 | n4321 ;
  assign n11788 = n11787 ^ n10745 ^ n6886 ;
  assign n11789 = n11786 & n11788 ;
  assign n11790 = n1348 | n7079 ;
  assign n11791 = n11789 | n11790 ;
  assign n11799 = n2829 ^ x111 ^ 1'b0 ;
  assign n11800 = n1400 & n11799 ;
  assign n11792 = n11514 ^ n4135 ^ 1'b0 ;
  assign n11793 = n920 & n11792 ;
  assign n11795 = x67 & ~n6290 ;
  assign n11796 = n11795 ^ n6196 ^ 1'b0 ;
  assign n11794 = n5868 & n9096 ;
  assign n11797 = n11796 ^ n11794 ^ 1'b0 ;
  assign n11798 = n11793 & ~n11797 ;
  assign n11801 = n11800 ^ n11798 ^ 1'b0 ;
  assign n11802 = n5112 | n6930 ;
  assign n11803 = n7270 & ~n11802 ;
  assign n11804 = n3482 | n6387 ;
  assign n11805 = ~n2353 & n5393 ;
  assign n11806 = n11805 ^ n9709 ^ 1'b0 ;
  assign n11807 = n249 & n7951 ;
  assign n11808 = n4633 & n7227 ;
  assign n11809 = ~n7113 & n8466 ;
  assign n11810 = n1950 & n11809 ;
  assign n11811 = ( n8702 & n11808 ) | ( n8702 & n11810 ) | ( n11808 & n11810 ) ;
  assign n11812 = ~n2176 & n2836 ;
  assign n11813 = n2404 & ~n7960 ;
  assign n11814 = n11384 ^ n5495 ^ 1'b0 ;
  assign n11815 = ( n3938 & ~n5705 ) | ( n3938 & n7369 ) | ( ~n5705 & n7369 ) ;
  assign n11816 = ~n8692 & n11815 ;
  assign n11817 = n11816 ^ n1381 ^ 1'b0 ;
  assign n11818 = n443 & n3001 ;
  assign n11819 = ~n5378 & n11818 ;
  assign n11820 = ( n1352 & ~n4753 ) | ( n1352 & n11819 ) | ( ~n4753 & n11819 ) ;
  assign n11821 = ( ~n1567 & n1809 ) | ( ~n1567 & n2456 ) | ( n1809 & n2456 ) ;
  assign n11822 = n7113 ^ n3898 ^ 1'b0 ;
  assign n11823 = n11822 ^ n9462 ^ n4465 ;
  assign n11824 = ( n744 & n11821 ) | ( n744 & n11823 ) | ( n11821 & n11823 ) ;
  assign n11826 = n4929 ^ n2041 ^ 1'b0 ;
  assign n11825 = n4124 | n4468 ;
  assign n11827 = n11826 ^ n11825 ^ 1'b0 ;
  assign n11828 = ( ~n601 & n4146 ) | ( ~n601 & n7147 ) | ( n4146 & n7147 ) ;
  assign n11829 = n9488 ^ n2055 ^ 1'b0 ;
  assign n11830 = n770 & n5322 ;
  assign n11831 = ~n1466 & n11830 ;
  assign n11833 = n4242 ^ n2047 ^ 1'b0 ;
  assign n11832 = ( n5104 & n7482 ) | ( n5104 & n9452 ) | ( n7482 & n9452 ) ;
  assign n11834 = n11833 ^ n11832 ^ n4794 ;
  assign n11835 = ( n3330 & n8023 ) | ( n3330 & ~n11030 ) | ( n8023 & ~n11030 ) ;
  assign n11836 = n5190 & n11037 ;
  assign n11837 = n7270 & ~n11836 ;
  assign n11838 = n11837 ^ n8159 ^ 1'b0 ;
  assign n11839 = n5883 ^ n2158 ^ 1'b0 ;
  assign n11840 = n1751 & n8345 ;
  assign n11841 = n11840 ^ n4695 ^ 1'b0 ;
  assign n11842 = x72 & n11841 ;
  assign n11843 = n11842 ^ n3991 ^ n1091 ;
  assign n11844 = n8084 & ~n11843 ;
  assign n11845 = n1712 ^ n1316 ^ 1'b0 ;
  assign n11846 = ( n6200 & n10006 ) | ( n6200 & n11845 ) | ( n10006 & n11845 ) ;
  assign n11847 = n7379 | n8334 ;
  assign n11852 = ~n4527 & n10299 ;
  assign n11853 = n11852 ^ n723 ^ 1'b0 ;
  assign n11854 = n11853 ^ n4265 ^ n1662 ;
  assign n11848 = x105 | n2066 ;
  assign n11849 = n1834 & ~n11848 ;
  assign n11850 = n11849 ^ n3277 ^ n606 ;
  assign n11851 = ( n169 & ~n8701 ) | ( n169 & n11850 ) | ( ~n8701 & n11850 ) ;
  assign n11855 = n11854 ^ n11851 ^ n4996 ;
  assign n11856 = ( ~n820 & n1199 ) | ( ~n820 & n2845 ) | ( n1199 & n2845 ) ;
  assign n11857 = ~n298 & n7369 ;
  assign n11858 = n1980 | n7204 ;
  assign n11859 = n11857 & ~n11858 ;
  assign n11860 = ( n5431 & n10762 ) | ( n5431 & n11859 ) | ( n10762 & n11859 ) ;
  assign n11861 = n11860 ^ n211 ^ 1'b0 ;
  assign n11862 = ~n11856 & n11861 ;
  assign n11863 = n240 | n11862 ;
  assign n11864 = ( n4039 & ~n8657 ) | ( n4039 & n10822 ) | ( ~n8657 & n10822 ) ;
  assign n11865 = n11864 ^ n6252 ^ 1'b0 ;
  assign n11866 = n3512 & ~n4533 ;
  assign n11867 = n7614 ^ n6998 ^ n4152 ;
  assign n11868 = n4610 ^ n3242 ^ 1'b0 ;
  assign n11869 = ~n3667 & n4035 ;
  assign n11870 = n5861 & n11869 ;
  assign n11871 = n11870 ^ n5810 ^ 1'b0 ;
  assign n11872 = n6335 & n11871 ;
  assign n11873 = n2698 | n11872 ;
  assign n11874 = n10544 | n11873 ;
  assign n11875 = x97 | n6289 ;
  assign n11876 = ( ~n5572 & n6625 ) | ( ~n5572 & n11875 ) | ( n6625 & n11875 ) ;
  assign n11877 = n11858 ^ x49 ^ 1'b0 ;
  assign n11878 = ~n2470 & n11877 ;
  assign n11882 = ~n987 & n6209 ;
  assign n11883 = n9004 & n11882 ;
  assign n11884 = n4669 & n11883 ;
  assign n11879 = ~x84 & n6718 ;
  assign n11880 = n5367 ^ n877 ^ 1'b0 ;
  assign n11881 = n11879 | n11880 ;
  assign n11885 = n11884 ^ n11881 ^ n5460 ;
  assign n11886 = n3967 & n5236 ;
  assign n11887 = n5013 ^ n4431 ^ 1'b0 ;
  assign n11888 = n11887 ^ n10492 ^ 1'b0 ;
  assign n11889 = n3863 & n11888 ;
  assign n11890 = x90 & n3563 ;
  assign n11891 = n3537 & n11890 ;
  assign n11892 = x89 & ~n366 ;
  assign n11893 = n11892 ^ n5161 ^ n3349 ;
  assign n11896 = n6497 ^ n6283 ^ 1'b0 ;
  assign n11897 = n6915 | n11896 ;
  assign n11898 = n3980 | n10822 ;
  assign n11899 = n11898 ^ n8786 ^ 1'b0 ;
  assign n11900 = n11897 | n11899 ;
  assign n11894 = n1202 & ~n2104 ;
  assign n11895 = n3777 & n11894 ;
  assign n11901 = n11900 ^ n11895 ^ 1'b0 ;
  assign n11905 = ~n3048 & n4743 ;
  assign n11906 = n11905 ^ n7602 ^ 1'b0 ;
  assign n11902 = n7324 ^ n2014 ^ 1'b0 ;
  assign n11903 = ~n1946 & n11902 ;
  assign n11904 = n7372 & n11903 ;
  assign n11907 = n11906 ^ n11904 ^ 1'b0 ;
  assign n11908 = n8231 ^ n2640 ^ 1'b0 ;
  assign n11909 = n11908 ^ n4461 ^ 1'b0 ;
  assign n11910 = n11909 ^ n4572 ^ n644 ;
  assign n11911 = n2038 ^ n1743 ^ 1'b0 ;
  assign n11912 = n9112 & ~n11911 ;
  assign n11913 = ~n11910 & n11912 ;
  assign n11914 = n6767 & ~n9665 ;
  assign n11915 = n11914 ^ n2100 ^ 1'b0 ;
  assign n11916 = n11915 ^ n5454 ^ n4712 ;
  assign n11917 = n10553 ^ n9996 ^ n4332 ;
  assign n11918 = n3598 | n6409 ;
  assign n11919 = n11918 ^ n4396 ^ 1'b0 ;
  assign n11920 = n1996 & ~n4533 ;
  assign n11921 = n3775 ^ n2125 ^ 1'b0 ;
  assign n11922 = n11920 & ~n11921 ;
  assign n11923 = ( n2106 & n2341 ) | ( n2106 & n4375 ) | ( n2341 & n4375 ) ;
  assign n11924 = n2841 ^ n2032 ^ 1'b0 ;
  assign n11925 = n11923 | n11924 ;
  assign n11926 = n4562 ^ n1990 ^ 1'b0 ;
  assign n11927 = ~n11925 & n11926 ;
  assign n11928 = n11927 ^ n10276 ^ n8904 ;
  assign n11931 = n5801 ^ n721 ^ 1'b0 ;
  assign n11932 = ( ~n1662 & n11631 ) | ( ~n1662 & n11931 ) | ( n11631 & n11931 ) ;
  assign n11929 = ( n210 & n2448 ) | ( n210 & n6885 ) | ( n2448 & n6885 ) ;
  assign n11930 = ~n5686 & n11929 ;
  assign n11933 = n11932 ^ n11930 ^ 1'b0 ;
  assign n11935 = ( x104 & n1459 ) | ( x104 & n1881 ) | ( n1459 & n1881 ) ;
  assign n11936 = n7033 | n11935 ;
  assign n11934 = n4160 ^ n3300 ^ n509 ;
  assign n11937 = n11936 ^ n11934 ^ 1'b0 ;
  assign n11938 = n11937 ^ n10011 ^ 1'b0 ;
  assign n11939 = ~n6835 & n11938 ;
  assign n11940 = ( n471 & n735 ) | ( n471 & n4434 ) | ( n735 & n4434 ) ;
  assign n11941 = n9533 ^ n3466 ^ 1'b0 ;
  assign n11942 = n3035 & ~n11941 ;
  assign n11943 = n11942 ^ n6271 ^ 1'b0 ;
  assign n11944 = n2633 & n11943 ;
  assign n11945 = n11944 ^ n2868 ^ 1'b0 ;
  assign n11946 = n7520 ^ n5855 ^ x1 ;
  assign n11947 = n2559 | n9296 ;
  assign n11948 = ( n1723 & ~n11946 ) | ( n1723 & n11947 ) | ( ~n11946 & n11947 ) ;
  assign n11949 = ~n11945 & n11948 ;
  assign n11951 = n11176 ^ n9524 ^ n8430 ;
  assign n11950 = n11719 ^ n6273 ^ 1'b0 ;
  assign n11952 = n11951 ^ n11950 ^ n7006 ;
  assign n11953 = x89 & n4265 ;
  assign n11954 = n11953 ^ n5168 ^ 1'b0 ;
  assign n11955 = n11954 ^ n6444 ^ n710 ;
  assign n11956 = n1053 | n1414 ;
  assign n11957 = n11956 ^ n9480 ^ 1'b0 ;
  assign n11958 = ( n2598 & n4245 ) | ( n2598 & n5477 ) | ( n4245 & n5477 ) ;
  assign n11959 = n11958 ^ n3674 ^ 1'b0 ;
  assign n11960 = n1485 | n11959 ;
  assign n11961 = n4906 | n6317 ;
  assign n11962 = n11960 & ~n11961 ;
  assign n11963 = n7774 & n11962 ;
  assign n11964 = n3187 ^ n761 ^ 1'b0 ;
  assign n11965 = ( n5113 & n5413 ) | ( n5113 & n7735 ) | ( n5413 & n7735 ) ;
  assign n11966 = n11965 ^ n6509 ^ 1'b0 ;
  assign n11967 = n3282 & ~n3784 ;
  assign n11968 = ~n3113 & n11967 ;
  assign n11969 = ~n11392 & n11968 ;
  assign n11970 = n2723 ^ n1702 ^ 1'b0 ;
  assign n11971 = n170 & ~n11970 ;
  assign n11972 = n11971 ^ n7276 ^ n3760 ;
  assign n11975 = n4641 ^ n1808 ^ 1'b0 ;
  assign n11973 = n7685 ^ n3837 ^ 1'b0 ;
  assign n11974 = n6849 | n11973 ;
  assign n11976 = n11975 ^ n11974 ^ x77 ;
  assign n11977 = ( n1284 & ~n1316 ) | ( n1284 & n3164 ) | ( ~n1316 & n3164 ) ;
  assign n11981 = n7869 ^ x86 ^ 1'b0 ;
  assign n11978 = n7342 | n8483 ;
  assign n11979 = n11978 ^ n254 ^ 1'b0 ;
  assign n11980 = n4231 & n11979 ;
  assign n11982 = n11981 ^ n11980 ^ 1'b0 ;
  assign n11983 = n3159 ^ n425 ^ 1'b0 ;
  assign n11984 = n1170 | n11983 ;
  assign n11985 = n2163 & ~n11984 ;
  assign n11986 = n10597 ^ n8979 ^ 1'b0 ;
  assign n11987 = ~n203 & n11986 ;
  assign n11988 = n3366 ^ n489 ^ 1'b0 ;
  assign n11989 = n143 & ~n7778 ;
  assign n11990 = n4249 | n9133 ;
  assign n11991 = ( n11854 & n11989 ) | ( n11854 & ~n11990 ) | ( n11989 & ~n11990 ) ;
  assign n11992 = n1458 & n4983 ;
  assign n11993 = n9609 ^ n6989 ^ n1392 ;
  assign n11995 = n6660 | n8752 ;
  assign n11996 = n3407 & ~n11995 ;
  assign n11994 = x19 & n3160 ;
  assign n11997 = n11996 ^ n11994 ^ 1'b0 ;
  assign n11998 = n5289 ^ n1138 ^ 1'b0 ;
  assign n11999 = n11998 ^ n5738 ^ 1'b0 ;
  assign n12001 = n816 & ~n11539 ;
  assign n12000 = ~n6596 & n10026 ;
  assign n12002 = n12001 ^ n12000 ^ 1'b0 ;
  assign n12003 = n10088 ^ n2741 ^ 1'b0 ;
  assign n12004 = ~n11038 & n12003 ;
  assign n12005 = n12004 ^ n5673 ^ 1'b0 ;
  assign n12006 = n9477 ^ n6433 ^ 1'b0 ;
  assign n12007 = n3713 ^ n1029 ^ 1'b0 ;
  assign n12008 = n12006 & ~n12007 ;
  assign n12009 = ( n3171 & ~n6335 ) | ( n3171 & n9630 ) | ( ~n6335 & n9630 ) ;
  assign n12010 = ( n526 & ~n7532 ) | ( n526 & n12009 ) | ( ~n7532 & n12009 ) ;
  assign n12011 = n4267 ^ n1093 ^ 1'b0 ;
  assign n12012 = ~n4738 & n12011 ;
  assign n12013 = n11446 | n12012 ;
  assign n12014 = ~n5771 & n6967 ;
  assign n12015 = n3701 | n4541 ;
  assign n12016 = n8345 | n12015 ;
  assign n12017 = n12016 ^ n8016 ^ 1'b0 ;
  assign n12018 = n1898 | n12017 ;
  assign n12019 = n6718 & ~n12018 ;
  assign n12020 = n12019 ^ n10152 ^ 1'b0 ;
  assign n12021 = n2724 | n12020 ;
  assign n12022 = ( ~n2196 & n3001 ) | ( ~n2196 & n3657 ) | ( n3001 & n3657 ) ;
  assign n12023 = n5467 ^ n3951 ^ 1'b0 ;
  assign n12024 = ~n7540 & n12023 ;
  assign n12025 = ~n5127 & n12024 ;
  assign n12026 = n950 | n4221 ;
  assign n12027 = n2435 | n12026 ;
  assign n12028 = n11024 & n12027 ;
  assign n12029 = ~n2944 & n12028 ;
  assign n12030 = n3986 | n4458 ;
  assign n12031 = n9569 & ~n12030 ;
  assign n12032 = n12031 ^ n10867 ^ 1'b0 ;
  assign n12033 = n7104 & n12032 ;
  assign n12034 = n377 & n2952 ;
  assign n12035 = ~x24 & n12034 ;
  assign n12036 = n12033 | n12035 ;
  assign n12037 = n10022 ^ n2934 ^ 1'b0 ;
  assign n12038 = n8949 & n12037 ;
  assign n12039 = n1694 & ~n5044 ;
  assign n12040 = n12039 ^ n8777 ^ n1175 ;
  assign n12041 = n4043 & n11515 ;
  assign n12042 = x70 & n4154 ;
  assign n12043 = n12042 ^ n5349 ^ 1'b0 ;
  assign n12044 = n12043 ^ n8192 ^ 1'b0 ;
  assign n12045 = n11095 ^ n2308 ^ 1'b0 ;
  assign n12046 = n10534 & ~n12045 ;
  assign n12047 = ~n6193 & n12046 ;
  assign n12048 = n12047 ^ n4708 ^ 1'b0 ;
  assign n12049 = n3383 ^ n685 ^ 1'b0 ;
  assign n12050 = ~n868 & n12049 ;
  assign n12051 = n3953 & n12050 ;
  assign n12052 = n4571 & n12051 ;
  assign n12053 = n12052 ^ n10436 ^ n8138 ;
  assign n12055 = n2141 ^ x8 ^ 1'b0 ;
  assign n12054 = n448 & n3316 ;
  assign n12056 = n12055 ^ n12054 ^ n1124 ;
  assign n12057 = n4132 | n12056 ;
  assign n12059 = n1136 & n4841 ;
  assign n12058 = n3844 | n5884 ;
  assign n12060 = n12059 ^ n12058 ^ 1'b0 ;
  assign n12061 = n3168 | n12060 ;
  assign n12062 = n3088 & ~n3209 ;
  assign n12063 = ~n4163 & n12062 ;
  assign n12064 = n6178 & n12063 ;
  assign n12065 = n6503 & ~n8903 ;
  assign n12066 = ( n3330 & n5088 ) | ( n3330 & n10920 ) | ( n5088 & n10920 ) ;
  assign n12067 = ~n9640 & n11802 ;
  assign n12068 = ~n2738 & n12067 ;
  assign n12069 = n12068 ^ n10503 ^ n10022 ;
  assign n12070 = n4181 ^ n1554 ^ 1'b0 ;
  assign n12071 = n7512 & n12070 ;
  assign n12072 = n12071 ^ n7682 ^ n3630 ;
  assign n12073 = n7260 ^ n1435 ^ 1'b0 ;
  assign n12074 = n1181 & n6522 ;
  assign n12075 = n247 & n12074 ;
  assign n12076 = ~n2086 & n11030 ;
  assign n12077 = n12076 ^ n3862 ^ 1'b0 ;
  assign n12078 = ( n1978 & n4180 ) | ( n1978 & n8737 ) | ( n4180 & n8737 ) ;
  assign n12080 = n2077 & ~n5284 ;
  assign n12081 = n3143 & n12080 ;
  assign n12079 = ~n1150 & n6784 ;
  assign n12082 = n12081 ^ n12079 ^ 1'b0 ;
  assign n12083 = n1284 | n1783 ;
  assign n12084 = n1283 | n3765 ;
  assign n12085 = n12083 | n12084 ;
  assign n12086 = n3391 & ~n12085 ;
  assign n12087 = n12086 ^ n6440 ^ 1'b0 ;
  assign n12088 = n2156 & n6668 ;
  assign n12089 = n12088 ^ n10168 ^ 1'b0 ;
  assign n12090 = ( n4605 & n5631 ) | ( n4605 & ~n12089 ) | ( n5631 & ~n12089 ) ;
  assign n12091 = n8429 ^ n4510 ^ 1'b0 ;
  assign n12094 = n2969 | n7834 ;
  assign n12095 = n6394 & ~n12094 ;
  assign n12093 = ~n298 & n10282 ;
  assign n12096 = n12095 ^ n12093 ^ 1'b0 ;
  assign n12097 = ~n1299 & n12096 ;
  assign n12098 = ~n5951 & n12097 ;
  assign n12092 = n9868 ^ n5747 ^ n4631 ;
  assign n12099 = n12098 ^ n12092 ^ 1'b0 ;
  assign n12100 = ( n2829 & n5669 ) | ( n2829 & ~n12099 ) | ( n5669 & ~n12099 ) ;
  assign n12101 = n7258 ^ n5399 ^ n2716 ;
  assign n12102 = n12101 ^ n9482 ^ 1'b0 ;
  assign n12103 = n5374 ^ n872 ^ 1'b0 ;
  assign n12104 = n12103 ^ n11434 ^ n7011 ;
  assign n12105 = n12104 ^ n2896 ^ 1'b0 ;
  assign n12106 = n3459 & n7328 ;
  assign n12108 = n8209 ^ n4388 ^ 1'b0 ;
  assign n12109 = n3614 & ~n12108 ;
  assign n12110 = n7339 ^ n2868 ^ 1'b0 ;
  assign n12111 = n12110 ^ n1837 ^ 1'b0 ;
  assign n12112 = n12109 & ~n12111 ;
  assign n12107 = x46 & ~n3779 ;
  assign n12113 = n12112 ^ n12107 ^ 1'b0 ;
  assign n12114 = n5058 | n8375 ;
  assign n12115 = n2252 & n5021 ;
  assign n12116 = ( n5032 & ~n9526 ) | ( n5032 & n12115 ) | ( ~n9526 & n12115 ) ;
  assign n12117 = n9273 ^ n2270 ^ 1'b0 ;
  assign n12118 = n447 & ~n12117 ;
  assign n12119 = x107 & n1947 ;
  assign n12120 = n906 & n12119 ;
  assign n12121 = n3721 & ~n11207 ;
  assign n12122 = n12120 & n12121 ;
  assign n12123 = n11804 | n12122 ;
  assign n12124 = n12118 | n12123 ;
  assign n12125 = ~n1447 & n2083 ;
  assign n12126 = ~n203 & n8492 ;
  assign n12127 = n12126 ^ n1055 ^ 1'b0 ;
  assign n12128 = n2014 & n7817 ;
  assign n12129 = ( n5291 & ~n12127 ) | ( n5291 & n12128 ) | ( ~n12127 & n12128 ) ;
  assign n12130 = n7284 & ~n9911 ;
  assign n12131 = ~x38 & n12130 ;
  assign n12132 = ( n5376 & n10061 ) | ( n5376 & ~n12131 ) | ( n10061 & ~n12131 ) ;
  assign n12133 = n211 & ~n9477 ;
  assign n12134 = ~n11881 & n12133 ;
  assign n12135 = n10985 & n11470 ;
  assign n12136 = ~n7675 & n8686 ;
  assign n12137 = ~n11233 & n12136 ;
  assign n12138 = n6507 | n12137 ;
  assign n12139 = n898 | n10115 ;
  assign n12140 = n10665 | n12139 ;
  assign n12141 = n5596 | n8892 ;
  assign n12142 = n2868 ^ n1215 ^ 1'b0 ;
  assign n12143 = n8687 & ~n12142 ;
  assign n12144 = ( ~n2197 & n5349 ) | ( ~n2197 & n12143 ) | ( n5349 & n12143 ) ;
  assign n12145 = n12144 ^ n7753 ^ 1'b0 ;
  assign n12146 = ~n3560 & n12145 ;
  assign n12147 = ( n1014 & ~n2265 ) | ( n1014 & n11824 ) | ( ~n2265 & n11824 ) ;
  assign n12148 = ~n3114 & n4369 ;
  assign n12149 = n9744 & n12148 ;
  assign n12150 = n11460 ^ n3352 ^ n853 ;
  assign n12151 = n8181 ^ n5811 ^ n3823 ;
  assign n12152 = n12151 ^ n7409 ^ 1'b0 ;
  assign n12153 = n6731 ^ n3748 ^ 1'b0 ;
  assign n12154 = ( n5130 & ~n9467 ) | ( n5130 & n12153 ) | ( ~n9467 & n12153 ) ;
  assign n12155 = n4164 & ~n12154 ;
  assign n12161 = n6121 & n10775 ;
  assign n12156 = n3698 & ~n12131 ;
  assign n12157 = n12156 ^ n4737 ^ 1'b0 ;
  assign n12158 = n12157 ^ n11911 ^ n7997 ;
  assign n12159 = n10284 ^ n9601 ^ 1'b0 ;
  assign n12160 = n12158 & ~n12159 ;
  assign n12162 = n12161 ^ n12160 ^ n4462 ;
  assign n12163 = n6812 & n7393 ;
  assign n12164 = ( n992 & n2997 ) | ( n992 & n12163 ) | ( n2997 & n12163 ) ;
  assign n12165 = n686 & n6003 ;
  assign n12166 = n11467 ^ n1046 ^ 1'b0 ;
  assign n12167 = n6439 & n12166 ;
  assign n12168 = n3772 | n3854 ;
  assign n12169 = n12168 ^ n1475 ^ n543 ;
  assign n12170 = n10264 ^ n7308 ^ 1'b0 ;
  assign n12171 = ~n8450 & n12170 ;
  assign n12172 = ( ~n10579 & n12169 ) | ( ~n10579 & n12171 ) | ( n12169 & n12171 ) ;
  assign n12173 = ( ~n2516 & n4593 ) | ( ~n2516 & n10284 ) | ( n4593 & n10284 ) ;
  assign n12174 = n12173 ^ n11293 ^ 1'b0 ;
  assign n12175 = n12174 ^ n3395 ^ 1'b0 ;
  assign n12176 = n4762 & n12175 ;
  assign n12177 = ~n421 & n10780 ;
  assign n12178 = ~n6040 & n12177 ;
  assign n12179 = ~n6132 & n8599 ;
  assign n12180 = ~n1272 & n12179 ;
  assign n12181 = n7766 & n9780 ;
  assign n12182 = n482 | n6462 ;
  assign n12183 = n12182 ^ n8982 ^ 1'b0 ;
  assign n12184 = n1700 ^ n740 ^ 1'b0 ;
  assign n12185 = ~n298 & n12184 ;
  assign n12186 = n4208 & ~n12185 ;
  assign n12193 = n4875 ^ n1507 ^ 1'b0 ;
  assign n12194 = n8730 ^ n5768 ^ 1'b0 ;
  assign n12195 = n12193 & ~n12194 ;
  assign n12191 = n10768 ^ n3023 ^ 1'b0 ;
  assign n12187 = n1378 & ~n3765 ;
  assign n12188 = ( n4382 & n5374 ) | ( n4382 & n12187 ) | ( n5374 & n12187 ) ;
  assign n12189 = ~n1264 & n12188 ;
  assign n12190 = n12189 ^ n8874 ^ 1'b0 ;
  assign n12192 = n12191 ^ n12190 ^ 1'b0 ;
  assign n12196 = n12195 ^ n12192 ^ n1331 ;
  assign n12197 = n597 ^ n173 ^ 1'b0 ;
  assign n12198 = n12040 ^ n4548 ^ 1'b0 ;
  assign n12199 = n6914 ^ n3946 ^ n1461 ;
  assign n12200 = n12199 ^ n5698 ^ 1'b0 ;
  assign n12201 = n566 | n12200 ;
  assign n12202 = ~n8031 & n10211 ;
  assign n12203 = n12131 & n12202 ;
  assign n12204 = ( ~n182 & n7789 ) | ( ~n182 & n12203 ) | ( n7789 & n12203 ) ;
  assign n12205 = n10807 ^ n7963 ^ 1'b0 ;
  assign n12206 = n8486 & ~n10769 ;
  assign n12207 = n4885 ^ n4150 ^ n1921 ;
  assign n12208 = ( x84 & n157 ) | ( x84 & n8130 ) | ( n157 & n8130 ) ;
  assign n12209 = n1078 & n1738 ;
  assign n12210 = n10461 & n12209 ;
  assign n12211 = ~n12208 & n12210 ;
  assign n12212 = n5189 ^ x51 ^ 1'b0 ;
  assign n12213 = n4695 & n12212 ;
  assign n12214 = n12213 ^ n6568 ^ 1'b0 ;
  assign n12215 = n4806 & n12214 ;
  assign n12216 = n2326 & ~n4951 ;
  assign n12217 = ~n1759 & n12216 ;
  assign n12218 = n12217 ^ n3023 ^ 1'b0 ;
  assign n12219 = ~n5423 & n12218 ;
  assign n12220 = n12219 ^ n9896 ^ 1'b0 ;
  assign n12221 = n12215 & ~n12220 ;
  assign n12222 = n7978 ^ n7852 ^ 1'b0 ;
  assign n12223 = ~n8735 & n12222 ;
  assign n12224 = n6665 | n9190 ;
  assign n12225 = n12223 | n12224 ;
  assign n12226 = n6261 | n10326 ;
  assign n12227 = n12226 ^ n6053 ^ 1'b0 ;
  assign n12228 = n12227 ^ n8504 ^ n773 ;
  assign n12229 = n3438 | n12228 ;
  assign n12230 = n3123 & ~n12229 ;
  assign n12231 = n7593 & ~n8777 ;
  assign n12233 = n286 & ~n1851 ;
  assign n12234 = n12233 ^ n1014 ^ 1'b0 ;
  assign n12235 = n5238 | n12234 ;
  assign n12232 = x111 & ~n6129 ;
  assign n12236 = n12235 ^ n12232 ^ 1'b0 ;
  assign n12237 = n1487 | n2837 ;
  assign n12238 = n6260 & ~n12237 ;
  assign n12239 = n440 & ~n11297 ;
  assign n12240 = n8125 ^ n4480 ^ 1'b0 ;
  assign n12241 = ~n6326 & n12240 ;
  assign n12242 = n12241 ^ n7462 ^ 1'b0 ;
  assign n12243 = ( ~n3426 & n5260 ) | ( ~n3426 & n12242 ) | ( n5260 & n12242 ) ;
  assign n12244 = n1686 & n12243 ;
  assign n12245 = ~n6395 & n12244 ;
  assign n12246 = ~n6752 & n12245 ;
  assign n12250 = n9412 ^ n6444 ^ 1'b0 ;
  assign n12247 = ~n210 & n5584 ;
  assign n12248 = n1887 & n12247 ;
  assign n12249 = n3397 & ~n12248 ;
  assign n12251 = n12250 ^ n12249 ^ 1'b0 ;
  assign n12252 = n3796 & n12251 ;
  assign n12253 = n11709 & n12252 ;
  assign n12254 = n4417 ^ n1203 ^ 1'b0 ;
  assign n12255 = ~n2139 & n2809 ;
  assign n12256 = n2186 & n12255 ;
  assign n12257 = n9837 ^ n6240 ^ 1'b0 ;
  assign n12258 = n3697 & ~n10446 ;
  assign n12259 = ~n940 & n12258 ;
  assign n12260 = n10888 ^ n4851 ^ n4726 ;
  assign n12261 = x107 & ~n12260 ;
  assign n12262 = n218 | n7017 ;
  assign n12263 = n9222 ^ n7947 ^ 1'b0 ;
  assign n12264 = n1384 | n2889 ;
  assign n12265 = n12264 ^ n6393 ^ n3221 ;
  assign n12266 = n10202 ^ n4010 ^ 1'b0 ;
  assign n12267 = ~n6537 & n12266 ;
  assign n12268 = n10235 ^ n5096 ^ 1'b0 ;
  assign n12269 = n11281 ^ n2773 ^ n1888 ;
  assign n12270 = ~n4425 & n4864 ;
  assign n12271 = n12270 ^ n1079 ^ 1'b0 ;
  assign n12272 = n2286 | n11465 ;
  assign n12273 = n12272 ^ n9298 ^ 1'b0 ;
  assign n12274 = n1744 ^ n249 ^ 1'b0 ;
  assign n12275 = n7400 ^ n4148 ^ 1'b0 ;
  assign n12276 = n5473 ^ n807 ^ 1'b0 ;
  assign n12277 = ~n4661 & n12276 ;
  assign n12278 = n3423 & n4027 ;
  assign n12279 = n12278 ^ x0 ^ 1'b0 ;
  assign n12280 = n877 | n8240 ;
  assign n12281 = n12280 ^ n4632 ^ 1'b0 ;
  assign n12282 = n4110 ^ n3721 ^ 1'b0 ;
  assign n12283 = ( ~n4691 & n9406 ) | ( ~n4691 & n12282 ) | ( n9406 & n12282 ) ;
  assign n12284 = x3 & ~n936 ;
  assign n12285 = n1696 & ~n2538 ;
  assign n12286 = n1256 & n12285 ;
  assign n12287 = n8892 ^ n3158 ^ 1'b0 ;
  assign n12288 = n2969 | n12287 ;
  assign n12289 = n7140 ^ n4598 ^ 1'b0 ;
  assign n12290 = n11500 ^ n6988 ^ 1'b0 ;
  assign n12291 = ~n2239 & n12290 ;
  assign n12292 = n1534 & n5337 ;
  assign n12293 = n1406 & n12292 ;
  assign n12295 = n334 | n8413 ;
  assign n12294 = ~n5689 & n6994 ;
  assign n12296 = n12295 ^ n12294 ^ 1'b0 ;
  assign n12297 = n339 & ~n6304 ;
  assign n12298 = n431 & ~n7301 ;
  assign n12299 = ~n12297 & n12298 ;
  assign n12300 = n12299 ^ n10264 ^ 1'b0 ;
  assign n12301 = ~n7713 & n12300 ;
  assign n12302 = n4726 ^ n2959 ^ 1'b0 ;
  assign n12303 = ( n4050 & n11911 ) | ( n4050 & n12302 ) | ( n11911 & n12302 ) ;
  assign n12305 = n5318 ^ n770 ^ 1'b0 ;
  assign n12306 = ~n339 & n12305 ;
  assign n12304 = n4446 & ~n4578 ;
  assign n12307 = n12306 ^ n12304 ^ 1'b0 ;
  assign n12308 = n12307 ^ n1720 ^ 1'b0 ;
  assign n12309 = n5982 & n12308 ;
  assign n12311 = n4236 ^ n1000 ^ 1'b0 ;
  assign n12310 = n823 & n2872 ;
  assign n12312 = n12311 ^ n12310 ^ 1'b0 ;
  assign n12313 = n11828 ^ n726 ^ 1'b0 ;
  assign n12314 = n12312 & ~n12313 ;
  assign n12317 = x58 & ~n5387 ;
  assign n12315 = n2599 & n6007 ;
  assign n12316 = n3734 & n12315 ;
  assign n12318 = n12317 ^ n12316 ^ n6462 ;
  assign n12319 = n12314 & n12318 ;
  assign n12320 = n10729 ^ n1653 ^ 1'b0 ;
  assign n12321 = n951 & n12320 ;
  assign n12322 = n11878 & n12321 ;
  assign n12323 = n2077 & n12322 ;
  assign n12324 = n2350 ^ n1427 ^ 1'b0 ;
  assign n12325 = ( ~n2879 & n5759 ) | ( ~n2879 & n12324 ) | ( n5759 & n12324 ) ;
  assign n12326 = n7473 & ~n12325 ;
  assign n12329 = n1196 & n4182 ;
  assign n12327 = ~n5057 & n5269 ;
  assign n12328 = ~n11802 & n12327 ;
  assign n12330 = n12329 ^ n12328 ^ 1'b0 ;
  assign n12331 = n9380 ^ n6641 ^ n5900 ;
  assign n12332 = n2466 & n3221 ;
  assign n12333 = ~n6875 & n12332 ;
  assign n12334 = n8374 | n12333 ;
  assign n12335 = n12334 ^ n9480 ^ 1'b0 ;
  assign n12336 = n965 ^ x104 ^ 1'b0 ;
  assign n12337 = n5447 & n12336 ;
  assign n12338 = n12337 ^ n1214 ^ 1'b0 ;
  assign n12339 = n3663 ^ n260 ^ 1'b0 ;
  assign n12342 = n146 | n1438 ;
  assign n12340 = n2709 | n8229 ;
  assign n12341 = n2413 & ~n12340 ;
  assign n12343 = n12342 ^ n12341 ^ n6724 ;
  assign n12344 = n12339 | n12343 ;
  assign n12345 = n12344 ^ x103 ^ 1'b0 ;
  assign n12346 = n12338 & n12345 ;
  assign n12347 = ~n7670 & n12346 ;
  assign n12348 = n7162 | n7918 ;
  assign n12349 = n289 | n2571 ;
  assign n12350 = n12349 ^ n5329 ^ 1'b0 ;
  assign n12351 = n8524 ^ n3382 ^ 1'b0 ;
  assign n12352 = n12351 ^ n4316 ^ n274 ;
  assign n12353 = n12155 ^ n7089 ^ 1'b0 ;
  assign n12354 = n6928 | n7254 ;
  assign n12355 = n1076 | n12354 ;
  assign n12356 = n3236 ^ x44 ^ 1'b0 ;
  assign n12357 = n4195 & n12356 ;
  assign n12358 = ~n12355 & n12357 ;
  assign n12359 = n915 ^ n820 ^ 1'b0 ;
  assign n12360 = n7987 & ~n12359 ;
  assign n12361 = n8860 ^ n8694 ^ n6060 ;
  assign n12362 = n12361 ^ n11908 ^ 1'b0 ;
  assign n12363 = n1068 | n12362 ;
  assign n12364 = ( ~n7068 & n10807 ) | ( ~n7068 & n12363 ) | ( n10807 & n12363 ) ;
  assign n12365 = n3610 & ~n3837 ;
  assign n12366 = ~n7302 & n12365 ;
  assign n12367 = ( n1435 & n7548 ) | ( n1435 & n12366 ) | ( n7548 & n12366 ) ;
  assign n12368 = n12364 | n12367 ;
  assign n12369 = n2134 & ~n12368 ;
  assign n12370 = n3972 | n6354 ;
  assign n12371 = n3011 | n12370 ;
  assign n12372 = n2390 | n12371 ;
  assign n12373 = n4328 & ~n12372 ;
  assign n12374 = n12373 ^ n1190 ^ 1'b0 ;
  assign n12375 = ~n3242 & n8013 ;
  assign n12376 = n12375 ^ n3196 ^ 1'b0 ;
  assign n12377 = ~n6295 & n12376 ;
  assign n12379 = ~n3315 & n8319 ;
  assign n12380 = n12379 ^ n12018 ^ 1'b0 ;
  assign n12378 = n3925 | n4993 ;
  assign n12381 = n12380 ^ n12378 ^ 1'b0 ;
  assign n12382 = n8159 ^ n5435 ^ n1475 ;
  assign n12383 = n9137 ^ n4798 ^ 1'b0 ;
  assign n12384 = n12383 ^ n2699 ^ n1130 ;
  assign n12386 = ~n985 & n10243 ;
  assign n12387 = n12386 ^ n9772 ^ 1'b0 ;
  assign n12388 = n12387 ^ n9651 ^ 1'b0 ;
  assign n12385 = ~n2460 & n8945 ;
  assign n12389 = n12388 ^ n12385 ^ 1'b0 ;
  assign n12392 = ~n661 & n5005 ;
  assign n12390 = n9630 | n11693 ;
  assign n12391 = n12390 ^ n5591 ^ 1'b0 ;
  assign n12393 = n12392 ^ n12391 ^ n2931 ;
  assign n12394 = n9730 ^ n4994 ^ n4074 ;
  assign n12395 = n6430 | n10431 ;
  assign n12396 = n12395 ^ n399 ^ 1'b0 ;
  assign n12397 = n12336 ^ n7718 ^ 1'b0 ;
  assign n12398 = n12396 & n12397 ;
  assign n12399 = n3666 | n11302 ;
  assign n12400 = ~n11953 & n12399 ;
  assign n12401 = n11137 | n12400 ;
  assign n12402 = n7923 ^ n1147 ^ 1'b0 ;
  assign n12403 = ~n3316 & n12402 ;
  assign n12404 = n12403 ^ n5912 ^ 1'b0 ;
  assign n12405 = ~n3390 & n12404 ;
  assign n12406 = ( n6928 & ~n8239 ) | ( n6928 & n12405 ) | ( ~n8239 & n12405 ) ;
  assign n12407 = n3803 | n4458 ;
  assign n12408 = n1521 & ~n12407 ;
  assign n12409 = n12408 ^ n5290 ^ 1'b0 ;
  assign n12410 = n4743 & n12409 ;
  assign n12411 = ~n8901 & n12410 ;
  assign n12412 = ( n5372 & n8052 ) | ( n5372 & n10613 ) | ( n8052 & n10613 ) ;
  assign n12416 = n12039 ^ n240 ^ 1'b0 ;
  assign n12417 = ~n3469 & n12416 ;
  assign n12413 = ~n2167 & n5460 ;
  assign n12414 = ~n9113 & n12413 ;
  assign n12415 = n1900 | n12414 ;
  assign n12418 = n12417 ^ n12415 ^ 1'b0 ;
  assign n12419 = n7437 ^ n6271 ^ n2028 ;
  assign n12420 = n12419 ^ n8229 ^ 1'b0 ;
  assign n12421 = n12418 & n12420 ;
  assign n12422 = n3802 & ~n9118 ;
  assign n12423 = n12422 ^ n6044 ^ n1582 ;
  assign n12424 = n9638 ^ n3162 ^ 1'b0 ;
  assign n12425 = n203 | n2991 ;
  assign n12426 = n3824 & ~n12425 ;
  assign n12427 = n8129 & n12426 ;
  assign n12428 = n3319 ^ x41 ^ 1'b0 ;
  assign n12429 = n5396 & n12428 ;
  assign n12430 = n12429 ^ n7725 ^ 1'b0 ;
  assign n12431 = ~n7934 & n9004 ;
  assign n12432 = ~n12430 & n12431 ;
  assign n12433 = ( n1046 & ~n2534 ) | ( n1046 & n12432 ) | ( ~n2534 & n12432 ) ;
  assign n12434 = n4999 & ~n7754 ;
  assign n12435 = n6381 & n12434 ;
  assign n12437 = n5313 ^ n3505 ^ 1'b0 ;
  assign n12438 = ~n7516 & n12437 ;
  assign n12439 = n12438 ^ n5977 ^ 1'b0 ;
  assign n12436 = n3880 & ~n8135 ;
  assign n12440 = n12439 ^ n12436 ^ 1'b0 ;
  assign n12441 = n4660 ^ n2347 ^ 1'b0 ;
  assign n12442 = n1888 & ~n12441 ;
  assign n12443 = ( n825 & n2301 ) | ( n825 & ~n12442 ) | ( n2301 & ~n12442 ) ;
  assign n12444 = n5578 ^ n4580 ^ 1'b0 ;
  assign n12445 = n12443 & n12444 ;
  assign n12446 = n5074 & ~n12149 ;
  assign n12447 = n8546 ^ n4973 ^ x8 ;
  assign n12448 = n2445 & ~n4844 ;
  assign n12449 = n11306 ^ n727 ^ 1'b0 ;
  assign n12450 = n1615 | n12449 ;
  assign n12451 = n12450 ^ n5746 ^ 1'b0 ;
  assign n12452 = n12451 ^ n2200 ^ n742 ;
  assign n12453 = n7989 | n8778 ;
  assign n12454 = ( n1317 & n4794 ) | ( n1317 & n7291 ) | ( n4794 & n7291 ) ;
  assign n12455 = n11730 & ~n12454 ;
  assign n12456 = ~n12453 & n12455 ;
  assign n12458 = ~n5552 & n9848 ;
  assign n12457 = n6426 ^ n4960 ^ n2366 ;
  assign n12459 = n12458 ^ n12457 ^ 1'b0 ;
  assign n12460 = ~n11376 & n12459 ;
  assign n12462 = n4041 ^ n625 ^ 1'b0 ;
  assign n12463 = n2500 & ~n12462 ;
  assign n12461 = n1741 & n9872 ;
  assign n12464 = n12463 ^ n12461 ^ n7788 ;
  assign n12465 = n12464 ^ n9802 ^ n9352 ;
  assign n12467 = n3503 & ~n9231 ;
  assign n12466 = ~n938 & n1542 ;
  assign n12468 = n12467 ^ n12466 ^ 1'b0 ;
  assign n12469 = ~n211 & n3964 ;
  assign n12470 = ~n870 & n12469 ;
  assign n12471 = x8 & ~n12470 ;
  assign n12472 = n12471 ^ n1860 ^ 1'b0 ;
  assign n12473 = ( n9036 & n10119 ) | ( n9036 & n12472 ) | ( n10119 & n12472 ) ;
  assign n12474 = n12473 ^ n161 ^ 1'b0 ;
  assign n12475 = n12468 & n12474 ;
  assign n12476 = n9303 ^ n5132 ^ 1'b0 ;
  assign n12477 = n7721 & n12476 ;
  assign n12478 = ( x92 & n2959 ) | ( x92 & ~n6461 ) | ( n2959 & ~n6461 ) ;
  assign n12479 = n1983 & n12478 ;
  assign n12480 = ~n12477 & n12479 ;
  assign n12481 = n10523 ^ n227 ^ n212 ;
  assign n12482 = n5973 ^ n3022 ^ 1'b0 ;
  assign n12483 = n12482 ^ n6004 ^ n2756 ;
  assign n12485 = n10057 ^ n9157 ^ n2456 ;
  assign n12484 = n7240 | n8448 ;
  assign n12486 = n12485 ^ n12484 ^ 1'b0 ;
  assign n12487 = n7463 & n11409 ;
  assign n12488 = n4169 ^ n1350 ^ 1'b0 ;
  assign n12489 = n5732 & ~n12488 ;
  assign n12490 = ~n12487 & n12489 ;
  assign n12491 = n3308 & ~n9503 ;
  assign n12492 = n12491 ^ n8084 ^ 1'b0 ;
  assign n12493 = ~n335 & n10918 ;
  assign n12494 = n12493 ^ n6195 ^ 1'b0 ;
  assign n12495 = ~n1422 & n12494 ;
  assign n12496 = ~n2228 & n6173 ;
  assign n12497 = n5552 ^ n4495 ^ n3978 ;
  assign n12499 = n6335 ^ n1567 ^ 1'b0 ;
  assign n12498 = n7083 & ~n11763 ;
  assign n12500 = n12499 ^ n12498 ^ 1'b0 ;
  assign n12501 = n2179 ^ n1148 ^ 1'b0 ;
  assign n12502 = ~n1767 & n12336 ;
  assign n12503 = ~n2021 & n12502 ;
  assign n12504 = n12503 ^ n7583 ^ n3968 ;
  assign n12507 = n1068 & ~n4645 ;
  assign n12506 = n4170 & n6581 ;
  assign n12508 = n12507 ^ n12506 ^ 1'b0 ;
  assign n12505 = n3479 & ~n6374 ;
  assign n12509 = n12508 ^ n12505 ^ 1'b0 ;
  assign n12510 = n1700 | n12509 ;
  assign n12511 = ~n2991 & n5569 ;
  assign n12512 = n2767 & ~n5186 ;
  assign n12513 = n2306 & ~n12512 ;
  assign n12514 = n4292 & ~n12513 ;
  assign n12515 = n3349 | n12514 ;
  assign n12516 = n10867 ^ n5614 ^ n3001 ;
  assign n12517 = n2776 & n12516 ;
  assign n12518 = n11356 & n12517 ;
  assign n12519 = n12518 ^ n9911 ^ 1'b0 ;
  assign n12520 = n12519 ^ n1510 ^ 1'b0 ;
  assign n12521 = ( n3612 & n3919 ) | ( n3612 & ~n12520 ) | ( n3919 & ~n12520 ) ;
  assign n12522 = n8818 & ~n12521 ;
  assign n12523 = n10406 ^ x61 ^ 1'b0 ;
  assign n12524 = n12523 ^ n9985 ^ n985 ;
  assign n12525 = n12440 ^ n12297 ^ n9726 ;
  assign n12526 = n3248 | n7839 ;
  assign n12527 = n12526 ^ n4483 ^ 1'b0 ;
  assign n12528 = ( n6258 & ~n7428 ) | ( n6258 & n7775 ) | ( ~n7428 & n7775 ) ;
  assign n12529 = ( n1527 & ~n4208 ) | ( n1527 & n5501 ) | ( ~n4208 & n5501 ) ;
  assign n12530 = n12529 ^ n2809 ^ 1'b0 ;
  assign n12531 = n8799 ^ n6407 ^ 1'b0 ;
  assign n12532 = ( n3781 & n5676 ) | ( n3781 & n7670 ) | ( n5676 & n7670 ) ;
  assign n12533 = n10958 ^ n7550 ^ 1'b0 ;
  assign n12534 = ~n1748 & n12533 ;
  assign n12535 = n12534 ^ n6646 ^ 1'b0 ;
  assign n12536 = n7994 & ~n12535 ;
  assign n12537 = n601 & ~n944 ;
  assign n12538 = n9200 ^ n4820 ^ 1'b0 ;
  assign n12539 = n12537 | n12538 ;
  assign n12540 = n2029 & n2420 ;
  assign n12541 = n2520 | n4855 ;
  assign n12542 = n12540 & ~n12541 ;
  assign n12543 = ~n685 & n12542 ;
  assign n12544 = n1493 & n12543 ;
  assign n12545 = n11215 & n12544 ;
  assign n12546 = n5543 & ~n7717 ;
  assign n12547 = n12546 ^ n10822 ^ 1'b0 ;
  assign n12548 = n1218 & ~n12547 ;
  assign n12549 = n4340 & n12548 ;
  assign n12550 = n2772 & n11870 ;
  assign n12551 = n12550 ^ n3150 ^ 1'b0 ;
  assign n12552 = n5703 & n12551 ;
  assign n12555 = x42 & n4210 ;
  assign n12553 = n7960 ^ n746 ^ n322 ;
  assign n12554 = n12553 ^ n9795 ^ n9544 ;
  assign n12556 = n12555 ^ n12554 ^ 1'b0 ;
  assign n12557 = n12552 & n12556 ;
  assign n12558 = n1725 & ~n12557 ;
  assign n12559 = n4646 ^ n1162 ^ 1'b0 ;
  assign n12560 = n2657 ^ n363 ^ 1'b0 ;
  assign n12561 = n770 & n12560 ;
  assign n12562 = n12561 ^ n886 ^ 1'b0 ;
  assign n12563 = n12559 & ~n12562 ;
  assign n12564 = ~n2124 & n12563 ;
  assign n12565 = n10960 ^ n10423 ^ n4662 ;
  assign n12566 = ( n980 & ~n11779 ) | ( n980 & n12565 ) | ( ~n11779 & n12565 ) ;
  assign n12567 = n6228 & n7269 ;
  assign n12568 = n12567 ^ n3054 ^ 1'b0 ;
  assign n12569 = n12568 ^ n4029 ^ n2124 ;
  assign n12570 = ~n8942 & n10076 ;
  assign n12571 = n5479 & n10107 ;
  assign n12572 = ( ~n950 & n9866 ) | ( ~n950 & n12571 ) | ( n9866 & n12571 ) ;
  assign n12573 = n6467 ^ n4166 ^ 1'b0 ;
  assign n12574 = n12573 ^ n5860 ^ n4993 ;
  assign n12575 = n2365 & ~n7956 ;
  assign n12576 = n8350 & n12575 ;
  assign n12577 = n9171 | n12576 ;
  assign n12578 = ~n982 & n1524 ;
  assign n12579 = n11412 | n12578 ;
  assign n12580 = n12579 ^ n9412 ^ n8854 ;
  assign n12581 = ~n2046 & n2731 ;
  assign n12582 = n4590 | n12581 ;
  assign n12583 = n12582 ^ n4452 ^ 1'b0 ;
  assign n12584 = n443 | n4669 ;
  assign n12585 = n12584 ^ n2641 ^ x106 ;
  assign n12586 = n1881 & ~n5765 ;
  assign n12587 = n12586 ^ n2763 ^ 1'b0 ;
  assign n12588 = ~n2898 & n3247 ;
  assign n12589 = n5384 & n8466 ;
  assign n12590 = n12589 ^ n6645 ^ 1'b0 ;
  assign n12592 = n2072 ^ n906 ^ 1'b0 ;
  assign n12593 = ~n1040 & n12592 ;
  assign n12591 = ~n1928 & n6756 ;
  assign n12594 = n12593 ^ n12591 ^ 1'b0 ;
  assign n12595 = n12594 ^ n9620 ^ 1'b0 ;
  assign n12596 = ~n12590 & n12595 ;
  assign n12597 = ( ~n1099 & n12588 ) | ( ~n1099 & n12596 ) | ( n12588 & n12596 ) ;
  assign n12598 = n6929 ^ n6496 ^ n285 ;
  assign n12599 = n12598 ^ n6860 ^ 1'b0 ;
  assign n12600 = ~n4942 & n7814 ;
  assign n12601 = n5425 & n9790 ;
  assign n12602 = n12601 ^ n6129 ^ 1'b0 ;
  assign n12604 = n1750 & n10260 ;
  assign n12603 = n1041 & n4945 ;
  assign n12605 = n12604 ^ n12603 ^ 1'b0 ;
  assign n12606 = n5442 ^ n3552 ^ 1'b0 ;
  assign n12607 = n7221 | n12606 ;
  assign n12610 = ( n3196 & ~n6013 ) | ( n3196 & n7548 ) | ( ~n6013 & n7548 ) ;
  assign n12611 = n12610 ^ n7648 ^ 1'b0 ;
  assign n12609 = n4271 ^ n2731 ^ 1'b0 ;
  assign n12608 = n3003 | n3953 ;
  assign n12612 = n12611 ^ n12609 ^ n12608 ;
  assign n12613 = n4584 | n5558 ;
  assign n12614 = n2756 & ~n12613 ;
  assign n12615 = n2597 & ~n12614 ;
  assign n12616 = ~n8786 & n10756 ;
  assign n12617 = ( ~x12 & n2488 ) | ( ~x12 & n7439 ) | ( n2488 & n7439 ) ;
  assign n12621 = n3974 ^ n2399 ^ 1'b0 ;
  assign n12620 = n5632 | n8240 ;
  assign n12622 = n12621 ^ n12620 ^ 1'b0 ;
  assign n12618 = ( n7402 & ~n7412 ) | ( n7402 & n9424 ) | ( ~n7412 & n9424 ) ;
  assign n12619 = n12618 ^ n4904 ^ n1880 ;
  assign n12623 = n12622 ^ n12619 ^ n1569 ;
  assign n12624 = n4938 & n12623 ;
  assign n12625 = ( n867 & n9860 ) | ( n867 & ~n11463 ) | ( n9860 & ~n11463 ) ;
  assign n12626 = n9955 ^ n8933 ^ 1'b0 ;
  assign n12627 = n3423 ^ n1611 ^ 1'b0 ;
  assign n12628 = n886 | n12627 ;
  assign n12629 = ~n968 & n12628 ;
  assign n12630 = n12626 | n12629 ;
  assign n12631 = n12625 | n12630 ;
  assign n12632 = ( n1637 & ~n2113 ) | ( n1637 & n4572 ) | ( ~n2113 & n4572 ) ;
  assign n12633 = n12632 ^ n5252 ^ 1'b0 ;
  assign n12634 = n8626 & ~n12633 ;
  assign n12635 = n4007 & ~n6076 ;
  assign n12636 = n12635 ^ n9668 ^ 1'b0 ;
  assign n12637 = n1273 ^ n256 ^ 1'b0 ;
  assign n12638 = n12637 ^ n6886 ^ n1819 ;
  assign n12639 = n12636 | n12638 ;
  assign n12640 = n2987 & ~n4433 ;
  assign n12641 = ~n193 & n9175 ;
  assign n12642 = n6834 & n12641 ;
  assign n12643 = n1308 & n12642 ;
  assign n12644 = ( n2055 & ~n3255 ) | ( n2055 & n4664 ) | ( ~n3255 & n4664 ) ;
  assign n12645 = n1069 & n12644 ;
  assign n12646 = n12645 ^ n4564 ^ 1'b0 ;
  assign n12647 = n12646 ^ n4925 ^ n3378 ;
  assign n12648 = n12647 ^ n9173 ^ n5815 ;
  assign n12650 = n10308 | n11748 ;
  assign n12651 = n12650 ^ n4426 ^ 1'b0 ;
  assign n12649 = n6009 & n9513 ;
  assign n12652 = n12651 ^ n12649 ^ 1'b0 ;
  assign n12653 = n12341 ^ n449 ^ 1'b0 ;
  assign n12654 = ~n3537 & n12653 ;
  assign n12655 = n11287 ^ n5737 ^ 1'b0 ;
  assign n12656 = n10413 & n12655 ;
  assign n12657 = n5870 ^ n470 ^ 1'b0 ;
  assign n12658 = n5984 | n9744 ;
  assign n12659 = n12657 & ~n12658 ;
  assign n12660 = n2125 | n10467 ;
  assign n12663 = ~n3169 & n6496 ;
  assign n12664 = ~n356 & n12663 ;
  assign n12665 = n1046 & n12664 ;
  assign n12666 = n5874 ^ n1441 ^ n1305 ;
  assign n12667 = n12665 & ~n12666 ;
  assign n12668 = n12667 ^ n1264 ^ 1'b0 ;
  assign n12661 = n1736 ^ n1470 ^ 1'b0 ;
  assign n12662 = ~n696 & n12661 ;
  assign n12669 = n12668 ^ n12662 ^ n8200 ;
  assign n12670 = n2969 ^ n2105 ^ 1'b0 ;
  assign n12671 = n4513 ^ n1523 ^ 1'b0 ;
  assign n12672 = n5132 | n12671 ;
  assign n12673 = n9406 ^ n5637 ^ n4733 ;
  assign n12674 = n8705 | n12673 ;
  assign n12675 = n12672 & ~n12674 ;
  assign n12676 = n798 & ~n6154 ;
  assign n12677 = n9921 & n12676 ;
  assign n12678 = n10887 ^ n9831 ^ n2061 ;
  assign n12679 = ( n5401 & ~n12677 ) | ( n5401 & n12678 ) | ( ~n12677 & n12678 ) ;
  assign n12681 = n5006 ^ n1748 ^ 1'b0 ;
  assign n12680 = n1417 & ~n3540 ;
  assign n12682 = n12681 ^ n12680 ^ 1'b0 ;
  assign n12683 = n8887 & n12682 ;
  assign n12684 = n12683 ^ n11737 ^ 1'b0 ;
  assign n12685 = n3037 | n12684 ;
  assign n12689 = n5623 & ~n7354 ;
  assign n12686 = n7749 ^ n6524 ^ n2834 ;
  assign n12687 = ~n9302 & n12686 ;
  assign n12688 = n10066 & n12687 ;
  assign n12690 = n12689 ^ n12688 ^ 1'b0 ;
  assign n12691 = n9825 ^ n9481 ^ 1'b0 ;
  assign n12692 = n7497 ^ n5818 ^ 1'b0 ;
  assign n12693 = n3669 & ~n12692 ;
  assign n12694 = n7807 & ~n12693 ;
  assign n12695 = n4289 ^ n2625 ^ 1'b0 ;
  assign n12696 = x111 & n2347 ;
  assign n12697 = ( ~n7829 & n12576 ) | ( ~n7829 & n12696 ) | ( n12576 & n12696 ) ;
  assign n12703 = ~n2296 & n4287 ;
  assign n12700 = n1947 & n9926 ;
  assign n12701 = ~n6722 & n12700 ;
  assign n12702 = n2872 & ~n12701 ;
  assign n12704 = n12703 ^ n12702 ^ 1'b0 ;
  assign n12698 = n5160 & n10723 ;
  assign n12699 = ~n1114 & n12698 ;
  assign n12705 = n12704 ^ n12699 ^ 1'b0 ;
  assign n12706 = n7610 & ~n7789 ;
  assign n12707 = ( n968 & n3958 ) | ( n968 & ~n5304 ) | ( n3958 & ~n5304 ) ;
  assign n12708 = n12707 ^ n9833 ^ n6409 ;
  assign n12709 = n7425 ^ n5717 ^ 1'b0 ;
  assign n12710 = ( n9952 & n10151 ) | ( n9952 & n11008 ) | ( n10151 & n11008 ) ;
  assign n12713 = ~x91 & n2534 ;
  assign n12711 = n2880 & n7488 ;
  assign n12712 = ~n1972 & n12711 ;
  assign n12714 = n12713 ^ n12712 ^ 1'b0 ;
  assign n12715 = n8483 | n12714 ;
  assign n12716 = n10969 ^ n2597 ^ 1'b0 ;
  assign n12717 = n6496 & n12716 ;
  assign n12718 = n2064 ^ n639 ^ 1'b0 ;
  assign n12719 = n9237 ^ n5180 ^ 1'b0 ;
  assign n12720 = n12718 & n12719 ;
  assign n12721 = n2316 & ~n12720 ;
  assign n12722 = ~n12717 & n12721 ;
  assign n12723 = n12722 ^ n11576 ^ n1231 ;
  assign n12727 = n3041 & n5822 ;
  assign n12725 = n1388 | n3796 ;
  assign n12724 = n12513 ^ n4341 ^ 1'b0 ;
  assign n12726 = n12725 ^ n12724 ^ n6673 ;
  assign n12728 = n12727 ^ n12726 ^ n819 ;
  assign n12729 = n7958 ^ n6354 ^ n5762 ;
  assign n12730 = ~n617 & n12729 ;
  assign n12731 = n12730 ^ n2259 ^ 1'b0 ;
  assign n12732 = n7484 ^ n4696 ^ 1'b0 ;
  assign n12733 = n6628 | n12732 ;
  assign n12734 = n1632 ^ n1376 ^ 1'b0 ;
  assign n12735 = n12734 ^ n8041 ^ 1'b0 ;
  assign n12736 = ~n862 & n10526 ;
  assign n12737 = ~n3834 & n12736 ;
  assign n12738 = n2660 | n12737 ;
  assign n12739 = n7886 | n12738 ;
  assign n12740 = n7511 & n11782 ;
  assign n12741 = n937 & ~n4387 ;
  assign n12742 = ~n790 & n12741 ;
  assign n12743 = ~n1406 & n8158 ;
  assign n12744 = n6216 & n12743 ;
  assign n12745 = n12744 ^ n11689 ^ 1'b0 ;
  assign n12746 = ~n12742 & n12745 ;
  assign n12747 = n7342 ^ n4774 ^ 1'b0 ;
  assign n12748 = x12 & ~n12747 ;
  assign n12749 = n1953 & n12748 ;
  assign n12751 = n4323 ^ n4103 ^ 1'b0 ;
  assign n12750 = n591 & n6631 ;
  assign n12752 = n12751 ^ n12750 ^ 1'b0 ;
  assign n12757 = n3279 ^ n1420 ^ n362 ;
  assign n12758 = x17 & ~n12757 ;
  assign n12759 = n12758 ^ n4645 ^ 1'b0 ;
  assign n12760 = ~n4703 & n12759 ;
  assign n12761 = ~n1273 & n12760 ;
  assign n12753 = n452 | n4618 ;
  assign n12754 = n139 | n12753 ;
  assign n12755 = n7021 & n12754 ;
  assign n12756 = n3122 & n12755 ;
  assign n12762 = n12761 ^ n12756 ^ n1491 ;
  assign n12763 = n9876 ^ n5788 ^ 1'b0 ;
  assign n12764 = n12039 | n12763 ;
  assign n12765 = ( n2475 & n7401 ) | ( n2475 & ~n7906 ) | ( n7401 & ~n7906 ) ;
  assign n12766 = n1545 | n12765 ;
  assign n12767 = n427 | n2404 ;
  assign n12768 = n12767 ^ n2383 ^ 1'b0 ;
  assign n12769 = n12768 ^ n8392 ^ 1'b0 ;
  assign n12773 = ( n158 & n422 ) | ( n158 & ~n12213 ) | ( n422 & ~n12213 ) ;
  assign n12774 = n12773 ^ n12115 ^ 1'b0 ;
  assign n12770 = n7077 ^ n802 ^ 1'b0 ;
  assign n12771 = n2769 & ~n12770 ;
  assign n12772 = n8994 & n12771 ;
  assign n12775 = n12774 ^ n12772 ^ 1'b0 ;
  assign n12776 = n5784 & n9268 ;
  assign n12777 = n4161 & n12776 ;
  assign n12779 = n240 & n2663 ;
  assign n12778 = n7258 ^ n3730 ^ 1'b0 ;
  assign n12780 = n12779 ^ n12778 ^ n9130 ;
  assign n12782 = ~n1743 & n3682 ;
  assign n12781 = n2809 & n10667 ;
  assign n12783 = n12782 ^ n12781 ^ 1'b0 ;
  assign n12784 = n5099 ^ n3441 ^ n1014 ;
  assign n12785 = n2939 ^ n560 ^ 1'b0 ;
  assign n12786 = ~n2350 & n12785 ;
  assign n12787 = n12786 ^ n5230 ^ 1'b0 ;
  assign n12789 = x112 | n2980 ;
  assign n12790 = n5244 ^ n307 ^ 1'b0 ;
  assign n12791 = n12789 & ~n12790 ;
  assign n12788 = n3614 | n10478 ;
  assign n12792 = n12791 ^ n12788 ^ n195 ;
  assign n12793 = n796 & ~n5800 ;
  assign n12794 = n2031 & n9465 ;
  assign n12795 = n9008 & n12794 ;
  assign n12796 = ~n453 & n2270 ;
  assign n12797 = n12796 ^ n5029 ^ n1773 ;
  assign n12798 = n12797 ^ n11903 ^ 1'b0 ;
  assign n12799 = n6128 | n12798 ;
  assign n12800 = ~n2250 & n11666 ;
  assign n12801 = n9609 & n12800 ;
  assign n12802 = ( n6019 & ~n6747 ) | ( n6019 & n12801 ) | ( ~n6747 & n12801 ) ;
  assign n12803 = n5399 ^ n3104 ^ 1'b0 ;
  assign n12804 = n9702 | n12803 ;
  assign n12805 = n10436 & ~n11136 ;
  assign n12806 = ~n2200 & n2417 ;
  assign n12807 = ~n3082 & n12806 ;
  assign n12808 = n12807 ^ n4641 ^ n526 ;
  assign n12809 = n12808 ^ n3689 ^ 1'b0 ;
  assign n12810 = n12809 ^ n9129 ^ n778 ;
  assign n12811 = ( n12804 & ~n12805 ) | ( n12804 & n12810 ) | ( ~n12805 & n12810 ) ;
  assign n12814 = n4207 ^ n2796 ^ 1'b0 ;
  assign n12815 = n3642 & n12814 ;
  assign n12812 = n5791 ^ n5595 ^ 1'b0 ;
  assign n12813 = n3505 & n12812 ;
  assign n12816 = n12815 ^ n12813 ^ 1'b0 ;
  assign n12817 = n12816 ^ n11741 ^ n4245 ;
  assign n12818 = n436 & n2256 ;
  assign n12819 = n7928 & ~n12818 ;
  assign n12820 = n4524 & n12819 ;
  assign n12821 = n1442 & n1917 ;
  assign n12822 = n12821 ^ n3090 ^ 1'b0 ;
  assign n12823 = n12822 ^ n5988 ^ n2524 ;
  assign n12824 = n10523 & ~n11702 ;
  assign n12825 = n12824 ^ n413 ^ 1'b0 ;
  assign n12826 = n1190 & ~n3663 ;
  assign n12827 = n8231 & n12826 ;
  assign n12828 = n12827 ^ n12578 ^ n606 ;
  assign n12829 = n4833 | n6717 ;
  assign n12830 = n9925 & ~n12829 ;
  assign n12831 = n4281 & ~n12830 ;
  assign n12832 = n2501 & ~n9145 ;
  assign n12833 = n12831 & n12832 ;
  assign n12834 = n5463 ^ n5314 ^ n4774 ;
  assign n12835 = n12834 ^ n9620 ^ 1'b0 ;
  assign n12836 = n2965 & ~n8864 ;
  assign n12837 = n12835 & n12836 ;
  assign n12839 = n849 | n7079 ;
  assign n12838 = n1556 & ~n4250 ;
  assign n12840 = n12839 ^ n12838 ^ 1'b0 ;
  assign n12841 = n2258 ^ n1770 ^ 1'b0 ;
  assign n12842 = n5436 | n11951 ;
  assign n12843 = n12842 ^ n7160 ^ 1'b0 ;
  assign n12844 = n6772 ^ n227 ^ 1'b0 ;
  assign n12845 = n12844 ^ n5423 ^ 1'b0 ;
  assign n12846 = n4849 ^ n3546 ^ 1'b0 ;
  assign n12847 = n12846 ^ n12317 ^ 1'b0 ;
  assign n12848 = ( ~n10076 & n11099 ) | ( ~n10076 & n12847 ) | ( n11099 & n12847 ) ;
  assign n12849 = n12848 ^ n10235 ^ n6664 ;
  assign n12850 = n1774 | n3739 ;
  assign n12851 = n5615 | n7350 ;
  assign n12852 = n1262 | n12851 ;
  assign n12853 = ( n3534 & ~n12850 ) | ( n3534 & n12852 ) | ( ~n12850 & n12852 ) ;
  assign n12858 = n4555 ^ n3521 ^ 1'b0 ;
  assign n12855 = n5854 ^ n1248 ^ 1'b0 ;
  assign n12856 = n1294 & n12855 ;
  assign n12854 = n8914 & n10270 ;
  assign n12857 = n12856 ^ n12854 ^ n1091 ;
  assign n12859 = n12858 ^ n12857 ^ n845 ;
  assign n12860 = n2391 | n8426 ;
  assign n12861 = ( n180 & n5500 ) | ( n180 & n12677 ) | ( n5500 & n12677 ) ;
  assign n12862 = n10960 & n12861 ;
  assign n12863 = n12862 ^ n8935 ^ 1'b0 ;
  assign n12864 = n9606 | n12863 ;
  assign n12867 = n1529 ^ n1375 ^ x126 ;
  assign n12868 = n1374 & n12867 ;
  assign n12869 = n12868 ^ n9497 ^ 1'b0 ;
  assign n12873 = n4329 ^ n3941 ^ n1542 ;
  assign n12874 = n12873 ^ n4079 ^ 1'b0 ;
  assign n12875 = ( n3413 & n4637 ) | ( n3413 & ~n12874 ) | ( n4637 & ~n12874 ) ;
  assign n12870 = ( n773 & ~n1619 ) | ( n773 & n4000 ) | ( ~n1619 & n4000 ) ;
  assign n12871 = n1876 & ~n12870 ;
  assign n12872 = n12512 & n12871 ;
  assign n12876 = n12875 ^ n12872 ^ 1'b0 ;
  assign n12877 = n12869 & ~n12876 ;
  assign n12865 = n1373 & n8024 ;
  assign n12866 = n1536 & n12865 ;
  assign n12878 = n12877 ^ n12866 ^ 1'b0 ;
  assign n12879 = n10048 & ~n12878 ;
  assign n12880 = n477 & ~n3024 ;
  assign n12881 = ~n1964 & n12880 ;
  assign n12882 = ( n2728 & n8298 ) | ( n2728 & ~n12881 ) | ( n8298 & ~n12881 ) ;
  assign n12883 = n4523 ^ n744 ^ 1'b0 ;
  assign n12884 = n12882 | n12883 ;
  assign n12885 = ( ~n1039 & n4167 ) | ( ~n1039 & n11182 ) | ( n4167 & n11182 ) ;
  assign n12886 = n12885 ^ n403 ^ 1'b0 ;
  assign n12887 = ~n452 & n4911 ;
  assign n12888 = n12887 ^ n1456 ^ 1'b0 ;
  assign n12889 = n12888 ^ n6946 ^ n4498 ;
  assign n12890 = n3541 ^ n3397 ^ 1'b0 ;
  assign n12891 = n2387 & ~n12890 ;
  assign n12892 = n1567 ^ n206 ^ 1'b0 ;
  assign n12893 = n878 & n12892 ;
  assign n12894 = n10343 | n12893 ;
  assign n12895 = n12891 | n12894 ;
  assign n12896 = ( ~n5164 & n6193 ) | ( ~n5164 & n11060 ) | ( n6193 & n11060 ) ;
  assign n12897 = ( n4463 & ~n6197 ) | ( n4463 & n12896 ) | ( ~n6197 & n12896 ) ;
  assign n12898 = n6273 | n12897 ;
  assign n12899 = n12898 ^ n8491 ^ 1'b0 ;
  assign n12908 = ~n1131 & n2567 ;
  assign n12909 = n12908 ^ n8961 ^ 1'b0 ;
  assign n12900 = n4070 ^ n3365 ^ x90 ;
  assign n12901 = n12900 ^ n4011 ^ 1'b0 ;
  assign n12905 = n2497 & ~n9303 ;
  assign n12902 = ~n1548 & n1674 ;
  assign n12903 = n475 | n9236 ;
  assign n12904 = n12902 & ~n12903 ;
  assign n12906 = n12905 ^ n12904 ^ n7854 ;
  assign n12907 = n12901 & ~n12906 ;
  assign n12910 = n12909 ^ n12907 ^ 1'b0 ;
  assign n12911 = n4447 ^ n867 ^ 1'b0 ;
  assign n12912 = n1381 | n2758 ;
  assign n12913 = n12911 | n12912 ;
  assign n12918 = n798 & n7327 ;
  assign n12914 = n3159 ^ x96 ^ 1'b0 ;
  assign n12915 = ~n4926 & n12914 ;
  assign n12916 = n7499 | n12915 ;
  assign n12917 = n8005 & n12916 ;
  assign n12919 = n12918 ^ n12917 ^ 1'b0 ;
  assign n12920 = n6143 ^ n6096 ^ 1'b0 ;
  assign n12921 = n5500 & ~n12920 ;
  assign n12922 = n11168 ^ n8255 ^ 1'b0 ;
  assign n12923 = n11469 ^ n3677 ^ n1415 ;
  assign n12924 = n12922 & n12923 ;
  assign n12925 = n12924 ^ n5235 ^ 1'b0 ;
  assign n12926 = n7520 & n12925 ;
  assign n12927 = ~n3890 & n7003 ;
  assign n12928 = n10919 ^ n4901 ^ 1'b0 ;
  assign n12929 = n2267 ^ n131 ^ 1'b0 ;
  assign n12930 = n7976 & n12929 ;
  assign n12931 = n397 | n947 ;
  assign n12932 = n12931 ^ n7730 ^ 1'b0 ;
  assign n12933 = n2965 | n12932 ;
  assign n12934 = n12933 ^ n1603 ^ 1'b0 ;
  assign n12935 = n10114 ^ n2349 ^ 1'b0 ;
  assign n12936 = ~n4753 & n6515 ;
  assign n12937 = n2565 ^ n1982 ^ 1'b0 ;
  assign n12938 = n12937 ^ n9673 ^ n410 ;
  assign n12939 = n2824 & n8272 ;
  assign n12940 = n12938 & ~n12939 ;
  assign n12941 = n1090 | n7610 ;
  assign n12944 = n1910 | n3106 ;
  assign n12945 = n12944 ^ n3828 ^ n755 ;
  assign n12946 = n12304 & n12945 ;
  assign n12943 = ~n1615 & n6178 ;
  assign n12947 = n12946 ^ n12943 ^ 1'b0 ;
  assign n12948 = ~n153 & n12947 ;
  assign n12942 = n356 & ~n11027 ;
  assign n12949 = n12948 ^ n12942 ^ 1'b0 ;
  assign n12950 = ( ~n1302 & n1445 ) | ( ~n1302 & n2089 ) | ( n1445 & n2089 ) ;
  assign n12951 = n6264 & n12950 ;
  assign n12952 = n6415 ^ n4887 ^ n2068 ;
  assign n12953 = n2981 & ~n9421 ;
  assign n12954 = n12953 ^ n4592 ^ 1'b0 ;
  assign n12955 = ~n12687 & n12954 ;
  assign n12956 = ~n3244 & n8924 ;
  assign n12957 = n12956 ^ n6663 ^ 1'b0 ;
  assign n12958 = ~n1366 & n12937 ;
  assign n12959 = n12958 ^ n7520 ^ 1'b0 ;
  assign n12960 = n12959 ^ n7774 ^ n6289 ;
  assign n12961 = ( n2241 & n4973 ) | ( n2241 & ~n8685 ) | ( n4973 & ~n8685 ) ;
  assign n12962 = ( n6208 & ~n10959 ) | ( n6208 & n12961 ) | ( ~n10959 & n12961 ) ;
  assign n12963 = ~n6730 & n8500 ;
  assign n12964 = n12963 ^ n4712 ^ 1'b0 ;
  assign n12965 = n11151 & n12964 ;
  assign n12966 = ~n5828 & n12965 ;
  assign n12967 = n2641 | n4917 ;
  assign n12968 = n3921 & ~n12967 ;
  assign n12969 = n12968 ^ x97 ^ 1'b0 ;
  assign n12970 = n5425 & ~n12969 ;
  assign n12971 = n12970 ^ n3615 ^ 1'b0 ;
  assign n12972 = n6537 & ~n12971 ;
  assign n12973 = ~n8690 & n12972 ;
  assign n12974 = n1550 ^ n936 ^ n425 ;
  assign n12975 = n3461 & n12974 ;
  assign n12976 = n12975 ^ n9705 ^ n218 ;
  assign n12977 = n3118 & n3758 ;
  assign n12978 = ( n634 & n5317 ) | ( n634 & n12977 ) | ( n5317 & n12977 ) ;
  assign n12979 = ( n5694 & ~n5698 ) | ( n5694 & n12350 ) | ( ~n5698 & n12350 ) ;
  assign n12980 = n2254 & ~n8522 ;
  assign n12981 = n12980 ^ n8763 ^ 1'b0 ;
  assign n12982 = n1163 | n12981 ;
  assign n12983 = ( ~n5421 & n11213 ) | ( ~n5421 & n12982 ) | ( n11213 & n12982 ) ;
  assign n12984 = ~x9 & n5151 ;
  assign n12985 = n1382 | n3928 ;
  assign n12986 = n4983 | n12985 ;
  assign n12987 = n6635 & ~n10485 ;
  assign n12988 = n2421 & n9889 ;
  assign n12989 = n11981 & n12988 ;
  assign n12992 = n4937 & ~n5952 ;
  assign n12993 = n12992 ^ n5380 ^ 1'b0 ;
  assign n12990 = n967 | n5093 ;
  assign n12991 = n2256 & ~n12990 ;
  assign n12994 = n12993 ^ n12991 ^ n4385 ;
  assign n12995 = n12388 ^ n8135 ^ n3552 ;
  assign n12996 = n5335 & n5955 ;
  assign n12997 = ~n1739 & n12996 ;
  assign n13000 = ( n3923 & n8955 ) | ( n3923 & n9670 ) | ( n8955 & n9670 ) ;
  assign n12998 = n325 | n1292 ;
  assign n12999 = n12998 ^ n11836 ^ 1'b0 ;
  assign n13001 = n13000 ^ n12999 ^ 1'b0 ;
  assign n13002 = n6512 ^ n794 ^ n252 ;
  assign n13003 = n3981 ^ n2917 ^ 1'b0 ;
  assign n13004 = n2829 & ~n13003 ;
  assign n13005 = n13002 & n13004 ;
  assign n13006 = n3023 & n10720 ;
  assign n13007 = n13006 ^ n4341 ^ n2321 ;
  assign n13008 = n7691 ^ n5431 ^ 1'b0 ;
  assign n13009 = ~n9220 & n13008 ;
  assign n13010 = n13007 & n13009 ;
  assign n13011 = n5775 ^ n1215 ^ 1'b0 ;
  assign n13012 = n2912 & n13011 ;
  assign n13013 = n6996 ^ n3199 ^ 1'b0 ;
  assign n13014 = n3059 & n13013 ;
  assign n13015 = ~n190 & n13014 ;
  assign n13016 = n13015 ^ n1173 ^ 1'b0 ;
  assign n13017 = n7221 ^ n6131 ^ 1'b0 ;
  assign n13018 = n8225 ^ n2078 ^ 1'b0 ;
  assign n13019 = n6681 & ~n6982 ;
  assign n13020 = n2633 & n13019 ;
  assign n13021 = ~n10416 & n13020 ;
  assign n13022 = n1910 ^ x57 ^ 1'b0 ;
  assign n13023 = n1695 | n13022 ;
  assign n13024 = ( n1226 & ~n1934 ) | ( n1226 & n8793 ) | ( ~n1934 & n8793 ) ;
  assign n13025 = n13024 ^ n8201 ^ n5258 ;
  assign n13026 = n13025 ^ n8662 ^ 1'b0 ;
  assign n13027 = n10753 ^ n969 ^ 1'b0 ;
  assign n13028 = ~n10618 & n13027 ;
  assign n13029 = n278 & n1621 ;
  assign n13030 = n381 | n13029 ;
  assign n13031 = n4071 & ~n13030 ;
  assign n13032 = n6220 ^ n4347 ^ 1'b0 ;
  assign n13033 = ~n1428 & n6924 ;
  assign n13034 = ~n13032 & n13033 ;
  assign n13035 = n1316 | n2306 ;
  assign n13036 = n13034 & ~n13035 ;
  assign n13037 = x51 | n8413 ;
  assign n13038 = n970 & n13037 ;
  assign n13039 = n1633 & n5060 ;
  assign n13040 = n711 & n13039 ;
  assign n13041 = n13040 ^ n9662 ^ n7473 ;
  assign n13042 = n9237 & n13041 ;
  assign n13043 = ( n452 & ~n5170 ) | ( n452 & n13042 ) | ( ~n5170 & n13042 ) ;
  assign n13044 = n9287 ^ n6472 ^ 1'b0 ;
  assign n13045 = n7852 ^ n701 ^ 1'b0 ;
  assign n13046 = n13045 ^ n3785 ^ n587 ;
  assign n13047 = n1358 | n6838 ;
  assign n13048 = n13046 & ~n13047 ;
  assign n13049 = n3040 & ~n4698 ;
  assign n13050 = ~n7133 & n12504 ;
  assign n13051 = n13049 & n13050 ;
  assign n13052 = n6758 ^ n1370 ^ 1'b0 ;
  assign n13053 = n9225 & ~n13052 ;
  assign n13054 = n13053 ^ n1181 ^ 1'b0 ;
  assign n13055 = n5366 | n13054 ;
  assign n13056 = n13055 ^ n6744 ^ 1'b0 ;
  assign n13057 = n2822 & ~n5153 ;
  assign n13058 = n4808 | n4847 ;
  assign n13059 = n13058 ^ n3428 ^ 1'b0 ;
  assign n13060 = n4570 ^ n1136 ^ n490 ;
  assign n13061 = n13060 ^ n4356 ^ 1'b0 ;
  assign n13062 = ( n681 & n13059 ) | ( n681 & ~n13061 ) | ( n13059 & ~n13061 ) ;
  assign n13063 = ~n9443 & n11873 ;
  assign n13064 = n167 | n6117 ;
  assign n13065 = n3741 ^ n1073 ^ n635 ;
  assign n13066 = n6207 ^ n2517 ^ 1'b0 ;
  assign n13067 = ~n13065 & n13066 ;
  assign n13068 = n218 | n7769 ;
  assign n13069 = n6567 ^ n3856 ^ n2072 ;
  assign n13070 = n13069 ^ n3136 ^ n673 ;
  assign n13071 = ( ~n932 & n3348 ) | ( ~n932 & n5823 ) | ( n3348 & n5823 ) ;
  assign n13072 = n8386 ^ n6247 ^ 1'b0 ;
  assign n13073 = ~n4486 & n13072 ;
  assign n13074 = n13073 ^ n9913 ^ 1'b0 ;
  assign n13075 = n2108 & n13074 ;
  assign n13076 = n1817 & n13075 ;
  assign n13077 = n402 & ~n8649 ;
  assign n13078 = ~n589 & n13077 ;
  assign n13079 = ( n4743 & ~n7726 ) | ( n4743 & n13078 ) | ( ~n7726 & n13078 ) ;
  assign n13080 = n982 | n5643 ;
  assign n13081 = n3533 & ~n13080 ;
  assign n13082 = n10164 & ~n13081 ;
  assign n13083 = ~n7730 & n13082 ;
  assign n13084 = n1064 | n5808 ;
  assign n13085 = ~n331 & n4035 ;
  assign n13086 = ~n3013 & n13085 ;
  assign n13087 = n13086 ^ n6603 ^ 1'b0 ;
  assign n13088 = n4539 ^ n3650 ^ 1'b0 ;
  assign n13089 = ( n3613 & ~n12818 ) | ( n3613 & n13088 ) | ( ~n12818 & n13088 ) ;
  assign n13090 = ( n2111 & n6447 ) | ( n2111 & n10793 ) | ( n6447 & n10793 ) ;
  assign n13091 = n10132 | n13090 ;
  assign n13092 = ( n2687 & n5986 ) | ( n2687 & ~n12470 ) | ( n5986 & ~n12470 ) ;
  assign n13093 = ~n484 & n6512 ;
  assign n13094 = n13093 ^ n420 ^ 1'b0 ;
  assign n13095 = n4633 ^ n3589 ^ n1470 ;
  assign n13099 = ( n172 & n770 ) | ( n172 & n9548 ) | ( n770 & n9548 ) ;
  assign n13096 = n3615 & ~n8318 ;
  assign n13097 = ( n138 & ~n1138 ) | ( n138 & n13096 ) | ( ~n1138 & n13096 ) ;
  assign n13098 = ~n1441 & n13097 ;
  assign n13100 = n13099 ^ n13098 ^ 1'b0 ;
  assign n13101 = n6550 ^ n4289 ^ 1'b0 ;
  assign n13102 = n4927 | n13101 ;
  assign n13103 = n13102 ^ n10341 ^ n3056 ;
  assign n13104 = ( x68 & n6740 ) | ( x68 & n13103 ) | ( n6740 & n13103 ) ;
  assign n13107 = n6803 | n10656 ;
  assign n13108 = n13107 ^ n1018 ^ 1'b0 ;
  assign n13105 = n2844 & ~n8231 ;
  assign n13106 = n3615 & n13105 ;
  assign n13109 = n13108 ^ n13106 ^ 1'b0 ;
  assign n13110 = ~n533 & n3859 ;
  assign n13111 = ( ~n1703 & n6565 ) | ( ~n1703 & n13110 ) | ( n6565 & n13110 ) ;
  assign n13112 = n7974 ^ n1291 ^ 1'b0 ;
  assign n13113 = n1908 | n13112 ;
  assign n13114 = n1720 | n13113 ;
  assign n13115 = n4467 & n13114 ;
  assign n13116 = n13111 & n13115 ;
  assign n13118 = n3007 ^ n2949 ^ 1'b0 ;
  assign n13119 = n13118 ^ n9912 ^ n1041 ;
  assign n13117 = n5376 | n7160 ;
  assign n13120 = n13119 ^ n13117 ^ 1'b0 ;
  assign n13121 = n3669 & ~n13120 ;
  assign n13122 = n1096 & n13121 ;
  assign n13123 = n13122 ^ n9028 ^ 1'b0 ;
  assign n13124 = n10629 & n13123 ;
  assign n13125 = ( n5214 & n5841 ) | ( n5214 & n13124 ) | ( n5841 & n13124 ) ;
  assign n13126 = ~n2100 & n2532 ;
  assign n13127 = n13126 ^ n990 ^ 1'b0 ;
  assign n13128 = ( n2417 & n3698 ) | ( n2417 & ~n10980 ) | ( n3698 & ~n10980 ) ;
  assign n13129 = n13128 ^ n726 ^ 1'b0 ;
  assign n13130 = n13129 ^ n12485 ^ 1'b0 ;
  assign n13131 = n13127 & ~n13130 ;
  assign n13132 = n7527 | n11389 ;
  assign n13133 = n2954 ^ n2829 ^ n773 ;
  assign n13134 = n10793 & ~n13133 ;
  assign n13135 = n13132 & n13134 ;
  assign n13138 = ( ~n788 & n2131 ) | ( ~n788 & n4913 ) | ( n2131 & n4913 ) ;
  assign n13136 = n6701 ^ n299 ^ 1'b0 ;
  assign n13137 = n5895 & n13136 ;
  assign n13139 = n13138 ^ n13137 ^ n979 ;
  assign n13142 = ( n5460 & ~n6585 ) | ( n5460 & n10464 ) | ( ~n6585 & n10464 ) ;
  assign n13143 = n13142 ^ n5754 ^ n3371 ;
  assign n13140 = n1788 | n3276 ;
  assign n13141 = n13140 ^ n2115 ^ 1'b0 ;
  assign n13144 = n13143 ^ n13141 ^ n6668 ;
  assign n13145 = n12371 ^ n5686 ^ 1'b0 ;
  assign n13146 = ( ~n3169 & n5572 ) | ( ~n3169 & n13145 ) | ( n5572 & n13145 ) ;
  assign n13147 = ~n6699 & n7457 ;
  assign n13148 = n13147 ^ n4589 ^ 1'b0 ;
  assign n13149 = n13148 ^ x71 ^ 1'b0 ;
  assign n13150 = n13146 & ~n13149 ;
  assign n13151 = ( n2599 & n10152 ) | ( n2599 & n10797 ) | ( n10152 & n10797 ) ;
  assign n13152 = ~n238 & n965 ;
  assign n13153 = n13152 ^ n1992 ^ 1'b0 ;
  assign n13154 = ( n11467 & ~n12399 ) | ( n11467 & n13153 ) | ( ~n12399 & n13153 ) ;
  assign n13155 = ( n827 & ~n6537 ) | ( n827 & n9441 ) | ( ~n6537 & n9441 ) ;
  assign n13156 = ~n4713 & n6513 ;
  assign n13157 = n13156 ^ n11229 ^ 1'b0 ;
  assign n13158 = n2986 | n5536 ;
  assign n13159 = n11397 & ~n13158 ;
  assign n13160 = ~n4146 & n6454 ;
  assign n13161 = n13160 ^ n12830 ^ n4219 ;
  assign n13162 = n9367 ^ n7209 ^ 1'b0 ;
  assign n13163 = n12349 & n13162 ;
  assign n13164 = n13161 & n13163 ;
  assign n13165 = n3794 & n12373 ;
  assign n13166 = ~n3403 & n13165 ;
  assign n13167 = n12757 ^ n4426 ^ 1'b0 ;
  assign n13168 = n3482 & n13167 ;
  assign n13169 = n13168 ^ n8438 ^ 1'b0 ;
  assign n13170 = n9520 | n10913 ;
  assign n13171 = n1769 | n13170 ;
  assign n13172 = n7618 ^ n3548 ^ 1'b0 ;
  assign n13173 = n4035 & n13172 ;
  assign n13174 = n13173 ^ n8430 ^ 1'b0 ;
  assign n13175 = n11797 | n13174 ;
  assign n13176 = ( ~n3523 & n3787 ) | ( ~n3523 & n11752 ) | ( n3787 & n11752 ) ;
  assign n13177 = n515 & ~n5499 ;
  assign n13179 = n13156 ^ n6242 ^ 1'b0 ;
  assign n13180 = n3821 & n13179 ;
  assign n13178 = n6442 & n7602 ;
  assign n13181 = n13180 ^ n13178 ^ 1'b0 ;
  assign n13182 = ( n5061 & ~n13177 ) | ( n5061 & n13181 ) | ( ~n13177 & n13181 ) ;
  assign n13183 = n387 | n7994 ;
  assign n13184 = n13183 ^ n4691 ^ 1'b0 ;
  assign n13185 = ( ~n331 & n1649 ) | ( ~n331 & n3679 ) | ( n1649 & n3679 ) ;
  assign n13186 = n9042 ^ n4088 ^ n3513 ;
  assign n13187 = n2750 & ~n3787 ;
  assign n13188 = ~n5611 & n13187 ;
  assign n13189 = ( n13185 & ~n13186 ) | ( n13185 & n13188 ) | ( ~n13186 & n13188 ) ;
  assign n13190 = n5294 & n7060 ;
  assign n13191 = n11428 & n13190 ;
  assign n13192 = n603 | n1181 ;
  assign n13193 = n295 | n7758 ;
  assign n13194 = n4123 & ~n9168 ;
  assign n13195 = n13194 ^ n6724 ^ 1'b0 ;
  assign n13196 = ( ~n313 & n5241 ) | ( ~n313 & n13195 ) | ( n5241 & n13195 ) ;
  assign n13197 = n2191 ^ n332 ^ 1'b0 ;
  assign n13198 = n6980 & ~n13197 ;
  assign n13199 = ~n1973 & n13198 ;
  assign n13200 = n13199 ^ n3734 ^ 1'b0 ;
  assign n13202 = n3965 ^ n730 ^ 1'b0 ;
  assign n13203 = n8900 & ~n13202 ;
  assign n13201 = ~n6647 & n9384 ;
  assign n13204 = n13203 ^ n13201 ^ 1'b0 ;
  assign n13205 = n2134 ^ n1179 ^ 1'b0 ;
  assign n13206 = n3884 & n13205 ;
  assign n13207 = ( n4326 & ~n5952 ) | ( n4326 & n8648 ) | ( ~n5952 & n8648 ) ;
  assign n13208 = n13207 ^ n3293 ^ 1'b0 ;
  assign n13209 = n1569 | n2544 ;
  assign n13210 = n10713 & ~n13209 ;
  assign n13211 = n13210 ^ n4445 ^ 1'b0 ;
  assign n13214 = n401 & n1037 ;
  assign n13215 = n13214 ^ n920 ^ 1'b0 ;
  assign n13216 = ( n8230 & n13138 ) | ( n8230 & ~n13215 ) | ( n13138 & ~n13215 ) ;
  assign n13212 = n1298 & n10549 ;
  assign n13213 = n13212 ^ n5406 ^ 1'b0 ;
  assign n13217 = n13216 ^ n13213 ^ n10039 ;
  assign n13218 = ~n148 & n2221 ;
  assign n13219 = n13218 ^ n822 ^ 1'b0 ;
  assign n13220 = n3814 ^ n1725 ^ 1'b0 ;
  assign n13221 = n13219 | n13220 ;
  assign n13222 = n8497 & ~n13221 ;
  assign n13223 = n4898 | n11539 ;
  assign n13224 = n13223 ^ n6457 ^ 1'b0 ;
  assign n13225 = n1311 & n4338 ;
  assign n13226 = ~x2 & n13225 ;
  assign n13227 = n5951 & ~n13226 ;
  assign n13228 = n13224 & n13227 ;
  assign n13229 = n10146 ^ n5305 ^ n1467 ;
  assign n13230 = n13229 ^ n5595 ^ 1'b0 ;
  assign n13231 = ( n7695 & n8185 ) | ( n7695 & n13230 ) | ( n8185 & n13230 ) ;
  assign n13232 = ( ~n4479 & n11323 ) | ( ~n4479 & n12486 ) | ( n11323 & n12486 ) ;
  assign n13236 = n1741 | n5587 ;
  assign n13237 = n2124 | n13236 ;
  assign n13238 = n3316 | n13237 ;
  assign n13233 = n3860 | n7803 ;
  assign n13234 = ( n399 & ~n12858 ) | ( n399 & n13233 ) | ( ~n12858 & n13233 ) ;
  assign n13235 = n4394 & ~n13234 ;
  assign n13239 = n13238 ^ n13235 ^ 1'b0 ;
  assign n13240 = n8417 ^ n4494 ^ n1584 ;
  assign n13241 = ~n6407 & n11653 ;
  assign n13242 = n12626 ^ n1723 ^ n298 ;
  assign n13243 = n2930 | n4267 ;
  assign n13244 = n13243 ^ n10732 ^ 1'b0 ;
  assign n13245 = ~n1008 & n5430 ;
  assign n13246 = n13245 ^ n2333 ^ 1'b0 ;
  assign n13247 = n7827 ^ n2708 ^ 1'b0 ;
  assign n13248 = n13246 & ~n13247 ;
  assign n13249 = n11010 & n13248 ;
  assign n13250 = n5043 & n13249 ;
  assign n13251 = n13244 | n13250 ;
  assign n13252 = ~n5178 & n10704 ;
  assign n13253 = ( ~n2842 & n4253 ) | ( ~n2842 & n10867 ) | ( n4253 & n10867 ) ;
  assign n13254 = n7803 ^ n2651 ^ 1'b0 ;
  assign n13255 = ~n5385 & n13254 ;
  assign n13256 = n9983 ^ n3237 ^ 1'b0 ;
  assign n13257 = ~n4590 & n6600 ;
  assign n13258 = ~n3247 & n13257 ;
  assign n13259 = n7649 | n13258 ;
  assign n13260 = n13256 | n13259 ;
  assign n13261 = n1895 | n8850 ;
  assign n13262 = n13261 ^ n340 ^ 1'b0 ;
  assign n13263 = n4440 & ~n4570 ;
  assign n13264 = n13263 ^ n5703 ^ 1'b0 ;
  assign n13265 = ( n1516 & n12403 ) | ( n1516 & n13264 ) | ( n12403 & n13264 ) ;
  assign n13266 = n13265 ^ n6651 ^ 1'b0 ;
  assign n13267 = n7829 & n13266 ;
  assign n13268 = n3494 & ~n5987 ;
  assign n13269 = ~n12968 & n13268 ;
  assign n13273 = n3032 ^ n2921 ^ n2740 ;
  assign n13270 = n2272 ^ n1764 ^ 1'b0 ;
  assign n13271 = n7035 & n13270 ;
  assign n13272 = ( ~n6150 & n6187 ) | ( ~n6150 & n13271 ) | ( n6187 & n13271 ) ;
  assign n13274 = n13273 ^ n13272 ^ 1'b0 ;
  assign n13275 = n12437 ^ n4476 ^ 1'b0 ;
  assign n13276 = ~n5764 & n13275 ;
  assign n13277 = n1084 & n10643 ;
  assign n13278 = n13277 ^ n10116 ^ 1'b0 ;
  assign n13279 = ( n13109 & ~n13276 ) | ( n13109 & n13278 ) | ( ~n13276 & n13278 ) ;
  assign n13282 = n2721 ^ n704 ^ 1'b0 ;
  assign n13280 = n8662 ^ n5033 ^ 1'b0 ;
  assign n13281 = n7179 | n13280 ;
  assign n13283 = n13282 ^ n13281 ^ 1'b0 ;
  assign n13286 = n9769 ^ n3548 ^ 1'b0 ;
  assign n13284 = n4195 & n6872 ;
  assign n13285 = n13284 ^ n5484 ^ 1'b0 ;
  assign n13287 = n13286 ^ n13285 ^ n11051 ;
  assign n13290 = ( n1895 & ~n2645 ) | ( n1895 & n2930 ) | ( ~n2645 & n2930 ) ;
  assign n13291 = n887 & n13290 ;
  assign n13288 = n10078 ^ n8955 ^ 1'b0 ;
  assign n13289 = n7388 | n13288 ;
  assign n13292 = n13291 ^ n13289 ^ 1'b0 ;
  assign n13293 = ~n8461 & n9985 ;
  assign n13295 = ~n4653 & n8853 ;
  assign n13296 = ~n4032 & n13295 ;
  assign n13294 = ~n5360 & n8486 ;
  assign n13297 = n13296 ^ n13294 ^ 1'b0 ;
  assign n13298 = n1236 & ~n7916 ;
  assign n13299 = n8658 ^ n8088 ^ 1'b0 ;
  assign n13300 = n10883 ^ n9078 ^ 1'b0 ;
  assign n13301 = n5890 | n6154 ;
  assign n13302 = n13301 ^ n941 ^ 1'b0 ;
  assign n13303 = ( n4342 & ~n6232 ) | ( n4342 & n13302 ) | ( ~n6232 & n13302 ) ;
  assign n13304 = n10519 ^ n8177 ^ 1'b0 ;
  assign n13307 = n3274 & n3771 ;
  assign n13308 = n1485 & n13307 ;
  assign n13309 = n7971 | n13308 ;
  assign n13310 = n13309 ^ n1560 ^ 1'b0 ;
  assign n13311 = n13310 ^ n7409 ^ n4864 ;
  assign n13305 = n6143 ^ n5907 ^ 1'b0 ;
  assign n13306 = n5561 & n13305 ;
  assign n13312 = n13311 ^ n13306 ^ n4866 ;
  assign n13313 = ( n1489 & n2598 ) | ( n1489 & ~n4144 ) | ( n2598 & ~n4144 ) ;
  assign n13314 = n6103 | n13313 ;
  assign n13315 = ( n11400 & n12439 ) | ( n11400 & ~n13314 ) | ( n12439 & ~n13314 ) ;
  assign n13316 = n9023 ^ x51 ^ 1'b0 ;
  assign n13317 = ~n10752 & n13316 ;
  assign n13318 = n4730 ^ n668 ^ 1'b0 ;
  assign n13319 = n13318 ^ n11329 ^ 1'b0 ;
  assign n13320 = ~n9927 & n13319 ;
  assign n13321 = n3908 & n13320 ;
  assign n13322 = n12610 ^ n4654 ^ n2100 ;
  assign n13323 = ( n1324 & n4113 ) | ( n1324 & ~n12193 ) | ( n4113 & ~n12193 ) ;
  assign n13324 = n13322 & ~n13323 ;
  assign n13325 = n4320 ^ n1327 ^ 1'b0 ;
  assign n13326 = n13325 ^ n5552 ^ 1'b0 ;
  assign n13327 = n8097 ^ n744 ^ 1'b0 ;
  assign n13328 = n10795 ^ n748 ^ 1'b0 ;
  assign n13329 = n4204 & n13328 ;
  assign n13330 = n11870 & ~n12846 ;
  assign n13338 = n1839 | n6216 ;
  assign n13339 = n1959 & ~n13338 ;
  assign n13336 = ( ~n606 & n3771 ) | ( ~n606 & n8335 ) | ( n3771 & n8335 ) ;
  assign n13337 = ~n7771 & n13336 ;
  assign n13340 = n13339 ^ n13337 ^ n5183 ;
  assign n13341 = n13340 ^ n3072 ^ 1'b0 ;
  assign n13331 = n4277 ^ n1398 ^ 1'b0 ;
  assign n13332 = n1685 & ~n13331 ;
  assign n13333 = ~n4712 & n13332 ;
  assign n13334 = n13333 ^ n8161 ^ 1'b0 ;
  assign n13335 = n10133 & n13334 ;
  assign n13342 = n13341 ^ n13335 ^ 1'b0 ;
  assign n13343 = n10715 & ~n12728 ;
  assign n13344 = n8662 & n13343 ;
  assign n13345 = ~n1817 & n12807 ;
  assign n13346 = n13345 ^ n744 ^ 1'b0 ;
  assign n13347 = n1222 & ~n13346 ;
  assign n13348 = n4914 ^ n2068 ^ 1'b0 ;
  assign n13349 = n6744 & n13348 ;
  assign n13350 = n1943 ^ n1720 ^ 1'b0 ;
  assign n13351 = n6087 & n13350 ;
  assign n13352 = n13349 & n13351 ;
  assign n13353 = ~n7297 & n13352 ;
  assign n13354 = n9388 & n9731 ;
  assign n13355 = n13353 & n13354 ;
  assign n13356 = n4650 & ~n6798 ;
  assign n13357 = ( ~n10224 & n12626 ) | ( ~n10224 & n13356 ) | ( n12626 & n13356 ) ;
  assign n13358 = ~n9212 & n13357 ;
  assign n13362 = ( n617 & ~n992 ) | ( n617 & n2163 ) | ( ~n992 & n2163 ) ;
  assign n13360 = n9212 ^ n4687 ^ n3884 ;
  assign n13361 = n13360 ^ n318 ^ 1'b0 ;
  assign n13359 = n4923 & ~n8875 ;
  assign n13363 = n13362 ^ n13361 ^ n13359 ;
  assign n13364 = n2102 & ~n3572 ;
  assign n13365 = n12893 & n13364 ;
  assign n13366 = ~x42 & n13365 ;
  assign n13368 = ( ~n2554 & n2947 ) | ( ~n2554 & n7689 ) | ( n2947 & n7689 ) ;
  assign n13369 = n2179 | n13368 ;
  assign n13370 = n13369 ^ n11163 ^ 1'b0 ;
  assign n13367 = ( n1199 & n1903 ) | ( n1199 & ~n4802 ) | ( n1903 & ~n4802 ) ;
  assign n13371 = n13370 ^ n13367 ^ 1'b0 ;
  assign n13372 = n9710 & n13371 ;
  assign n13375 = n6630 ^ n866 ^ 1'b0 ;
  assign n13373 = ~n7856 & n8788 ;
  assign n13374 = ~n5880 & n13373 ;
  assign n13376 = n13375 ^ n13374 ^ n1121 ;
  assign n13378 = n1137 ^ n732 ^ 1'b0 ;
  assign n13377 = ~n2318 & n5620 ;
  assign n13379 = n13378 ^ n13377 ^ 1'b0 ;
  assign n13380 = ( ~n579 & n5577 ) | ( ~n579 & n8673 ) | ( n5577 & n8673 ) ;
  assign n13381 = n3923 & n13380 ;
  assign n13382 = n13381 ^ n5110 ^ 1'b0 ;
  assign n13383 = n6422 ^ n667 ^ 1'b0 ;
  assign n13384 = n1851 | n11570 ;
  assign n13385 = n6645 ^ n2059 ^ 1'b0 ;
  assign n13386 = n4163 | n13385 ;
  assign n13387 = n7137 ^ n3775 ^ 1'b0 ;
  assign n13388 = ~n1795 & n13387 ;
  assign n13389 = n13388 ^ n9609 ^ 1'b0 ;
  assign n13390 = ~n4863 & n13389 ;
  assign n13391 = n2976 & n13390 ;
  assign n13392 = ( ~n6519 & n8787 ) | ( ~n6519 & n13391 ) | ( n8787 & n13391 ) ;
  assign n13393 = n7204 | n11586 ;
  assign n13394 = n13393 ^ n4190 ^ 1'b0 ;
  assign n13395 = n7137 ^ n6361 ^ n3120 ;
  assign n13396 = n13395 ^ n6744 ^ 1'b0 ;
  assign n13397 = n1976 | n4712 ;
  assign n13398 = n5164 ^ n3907 ^ 1'b0 ;
  assign n13399 = n13398 ^ n8744 ^ n4646 ;
  assign n13400 = n2528 & n3731 ;
  assign n13401 = n13400 ^ n7862 ^ 1'b0 ;
  assign n13402 = ( n257 & n7610 ) | ( n257 & ~n13401 ) | ( n7610 & ~n13401 ) ;
  assign n13403 = n13402 ^ n12553 ^ 1'b0 ;
  assign n13404 = n6507 ^ n784 ^ 1'b0 ;
  assign n13405 = n5670 & ~n13404 ;
  assign n13406 = n13405 ^ n2686 ^ 1'b0 ;
  assign n13407 = n3642 & n13406 ;
  assign n13408 = ~n5669 & n13407 ;
  assign n13413 = ~n3486 & n4294 ;
  assign n13411 = x89 & n1343 ;
  assign n13412 = n779 & n13411 ;
  assign n13414 = n13413 ^ n13412 ^ n1840 ;
  assign n13415 = n2679 & n13414 ;
  assign n13416 = n9651 & n13415 ;
  assign n13409 = n9528 ^ n6818 ^ 1'b0 ;
  assign n13410 = n13409 ^ n1895 ^ n801 ;
  assign n13417 = n13416 ^ n13410 ^ 1'b0 ;
  assign n13418 = ~n9599 & n13417 ;
  assign n13419 = ~n3237 & n13418 ;
  assign n13420 = n12703 ^ n6060 ^ 1'b0 ;
  assign n13421 = n5347 & n7054 ;
  assign n13422 = ( ~n4149 & n4267 ) | ( ~n4149 & n7905 ) | ( n4267 & n7905 ) ;
  assign n13423 = n13422 ^ n9033 ^ 1'b0 ;
  assign n13424 = n2879 ^ n1305 ^ 1'b0 ;
  assign n13425 = n295 | n13424 ;
  assign n13426 = n13425 ^ n3382 ^ n1266 ;
  assign n13427 = ~n5422 & n13426 ;
  assign n13428 = n2635 & n13336 ;
  assign n13429 = n13428 ^ n4124 ^ 1'b0 ;
  assign n13432 = n3265 ^ n2149 ^ 1'b0 ;
  assign n13433 = n4085 & n13432 ;
  assign n13434 = n13433 ^ n8119 ^ 1'b0 ;
  assign n13435 = n7945 | n13434 ;
  assign n13430 = n1700 | n4665 ;
  assign n13431 = ~n591 & n13430 ;
  assign n13436 = n13435 ^ n13431 ^ 1'b0 ;
  assign n13437 = n8327 ^ n5006 ^ 1'b0 ;
  assign n13438 = n8178 ^ n6285 ^ 1'b0 ;
  assign n13439 = n1086 | n7834 ;
  assign n13440 = n13438 & ~n13439 ;
  assign n13441 = ~n13437 & n13440 ;
  assign n13442 = n13441 ^ n6483 ^ n6271 ;
  assign n13443 = n4633 & ~n13442 ;
  assign n13444 = ( n8691 & ~n9538 ) | ( n8691 & n12554 ) | ( ~n9538 & n12554 ) ;
  assign n13445 = ~n11692 & n13444 ;
  assign n13446 = ( ~n2167 & n5223 ) | ( ~n2167 & n7750 ) | ( n5223 & n7750 ) ;
  assign n13447 = ~n11579 & n13446 ;
  assign n13448 = n13447 ^ n11206 ^ 1'b0 ;
  assign n13449 = n8523 & ~n11389 ;
  assign n13450 = n5867 & n11015 ;
  assign n13451 = ~n4455 & n8265 ;
  assign n13452 = n7292 ^ n885 ^ 1'b0 ;
  assign n13453 = n13451 & ~n13452 ;
  assign n13455 = ~n1002 & n11958 ;
  assign n13454 = n593 | n13268 ;
  assign n13456 = n13455 ^ n13454 ^ 1'b0 ;
  assign n13457 = n880 & ~n8410 ;
  assign n13458 = n13457 ^ n6341 ^ n3212 ;
  assign n13459 = x106 | n319 ;
  assign n13460 = n8675 & ~n13459 ;
  assign n13461 = n13460 ^ n12587 ^ n5458 ;
  assign n13462 = n416 | n5168 ;
  assign n13463 = n6671 & ~n13462 ;
  assign n13464 = ~n10088 & n10969 ;
  assign n13465 = n13464 ^ n10881 ^ 1'b0 ;
  assign n13466 = n10005 & ~n13465 ;
  assign n13467 = n6695 ^ n2413 ^ 1'b0 ;
  assign n13468 = n13467 ^ n10460 ^ 1'b0 ;
  assign n13478 = n2099 ^ n1761 ^ 1'b0 ;
  assign n13472 = n4908 ^ n3056 ^ n831 ;
  assign n13473 = n7771 ^ n2657 ^ 1'b0 ;
  assign n13474 = ~n3353 & n10080 ;
  assign n13475 = ~n4298 & n13474 ;
  assign n13476 = ( ~n13472 & n13473 ) | ( ~n13472 & n13475 ) | ( n13473 & n13475 ) ;
  assign n13477 = n13476 ^ n12031 ^ n599 ;
  assign n13469 = ( n8022 & n9160 ) | ( n8022 & n10777 ) | ( n9160 & n10777 ) ;
  assign n13470 = ~n1776 & n6498 ;
  assign n13471 = ~n13469 & n13470 ;
  assign n13479 = n13478 ^ n13477 ^ n13471 ;
  assign n13480 = n3050 ^ n2952 ^ 1'b0 ;
  assign n13481 = n9424 ^ n490 ^ 1'b0 ;
  assign n13482 = n13480 | n13481 ;
  assign n13483 = n13482 ^ n12703 ^ 1'b0 ;
  assign n13484 = n7965 ^ n7182 ^ n2604 ;
  assign n13485 = n7116 | n13484 ;
  assign n13486 = n13485 ^ n9070 ^ 1'b0 ;
  assign n13487 = n181 & n5187 ;
  assign n13488 = n13487 ^ n3943 ^ 1'b0 ;
  assign n13489 = n10304 ^ n7543 ^ 1'b0 ;
  assign n13490 = n13488 | n13489 ;
  assign n13491 = n3011 & ~n13490 ;
  assign n13492 = n701 & n13491 ;
  assign n13493 = n7245 ^ n4013 ^ 1'b0 ;
  assign n13494 = n7793 & n13493 ;
  assign n13495 = n13494 ^ n6138 ^ n4492 ;
  assign n13496 = ~n1660 & n7420 ;
  assign n13497 = n13496 ^ n9579 ^ x0 ;
  assign n13498 = ~n4940 & n13497 ;
  assign n13499 = ~n8056 & n13498 ;
  assign n13500 = n12382 ^ n10235 ^ 1'b0 ;
  assign n13501 = ~n13499 & n13500 ;
  assign n13502 = n4809 ^ n2519 ^ 1'b0 ;
  assign n13503 = n3608 & ~n13502 ;
  assign n13504 = n5773 ^ n1008 ^ 1'b0 ;
  assign n13505 = n700 | n13504 ;
  assign n13506 = n10515 | n13505 ;
  assign n13507 = n13503 & ~n13506 ;
  assign n13508 = n3642 ^ n2699 ^ n2645 ;
  assign n13509 = n13508 ^ n247 ^ 1'b0 ;
  assign n13510 = n1230 & ~n13509 ;
  assign n13511 = n3731 & n13510 ;
  assign n13512 = n13511 ^ n2638 ^ 1'b0 ;
  assign n13513 = ~n7766 & n11468 ;
  assign n13514 = n13513 ^ n3173 ^ 1'b0 ;
  assign n13515 = n1334 ^ n844 ^ 1'b0 ;
  assign n13516 = n9089 & n13515 ;
  assign n13517 = ~n13514 & n13516 ;
  assign n13518 = n1294 ^ n1049 ^ 1'b0 ;
  assign n13519 = ~n1992 & n13518 ;
  assign n13520 = n10699 & n13519 ;
  assign n13521 = n13517 & n13520 ;
  assign n13522 = ~n584 & n11954 ;
  assign n13523 = n13521 & ~n13522 ;
  assign n13524 = n7932 ^ n7482 ^ 1'b0 ;
  assign n13525 = ~n3522 & n13524 ;
  assign n13526 = ~n6915 & n13525 ;
  assign n13527 = ~n6003 & n13526 ;
  assign n13528 = n4378 & n7152 ;
  assign n13529 = n5351 ^ n3428 ^ 1'b0 ;
  assign n13530 = n13528 & ~n13529 ;
  assign n13531 = n5817 ^ n2653 ^ 1'b0 ;
  assign n13532 = n2507 & n13531 ;
  assign n13533 = n13532 ^ n2971 ^ 1'b0 ;
  assign n13534 = n13533 ^ n9427 ^ 1'b0 ;
  assign n13536 = ( n298 & n914 ) | ( n298 & n2435 ) | ( n914 & n2435 ) ;
  assign n13535 = n1895 & n12540 ;
  assign n13537 = n13536 ^ n13535 ^ n5599 ;
  assign n13538 = n9995 ^ n2660 ^ 1'b0 ;
  assign n13544 = n9921 ^ x39 ^ 1'b0 ;
  assign n13541 = n10903 ^ n6200 ^ 1'b0 ;
  assign n13539 = n5008 ^ n4434 ^ n2638 ;
  assign n13540 = n13539 ^ n6243 ^ n3661 ;
  assign n13542 = n13541 ^ n13540 ^ n2740 ;
  assign n13543 = n13542 ^ n4343 ^ n1381 ;
  assign n13545 = n13544 ^ n13543 ^ 1'b0 ;
  assign n13546 = n11354 | n13545 ;
  assign n13547 = ( ~n2042 & n10056 ) | ( ~n2042 & n13141 ) | ( n10056 & n13141 ) ;
  assign n13548 = n9300 & n11069 ;
  assign n13549 = n4132 ^ n1888 ^ n831 ;
  assign n13550 = n1365 | n13549 ;
  assign n13551 = n2905 | n5305 ;
  assign n13552 = n4798 & ~n13551 ;
  assign n13553 = n13552 ^ n9759 ^ n6274 ;
  assign n13554 = n8626 ^ n8487 ^ 1'b0 ;
  assign n13555 = n13553 | n13554 ;
  assign n13556 = n3118 ^ n2278 ^ 1'b0 ;
  assign n13557 = n10275 | n13556 ;
  assign n13558 = n5788 & ~n13557 ;
  assign n13559 = ~n9105 & n12412 ;
  assign n13560 = n4983 & n13559 ;
  assign n13561 = n13560 ^ n4054 ^ 1'b0 ;
  assign n13562 = n2715 | n13561 ;
  assign n13563 = n6628 & ~n13562 ;
  assign n13564 = ~n1521 & n6186 ;
  assign n13565 = n8845 ^ n935 ^ 1'b0 ;
  assign n13566 = ( ~n3533 & n13564 ) | ( ~n3533 & n13565 ) | ( n13564 & n13565 ) ;
  assign n13567 = n6705 ^ n5540 ^ 1'b0 ;
  assign n13568 = n940 | n13567 ;
  assign n13569 = n13568 ^ n9421 ^ 1'b0 ;
  assign n13570 = n13566 | n13569 ;
  assign n13572 = n1046 | n4431 ;
  assign n13573 = n13572 ^ n1594 ^ 1'b0 ;
  assign n13571 = ~n7059 & n10501 ;
  assign n13574 = n13573 ^ n13571 ^ 1'b0 ;
  assign n13575 = n9955 ^ n7911 ^ n7369 ;
  assign n13576 = ( n1759 & n2886 ) | ( n1759 & n6452 ) | ( n2886 & n6452 ) ;
  assign n13577 = n6633 & n13576 ;
  assign n13578 = ( n3758 & ~n13575 ) | ( n3758 & n13577 ) | ( ~n13575 & n13577 ) ;
  assign n13579 = n5939 ^ n2450 ^ n1470 ;
  assign n13580 = ~n12452 & n13283 ;
  assign n13581 = n9709 ^ n131 ^ 1'b0 ;
  assign n13582 = x106 & n13581 ;
  assign n13583 = x6 & n818 ;
  assign n13584 = n13583 ^ n867 ^ 1'b0 ;
  assign n13585 = n8543 & ~n13584 ;
  assign n13586 = n7839 & n13585 ;
  assign n13587 = n13586 ^ n12325 ^ 1'b0 ;
  assign n13588 = ~n13582 & n13587 ;
  assign n13589 = n9135 ^ n5801 ^ 1'b0 ;
  assign n13590 = n4173 ^ n3180 ^ 1'b0 ;
  assign n13591 = n870 & ~n13590 ;
  assign n13592 = n10815 ^ n2811 ^ 1'b0 ;
  assign n13593 = n11007 & n13592 ;
  assign n13594 = ( n5149 & n6286 ) | ( n5149 & ~n11232 ) | ( n6286 & ~n11232 ) ;
  assign n13595 = ( ~n2582 & n8801 ) | ( ~n2582 & n13594 ) | ( n8801 & n13594 ) ;
  assign n13596 = n11694 ^ x74 ^ 1'b0 ;
  assign n13597 = n3199 & ~n4563 ;
  assign n13598 = n7030 & n10117 ;
  assign n13599 = n10992 ^ n10520 ^ 1'b0 ;
  assign n13600 = n1985 | n8840 ;
  assign n13601 = n10045 ^ n9392 ^ 1'b0 ;
  assign n13602 = n13600 | n13601 ;
  assign n13603 = n10567 ^ n4182 ^ 1'b0 ;
  assign n13604 = n2635 & n5032 ;
  assign n13606 = n3262 ^ n1532 ^ 1'b0 ;
  assign n13605 = n8712 ^ n7760 ^ 1'b0 ;
  assign n13607 = n13606 ^ n13605 ^ 1'b0 ;
  assign n13608 = n13604 | n13607 ;
  assign n13609 = ~n5224 & n6143 ;
  assign n13610 = n13609 ^ n2028 ^ 1'b0 ;
  assign n13611 = n1257 & n11430 ;
  assign n13612 = n13611 ^ n3187 ^ 1'b0 ;
  assign n13613 = n8359 | n13612 ;
  assign n13615 = ( n1639 & n4521 ) | ( n1639 & n6591 ) | ( n4521 & n6591 ) ;
  assign n13614 = ~x13 & n7455 ;
  assign n13616 = n13615 ^ n13614 ^ 1'b0 ;
  assign n13617 = ~n2660 & n13616 ;
  assign n13619 = n1256 | n9601 ;
  assign n13620 = n351 & ~n13619 ;
  assign n13618 = ( ~n4182 & n5928 ) | ( ~n4182 & n9042 ) | ( n5928 & n9042 ) ;
  assign n13621 = n13620 ^ n13618 ^ 1'b0 ;
  assign n13622 = n13621 ^ n6701 ^ n4753 ;
  assign n13623 = n4221 ^ n1542 ^ n905 ;
  assign n13624 = n1345 | n13623 ;
  assign n13625 = ( n4830 & n8283 ) | ( n4830 & n13460 ) | ( n8283 & n13460 ) ;
  assign n13626 = ~n2288 & n13625 ;
  assign n13627 = n4069 ^ n3139 ^ n210 ;
  assign n13628 = n8778 & n13627 ;
  assign n13629 = ( ~n3177 & n13626 ) | ( ~n3177 & n13628 ) | ( n13626 & n13628 ) ;
  assign n13630 = x78 & n5850 ;
  assign n13631 = n10116 & n13630 ;
  assign n13632 = ~n2863 & n5921 ;
  assign n13633 = n2408 & ~n13632 ;
  assign n13634 = n13631 & n13633 ;
  assign n13635 = n8253 | n11134 ;
  assign n13636 = n4235 | n7923 ;
  assign n13637 = n5868 ^ n5283 ^ 1'b0 ;
  assign n13638 = n3953 & n12734 ;
  assign n13639 = n7871 & ~n13638 ;
  assign n13640 = ~n10925 & n13639 ;
  assign n13642 = n1953 | n10531 ;
  assign n13643 = n10348 & n13642 ;
  assign n13641 = n3726 & ~n9345 ;
  assign n13644 = n13643 ^ n13641 ^ 1'b0 ;
  assign n13645 = n12628 ^ n11560 ^ n551 ;
  assign n13646 = n5720 & ~n13645 ;
  assign n13647 = n2435 ^ n1898 ^ 1'b0 ;
  assign n13648 = n3046 ^ n828 ^ 1'b0 ;
  assign n13649 = n11460 & n13648 ;
  assign n13650 = ( n2738 & n7038 ) | ( n2738 & ~n8936 ) | ( n7038 & ~n8936 ) ;
  assign n13652 = n5291 | n11368 ;
  assign n13653 = ( n4247 & n6928 ) | ( n4247 & n13652 ) | ( n6928 & n13652 ) ;
  assign n13651 = n3530 | n6976 ;
  assign n13654 = n13653 ^ n13651 ^ 1'b0 ;
  assign n13655 = ( n10165 & n13650 ) | ( n10165 & ~n13654 ) | ( n13650 & ~n13654 ) ;
  assign n13660 = n3564 | n5804 ;
  assign n13657 = n3196 ^ n1853 ^ 1'b0 ;
  assign n13658 = x25 & n13657 ;
  assign n13656 = n4159 & ~n4415 ;
  assign n13659 = n13658 ^ n13656 ^ 1'b0 ;
  assign n13661 = n13660 ^ n13659 ^ n968 ;
  assign n13665 = n9427 ^ n1355 ^ 1'b0 ;
  assign n13662 = n6785 & n9688 ;
  assign n13663 = ~n1020 & n13662 ;
  assign n13664 = n10643 & ~n13663 ;
  assign n13666 = n13665 ^ n13664 ^ 1'b0 ;
  assign n13667 = n2000 & n13666 ;
  assign n13668 = ~n5752 & n13667 ;
  assign n13669 = n2155 | n2200 ;
  assign n13670 = n13669 ^ n139 ^ 1'b0 ;
  assign n13671 = n199 & n4170 ;
  assign n13672 = ~n13670 & n13671 ;
  assign n13673 = n10784 & n13672 ;
  assign n13674 = n1802 & ~n3561 ;
  assign n13675 = n13674 ^ n3819 ^ 1'b0 ;
  assign n13676 = n9883 ^ n8575 ^ 1'b0 ;
  assign n13677 = n1933 & n8507 ;
  assign n13678 = ~n6811 & n13677 ;
  assign n13679 = n7750 ^ n6191 ^ 1'b0 ;
  assign n13680 = ( n3371 & ~n3828 ) | ( n3371 & n13679 ) | ( ~n3828 & n13679 ) ;
  assign n13681 = n6415 & n6645 ;
  assign n13682 = n13681 ^ n8020 ^ 1'b0 ;
  assign n13683 = n1739 | n3506 ;
  assign n13684 = n10833 & ~n13683 ;
  assign n13685 = n13684 ^ n11891 ^ 1'b0 ;
  assign n13686 = n2822 & n13685 ;
  assign n13687 = n10429 ^ n5599 ^ 1'b0 ;
  assign n13688 = n1812 & n13687 ;
  assign n13689 = n12619 ^ n6591 ^ n432 ;
  assign n13690 = n12358 ^ n351 ^ 1'b0 ;
  assign n13691 = ~n5885 & n9131 ;
  assign n13692 = n2150 ^ n1691 ^ 1'b0 ;
  assign n13693 = n9445 | n13692 ;
  assign n13694 = ( n855 & n3878 ) | ( n855 & ~n7906 ) | ( n3878 & ~n7906 ) ;
  assign n13695 = ( n13691 & n13693 ) | ( n13691 & ~n13694 ) | ( n13693 & ~n13694 ) ;
  assign n13696 = ~n2898 & n4204 ;
  assign n13697 = n3160 ^ x78 ^ 1'b0 ;
  assign n13698 = ~n13696 & n13697 ;
  assign n13705 = n6042 & n7121 ;
  assign n13699 = n6838 ^ n4498 ^ 1'b0 ;
  assign n13700 = n7064 ^ n3302 ^ n2411 ;
  assign n13701 = n10440 & ~n13700 ;
  assign n13702 = n8846 & n13701 ;
  assign n13703 = n5974 | n13702 ;
  assign n13704 = n13699 | n13703 ;
  assign n13706 = n13705 ^ n13704 ^ n2510 ;
  assign n13707 = n6288 ^ n5680 ^ n1190 ;
  assign n13708 = ( n7287 & ~n11514 ) | ( n7287 & n13707 ) | ( ~n11514 & n13707 ) ;
  assign n13710 = n5741 ^ n2070 ^ 1'b0 ;
  assign n13709 = n1233 ^ n710 ^ 1'b0 ;
  assign n13711 = n13710 ^ n13709 ^ 1'b0 ;
  assign n13712 = ( n7116 & n12410 ) | ( n7116 & ~n13711 ) | ( n12410 & ~n13711 ) ;
  assign n13713 = n2198 & n11998 ;
  assign n13714 = ( n795 & ~n7266 ) | ( n795 & n7349 ) | ( ~n7266 & n7349 ) ;
  assign n13715 = n13714 ^ n3486 ^ 1'b0 ;
  assign n13716 = n9465 & n13715 ;
  assign n13717 = ~n6111 & n8458 ;
  assign n13718 = n13717 ^ n9760 ^ 1'b0 ;
  assign n13722 = n8969 & ~n11763 ;
  assign n13723 = n13722 ^ x12 ^ 1'b0 ;
  assign n13724 = n13723 ^ n4054 ^ n3318 ;
  assign n13719 = n11653 ^ n6271 ^ 1'b0 ;
  assign n13720 = n12852 ^ n2002 ^ 1'b0 ;
  assign n13721 = n13719 | n13720 ;
  assign n13725 = n13724 ^ n13721 ^ 1'b0 ;
  assign n13726 = n13718 & n13725 ;
  assign n13727 = n3228 ^ n1192 ^ n216 ;
  assign n13728 = n11294 ^ n285 ^ 1'b0 ;
  assign n13729 = n13727 & n13728 ;
  assign n13730 = ~n10883 & n13729 ;
  assign n13731 = n3310 & n13730 ;
  assign n13732 = ( n259 & n1257 ) | ( n259 & n7977 ) | ( n1257 & n7977 ) ;
  assign n13733 = n2601 & n6845 ;
  assign n13734 = n13733 ^ n4191 ^ 1'b0 ;
  assign n13735 = n13732 & ~n13734 ;
  assign n13736 = n368 & n13326 ;
  assign n13737 = ~n1720 & n13736 ;
  assign n13738 = n825 & ~n1800 ;
  assign n13739 = n7663 ^ n3660 ^ n2338 ;
  assign n13740 = n13739 ^ n10184 ^ 1'b0 ;
  assign n13741 = n5936 | n13740 ;
  assign n13742 = n13741 ^ n843 ^ 1'b0 ;
  assign n13743 = ( n4570 & n13738 ) | ( n4570 & ~n13742 ) | ( n13738 & ~n13742 ) ;
  assign n13744 = n11115 ^ n7241 ^ 1'b0 ;
  assign n13745 = ~n4859 & n11616 ;
  assign n13746 = n13745 ^ n12318 ^ 1'b0 ;
  assign n13747 = n4090 & ~n13746 ;
  assign n13748 = n2554 & ~n9121 ;
  assign n13749 = ~n5297 & n13748 ;
  assign n13750 = n10972 | n13749 ;
  assign n13751 = n7546 ^ n6938 ^ 1'b0 ;
  assign n13752 = ( ~n781 & n13750 ) | ( ~n781 & n13751 ) | ( n13750 & n13751 ) ;
  assign n13753 = n7604 ^ n6855 ^ n1797 ;
  assign n13754 = n10383 ^ n3739 ^ n1772 ;
  assign n13755 = ( n6365 & n10833 ) | ( n6365 & n13754 ) | ( n10833 & n13754 ) ;
  assign n13756 = n670 & ~n5393 ;
  assign n13757 = ~n2723 & n7030 ;
  assign n13758 = n13756 & n13757 ;
  assign n13759 = n13758 ^ n9968 ^ 1'b0 ;
  assign n13760 = n13755 & n13759 ;
  assign n13761 = ( n1215 & ~n3044 ) | ( n1215 & n10804 ) | ( ~n3044 & n10804 ) ;
  assign n13762 = ~n8651 & n13761 ;
  assign n13763 = n1767 & n13762 ;
  assign n13764 = n13763 ^ n3070 ^ 1'b0 ;
  assign n13765 = n232 & n710 ;
  assign n13766 = n13765 ^ n8255 ^ 1'b0 ;
  assign n13767 = ~n1452 & n7405 ;
  assign n13768 = n13767 ^ n12127 ^ 1'b0 ;
  assign n13769 = n11446 | n13768 ;
  assign n13770 = n1200 & n3237 ;
  assign n13771 = n13770 ^ n344 ^ 1'b0 ;
  assign n13772 = ( ~n4163 & n13769 ) | ( ~n4163 & n13771 ) | ( n13769 & n13771 ) ;
  assign n13773 = n2590 & ~n12009 ;
  assign n13774 = n12977 ^ n6772 ^ 1'b0 ;
  assign n13775 = ~n6764 & n13437 ;
  assign n13776 = n13545 ^ n3173 ^ 1'b0 ;
  assign n13777 = n13775 & n13776 ;
  assign n13778 = n13777 ^ n11310 ^ 1'b0 ;
  assign n13779 = n1710 | n12236 ;
  assign n13780 = n8256 & ~n10687 ;
  assign n13781 = n7204 | n13412 ;
  assign n13782 = n8278 | n13781 ;
  assign n13783 = ( n12452 & n13195 ) | ( n12452 & n13782 ) | ( n13195 & n13782 ) ;
  assign n13784 = ( ~n5332 & n5665 ) | ( ~n5332 & n7438 ) | ( n5665 & n7438 ) ;
  assign n13785 = n5093 | n10375 ;
  assign n13786 = n13430 | n13785 ;
  assign n13787 = n3652 & n8702 ;
  assign n13788 = n13115 & n13787 ;
  assign n13789 = n13788 ^ n872 ^ 1'b0 ;
  assign n13790 = n1928 | n13449 ;
  assign n13791 = n13790 ^ n708 ^ 1'b0 ;
  assign n13792 = n427 | n11999 ;
  assign n13793 = ( ~n4735 & n6743 ) | ( ~n4735 & n8444 ) | ( n6743 & n8444 ) ;
  assign n13794 = n13793 ^ n4511 ^ 1'b0 ;
  assign n13795 = n1649 & n13794 ;
  assign n13796 = n13795 ^ n2628 ^ 1'b0 ;
  assign n13797 = ( n917 & n3396 ) | ( n917 & ~n13796 ) | ( n3396 & ~n13796 ) ;
  assign n13798 = n4364 ^ n2760 ^ 1'b0 ;
  assign n13799 = ~n3217 & n13798 ;
  assign n13800 = n9742 ^ n7274 ^ 1'b0 ;
  assign n13801 = n13799 & ~n13800 ;
  assign n13802 = n13801 ^ n9455 ^ n6381 ;
  assign n13803 = n4781 & ~n4958 ;
  assign n13804 = n7939 & n13803 ;
  assign n13805 = n12891 ^ n8047 ^ 1'b0 ;
  assign n13806 = n12681 & ~n13805 ;
  assign n13807 = ( ~n2797 & n2897 ) | ( ~n2797 & n4512 ) | ( n2897 & n4512 ) ;
  assign n13808 = ~n1000 & n13807 ;
  assign n13809 = n13808 ^ n3559 ^ n773 ;
  assign n13810 = n2607 | n4632 ;
  assign n13811 = n12778 ^ n1871 ^ 1'b0 ;
  assign n13812 = n11155 & ~n13811 ;
  assign n13813 = n2580 ^ n1818 ^ 1'b0 ;
  assign n13814 = ~n2074 & n13813 ;
  assign n13815 = n9992 & ~n13494 ;
  assign n13816 = n2203 ^ n2195 ^ n843 ;
  assign n13823 = n7590 & ~n8018 ;
  assign n13824 = ( n3172 & n12881 ) | ( n3172 & ~n13823 ) | ( n12881 & ~n13823 ) ;
  assign n13819 = n4193 ^ n2494 ^ 1'b0 ;
  assign n13820 = n13819 ^ n3076 ^ 1'b0 ;
  assign n13821 = n4029 & ~n13820 ;
  assign n13817 = ( ~n9971 & n11148 ) | ( ~n9971 & n11357 ) | ( n11148 & n11357 ) ;
  assign n13818 = ~n6655 & n13817 ;
  assign n13822 = n13821 ^ n13818 ^ 1'b0 ;
  assign n13825 = n13824 ^ n13822 ^ n6158 ;
  assign n13826 = n7832 & ~n9655 ;
  assign n13827 = n5123 & n8783 ;
  assign n13828 = n13827 ^ n12875 ^ n6551 ;
  assign n13829 = n2260 ^ n545 ^ 1'b0 ;
  assign n13830 = n416 | n13829 ;
  assign n13831 = n2361 | n13830 ;
  assign n13832 = n13828 & n13831 ;
  assign n13833 = n138 | n3279 ;
  assign n13834 = n4461 & n4641 ;
  assign n13835 = n4572 & n13834 ;
  assign n13836 = n13835 ^ n7740 ^ 1'b0 ;
  assign n13837 = n5958 | n13836 ;
  assign n13838 = n6986 & n13205 ;
  assign n13839 = ~n4895 & n13838 ;
  assign n13840 = n13839 ^ n8833 ^ n2187 ;
  assign n13841 = n3975 ^ n2517 ^ n293 ;
  assign n13842 = x119 & ~n8482 ;
  assign n13843 = n13842 ^ n5823 ^ 1'b0 ;
  assign n13844 = n7721 & n13843 ;
  assign n13845 = ~n13841 & n13844 ;
  assign n13846 = n9764 & n13845 ;
  assign n13847 = n3974 ^ n820 ^ 1'b0 ;
  assign n13848 = n4586 & n13847 ;
  assign n13849 = n3231 & n13848 ;
  assign n13853 = n2261 | n3160 ;
  assign n13850 = n693 | n11967 ;
  assign n13851 = n13019 ^ n1671 ^ 1'b0 ;
  assign n13852 = n13850 & n13851 ;
  assign n13854 = n13853 ^ n13852 ^ 1'b0 ;
  assign n13855 = n13854 ^ n11699 ^ n6810 ;
  assign n13859 = ~n2183 & n11833 ;
  assign n13856 = ( n3117 & ~n4219 ) | ( n3117 & n6131 ) | ( ~n4219 & n6131 ) ;
  assign n13857 = ( n5178 & n12050 ) | ( n5178 & ~n13856 ) | ( n12050 & ~n13856 ) ;
  assign n13858 = ~n2275 & n13857 ;
  assign n13860 = n13859 ^ n13858 ^ 1'b0 ;
  assign n13861 = n13860 ^ n8131 ^ n1715 ;
  assign n13862 = n8583 ^ n3574 ^ 1'b0 ;
  assign n13863 = ( n5956 & ~n6673 ) | ( n5956 & n13862 ) | ( ~n6673 & n13862 ) ;
  assign n13864 = n13292 & n13863 ;
  assign n13865 = n6601 ^ n358 ^ 1'b0 ;
  assign n13866 = n9623 | n13865 ;
  assign n13867 = n3741 & n10173 ;
  assign n13869 = n1548 ^ n589 ^ 1'b0 ;
  assign n13870 = n9616 & n10667 ;
  assign n13871 = n1818 & n13870 ;
  assign n13872 = n13869 & n13871 ;
  assign n13868 = n11055 ^ n10180 ^ n9247 ;
  assign n13873 = n13872 ^ n13868 ^ n9458 ;
  assign n13874 = n13873 ^ n13296 ^ 1'b0 ;
  assign n13875 = ~n8513 & n9456 ;
  assign n13876 = n10630 ^ n6407 ^ n3791 ;
  assign n13877 = n2783 ^ n1179 ^ 1'b0 ;
  assign n13878 = n4316 & n13877 ;
  assign n13879 = n13878 ^ n9090 ^ 1'b0 ;
  assign n13885 = n5080 & n6824 ;
  assign n13886 = ( n1383 & n7894 ) | ( n1383 & n13885 ) | ( n7894 & n13885 ) ;
  assign n13882 = n2984 ^ n2573 ^ 1'b0 ;
  assign n13880 = n2954 ^ n370 ^ 1'b0 ;
  assign n13881 = n12188 & n13880 ;
  assign n13883 = n13882 ^ n13881 ^ n13621 ;
  assign n13884 = ~n13437 & n13883 ;
  assign n13887 = n13886 ^ n13884 ^ 1'b0 ;
  assign n13889 = n927 | n1545 ;
  assign n13888 = n2371 | n7343 ;
  assign n13890 = n13889 ^ n13888 ^ 1'b0 ;
  assign n13896 = n7621 ^ n5259 ^ 1'b0 ;
  assign n13897 = n8510 & n13896 ;
  assign n13891 = n13152 ^ n1543 ^ 1'b0 ;
  assign n13892 = n261 & n13891 ;
  assign n13893 = ~n9157 & n13892 ;
  assign n13894 = n13893 ^ n923 ^ 1'b0 ;
  assign n13895 = n13894 ^ n11389 ^ n7170 ;
  assign n13898 = n13897 ^ n13895 ^ 1'b0 ;
  assign n13899 = ( n4044 & n13360 ) | ( n4044 & n13898 ) | ( n13360 & n13898 ) ;
  assign n13900 = ( n1392 & n2282 ) | ( n1392 & ~n9729 ) | ( n2282 & ~n9729 ) ;
  assign n13901 = ( n1556 & ~n1817 ) | ( n1556 & n6524 ) | ( ~n1817 & n6524 ) ;
  assign n13902 = n5546 & n9831 ;
  assign n13903 = n3720 | n13902 ;
  assign n13904 = n725 | n13903 ;
  assign n13905 = ~n13901 & n13904 ;
  assign n13906 = n13905 ^ n1035 ^ 1'b0 ;
  assign n13907 = n1552 | n10722 ;
  assign n13908 = n7670 ^ n1983 ^ 1'b0 ;
  assign n13909 = ~n1353 & n13908 ;
  assign n13910 = n13909 ^ n2419 ^ 1'b0 ;
  assign n13911 = n1342 | n1674 ;
  assign n13912 = n13910 & ~n13911 ;
  assign n13913 = ( n5138 & n10057 ) | ( n5138 & n13912 ) | ( n10057 & n13912 ) ;
  assign n13914 = n6380 ^ n4803 ^ n1150 ;
  assign n13915 = ( n3324 & n7082 ) | ( n3324 & n13914 ) | ( n7082 & n13914 ) ;
  assign n13916 = ~n3472 & n4664 ;
  assign n13917 = n1036 & n8875 ;
  assign n13918 = n13916 & n13917 ;
  assign n13919 = n968 & n6844 ;
  assign n13920 = n250 & ~n1473 ;
  assign n13921 = ~n6543 & n13414 ;
  assign n13922 = n3591 | n5956 ;
  assign n13923 = n13922 ^ n1353 ^ 1'b0 ;
  assign n13924 = ( ~n5594 & n13040 ) | ( ~n5594 & n13727 ) | ( n13040 & n13727 ) ;
  assign n13925 = n3348 | n13924 ;
  assign n13926 = n9648 ^ n3080 ^ 1'b0 ;
  assign n13927 = n13926 ^ n11916 ^ n1803 ;
  assign n13928 = n893 & ~n2862 ;
  assign n13929 = n12392 ^ n496 ^ 1'b0 ;
  assign n13930 = ( ~n2559 & n6591 ) | ( ~n2559 & n8957 ) | ( n6591 & n8957 ) ;
  assign n13931 = n509 & ~n9956 ;
  assign n13933 = ~n8829 & n10775 ;
  assign n13932 = n12636 ^ n5872 ^ 1'b0 ;
  assign n13934 = n13933 ^ n13932 ^ n9309 ;
  assign n13935 = n7274 ^ n2389 ^ 1'b0 ;
  assign n13936 = n5213 & ~n13935 ;
  assign n13937 = n6372 ^ n5807 ^ n1269 ;
  assign n13938 = n6772 ^ n6335 ^ 1'b0 ;
  assign n13939 = n5151 & n13938 ;
  assign n13940 = n7316 | n7593 ;
  assign n13941 = n10173 | n13940 ;
  assign n13942 = n13097 ^ n12366 ^ n10790 ;
  assign n13943 = n4271 ^ n608 ^ 1'b0 ;
  assign n13944 = n13943 ^ n5302 ^ n4795 ;
  assign n13945 = ( n3720 & n5178 ) | ( n3720 & ~n13944 ) | ( n5178 & ~n13944 ) ;
  assign n13946 = n8970 ^ x54 ^ 1'b0 ;
  assign n13947 = n13946 ^ n12563 ^ n4436 ;
  assign n13948 = ( n7425 & n13945 ) | ( n7425 & ~n13947 ) | ( n13945 & ~n13947 ) ;
  assign n13949 = n1758 ^ n1355 ^ 1'b0 ;
  assign n13950 = n3652 | n7462 ;
  assign n13951 = n13950 ^ n8367 ^ 1'b0 ;
  assign n13952 = ~n10343 & n13951 ;
  assign n13953 = n9223 & n13952 ;
  assign n13954 = n13953 ^ n866 ^ 1'b0 ;
  assign n13955 = n13949 | n13954 ;
  assign n13956 = n4901 ^ n1781 ^ 1'b0 ;
  assign n13957 = n6736 ^ n822 ^ 1'b0 ;
  assign n13958 = n13957 ^ n2514 ^ 1'b0 ;
  assign n13959 = n4223 | n13958 ;
  assign n13966 = ( ~n4281 & n6273 ) | ( ~n4281 & n7505 ) | ( n6273 & n7505 ) ;
  assign n13960 = n1853 | n6489 ;
  assign n13961 = n13960 ^ n7407 ^ 1'b0 ;
  assign n13962 = ( ~n975 & n7955 ) | ( ~n975 & n13961 ) | ( n7955 & n13961 ) ;
  assign n13963 = n2041 | n13962 ;
  assign n13964 = n13963 ^ n2761 ^ 1'b0 ;
  assign n13965 = n2197 & n13964 ;
  assign n13967 = n13966 ^ n13965 ^ 1'b0 ;
  assign n13968 = n356 & ~n13967 ;
  assign n13969 = n7079 ^ n1739 ^ 1'b0 ;
  assign n13970 = ~n12779 & n13969 ;
  assign n13971 = ~n4868 & n10991 ;
  assign n13972 = n2382 & n13971 ;
  assign n13973 = n13972 ^ n12402 ^ n4183 ;
  assign n13974 = ( n8735 & n13970 ) | ( n8735 & ~n13973 ) | ( n13970 & ~n13973 ) ;
  assign n13975 = n9231 & ~n13974 ;
  assign n13976 = n7841 & n13975 ;
  assign n13977 = n4958 ^ n3961 ^ 1'b0 ;
  assign n13978 = n1695 | n13977 ;
  assign n13979 = ~n9119 & n11377 ;
  assign n13980 = n8988 ^ n3093 ^ 1'b0 ;
  assign n13981 = n639 & n8807 ;
  assign n13982 = n6520 | n11842 ;
  assign n13983 = n1170 & ~n13982 ;
  assign n13984 = n9925 ^ n2358 ^ n234 ;
  assign n13985 = n3150 | n13984 ;
  assign n13986 = n13985 ^ n3915 ^ 1'b0 ;
  assign n13987 = ~n3722 & n13986 ;
  assign n13988 = n13987 ^ n214 ^ 1'b0 ;
  assign n13989 = ~n2728 & n5648 ;
  assign n13990 = ~n6410 & n13989 ;
  assign n13991 = ( n1719 & n4917 ) | ( n1719 & n12682 ) | ( n4917 & n12682 ) ;
  assign n13992 = n1784 & n6203 ;
  assign n13993 = n13992 ^ n8375 ^ 1'b0 ;
  assign n13994 = n6503 & ~n6976 ;
  assign n13995 = n13994 ^ n3158 ^ 1'b0 ;
  assign n13997 = ~n993 & n1067 ;
  assign n13996 = n1855 | n2340 ;
  assign n13998 = n13997 ^ n13996 ^ 1'b0 ;
  assign n13999 = n4934 | n13998 ;
  assign n14000 = ( n4701 & ~n11061 ) | ( n4701 & n13999 ) | ( ~n11061 & n13999 ) ;
  assign n14001 = ~n356 & n1689 ;
  assign n14002 = n14001 ^ n915 ^ 1'b0 ;
  assign n14003 = n13631 & ~n14002 ;
  assign n14004 = n5514 | n13813 ;
  assign n14005 = ( ~n1159 & n4152 ) | ( ~n1159 & n6420 ) | ( n4152 & n6420 ) ;
  assign n14006 = n4636 & ~n14005 ;
  assign n14007 = n4287 ^ n3417 ^ 1'b0 ;
  assign n14008 = n5297 & ~n14007 ;
  assign n14009 = ~n3271 & n8233 ;
  assign n14010 = n12882 ^ n4039 ^ 1'b0 ;
  assign n14011 = n1558 & n14010 ;
  assign n14012 = ( n4856 & n5337 ) | ( n4856 & ~n14011 ) | ( n5337 & ~n14011 ) ;
  assign n14013 = n14012 ^ n4952 ^ n990 ;
  assign n14014 = n10847 ^ n4475 ^ n1577 ;
  assign n14015 = n14014 ^ n4855 ^ n3634 ;
  assign n14016 = n14015 ^ n2488 ^ 1'b0 ;
  assign n14017 = ~n480 & n13761 ;
  assign n14018 = ~n13761 & n14017 ;
  assign n14019 = n6458 | n14018 ;
  assign n14020 = n14018 & ~n14019 ;
  assign n14021 = n14016 & ~n14020 ;
  assign n14022 = ~n14016 & n14021 ;
  assign n14023 = x92 & n9144 ;
  assign n14024 = n14023 ^ n2874 ^ 1'b0 ;
  assign n14025 = n2758 | n12085 ;
  assign n14026 = ( n2181 & n5135 ) | ( n2181 & n7401 ) | ( n5135 & n7401 ) ;
  assign n14027 = n14026 ^ n5864 ^ 1'b0 ;
  assign n14028 = n4964 & ~n8773 ;
  assign n14029 = n14028 ^ n7634 ^ 1'b0 ;
  assign n14030 = n12693 & ~n14029 ;
  assign n14031 = n12825 ^ n10504 ^ n4687 ;
  assign n14032 = n2597 | n7460 ;
  assign n14033 = n14032 ^ n13008 ^ 1'b0 ;
  assign n14034 = ~n1368 & n2455 ;
  assign n14035 = ~n12504 & n14034 ;
  assign n14036 = ( ~n3578 & n4647 ) | ( ~n3578 & n11998 ) | ( n4647 & n11998 ) ;
  assign n14037 = n1833 ^ n1133 ^ 1'b0 ;
  assign n14038 = ( n5393 & ~n10926 ) | ( n5393 & n14037 ) | ( ~n10926 & n14037 ) ;
  assign n14049 = n8060 & n9669 ;
  assign n14050 = n1353 & n14049 ;
  assign n14046 = n205 & ~n4653 ;
  assign n14047 = n6628 & n14046 ;
  assign n14048 = n14047 ^ n10558 ^ n4810 ;
  assign n14042 = n9504 ^ n6404 ^ n3491 ;
  assign n14039 = n2282 | n9014 ;
  assign n14040 = n11734 & ~n14039 ;
  assign n14041 = n14040 ^ n421 ^ 1'b0 ;
  assign n14043 = n14042 ^ n14041 ^ 1'b0 ;
  assign n14044 = n11685 | n14043 ;
  assign n14045 = n14044 ^ n4915 ^ n1390 ;
  assign n14051 = n14050 ^ n14048 ^ n14045 ;
  assign n14052 = n7929 & ~n10309 ;
  assign n14053 = n9228 ^ n2411 ^ n2131 ;
  assign n14054 = n13618 ^ n3459 ^ 1'b0 ;
  assign n14055 = n14053 & n14054 ;
  assign n14056 = n1440 ^ n1282 ^ 1'b0 ;
  assign n14057 = n2077 & ~n14056 ;
  assign n14058 = n2285 & ~n3989 ;
  assign n14059 = n14058 ^ n7339 ^ 1'b0 ;
  assign n14060 = ~n1810 & n14059 ;
  assign n14061 = ( n1979 & n3988 ) | ( n1979 & ~n14060 ) | ( n3988 & ~n14060 ) ;
  assign n14064 = n8590 ^ n2785 ^ 1'b0 ;
  assign n14065 = n9499 & ~n14064 ;
  assign n14062 = n1921 & n8295 ;
  assign n14063 = n5582 & n14062 ;
  assign n14066 = n14065 ^ n14063 ^ 1'b0 ;
  assign n14072 = n958 & ~n3503 ;
  assign n14068 = ~n491 & n1158 ;
  assign n14069 = n14068 ^ n4444 ^ 1'b0 ;
  assign n14070 = n14069 ^ n8099 ^ n5737 ;
  assign n14071 = n5377 | n14070 ;
  assign n14073 = n14072 ^ n14071 ^ 1'b0 ;
  assign n14067 = n12911 ^ n6261 ^ n438 ;
  assign n14074 = n14073 ^ n14067 ^ 1'b0 ;
  assign n14075 = n6515 | n14074 ;
  assign n14076 = ~n866 & n932 ;
  assign n14077 = n5446 & ~n13426 ;
  assign n14078 = n2926 & n14077 ;
  assign n14079 = ( n4271 & ~n5072 ) | ( n4271 & n14078 ) | ( ~n5072 & n14078 ) ;
  assign n14080 = ( ~n1545 & n4392 ) | ( ~n1545 & n14079 ) | ( n4392 & n14079 ) ;
  assign n14081 = n3664 ^ n2145 ^ 1'b0 ;
  assign n14082 = n12968 ^ n10649 ^ 1'b0 ;
  assign n14083 = ~n950 & n14082 ;
  assign n14084 = ( n11627 & n12188 ) | ( n11627 & ~n14083 ) | ( n12188 & ~n14083 ) ;
  assign n14085 = n3704 ^ n1649 ^ 1'b0 ;
  assign n14086 = n10180 & ~n14085 ;
  assign n14087 = n2308 & n9619 ;
  assign n14088 = ~n14086 & n14087 ;
  assign n14089 = n7265 & n14088 ;
  assign n14090 = ~n637 & n7491 ;
  assign n14091 = n9476 ^ n8936 ^ 1'b0 ;
  assign n14092 = n6067 | n14091 ;
  assign n14093 = n14092 ^ n6145 ^ 1'b0 ;
  assign n14094 = n8984 & n14093 ;
  assign n14095 = ( n1076 & n3299 ) | ( n1076 & n5788 ) | ( n3299 & n5788 ) ;
  assign n14096 = ~n1686 & n14095 ;
  assign n14097 = n8995 ^ n2296 ^ 1'b0 ;
  assign n14098 = n5226 & ~n14097 ;
  assign n14099 = ~n5591 & n7902 ;
  assign n14100 = n13582 ^ n944 ^ 1'b0 ;
  assign n14102 = n5003 & ~n6907 ;
  assign n14101 = n4231 & ~n8129 ;
  assign n14103 = n14102 ^ n14101 ^ 1'b0 ;
  assign n14104 = n3383 & ~n8961 ;
  assign n14105 = n270 & ~n4927 ;
  assign n14108 = n2879 ^ n765 ^ 1'b0 ;
  assign n14109 = n1626 | n14108 ;
  assign n14106 = n9526 ^ n1985 ^ 1'b0 ;
  assign n14107 = ~n9130 & n14106 ;
  assign n14110 = n14109 ^ n14107 ^ 1'b0 ;
  assign n14111 = ( n3834 & n4202 ) | ( n3834 & n7530 ) | ( n4202 & n7530 ) ;
  assign n14112 = n8717 & n14111 ;
  assign n14113 = n9064 ^ n4803 ^ 1'b0 ;
  assign n14114 = n14113 ^ n5198 ^ 1'b0 ;
  assign n14115 = n3136 & ~n14114 ;
  assign n14116 = ( n7217 & n12547 ) | ( n7217 & ~n14115 ) | ( n12547 & ~n14115 ) ;
  assign n14117 = n11193 ^ n7781 ^ n379 ;
  assign n14122 = ( n2375 & n3517 ) | ( n2375 & n5002 ) | ( n3517 & n5002 ) ;
  assign n14118 = n4637 ^ n2448 ^ 1'b0 ;
  assign n14119 = n366 & n14118 ;
  assign n14120 = ~n295 & n14119 ;
  assign n14121 = n14120 ^ n1150 ^ 1'b0 ;
  assign n14123 = n14122 ^ n14121 ^ n6159 ;
  assign n14124 = n14123 ^ n1971 ^ 1'b0 ;
  assign n14125 = n14124 ^ n14111 ^ 1'b0 ;
  assign n14126 = n9826 ^ n7007 ^ 1'b0 ;
  assign n14129 = ~n381 & n10413 ;
  assign n14130 = ~n5783 & n14129 ;
  assign n14131 = n14130 ^ n13985 ^ n9039 ;
  assign n14127 = n14037 ^ n9963 ^ n6819 ;
  assign n14128 = n12065 & n14127 ;
  assign n14132 = n14131 ^ n14128 ^ 1'b0 ;
  assign n14133 = n6741 | n9482 ;
  assign n14135 = ( x61 & n3239 ) | ( x61 & n4029 ) | ( n3239 & n4029 ) ;
  assign n14136 = n402 & n14135 ;
  assign n14137 = n14136 ^ n312 ^ 1'b0 ;
  assign n14134 = ~n6976 & n12100 ;
  assign n14138 = n14137 ^ n14134 ^ 1'b0 ;
  assign n14139 = n11115 ^ n10290 ^ n8366 ;
  assign n14140 = n8677 ^ n3388 ^ x62 ;
  assign n14141 = n4051 ^ n2999 ^ 1'b0 ;
  assign n14142 = n14141 ^ n2654 ^ n1999 ;
  assign n14143 = ~n2171 & n13077 ;
  assign n14144 = n7231 ^ n5902 ^ n330 ;
  assign n14145 = n3560 ^ n1246 ^ n913 ;
  assign n14146 = n14145 ^ n6295 ^ 1'b0 ;
  assign n14147 = n14144 & ~n14146 ;
  assign n14148 = ( n5664 & n5828 ) | ( n5664 & ~n10305 ) | ( n5828 & ~n10305 ) ;
  assign n14149 = ( n3932 & n6522 ) | ( n3932 & ~n14148 ) | ( n6522 & ~n14148 ) ;
  assign n14150 = n5665 ^ n5141 ^ n3430 ;
  assign n14151 = n14149 & ~n14150 ;
  assign n14152 = n7565 ^ n6070 ^ n1712 ;
  assign n14153 = ( n4261 & ~n8572 ) | ( n4261 & n12053 ) | ( ~n8572 & n12053 ) ;
  assign n14154 = n9747 ^ n3731 ^ n344 ;
  assign n14155 = n14009 & ~n14154 ;
  assign n14156 = n8447 ^ n5499 ^ 1'b0 ;
  assign n14157 = n4994 ^ n2570 ^ 1'b0 ;
  assign n14158 = ~n6828 & n14157 ;
  assign n14159 = ~n3971 & n14158 ;
  assign n14160 = n6382 ^ n4261 ^ 1'b0 ;
  assign n14161 = n10160 & n14160 ;
  assign n14162 = n1057 & ~n11256 ;
  assign n14163 = n8769 ^ n429 ^ 1'b0 ;
  assign n14164 = n6050 ^ n4638 ^ 1'b0 ;
  assign n14165 = ~n14163 & n14164 ;
  assign n14166 = n1250 & ~n2748 ;
  assign n14167 = n14166 ^ n9678 ^ 1'b0 ;
  assign n14168 = n5495 | n6227 ;
  assign n14169 = n14168 ^ n5702 ^ 1'b0 ;
  assign n14170 = n14169 ^ n9400 ^ n6003 ;
  assign n14171 = ( n10087 & ~n14167 ) | ( n10087 & n14170 ) | ( ~n14167 & n14170 ) ;
  assign n14172 = n11310 & ~n13325 ;
  assign n14173 = n14172 ^ n10515 ^ 1'b0 ;
  assign n14174 = ~n2163 & n5970 ;
  assign n14175 = n14174 ^ n4396 ^ 1'b0 ;
  assign n14176 = ( ~n6346 & n7565 ) | ( ~n6346 & n14175 ) | ( n7565 & n14175 ) ;
  assign n14177 = n1347 | n5617 ;
  assign n14178 = n6404 ^ n5880 ^ 1'b0 ;
  assign n14179 = ~n14177 & n14178 ;
  assign n14180 = n14176 & n14179 ;
  assign n14181 = n6298 | n12254 ;
  assign n14182 = n11061 & ~n14181 ;
  assign n14183 = n11070 ^ n5308 ^ 1'b0 ;
  assign n14184 = n6339 ^ n5139 ^ 1'b0 ;
  assign n14185 = n14184 ^ n7117 ^ n142 ;
  assign n14186 = ( n1608 & n7103 ) | ( n1608 & n10498 ) | ( n7103 & n10498 ) ;
  assign n14187 = n8869 ^ n2801 ^ n580 ;
  assign n14188 = ( n1996 & n9345 ) | ( n1996 & ~n12818 ) | ( n9345 & ~n12818 ) ;
  assign n14189 = n1200 & ~n1450 ;
  assign n14190 = n6247 ^ n5103 ^ 1'b0 ;
  assign n14191 = ( ~n210 & n14189 ) | ( ~n210 & n14190 ) | ( n14189 & n14190 ) ;
  assign n14192 = n7073 & n10183 ;
  assign n14193 = n10337 ^ n7506 ^ 1'b0 ;
  assign n14194 = ~n2382 & n5571 ;
  assign n14197 = n6803 ^ n6288 ^ n819 ;
  assign n14198 = n1168 & ~n14197 ;
  assign n14195 = n1763 ^ n1186 ^ n586 ;
  assign n14196 = n14195 ^ n1188 ^ 1'b0 ;
  assign n14199 = n14198 ^ n14196 ^ n12768 ;
  assign n14205 = n10387 ^ n5392 ^ 1'b0 ;
  assign n14204 = ~x6 & n4376 ;
  assign n14200 = n349 & ~n4269 ;
  assign n14201 = ~n11204 & n14200 ;
  assign n14202 = n9111 ^ n8987 ^ 1'b0 ;
  assign n14203 = ~n14201 & n14202 ;
  assign n14206 = n14205 ^ n14204 ^ n14203 ;
  assign n14210 = n3610 | n11841 ;
  assign n14211 = n4515 & n14210 ;
  assign n14212 = n14211 ^ n3002 ^ 1'b0 ;
  assign n14207 = n7513 ^ n5205 ^ 1'b0 ;
  assign n14208 = n5928 & ~n14207 ;
  assign n14209 = n14208 ^ n8216 ^ n2599 ;
  assign n14213 = n14212 ^ n14209 ^ n4261 ;
  assign n14214 = n6775 ^ n1186 ^ 1'b0 ;
  assign n14215 = ~n1815 & n14214 ;
  assign n14216 = n14215 ^ n11612 ^ 1'b0 ;
  assign n14217 = n9192 ^ n3100 ^ 1'b0 ;
  assign n14218 = n1473 | n5754 ;
  assign n14219 = n7006 | n14218 ;
  assign n14220 = n6620 | n8580 ;
  assign n14221 = n4463 & ~n14220 ;
  assign n14222 = n3255 | n14221 ;
  assign n14223 = n14222 ^ n6781 ^ 1'b0 ;
  assign n14224 = n8194 ^ n5635 ^ n1334 ;
  assign n14225 = ( n3967 & ~n4962 ) | ( n3967 & n14224 ) | ( ~n4962 & n14224 ) ;
  assign n14226 = ~n165 & n14225 ;
  assign n14227 = n1501 & ~n5367 ;
  assign n14228 = n3177 & n14227 ;
  assign n14231 = n1855 & n2795 ;
  assign n14232 = n14231 ^ n3186 ^ 1'b0 ;
  assign n14229 = ~n5170 & n7143 ;
  assign n14230 = ~n3056 & n14229 ;
  assign n14233 = n14232 ^ n14230 ^ n10598 ;
  assign n14234 = ( x17 & n2353 ) | ( x17 & ~n9228 ) | ( n2353 & ~n9228 ) ;
  assign n14235 = n14234 ^ n11763 ^ 1'b0 ;
  assign n14236 = n14233 | n14235 ;
  assign n14237 = n5558 | n13131 ;
  assign n14238 = n10021 ^ n8933 ^ 1'b0 ;
  assign n14239 = n11307 & ~n14238 ;
  assign n14240 = ( ~n1795 & n6867 ) | ( ~n1795 & n14239 ) | ( n6867 & n14239 ) ;
  assign n14241 = n2155 & n14240 ;
  assign n14242 = n5552 | n6052 ;
  assign n14243 = n14242 ^ n1607 ^ 1'b0 ;
  assign n14246 = n2993 | n7984 ;
  assign n14244 = n11524 ^ n4052 ^ 1'b0 ;
  assign n14245 = n8926 | n14244 ;
  assign n14247 = n14246 ^ n14245 ^ 1'b0 ;
  assign n14248 = n6164 | n6939 ;
  assign n14249 = n4671 & ~n14248 ;
  assign n14250 = n14249 ^ n2397 ^ 1'b0 ;
  assign n14251 = n14247 | n14250 ;
  assign n14252 = n3043 & ~n14251 ;
  assign n14253 = n14252 ^ n11038 ^ 1'b0 ;
  assign n14254 = n9876 ^ n8697 ^ n1139 ;
  assign n14255 = n5664 ^ n3949 ^ 1'b0 ;
  assign n14256 = ~n339 & n14255 ;
  assign n14257 = n14256 ^ n5865 ^ 1'b0 ;
  assign n14258 = n14257 ^ n2772 ^ 1'b0 ;
  assign n14259 = ~n14254 & n14258 ;
  assign n14260 = ~n2345 & n9495 ;
  assign n14261 = n2357 & n14260 ;
  assign n14262 = n14261 ^ n9283 ^ n2212 ;
  assign n14263 = n3149 & ~n4664 ;
  assign n14264 = n14263 ^ n9693 ^ 1'b0 ;
  assign n14265 = n12534 & ~n14264 ;
  assign n14266 = n1461 & n2733 ;
  assign n14267 = ( ~n2944 & n4738 ) | ( ~n2944 & n14266 ) | ( n4738 & n14266 ) ;
  assign n14268 = n12852 ^ n9492 ^ 1'b0 ;
  assign n14269 = ~n14267 & n14268 ;
  assign n14270 = n1702 & n14269 ;
  assign n14271 = n14270 ^ n8016 ^ 1'b0 ;
  assign n14272 = n6208 ^ n3729 ^ 1'b0 ;
  assign n14273 = n3023 | n10114 ;
  assign n14274 = n14273 ^ n5546 ^ 1'b0 ;
  assign n14275 = ( n410 & ~n5902 ) | ( n410 & n6300 ) | ( ~n5902 & n6300 ) ;
  assign n14276 = n14275 ^ n13251 ^ n5613 ;
  assign n14277 = ( ~n2042 & n6342 ) | ( ~n2042 & n10372 ) | ( n6342 & n10372 ) ;
  assign n14278 = n14277 ^ n1853 ^ 1'b0 ;
  assign n14279 = ( n4498 & ~n6653 ) | ( n4498 & n9591 ) | ( ~n6653 & n9591 ) ;
  assign n14280 = n11304 | n14279 ;
  assign n14281 = n14280 ^ x9 ^ 1'b0 ;
  assign n14282 = n4783 & ~n14281 ;
  assign n14283 = n2254 & ~n14282 ;
  assign n14284 = n13799 ^ n7638 ^ 1'b0 ;
  assign n14285 = ( n595 & ~n2930 ) | ( n595 & n9398 ) | ( ~n2930 & n9398 ) ;
  assign n14286 = ( n478 & n8824 ) | ( n478 & n13549 ) | ( n8824 & n13549 ) ;
  assign n14287 = x8 & n12789 ;
  assign n14288 = ~n14286 & n14287 ;
  assign n14289 = ~n6508 & n14288 ;
  assign n14290 = n13090 ^ n8151 ^ n296 ;
  assign n14291 = ~n14289 & n14290 ;
  assign n14292 = n4621 & n14291 ;
  assign n14293 = n2334 & n5171 ;
  assign n14294 = n9569 ^ n3888 ^ n685 ;
  assign n14295 = ~n14221 & n14294 ;
  assign n14296 = n14295 ^ n5931 ^ 1'b0 ;
  assign n14297 = n8995 & n14296 ;
  assign n14298 = ~n14293 & n14297 ;
  assign n14299 = n13567 ^ n4094 ^ 1'b0 ;
  assign n14300 = n6571 | n12052 ;
  assign n14301 = n9037 ^ n4382 ^ 1'b0 ;
  assign n14302 = n6598 | n14301 ;
  assign n14303 = ~n3284 & n14302 ;
  assign n14304 = n160 & ~n3027 ;
  assign n14305 = ~n3212 & n14304 ;
  assign n14306 = n1067 & n4344 ;
  assign n14307 = ~n6550 & n14306 ;
  assign n14308 = n11591 | n14307 ;
  assign n14309 = n14305 & ~n14308 ;
  assign n14310 = n14309 ^ n7738 ^ 1'b0 ;
  assign n14316 = n5620 ^ n1894 ^ 1'b0 ;
  assign n14314 = n12333 & n13885 ;
  assign n14311 = n5169 ^ n5026 ^ 1'b0 ;
  assign n14312 = n6508 & ~n7625 ;
  assign n14313 = ( ~n4367 & n14311 ) | ( ~n4367 & n14312 ) | ( n14311 & n14312 ) ;
  assign n14315 = n14314 ^ n14313 ^ n4703 ;
  assign n14317 = n14316 ^ n14315 ^ 1'b0 ;
  assign n14324 = n1116 ^ n958 ^ n878 ;
  assign n14323 = n6066 ^ n1381 ^ 1'b0 ;
  assign n14318 = n3342 & ~n5512 ;
  assign n14319 = ~n2915 & n14318 ;
  assign n14320 = n6076 | n10098 ;
  assign n14321 = n14319 & ~n14320 ;
  assign n14322 = n14321 ^ n2534 ^ 1'b0 ;
  assign n14325 = n14324 ^ n14323 ^ n14322 ;
  assign n14326 = n4954 ^ x95 ^ 1'b0 ;
  assign n14327 = n14326 ^ n3758 ^ n2745 ;
  assign n14328 = n11962 ^ n2218 ^ 1'b0 ;
  assign n14329 = ( n1470 & ~n9231 ) | ( n1470 & n10827 ) | ( ~n9231 & n10827 ) ;
  assign n14330 = n4756 & ~n7880 ;
  assign n14331 = n14329 & n14330 ;
  assign n14332 = n7404 | n14122 ;
  assign n14333 = ( n4961 & n6630 ) | ( n4961 & n14332 ) | ( n6630 & n14332 ) ;
  assign n14334 = n10165 ^ n5937 ^ n5561 ;
  assign n14335 = ( n1383 & ~n4973 ) | ( n1383 & n14334 ) | ( ~n4973 & n14334 ) ;
  assign n14336 = n6641 ^ n1642 ^ 1'b0 ;
  assign n14337 = n804 & n14336 ;
  assign n14338 = n7091 ^ n3503 ^ 1'b0 ;
  assign n14339 = n14338 ^ n4452 ^ 1'b0 ;
  assign n14340 = n7563 ^ n850 ^ 1'b0 ;
  assign n14341 = n191 & n14340 ;
  assign n14342 = ( ~n3279 & n4273 ) | ( ~n3279 & n14341 ) | ( n4273 & n14341 ) ;
  assign n14343 = n8786 & n14342 ;
  assign n14344 = n9744 | n14343 ;
  assign n14345 = n4472 | n5421 ;
  assign n14346 = n11826 ^ n10851 ^ 1'b0 ;
  assign n14347 = ~n4656 & n13614 ;
  assign n14348 = ( ~n2104 & n8311 ) | ( ~n2104 & n14347 ) | ( n8311 & n14347 ) ;
  assign n14349 = ( n1512 & n10309 ) | ( n1512 & n12099 ) | ( n10309 & n12099 ) ;
  assign n14350 = ~n5088 & n6158 ;
  assign n14351 = n14350 ^ n6509 ^ 1'b0 ;
  assign n14352 = n7571 | n10027 ;
  assign n14353 = ( n1567 & n4492 ) | ( n1567 & ~n8049 ) | ( n4492 & ~n8049 ) ;
  assign n14354 = n14353 ^ n13008 ^ 1'b0 ;
  assign n14355 = n2560 & n6228 ;
  assign n14356 = n10326 & n14355 ;
  assign n14357 = ( n3999 & n7017 ) | ( n3999 & ~n7318 ) | ( n7017 & ~n7318 ) ;
  assign n14358 = n14357 ^ n8075 ^ 1'b0 ;
  assign n14359 = ~n591 & n5791 ;
  assign n14360 = ~n2473 & n11347 ;
  assign n14361 = n11153 & n14360 ;
  assign n14362 = n1776 | n7603 ;
  assign n14363 = n14362 ^ n10202 ^ 1'b0 ;
  assign n14364 = n2092 ^ n1713 ^ 1'b0 ;
  assign n14365 = n14164 & ~n14364 ;
  assign n14366 = n14363 & n14365 ;
  assign n14367 = n2034 & n2843 ;
  assign n14368 = ~n14275 & n14367 ;
  assign n14369 = n14368 ^ n11389 ^ n2213 ;
  assign n14370 = n5811 ^ n1585 ^ 1'b0 ;
  assign n14371 = ~n12452 & n14370 ;
  assign n14372 = n14371 ^ n1262 ^ 1'b0 ;
  assign n14373 = n2687 ^ n927 ^ 1'b0 ;
  assign n14374 = n10433 & ~n14373 ;
  assign n14375 = ( n1287 & n3645 ) | ( n1287 & ~n4833 ) | ( n3645 & ~n4833 ) ;
  assign n14376 = x108 & n9743 ;
  assign n14377 = n5137 & n14376 ;
  assign n14378 = ~n194 & n7403 ;
  assign n14379 = ( ~n11679 & n12970 ) | ( ~n11679 & n14378 ) | ( n12970 & n14378 ) ;
  assign n14380 = n14379 ^ n6230 ^ 1'b0 ;
  assign n14381 = ~n13983 & n14380 ;
  assign n14382 = n14381 ^ n14267 ^ 1'b0 ;
  assign n14390 = ~n5135 & n5413 ;
  assign n14383 = n586 & n940 ;
  assign n14384 = ~n586 & n14383 ;
  assign n14385 = n14384 ^ n7200 ^ n1480 ;
  assign n14386 = n5834 & n14385 ;
  assign n14387 = ~n448 & n14386 ;
  assign n14388 = n9121 | n14387 ;
  assign n14389 = n6653 & ~n14388 ;
  assign n14391 = n14390 ^ n14389 ^ n6857 ;
  assign n14392 = ( n1199 & n3598 ) | ( n1199 & n5174 ) | ( n3598 & n5174 ) ;
  assign n14393 = n14392 ^ n10873 ^ n8817 ;
  assign n14394 = n14393 ^ n3995 ^ 1'b0 ;
  assign n14395 = n5180 | n14394 ;
  assign n14396 = ( n6198 & ~n6247 ) | ( n6198 & n6424 ) | ( ~n6247 & n6424 ) ;
  assign n14397 = n13239 ^ n4236 ^ 1'b0 ;
  assign n14398 = n5126 & ~n14052 ;
  assign n14399 = n12618 ^ n3463 ^ x53 ;
  assign n14400 = n13714 ^ n12173 ^ 1'b0 ;
  assign n14402 = ~n2607 & n4950 ;
  assign n14403 = n4745 & n14402 ;
  assign n14401 = ( n246 & n1010 ) | ( n246 & n13819 ) | ( n1010 & n13819 ) ;
  assign n14404 = n14403 ^ n14401 ^ n8350 ;
  assign n14405 = n13915 ^ n7782 ^ 1'b0 ;
  assign n14406 = n6810 & n14405 ;
  assign n14407 = n250 | n9293 ;
  assign n14408 = n14407 ^ n6922 ^ 1'b0 ;
  assign n14409 = n11764 & ~n14408 ;
  assign n14410 = n11032 ^ n2483 ^ 1'b0 ;
  assign n14411 = n5070 & n11676 ;
  assign n14412 = n8706 & n14411 ;
  assign n14413 = ~n1600 & n8159 ;
  assign n14414 = n14413 ^ n7170 ^ n3928 ;
  assign n14415 = n5700 ^ n5449 ^ 1'b0 ;
  assign n14416 = n2197 ^ n1619 ^ n372 ;
  assign n14417 = ( n3237 & n4431 ) | ( n3237 & ~n6169 ) | ( n4431 & ~n6169 ) ;
  assign n14418 = ( n1313 & n14416 ) | ( n1313 & ~n14417 ) | ( n14416 & ~n14417 ) ;
  assign n14419 = n14415 | n14418 ;
  assign n14420 = n14419 ^ n13503 ^ n3983 ;
  assign n14423 = x119 & ~n2384 ;
  assign n14424 = ~n3181 & n14423 ;
  assign n14421 = ( ~n6201 & n8021 ) | ( ~n6201 & n9406 ) | ( n8021 & n9406 ) ;
  assign n14422 = ~n9626 & n14421 ;
  assign n14425 = n14424 ^ n14422 ^ 1'b0 ;
  assign n14426 = n5337 ^ n4442 ^ 1'b0 ;
  assign n14427 = n654 & ~n6017 ;
  assign n14428 = n14427 ^ n4308 ^ 1'b0 ;
  assign n14429 = ~n491 & n14428 ;
  assign n14430 = ~n12180 & n12564 ;
  assign n14431 = ~n14429 & n14430 ;
  assign n14432 = n1260 & n14011 ;
  assign n14433 = n10050 ^ n9107 ^ n6668 ;
  assign n14434 = x7 & n3828 ;
  assign n14435 = n8126 & n14434 ;
  assign n14436 = n14435 ^ n2796 ^ n339 ;
  assign n14437 = n8922 & n14436 ;
  assign n14438 = n7082 ^ n4424 ^ n2106 ;
  assign n14439 = n6425 | n14438 ;
  assign n14440 = n2976 & ~n14439 ;
  assign n14441 = ~n10145 & n14440 ;
  assign n14443 = ~n5172 & n10398 ;
  assign n14444 = n14443 ^ n6432 ^ 1'b0 ;
  assign n14442 = n5719 & ~n6763 ;
  assign n14445 = n14444 ^ n14442 ^ 1'b0 ;
  assign n14447 = n1723 & ~n8130 ;
  assign n14448 = n1935 & n14447 ;
  assign n14446 = n404 & ~n3234 ;
  assign n14449 = n14448 ^ n14446 ^ 1'b0 ;
  assign n14450 = n11957 | n14449 ;
  assign n14453 = ~n13693 & n14418 ;
  assign n14454 = n1809 & n14453 ;
  assign n14451 = ~n2879 & n9392 ;
  assign n14452 = n7975 & n14451 ;
  assign n14455 = n14454 ^ n14452 ^ 1'b0 ;
  assign n14456 = n1441 & ~n2222 ;
  assign n14457 = n14456 ^ n8668 ^ 1'b0 ;
  assign n14462 = ( n923 & ~n5360 ) | ( n923 & n8617 ) | ( ~n5360 & n8617 ) ;
  assign n14459 = ~x98 & n5561 ;
  assign n14458 = n3342 & n8855 ;
  assign n14460 = n14459 ^ n14458 ^ 1'b0 ;
  assign n14461 = n13508 & ~n14460 ;
  assign n14463 = n14462 ^ n14461 ^ 1'b0 ;
  assign n14464 = ( n3978 & n6509 ) | ( n3978 & n9638 ) | ( n6509 & n9638 ) ;
  assign n14465 = ( ~x92 & n523 ) | ( ~x92 & n2092 ) | ( n523 & n2092 ) ;
  assign n14466 = ( n3241 & ~n14464 ) | ( n3241 & n14465 ) | ( ~n14464 & n14465 ) ;
  assign n14467 = n14466 ^ n210 ^ 1'b0 ;
  assign n14468 = n8787 ^ n1878 ^ 1'b0 ;
  assign n14469 = n6693 | n14468 ;
  assign n14470 = n14469 ^ n152 ^ 1'b0 ;
  assign n14471 = n914 | n9020 ;
  assign n14472 = n13383 & n14471 ;
  assign n14473 = n1924 & n14472 ;
  assign n14475 = ( ~n303 & n665 ) | ( ~n303 & n10076 ) | ( n665 & n10076 ) ;
  assign n14474 = n1997 & n4445 ;
  assign n14476 = n14475 ^ n14474 ^ 1'b0 ;
  assign n14477 = n2648 | n14476 ;
  assign n14478 = n10241 & n10998 ;
  assign n14479 = n14478 ^ n7607 ^ 1'b0 ;
  assign n14480 = n10731 & n14479 ;
  assign n14481 = n14480 ^ n13480 ^ 1'b0 ;
  assign n14482 = n12850 ^ n1683 ^ 1'b0 ;
  assign n14483 = n14482 ^ n6195 ^ 1'b0 ;
  assign n14486 = n3964 ^ n3903 ^ n2898 ;
  assign n14484 = n2415 & n9539 ;
  assign n14485 = n9169 & ~n14484 ;
  assign n14487 = n14486 ^ n14485 ^ n8412 ;
  assign n14488 = n11259 ^ n5772 ^ 1'b0 ;
  assign n14489 = n9532 & n14204 ;
  assign n14490 = ~n3734 & n4914 ;
  assign n14491 = n11579 ^ n8939 ^ 1'b0 ;
  assign n14492 = n14490 | n14491 ;
  assign n14493 = n3674 ^ n1914 ^ 1'b0 ;
  assign n14494 = n8426 ^ n4919 ^ 1'b0 ;
  assign n14495 = n14494 ^ n8645 ^ n1882 ;
  assign n14496 = n14495 ^ n4600 ^ 1'b0 ;
  assign n14497 = n14493 & n14496 ;
  assign n14498 = n453 & n14289 ;
  assign n14499 = n8978 ^ n4597 ^ 1'b0 ;
  assign n14500 = n572 | n14499 ;
  assign n14501 = n12199 ^ n3862 ^ 1'b0 ;
  assign n14502 = n14500 | n14501 ;
  assign n14503 = n5438 & ~n14502 ;
  assign n14504 = n14503 ^ n8958 ^ n4793 ;
  assign n14505 = ~n4246 & n5171 ;
  assign n14506 = n3323 ^ n2933 ^ 1'b0 ;
  assign n14507 = ( n986 & n14505 ) | ( n986 & ~n14506 ) | ( n14505 & ~n14506 ) ;
  assign n14508 = n3484 & n14507 ;
  assign n14509 = n14508 ^ n14395 ^ 1'b0 ;
  assign n14510 = n12719 ^ n5384 ^ n242 ;
  assign n14511 = n3809 | n4175 ;
  assign n14512 = ( ~n1107 & n14510 ) | ( ~n1107 & n14511 ) | ( n14510 & n14511 ) ;
  assign n14513 = n181 & ~n11547 ;
  assign n14514 = ~n5403 & n14513 ;
  assign n14515 = n1897 & ~n14514 ;
  assign n14516 = ~n12709 & n14515 ;
  assign n14517 = n2447 & n5781 ;
  assign n14518 = n14517 ^ n13899 ^ n9476 ;
  assign n14519 = ( n2520 & n3436 ) | ( n2520 & ~n5357 ) | ( n3436 & ~n5357 ) ;
  assign n14520 = n12621 ^ n3747 ^ 1'b0 ;
  assign n14521 = n14519 & n14520 ;
  assign n14522 = n6908 & n14521 ;
  assign n14523 = n14522 ^ n6243 ^ 1'b0 ;
  assign n14524 = n5717 ^ n4103 ^ 1'b0 ;
  assign n14525 = ~n929 & n1956 ;
  assign n14526 = n6187 & n14525 ;
  assign n14527 = n14524 & ~n14526 ;
  assign n14528 = ~n14523 & n14527 ;
  assign n14529 = ( ~n9421 & n12338 ) | ( ~n9421 & n12572 ) | ( n12338 & n12572 ) ;
  assign n14530 = n420 & n7592 ;
  assign n14531 = n5587 & n14530 ;
  assign n14532 = n9049 ^ n6965 ^ n1470 ;
  assign n14533 = n8383 & ~n14532 ;
  assign n14534 = n14531 & n14533 ;
  assign n14535 = n14534 ^ n5338 ^ 1'b0 ;
  assign n14536 = ~n4669 & n6537 ;
  assign n14537 = n14536 ^ n3024 ^ 1'b0 ;
  assign n14538 = n14537 ^ n14390 ^ 1'b0 ;
  assign n14539 = n8205 | n14538 ;
  assign n14540 = n673 & ~n14539 ;
  assign n14541 = ~n1113 & n3995 ;
  assign n14542 = n14541 ^ n7087 ^ 1'b0 ;
  assign n14545 = n6058 ^ n2296 ^ 1'b0 ;
  assign n14546 = ~n12341 & n14545 ;
  assign n14543 = n4592 ^ n2167 ^ 1'b0 ;
  assign n14544 = n3637 & ~n14543 ;
  assign n14547 = n14546 ^ n14544 ^ n1023 ;
  assign n14548 = n1626 & n14547 ;
  assign n14549 = n14548 ^ n5689 ^ 1'b0 ;
  assign n14550 = n4248 ^ n3769 ^ n3293 ;
  assign n14551 = n2331 ^ n2155 ^ n1554 ;
  assign n14552 = n1291 & n10049 ;
  assign n14553 = n14551 & n14552 ;
  assign n14554 = n14553 ^ n14095 ^ 1'b0 ;
  assign n14555 = n9945 ^ n7392 ^ 1'b0 ;
  assign n14556 = n3905 | n14555 ;
  assign n14557 = n6013 | n14556 ;
  assign n14558 = n14557 ^ n5696 ^ 1'b0 ;
  assign n14559 = ( n14550 & n14554 ) | ( n14550 & n14558 ) | ( n14554 & n14558 ) ;
  assign n14560 = n4714 ^ n319 ^ 1'b0 ;
  assign n14561 = n14560 ^ n3187 ^ n1041 ;
  assign n14562 = n10978 & n14561 ;
  assign n14563 = n8939 & n10966 ;
  assign n14564 = n11616 ^ n5433 ^ 1'b0 ;
  assign n14565 = n325 | n593 ;
  assign n14566 = n1939 | n14565 ;
  assign n14567 = n9794 ^ n565 ^ 1'b0 ;
  assign n14568 = n5159 & ~n14567 ;
  assign n14569 = n13822 | n14568 ;
  assign n14570 = n11498 ^ n9795 ^ 1'b0 ;
  assign n14571 = n1515 & ~n2195 ;
  assign n14572 = n4215 & n14571 ;
  assign n14573 = n14570 | n14572 ;
  assign n14574 = n5586 & ~n14573 ;
  assign n14575 = n6333 & n14574 ;
  assign n14576 = ( n3552 & n11343 ) | ( n3552 & ~n14575 ) | ( n11343 & ~n14575 ) ;
  assign n14579 = n424 & ~n10366 ;
  assign n14580 = n14579 ^ n6730 ^ 1'b0 ;
  assign n14577 = ~n1381 & n5533 ;
  assign n14578 = n240 & n14577 ;
  assign n14581 = n14580 ^ n14578 ^ n5634 ;
  assign n14582 = ( ~n1126 & n1714 ) | ( ~n1126 & n9620 ) | ( n1714 & n9620 ) ;
  assign n14586 = n14314 ^ n11858 ^ 1'b0 ;
  assign n14587 = ~n13075 & n14586 ;
  assign n14584 = n4233 ^ n2535 ^ 1'b0 ;
  assign n14585 = n14584 ^ n6083 ^ n258 ;
  assign n14583 = ( n2070 & n8756 ) | ( n2070 & ~n10909 ) | ( n8756 & ~n10909 ) ;
  assign n14588 = n14587 ^ n14585 ^ n14583 ;
  assign n14589 = n14582 & n14588 ;
  assign n14590 = n8425 & ~n11321 ;
  assign n14591 = n650 & ~n12161 ;
  assign n14592 = n14591 ^ n6917 ^ 1'b0 ;
  assign n14593 = ~n14590 & n14592 ;
  assign n14594 = n133 & ~n911 ;
  assign n14595 = n2779 & n14594 ;
  assign n14596 = n14595 ^ n1712 ^ 1'b0 ;
  assign n14597 = n14593 & n14596 ;
  assign n14601 = n155 | n5016 ;
  assign n14598 = n6484 ^ n4834 ^ 1'b0 ;
  assign n14599 = n14598 ^ n2536 ^ n1685 ;
  assign n14600 = n14599 ^ n8440 ^ n3448 ;
  assign n14602 = n14601 ^ n14600 ^ 1'b0 ;
  assign n14603 = ~n1748 & n14602 ;
  assign n14604 = n8193 ^ n6768 ^ 1'b0 ;
  assign n14605 = n6620 | n14604 ;
  assign n14606 = ( n4700 & n8900 ) | ( n4700 & n14605 ) | ( n8900 & n14605 ) ;
  assign n14607 = n8271 ^ n1669 ^ 1'b0 ;
  assign n14608 = ~n11632 & n14607 ;
  assign n14609 = n3770 ^ n2328 ^ 1'b0 ;
  assign n14610 = n8676 & ~n14609 ;
  assign n14611 = n1353 & n14610 ;
  assign n14612 = n471 & ~n3830 ;
  assign n14613 = n9591 ^ n331 ^ 1'b0 ;
  assign n14614 = ~n14612 & n14613 ;
  assign n14617 = ~n2651 & n11442 ;
  assign n14618 = n14617 ^ n6232 ^ 1'b0 ;
  assign n14615 = ( n4035 & n5499 ) | ( n4035 & ~n9904 ) | ( n5499 & ~n9904 ) ;
  assign n14616 = ~n3694 & n14615 ;
  assign n14619 = n14618 ^ n14616 ^ 1'b0 ;
  assign n14621 = ~n2837 & n4978 ;
  assign n14622 = n14621 ^ n8649 ^ 1'b0 ;
  assign n14620 = ( n3060 & n4743 ) | ( n3060 & ~n10166 ) | ( n4743 & ~n10166 ) ;
  assign n14623 = n14622 ^ n14620 ^ 1'b0 ;
  assign n14624 = n8112 ^ n3236 ^ 1'b0 ;
  assign n14625 = n14624 ^ n8438 ^ 1'b0 ;
  assign n14626 = n2611 & ~n2933 ;
  assign n14627 = n14626 ^ n3681 ^ 1'b0 ;
  assign n14628 = n14627 ^ n9402 ^ n3686 ;
  assign n14629 = ( ~n10643 & n14625 ) | ( ~n10643 & n14628 ) | ( n14625 & n14628 ) ;
  assign n14630 = n2630 & n4542 ;
  assign n14631 = ( ~n1470 & n7229 ) | ( ~n1470 & n14630 ) | ( n7229 & n14630 ) ;
  assign n14632 = n14631 ^ n11987 ^ n5131 ;
  assign n14633 = ~n5005 & n14632 ;
  assign n14634 = n14633 ^ n8751 ^ 1'b0 ;
  assign n14635 = n3660 & n7794 ;
  assign n14636 = ~n8780 & n9271 ;
  assign n14637 = n14636 ^ n1615 ^ 1'b0 ;
  assign n14638 = ~n1020 & n10974 ;
  assign n14639 = n2710 & n14638 ;
  assign n14640 = n14639 ^ n6876 ^ 1'b0 ;
  assign n14641 = ( n4589 & ~n14637 ) | ( n4589 & n14640 ) | ( ~n14637 & n14640 ) ;
  assign n14642 = n905 & ~n8149 ;
  assign n14643 = n14642 ^ n3776 ^ 1'b0 ;
  assign n14644 = n8824 & ~n8837 ;
  assign n14645 = ~n6913 & n14644 ;
  assign n14646 = n2120 ^ n1084 ^ 1'b0 ;
  assign n14647 = n6702 & ~n14646 ;
  assign n14648 = n14647 ^ n2576 ^ 1'b0 ;
  assign n14649 = n2139 | n11365 ;
  assign n14650 = n14649 ^ n12942 ^ 1'b0 ;
  assign n14651 = n6025 ^ n3930 ^ 1'b0 ;
  assign n14652 = n6333 ^ n4858 ^ 1'b0 ;
  assign n14653 = n1295 & n10297 ;
  assign n14654 = n14653 ^ n8952 ^ 1'b0 ;
  assign n14655 = n12100 ^ n1114 ^ 1'b0 ;
  assign n14656 = n7992 | n12052 ;
  assign n14657 = n597 & ~n14656 ;
  assign n14658 = n3545 ^ n3179 ^ 1'b0 ;
  assign n14659 = n14657 | n14658 ;
  assign n14660 = n14659 ^ n477 ^ 1'b0 ;
  assign n14661 = ( n4463 & n4884 ) | ( n4463 & ~n6426 ) | ( n4884 & ~n6426 ) ;
  assign n14662 = ( n6137 & ~n6221 ) | ( n6137 & n14661 ) | ( ~n6221 & n14661 ) ;
  assign n14663 = n10780 ^ n944 ^ 1'b0 ;
  assign n14664 = n5387 & ~n5979 ;
  assign n14665 = n5181 ^ n1552 ^ x0 ;
  assign n14666 = n14665 ^ n6891 ^ n3349 ;
  assign n14667 = ( n1025 & n1156 ) | ( n1025 & ~n1349 ) | ( n1156 & ~n1349 ) ;
  assign n14668 = n4549 | n14667 ;
  assign n14669 = n14668 ^ n1242 ^ 1'b0 ;
  assign n14670 = n13423 ^ n1383 ^ 1'b0 ;
  assign n14671 = ( ~n2500 & n4120 ) | ( ~n2500 & n7034 ) | ( n4120 & n7034 ) ;
  assign n14672 = n1868 | n14671 ;
  assign n14673 = n1485 & ~n14672 ;
  assign n14674 = n6768 ^ n3123 ^ 1'b0 ;
  assign n14676 = n1011 | n11465 ;
  assign n14675 = n7133 ^ n4005 ^ n2422 ;
  assign n14677 = n14676 ^ n14675 ^ n14627 ;
  assign n14678 = ~n2695 & n5895 ;
  assign n14679 = n14678 ^ n7103 ^ 1'b0 ;
  assign n14680 = n11015 & n13300 ;
  assign n14681 = ~n819 & n10499 ;
  assign n14682 = n14681 ^ n10599 ^ 1'b0 ;
  assign n14683 = n14682 ^ n11829 ^ 1'b0 ;
  assign n14684 = n1300 & ~n14683 ;
  assign n14685 = ( ~n279 & n9090 ) | ( ~n279 & n13413 ) | ( n9090 & n13413 ) ;
  assign n14686 = n6930 ^ n6316 ^ 1'b0 ;
  assign n14687 = n4206 & n14686 ;
  assign n14688 = n7794 ^ n7415 ^ 1'b0 ;
  assign n14689 = n8438 ^ n3342 ^ 1'b0 ;
  assign n14690 = n1648 & n14689 ;
  assign n14694 = n14465 ^ n5269 ^ 1'b0 ;
  assign n14691 = n9162 ^ n1136 ^ n509 ;
  assign n14692 = n14691 ^ n8599 ^ n6859 ;
  assign n14693 = n14664 | n14692 ;
  assign n14695 = n14694 ^ n14693 ^ 1'b0 ;
  assign n14696 = ~n180 & n8700 ;
  assign n14698 = n8801 ^ n8099 ^ n4574 ;
  assign n14697 = n12727 ^ n4088 ^ 1'b0 ;
  assign n14699 = n14698 ^ n14697 ^ 1'b0 ;
  assign n14700 = n14696 & n14699 ;
  assign n14701 = n9605 & n13933 ;
  assign n14702 = ~n12937 & n14701 ;
  assign n14703 = n461 | n8550 ;
  assign n14704 = ( ~x0 & n7392 ) | ( ~x0 & n11323 ) | ( n7392 & n11323 ) ;
  assign n14705 = n14703 & n14704 ;
  assign n14706 = n14705 ^ n8835 ^ 1'b0 ;
  assign n14707 = n8258 | n14706 ;
  assign n14708 = ( n5800 & n14702 ) | ( n5800 & ~n14707 ) | ( n14702 & ~n14707 ) ;
  assign n14709 = n366 | n3665 ;
  assign n14710 = n3558 & n14709 ;
  assign n14711 = ~n4380 & n14710 ;
  assign n14712 = ( ~n423 & n10036 ) | ( ~n423 & n14711 ) | ( n10036 & n14711 ) ;
  assign n14713 = n8910 ^ n6522 ^ 1'b0 ;
  assign n14714 = ( n793 & n1914 ) | ( n793 & ~n14713 ) | ( n1914 & ~n14713 ) ;
  assign n14715 = n10894 ^ n1485 ^ 1'b0 ;
  assign n14716 = n10033 & n14715 ;
  assign n14717 = n1929 | n11891 ;
  assign n14718 = n14717 ^ n5689 ^ 1'b0 ;
  assign n14719 = n13813 ^ n862 ^ 1'b0 ;
  assign n14720 = n356 & n10974 ;
  assign n14721 = n14720 ^ n9357 ^ 1'b0 ;
  assign n14724 = ~n8268 & n10824 ;
  assign n14725 = n14724 ^ x20 ^ 1'b0 ;
  assign n14722 = n14312 ^ n8762 ^ n7133 ;
  assign n14723 = n1216 | n14722 ;
  assign n14726 = n14725 ^ n14723 ^ 1'b0 ;
  assign n14727 = ~n1815 & n13957 ;
  assign n14728 = ~n5854 & n7323 ;
  assign n14729 = ~n773 & n14728 ;
  assign n14730 = n146 | n11301 ;
  assign n14731 = ( n1584 & ~n2011 ) | ( n1584 & n3686 ) | ( ~n2011 & n3686 ) ;
  assign n14732 = n14731 ^ n10640 ^ 1'b0 ;
  assign n14733 = n11860 ^ n5661 ^ 1'b0 ;
  assign n14734 = ( n8533 & n14732 ) | ( n8533 & n14733 ) | ( n14732 & n14733 ) ;
  assign n14735 = n6440 ^ n2778 ^ 1'b0 ;
  assign n14736 = ~n8365 & n14735 ;
  assign n14737 = n14736 ^ n11470 ^ 1'b0 ;
  assign n14738 = n3271 | n9524 ;
  assign n14739 = ( n6199 & ~n14737 ) | ( n6199 & n14738 ) | ( ~n14737 & n14738 ) ;
  assign n14740 = n5677 & ~n10834 ;
  assign n14741 = n14740 ^ n6580 ^ 1'b0 ;
  assign n14742 = n14741 ^ n10233 ^ 1'b0 ;
  assign n14743 = ~n2344 & n14742 ;
  assign n14744 = ( n5595 & n6041 ) | ( n5595 & ~n7051 ) | ( n6041 & ~n7051 ) ;
  assign n14745 = n14744 ^ n9586 ^ 1'b0 ;
  assign n14746 = n9619 ^ n6899 ^ 1'b0 ;
  assign n14747 = n14745 | n14746 ;
  assign n14748 = n2124 | n5313 ;
  assign n14749 = n9038 ^ n8400 ^ 1'b0 ;
  assign n14750 = n14748 & ~n14749 ;
  assign n14751 = n484 | n7116 ;
  assign n14752 = n11230 & ~n14751 ;
  assign n14755 = n6312 ^ n4456 ^ 1'b0 ;
  assign n14753 = n1929 & n4904 ;
  assign n14754 = n14753 ^ n10393 ^ 1'b0 ;
  assign n14756 = n14755 ^ n14754 ^ n9441 ;
  assign n14757 = n12277 ^ n7737 ^ n868 ;
  assign n14758 = n1882 ^ n459 ^ 1'b0 ;
  assign n14759 = n3189 & ~n14758 ;
  assign n14760 = n14759 ^ n8144 ^ n3772 ;
  assign n14761 = n14757 & n14760 ;
  assign n14762 = ~n4103 & n5555 ;
  assign n14763 = n7316 | n11342 ;
  assign n14764 = ~n5750 & n14763 ;
  assign n14765 = ~n14762 & n14764 ;
  assign n14766 = n11402 | n11458 ;
  assign n14767 = n12814 & ~n14766 ;
  assign n14768 = n2163 | n3389 ;
  assign n14769 = n14768 ^ n10777 ^ 1'b0 ;
  assign n14770 = n4373 & ~n9160 ;
  assign n14771 = n10300 | n14770 ;
  assign n14772 = n14769 & ~n14771 ;
  assign n14773 = n1712 | n11609 ;
  assign n14774 = ( n8411 & n13833 ) | ( n8411 & ~n14773 ) | ( n13833 & ~n14773 ) ;
  assign n14775 = n5732 & n11304 ;
  assign n14776 = n7350 | n14775 ;
  assign n14777 = n14595 ^ n4714 ^ 1'b0 ;
  assign n14778 = n5910 & n14777 ;
  assign n14779 = x119 & n14778 ;
  assign n14780 = n14779 ^ n1428 ^ 1'b0 ;
  assign n14781 = ( n3858 & ~n8539 ) | ( n3858 & n14780 ) | ( ~n8539 & n14780 ) ;
  assign n14782 = n14781 ^ n14119 ^ 1'b0 ;
  assign n14783 = ( ~n5514 & n8198 ) | ( ~n5514 & n10036 ) | ( n8198 & n10036 ) ;
  assign n14784 = n14783 ^ n3359 ^ 1'b0 ;
  assign n14785 = n14782 & ~n14784 ;
  assign n14786 = n7778 | n10027 ;
  assign n14787 = n14786 ^ n4078 ^ 1'b0 ;
  assign n14788 = n11068 | n14787 ;
  assign n14789 = n14788 ^ n13899 ^ 1'b0 ;
  assign n14790 = ~n2066 & n14789 ;
  assign n14791 = n5003 ^ n2169 ^ 1'b0 ;
  assign n14796 = n946 | n2512 ;
  assign n14797 = n14796 ^ n2275 ^ 1'b0 ;
  assign n14798 = n14797 ^ n6885 ^ n2633 ;
  assign n14795 = n1803 & n13142 ;
  assign n14792 = n2948 & n10164 ;
  assign n14793 = n14792 ^ n8504 ^ 1'b0 ;
  assign n14794 = ( n3819 & ~n5958 ) | ( n3819 & n14793 ) | ( ~n5958 & n14793 ) ;
  assign n14799 = n14798 ^ n14795 ^ n14794 ;
  assign n14800 = ( x120 & n9093 ) | ( x120 & n9424 ) | ( n9093 & n9424 ) ;
  assign n14801 = n429 ^ n203 ^ 1'b0 ;
  assign n14802 = n5460 | n14801 ;
  assign n14803 = n8576 & n14802 ;
  assign n14804 = n2891 & n8426 ;
  assign n14805 = n7699 & n14804 ;
  assign n14806 = n6186 & ~n14805 ;
  assign n14807 = n14806 ^ n964 ^ 1'b0 ;
  assign n14809 = n7180 & ~n8812 ;
  assign n14810 = ~n6092 & n14809 ;
  assign n14808 = n3035 & n12244 ;
  assign n14811 = n14810 ^ n14808 ^ 1'b0 ;
  assign n14815 = n4369 ^ n4193 ^ n1984 ;
  assign n14812 = ( n4374 & n12945 ) | ( n4374 & n14047 ) | ( n12945 & n14047 ) ;
  assign n14813 = ( n2150 & n10605 ) | ( n2150 & n14812 ) | ( n10605 & n14812 ) ;
  assign n14814 = n14813 ^ n10502 ^ 1'b0 ;
  assign n14816 = n14815 ^ n14814 ^ 1'b0 ;
  assign n14817 = n184 & n9499 ;
  assign n14820 = n13926 ^ n12366 ^ n5397 ;
  assign n14818 = ~n2930 & n10224 ;
  assign n14819 = n453 & ~n14818 ;
  assign n14821 = n14820 ^ n14819 ^ 1'b0 ;
  assign n14823 = ( n5725 & ~n5783 ) | ( n5725 & n7212 ) | ( ~n5783 & n7212 ) ;
  assign n14822 = n13510 ^ n6880 ^ n1108 ;
  assign n14824 = n14823 ^ n14822 ^ n274 ;
  assign n14825 = n10110 ^ n6269 ^ n5533 ;
  assign n14826 = n14825 ^ n8033 ^ 1'b0 ;
  assign n14827 = n14826 ^ n6198 ^ n2521 ;
  assign n14828 = n4574 & n14775 ;
  assign n14829 = ~n14827 & n14828 ;
  assign n14830 = n6533 ^ n6166 ^ 1'b0 ;
  assign n14831 = n5037 & n13713 ;
  assign n14832 = n7206 & n14831 ;
  assign n14833 = n10352 ^ n2682 ^ 1'b0 ;
  assign n14834 = ~n8598 & n14833 ;
  assign n14835 = n421 | n7137 ;
  assign n14836 = n8839 & ~n14835 ;
  assign n14837 = n14836 ^ n4206 ^ n4059 ;
  assign n14842 = n3359 | n5016 ;
  assign n14843 = n14842 ^ n7308 ^ 1'b0 ;
  assign n14841 = n4896 & ~n6619 ;
  assign n14844 = n14843 ^ n14841 ^ 1'b0 ;
  assign n14838 = ( n2755 & n8447 ) | ( n2755 & n12626 ) | ( n8447 & n12626 ) ;
  assign n14839 = n8312 | n14838 ;
  assign n14840 = n14839 ^ n1655 ^ 1'b0 ;
  assign n14845 = n14844 ^ n14840 ^ 1'b0 ;
  assign n14846 = n7984 & n10487 ;
  assign n14847 = n14846 ^ n787 ^ 1'b0 ;
  assign n14848 = n5539 & n14847 ;
  assign n14849 = ~n14845 & n14848 ;
  assign n14850 = n6758 ^ n5784 ^ 1'b0 ;
  assign n14852 = n259 | n2259 ;
  assign n14853 = n14852 ^ n10965 ^ n6984 ;
  assign n14851 = n8990 | n9238 ;
  assign n14854 = n14853 ^ n14851 ^ 1'b0 ;
  assign n14855 = n9703 ^ n7686 ^ n3025 ;
  assign n14856 = n8757 & ~n14855 ;
  assign n14857 = n14856 ^ n14143 ^ 1'b0 ;
  assign n14858 = ~n1888 & n3479 ;
  assign n14859 = ~n9575 & n14858 ;
  assign n14860 = n5890 | n13374 ;
  assign n14861 = ~n386 & n1986 ;
  assign n14862 = n14861 ^ n3323 ^ 1'b0 ;
  assign n14863 = n5131 & ~n8314 ;
  assign n14864 = ~n14862 & n14863 ;
  assign n14865 = x105 & n2686 ;
  assign n14866 = n14865 ^ n3523 ^ 1'b0 ;
  assign n14867 = n3655 & n10015 ;
  assign n14868 = n14866 & n14867 ;
  assign n14869 = n14122 ^ n5815 ^ n1748 ;
  assign n14870 = n370 | n8154 ;
  assign n14871 = n2709 ^ n2494 ^ 1'b0 ;
  assign n14872 = ~n7716 & n14871 ;
  assign n14873 = n14872 ^ n5954 ^ 1'b0 ;
  assign n14874 = ~n10476 & n14873 ;
  assign n14875 = n246 & ~n1096 ;
  assign n14876 = ~n4512 & n14875 ;
  assign n14877 = n11078 ^ n403 ^ 1'b0 ;
  assign n14878 = n14877 ^ n11935 ^ n4342 ;
  assign n14879 = n14876 | n14878 ;
  assign n14880 = n11282 | n14879 ;
  assign n14881 = n13478 | n14495 ;
  assign n14882 = n2273 | n14881 ;
  assign n14883 = n7176 ^ n523 ^ 1'b0 ;
  assign n14884 = n9586 ^ n4607 ^ 1'b0 ;
  assign n14885 = n5984 & n14884 ;
  assign n14886 = n9409 ^ n4722 ^ 1'b0 ;
  assign n14887 = ~n1623 & n14886 ;
  assign n14888 = n1496 | n10847 ;
  assign n14889 = n14888 ^ n822 ^ 1'b0 ;
  assign n14890 = n4263 ^ n1216 ^ 1'b0 ;
  assign n14891 = ~n2173 & n14890 ;
  assign n14892 = n14891 ^ n1218 ^ 1'b0 ;
  assign n14893 = ~n11153 & n14892 ;
  assign n14894 = ~n10644 & n14893 ;
  assign n14895 = n3559 & n14894 ;
  assign n14896 = ~n898 & n8824 ;
  assign n14897 = n14896 ^ n718 ^ 1'b0 ;
  assign n14898 = n14897 ^ n6196 ^ n295 ;
  assign n14899 = n2954 & n8406 ;
  assign n14900 = n14899 ^ n5340 ^ 1'b0 ;
  assign n14901 = ~n5915 & n7557 ;
  assign n14902 = n6909 & n14901 ;
  assign n14903 = n12341 | n14902 ;
  assign n14904 = n14900 & ~n14903 ;
  assign n14905 = n5784 & n10168 ;
  assign n14906 = ~n4658 & n14905 ;
  assign n14907 = n1478 & n6374 ;
  assign n14908 = n14907 ^ n11665 ^ 1'b0 ;
  assign n14909 = n14908 ^ n1190 ^ 1'b0 ;
  assign n14910 = n10673 ^ n5808 ^ 1'b0 ;
  assign n14911 = ~n8257 & n10967 ;
  assign n14912 = n14911 ^ n3001 ^ 1'b0 ;
  assign n14913 = n715 & n10597 ;
  assign n14914 = n11946 ^ n9132 ^ 1'b0 ;
  assign n14915 = n8494 ^ n7534 ^ n984 ;
  assign n14916 = ( ~n2737 & n2833 ) | ( ~n2737 & n7339 ) | ( n2833 & n7339 ) ;
  assign n14917 = n2808 & ~n8759 ;
  assign n14918 = ~n14916 & n14917 ;
  assign n14919 = ( n1240 & n14915 ) | ( n1240 & ~n14918 ) | ( n14915 & ~n14918 ) ;
  assign n14922 = n5904 ^ n4645 ^ n1539 ;
  assign n14923 = n14922 ^ n11808 ^ 1'b0 ;
  assign n14920 = n1517 & n2028 ;
  assign n14921 = n6889 | n14920 ;
  assign n14924 = n14923 ^ n14921 ^ n11001 ;
  assign n14927 = ~n3319 & n8241 ;
  assign n14925 = n3102 | n10592 ;
  assign n14926 = n10193 | n14925 ;
  assign n14928 = n14927 ^ n14926 ^ 1'b0 ;
  assign n14929 = n13970 ^ n9801 ^ 1'b0 ;
  assign n14930 = n4078 & ~n14929 ;
  assign n14931 = n14136 ^ n11207 ^ 1'b0 ;
  assign n14932 = n14930 & n14931 ;
  assign n14933 = n4288 | n5522 ;
  assign n14934 = ( n438 & ~n4664 ) | ( n438 & n14933 ) | ( ~n4664 & n14933 ) ;
  assign n14935 = n7094 & ~n14934 ;
  assign n14936 = n14934 & n14935 ;
  assign n14937 = n9848 ^ n5963 ^ n3281 ;
  assign n14938 = n3169 | n9369 ;
  assign n14939 = n14938 ^ n3126 ^ 1'b0 ;
  assign n14940 = ( n1936 & n11420 ) | ( n1936 & ~n14939 ) | ( n11420 & ~n14939 ) ;
  assign n14941 = ( n3330 & n3816 ) | ( n3330 & ~n6585 ) | ( n3816 & ~n6585 ) ;
  assign n14942 = n501 & n14941 ;
  assign n14943 = n14942 ^ n9933 ^ 1'b0 ;
  assign n14944 = n4578 ^ n1659 ^ n477 ;
  assign n14945 = ( n6396 & n7593 ) | ( n6396 & n14944 ) | ( n7593 & n14944 ) ;
  assign n14946 = n9203 & n10181 ;
  assign n14947 = n14945 & n14946 ;
  assign n14948 = n5859 | n8130 ;
  assign n14949 = n14948 ^ x13 ^ 1'b0 ;
  assign n14950 = ( n7016 & ~n8845 ) | ( n7016 & n11944 ) | ( ~n8845 & n11944 ) ;
  assign n14951 = n7543 & n14950 ;
  assign n14952 = ( ~n2930 & n3583 ) | ( ~n2930 & n7932 ) | ( n3583 & n7932 ) ;
  assign n14953 = n13133 ^ n9619 ^ 1'b0 ;
  assign n14954 = n13670 ^ n716 ^ 1'b0 ;
  assign n14955 = n2399 & n14954 ;
  assign n14956 = ~n1779 & n14955 ;
  assign n14957 = n4186 & n14956 ;
  assign n14958 = n12786 | n14957 ;
  assign n14959 = n14958 ^ n5692 ^ 1'b0 ;
  assign n14960 = n14814 & ~n14959 ;
  assign n14961 = n12933 ^ n1222 ^ 1'b0 ;
  assign n14962 = n6645 & ~n14961 ;
  assign n14963 = ( ~n9445 & n12299 ) | ( ~n9445 & n14962 ) | ( n12299 & n14962 ) ;
  assign n14964 = ( n5734 & ~n9018 ) | ( n5734 & n11394 ) | ( ~n9018 & n11394 ) ;
  assign n14965 = n6794 & n10429 ;
  assign n14966 = n4596 ^ n3519 ^ 1'b0 ;
  assign n14967 = ~n992 & n14966 ;
  assign n14968 = n14967 ^ n8163 ^ 1'b0 ;
  assign n14969 = n1311 & n14968 ;
  assign n14970 = n10541 & n14969 ;
  assign n14971 = n7237 ^ n207 ^ 1'b0 ;
  assign n14972 = n6766 & ~n14971 ;
  assign n14973 = n14972 ^ n2221 ^ 1'b0 ;
  assign n14974 = n11368 ^ n6609 ^ n2458 ;
  assign n14975 = n14974 ^ n7707 ^ n5652 ;
  assign n14977 = ~n1729 & n7807 ;
  assign n14978 = n14977 ^ n12714 ^ 1'b0 ;
  assign n14976 = n2860 & ~n7916 ;
  assign n14979 = n14978 ^ n14976 ^ 1'b0 ;
  assign n14980 = n14587 & ~n14979 ;
  assign n14981 = n6772 ^ n5401 ^ n4689 ;
  assign n14982 = n12662 & ~n14981 ;
  assign n14983 = n14982 ^ n4669 ^ 1'b0 ;
  assign n14984 = n14249 ^ n3449 ^ 1'b0 ;
  assign n14985 = ~n9528 & n14984 ;
  assign n14986 = n2536 & n14985 ;
  assign n14987 = n5515 & n14986 ;
  assign n14988 = n6282 & n8478 ;
  assign n14989 = n14988 ^ n3811 ^ 1'b0 ;
  assign n14990 = n2687 & n14989 ;
  assign n14991 = n14990 ^ n1931 ^ 1'b0 ;
  assign n14992 = n11088 ^ n1503 ^ 1'b0 ;
  assign n14993 = n11784 ^ n11255 ^ 1'b0 ;
  assign n14994 = n6668 ^ n1006 ^ 1'b0 ;
  assign n14995 = n1596 | n8767 ;
  assign n14996 = n7618 | n14995 ;
  assign n14997 = n6053 | n14996 ;
  assign n14998 = n6527 & n14997 ;
  assign n14999 = n3463 & n6214 ;
  assign n15000 = n4584 & n14999 ;
  assign n15001 = ( n14994 & ~n14998 ) | ( n14994 & n15000 ) | ( ~n14998 & n15000 ) ;
  assign n15002 = n15001 ^ n12816 ^ n12201 ;
  assign n15008 = ~n6232 & n10620 ;
  assign n15003 = ( ~n1305 & n8298 ) | ( ~n1305 & n13332 ) | ( n8298 & n13332 ) ;
  assign n15004 = n15003 ^ n5522 ^ 1'b0 ;
  assign n15005 = ~n6897 & n15004 ;
  assign n15006 = n2598 & n15005 ;
  assign n15007 = n15006 ^ n927 ^ 1'b0 ;
  assign n15009 = n15008 ^ n15007 ^ 1'b0 ;
  assign n15010 = n6254 & ~n15009 ;
  assign n15011 = n9226 ^ n606 ^ 1'b0 ;
  assign n15012 = ~x20 & n5147 ;
  assign n15013 = n15012 ^ n6686 ^ n5933 ;
  assign n15014 = n3403 ^ n2905 ^ n985 ;
  assign n15015 = n4246 ^ n730 ^ 1'b0 ;
  assign n15019 = n3593 ^ n3240 ^ 1'b0 ;
  assign n15016 = n7341 & n13102 ;
  assign n15017 = n15016 ^ n1558 ^ n646 ;
  assign n15018 = n9903 | n15017 ;
  assign n15020 = n15019 ^ n15018 ^ 1'b0 ;
  assign n15021 = n4342 | n9362 ;
  assign n15022 = n9236 | n11841 ;
  assign n15023 = n15022 ^ n7958 ^ 1'b0 ;
  assign n15024 = ( n846 & n3883 ) | ( n846 & ~n15023 ) | ( n3883 & ~n15023 ) ;
  assign n15025 = n13029 ^ n5962 ^ 1'b0 ;
  assign n15026 = ~n1317 & n15025 ;
  assign n15027 = ( n918 & n1554 ) | ( n918 & ~n15026 ) | ( n1554 & ~n15026 ) ;
  assign n15028 = n15027 ^ n9613 ^ 1'b0 ;
  assign n15029 = n11574 | n15028 ;
  assign n15030 = n10699 | n15029 ;
  assign n15035 = n2409 ^ n1756 ^ 1'b0 ;
  assign n15032 = n4691 & n10309 ;
  assign n15033 = n9526 & n15032 ;
  assign n15034 = n6477 & ~n15033 ;
  assign n15036 = n15035 ^ n15034 ^ 1'b0 ;
  assign n15031 = n7732 | n14981 ;
  assign n15037 = n15036 ^ n15031 ^ 1'b0 ;
  assign n15038 = n15037 ^ n8929 ^ 1'b0 ;
  assign n15039 = n7859 ^ n1470 ^ 1'b0 ;
  assign n15040 = ~n13065 & n15039 ;
  assign n15041 = ~n5987 & n15040 ;
  assign n15042 = n15041 ^ n5548 ^ 1'b0 ;
  assign n15043 = n5011 | n5958 ;
  assign n15044 = n9464 ^ n4077 ^ 1'b0 ;
  assign n15045 = ~n3134 & n15044 ;
  assign n15046 = n13556 ^ n12726 ^ 1'b0 ;
  assign n15048 = n6668 ^ n5786 ^ 1'b0 ;
  assign n15049 = ( ~n7828 & n9553 ) | ( ~n7828 & n15048 ) | ( n9553 & n15048 ) ;
  assign n15047 = n2859 & ~n6380 ;
  assign n15050 = n15049 ^ n15047 ^ 1'b0 ;
  assign n15051 = n15050 ^ n12611 ^ n2456 ;
  assign n15052 = ( ~n6136 & n11297 ) | ( ~n6136 & n15051 ) | ( n11297 & n15051 ) ;
  assign n15053 = n4095 ^ n2910 ^ 1'b0 ;
  assign n15054 = n15053 ^ n8184 ^ n3403 ;
  assign n15055 = n4854 ^ n368 ^ 1'b0 ;
  assign n15056 = n13173 & n15055 ;
  assign n15057 = n2988 & ~n5243 ;
  assign n15058 = n15057 ^ n14037 ^ 1'b0 ;
  assign n15059 = n6161 ^ n1212 ^ 1'b0 ;
  assign n15060 = n496 | n15059 ;
  assign n15061 = ( n148 & n1656 ) | ( n148 & ~n2982 ) | ( n1656 & ~n2982 ) ;
  assign n15062 = ~n14843 & n15061 ;
  assign n15063 = ~n15060 & n15062 ;
  assign n15064 = ( n3392 & n9371 ) | ( n3392 & ~n10129 ) | ( n9371 & ~n10129 ) ;
  assign n15065 = ~n2025 & n5143 ;
  assign n15066 = n685 | n11454 ;
  assign n15067 = n10066 | n15066 ;
  assign n15069 = n290 & ~n6959 ;
  assign n15070 = n15069 ^ n4717 ^ 1'b0 ;
  assign n15068 = ( n286 & n2660 ) | ( n286 & n3368 ) | ( n2660 & n3368 ) ;
  assign n15071 = n15070 ^ n15068 ^ n12509 ;
  assign n15074 = ~n2345 & n3474 ;
  assign n15075 = n4792 & n15074 ;
  assign n15072 = ~n274 & n2370 ;
  assign n15073 = n15072 ^ n796 ^ 1'b0 ;
  assign n15076 = n15075 ^ n15073 ^ n4546 ;
  assign n15077 = n15076 ^ n6612 ^ 1'b0 ;
  assign n15078 = n15071 & n15077 ;
  assign n15079 = n1868 & ~n6043 ;
  assign n15080 = n6398 & n14092 ;
  assign n15081 = ( ~n10259 & n10376 ) | ( ~n10259 & n14424 ) | ( n10376 & n14424 ) ;
  assign n15082 = n1542 ^ n1463 ^ 1'b0 ;
  assign n15083 = ~n15081 & n15082 ;
  assign n15084 = n2653 & n9310 ;
  assign n15085 = ~n15083 & n15084 ;
  assign n15086 = n7968 ^ n5745 ^ 1'b0 ;
  assign n15087 = n786 & n15086 ;
  assign n15088 = n15087 ^ n11821 ^ 1'b0 ;
  assign n15089 = n5278 ^ n4891 ^ n395 ;
  assign n15090 = n4290 & n15089 ;
  assign n15091 = n15088 & n15090 ;
  assign n15092 = ~n732 & n8854 ;
  assign n15093 = n13198 & ~n15092 ;
  assign n15094 = n7834 ^ x118 ^ 1'b0 ;
  assign n15095 = n15093 & ~n15094 ;
  assign n15096 = n15095 ^ n10259 ^ n4032 ;
  assign n15097 = ( x38 & n3533 ) | ( x38 & ~n15096 ) | ( n3533 & ~n15096 ) ;
  assign n15098 = n13847 ^ n4073 ^ 1'b0 ;
  assign n15099 = n15097 & n15098 ;
  assign n15100 = n2083 | n12517 ;
  assign n15101 = ( n5502 & n5514 ) | ( n5502 & ~n8626 ) | ( n5514 & ~n8626 ) ;
  assign n15102 = n15101 ^ n5494 ^ n2730 ;
  assign n15103 = ~n7572 & n8872 ;
  assign n15104 = n15103 ^ n4224 ^ 1'b0 ;
  assign n15105 = n1876 & ~n14551 ;
  assign n15106 = ~n9527 & n15105 ;
  assign n15107 = n5259 ^ n3792 ^ n1680 ;
  assign n15108 = ~n15106 & n15107 ;
  assign n15109 = n15108 ^ n143 ^ 1'b0 ;
  assign n15110 = ~n10009 & n12024 ;
  assign n15111 = ( ~n2903 & n12209 ) | ( ~n2903 & n15110 ) | ( n12209 & n15110 ) ;
  assign n15112 = n1564 & n10180 ;
  assign n15113 = ~x79 & n3334 ;
  assign n15114 = n15113 ^ n12405 ^ 1'b0 ;
  assign n15115 = n3991 | n5079 ;
  assign n15116 = n3876 & ~n15115 ;
  assign n15117 = n627 & n15116 ;
  assign n15118 = n10271 & n15117 ;
  assign n15119 = n1819 | n11963 ;
  assign n15120 = n320 | n15119 ;
  assign n15121 = ( n324 & n3358 ) | ( n324 & ~n4779 ) | ( n3358 & ~n4779 ) ;
  assign n15122 = n15121 ^ n4478 ^ 1'b0 ;
  assign n15123 = n6009 & n15122 ;
  assign n15124 = n13388 & n15123 ;
  assign n15125 = n15124 ^ n1435 ^ 1'b0 ;
  assign n15126 = n15125 ^ n3109 ^ 1'b0 ;
  assign n15127 = n6889 ^ n6444 ^ 1'b0 ;
  assign n15128 = n9838 | n15127 ;
  assign n15129 = n4172 | n4264 ;
  assign n15130 = n1890 | n13112 ;
  assign n15131 = n15129 & ~n15130 ;
  assign n15132 = n15131 ^ n13006 ^ n8667 ;
  assign n15134 = x99 & ~n660 ;
  assign n15135 = n15134 ^ n9441 ^ 1'b0 ;
  assign n15136 = n15135 ^ n289 ^ 1'b0 ;
  assign n15137 = n9233 & ~n15136 ;
  assign n15133 = n6157 ^ n947 ^ n803 ;
  assign n15138 = n15137 ^ n15133 ^ 1'b0 ;
  assign n15139 = n3699 | n15138 ;
  assign n15140 = ( n3488 & n3880 ) | ( n3488 & ~n7549 ) | ( n3880 & ~n7549 ) ;
  assign n15141 = n15140 ^ n2469 ^ 1'b0 ;
  assign n15142 = n8813 ^ n1919 ^ 1'b0 ;
  assign n15143 = n6444 | n15142 ;
  assign n15144 = n10031 | n15143 ;
  assign n15145 = ~n15141 & n15144 ;
  assign n15146 = n7744 | n14578 ;
  assign n15147 = n15146 ^ n3971 ^ 1'b0 ;
  assign n15148 = ( n2512 & n8355 ) | ( n2512 & ~n12552 ) | ( n8355 & ~n12552 ) ;
  assign n15150 = ~n781 & n2815 ;
  assign n15149 = n10640 ^ n4184 ^ n1767 ;
  assign n15151 = n15150 ^ n15149 ^ n7892 ;
  assign n15152 = ( n4714 & n15148 ) | ( n4714 & n15151 ) | ( n15148 & n15151 ) ;
  assign n15156 = ~n2246 & n2804 ;
  assign n15157 = ~n4656 & n15156 ;
  assign n15158 = n307 | n15157 ;
  assign n15159 = n15158 ^ n6586 ^ 1'b0 ;
  assign n15160 = n15159 ^ n3029 ^ 1'b0 ;
  assign n15153 = ( ~n2126 & n3442 ) | ( ~n2126 & n7711 ) | ( n3442 & n7711 ) ;
  assign n15154 = n15153 ^ n2780 ^ 1'b0 ;
  assign n15155 = ~n784 & n15154 ;
  assign n15161 = n15160 ^ n15155 ^ n14853 ;
  assign n15164 = n13052 ^ n9837 ^ 1'b0 ;
  assign n15165 = n3545 | n15164 ;
  assign n15162 = n10969 & n12477 ;
  assign n15163 = n15162 ^ n11811 ^ x17 ;
  assign n15166 = n15165 ^ n15163 ^ 1'b0 ;
  assign n15167 = n8489 & ~n9482 ;
  assign n15168 = n15167 ^ n1763 ^ 1'b0 ;
  assign n15169 = n15168 ^ n4636 ^ n2760 ;
  assign n15170 = n8502 ^ n5079 ^ 1'b0 ;
  assign n15171 = n9588 ^ n3923 ^ 1'b0 ;
  assign n15172 = ~n9308 & n15171 ;
  assign n15173 = n15172 ^ n5096 ^ n3582 ;
  assign n15174 = ( n606 & ~n5634 ) | ( n606 & n5919 ) | ( ~n5634 & n5919 ) ;
  assign n15175 = n1104 & n5417 ;
  assign n15176 = n15174 & n15175 ;
  assign n15177 = n15176 ^ n5571 ^ n4946 ;
  assign n15178 = n8974 ^ n2741 ^ 1'b0 ;
  assign n15179 = n4219 ^ n2247 ^ 1'b0 ;
  assign n15180 = n15179 ^ n397 ^ 1'b0 ;
  assign n15181 = n6668 | n15180 ;
  assign n15182 = ( n5092 & n9225 ) | ( n5092 & n11666 ) | ( n9225 & n11666 ) ;
  assign n15183 = n15182 ^ n8099 ^ 1'b0 ;
  assign n15184 = ~n1159 & n3792 ;
  assign n15185 = n15035 ^ n4103 ^ 1'b0 ;
  assign n15186 = n4716 & n12612 ;
  assign n15187 = n8785 | n10323 ;
  assign n15188 = n2138 | n2411 ;
  assign n15189 = n2025 & ~n15188 ;
  assign n15190 = n15189 ^ n7219 ^ 1'b0 ;
  assign n15191 = ~n10024 & n15190 ;
  assign n15192 = n629 & n10148 ;
  assign n15193 = n15192 ^ n5379 ^ 1'b0 ;
  assign n15194 = ( ~n1417 & n6066 ) | ( ~n1417 & n15193 ) | ( n6066 & n15193 ) ;
  assign n15195 = n15191 & ~n15194 ;
  assign n15196 = ( n3182 & n4404 ) | ( n3182 & ~n15195 ) | ( n4404 & ~n15195 ) ;
  assign n15197 = n15196 ^ n9018 ^ 1'b0 ;
  assign n15198 = n15187 | n15197 ;
  assign n15199 = n1322 & n1450 ;
  assign n15200 = n15198 & n15199 ;
  assign n15201 = n8634 & ~n14152 ;
  assign n15202 = n6605 & ~n11725 ;
  assign n15203 = n8499 ^ n1260 ^ 1'b0 ;
  assign n15204 = ( n2034 & ~n2196 ) | ( n2034 & n15203 ) | ( ~n2196 & n15203 ) ;
  assign n15205 = n2217 & n15204 ;
  assign n15206 = n7354 & ~n15205 ;
  assign n15207 = n1726 & n2813 ;
  assign n15208 = n12231 | n15207 ;
  assign n15209 = n15208 ^ n2344 ^ 1'b0 ;
  assign n15210 = ~n4430 & n12109 ;
  assign n15211 = ~n2721 & n15210 ;
  assign n15212 = ~n2107 & n5395 ;
  assign n15213 = ~n6264 & n15212 ;
  assign n15214 = ~n10678 & n15213 ;
  assign n15215 = n10231 ^ n935 ^ 1'b0 ;
  assign n15216 = ~n11448 & n13658 ;
  assign n15217 = ~n4281 & n15216 ;
  assign n15218 = n15217 ^ n10509 ^ n5910 ;
  assign n15219 = n154 & ~n2180 ;
  assign n15220 = n7213 | n15219 ;
  assign n15224 = n5495 ^ n1362 ^ 1'b0 ;
  assign n15225 = ( ~n767 & n1636 ) | ( ~n767 & n15224 ) | ( n1636 & n15224 ) ;
  assign n15226 = n15225 ^ n7276 ^ 1'b0 ;
  assign n15221 = ( n4269 & n4678 ) | ( n4269 & ~n12779 ) | ( n4678 & ~n12779 ) ;
  assign n15222 = n15221 ^ n12085 ^ 1'b0 ;
  assign n15223 = ~n7642 & n15222 ;
  assign n15227 = n15226 ^ n15223 ^ 1'b0 ;
  assign n15233 = ~n2477 & n12873 ;
  assign n15234 = n15233 ^ x6 ^ 1'b0 ;
  assign n15235 = n15234 ^ n12428 ^ 1'b0 ;
  assign n15236 = n309 & ~n15235 ;
  assign n15228 = n7965 ^ n5235 ^ 1'b0 ;
  assign n15229 = ( n1329 & n1791 ) | ( n1329 & ~n6419 ) | ( n1791 & ~n6419 ) ;
  assign n15230 = ~n360 & n15229 ;
  assign n15231 = n15230 ^ n8158 ^ 1'b0 ;
  assign n15232 = n15228 & ~n15231 ;
  assign n15237 = n15236 ^ n15232 ^ 1'b0 ;
  assign n15238 = ( n5337 & ~n10412 ) | ( n5337 & n15123 ) | ( ~n10412 & n15123 ) ;
  assign n15242 = n13060 ^ n8294 ^ 1'b0 ;
  assign n15239 = n6471 | n10044 ;
  assign n15240 = ~n2715 & n2808 ;
  assign n15241 = n15239 & n15240 ;
  assign n15243 = n15242 ^ n15241 ^ n9982 ;
  assign n15244 = ( n10745 & n15238 ) | ( n10745 & n15243 ) | ( n15238 & n15243 ) ;
  assign n15245 = n927 | n2736 ;
  assign n15246 = n15245 ^ n2189 ^ 1'b0 ;
  assign n15247 = n6114 ^ n4495 ^ 1'b0 ;
  assign n15248 = ( n5126 & n8441 ) | ( n5126 & ~n15247 ) | ( n8441 & ~n15247 ) ;
  assign n15249 = n7577 | n13560 ;
  assign n15250 = n10340 ^ n6171 ^ 1'b0 ;
  assign n15251 = n2811 & ~n15250 ;
  assign n15252 = ~x54 & n2703 ;
  assign n15253 = n5762 ^ n3113 ^ 1'b0 ;
  assign n15254 = n12961 ^ n788 ^ 1'b0 ;
  assign n15255 = n15254 ^ n6092 ^ 1'b0 ;
  assign n15256 = n7338 ^ n5008 ^ 1'b0 ;
  assign n15257 = ( n3616 & ~n7448 ) | ( n3616 & n13576 ) | ( ~n7448 & n13576 ) ;
  assign n15258 = n7980 ^ n7890 ^ n6830 ;
  assign n15259 = n15005 ^ n8209 ^ 1'b0 ;
  assign n15260 = n7277 & n9736 ;
  assign n15262 = n2481 ^ n1410 ^ 1'b0 ;
  assign n15261 = n8483 | n14026 ;
  assign n15263 = n15262 ^ n15261 ^ 1'b0 ;
  assign n15264 = n3647 & ~n15263 ;
  assign n15265 = ~n5003 & n15264 ;
  assign n15266 = n5755 | n11432 ;
  assign n15267 = n15266 ^ n11945 ^ 1'b0 ;
  assign n15268 = n15267 ^ n4021 ^ 1'b0 ;
  assign n15271 = n5823 ^ n3408 ^ 1'b0 ;
  assign n15269 = n945 | n3650 ;
  assign n15270 = ( n4584 & ~n11158 ) | ( n4584 & n15269 ) | ( ~n11158 & n15269 ) ;
  assign n15272 = n15271 ^ n15270 ^ n9790 ;
  assign n15273 = n8086 ^ n2923 ^ 1'b0 ;
  assign n15274 = n7227 & n15273 ;
  assign n15275 = n15274 ^ n5387 ^ n4658 ;
  assign n15276 = n6137 | n11936 ;
  assign n15277 = n15276 ^ n10381 ^ 1'b0 ;
  assign n15278 = ~n2296 & n15277 ;
  assign n15279 = n4107 & ~n10176 ;
  assign n15280 = n15279 ^ n8500 ^ 1'b0 ;
  assign n15281 = n10010 & n13901 ;
  assign n15282 = ~n701 & n15281 ;
  assign n15283 = ( n181 & n1554 ) | ( n181 & n12096 ) | ( n1554 & n12096 ) ;
  assign n15284 = ( n236 & n1029 ) | ( n236 & n15283 ) | ( n1029 & n15283 ) ;
  assign n15285 = ~n15282 & n15284 ;
  assign n15286 = n1910 ^ n799 ^ 1'b0 ;
  assign n15287 = ( n173 & ~n9887 ) | ( n173 & n15286 ) | ( ~n9887 & n15286 ) ;
  assign n15288 = n2159 ^ n2070 ^ 1'b0 ;
  assign n15289 = n10549 & n15288 ;
  assign n15290 = n9940 & n15289 ;
  assign n15291 = ~n3865 & n15290 ;
  assign n15292 = n7691 | n15291 ;
  assign n15293 = n1362 & ~n15292 ;
  assign n15294 = ( ~n15285 & n15287 ) | ( ~n15285 & n15293 ) | ( n15287 & n15293 ) ;
  assign n15295 = ~n1423 & n7234 ;
  assign n15296 = n2149 ^ n1470 ^ 1'b0 ;
  assign n15297 = n2326 & n13796 ;
  assign n15298 = ~n9988 & n15297 ;
  assign n15299 = ( ~n1331 & n15296 ) | ( ~n1331 & n15298 ) | ( n15296 & n15298 ) ;
  assign n15300 = ~n2487 & n6203 ;
  assign n15301 = ~n15299 & n15300 ;
  assign n15302 = ~n2889 & n3236 ;
  assign n15303 = ~n9697 & n15302 ;
  assign n15304 = n15303 ^ n4504 ^ n3381 ;
  assign n15305 = n357 & ~n10046 ;
  assign n15306 = x49 | n938 ;
  assign n15307 = n15306 ^ n7923 ^ 1'b0 ;
  assign n15308 = n12451 | n12709 ;
  assign n15309 = ~n10451 & n13065 ;
  assign n15311 = n2177 & n3709 ;
  assign n15312 = n15311 ^ n7172 ^ 1'b0 ;
  assign n15313 = n8014 ^ n3091 ^ 1'b0 ;
  assign n15314 = n15312 | n15313 ;
  assign n15310 = n4131 ^ n668 ^ 1'b0 ;
  assign n15315 = n15314 ^ n15310 ^ n9781 ;
  assign n15316 = n6537 & n7532 ;
  assign n15317 = n6888 & n7794 ;
  assign n15318 = ~n1402 & n6628 ;
  assign n15319 = n15318 ^ n4255 ^ n977 ;
  assign n15320 = n14187 ^ n4737 ^ 1'b0 ;
  assign n15321 = n193 & ~n15320 ;
  assign n15322 = n9091 & n15321 ;
  assign n15323 = n15319 & n15322 ;
  assign n15324 = n2839 | n15323 ;
  assign n15325 = n915 | n15324 ;
  assign n15326 = n9833 ^ n1487 ^ 1'b0 ;
  assign n15327 = ~n12664 & n15326 ;
  assign n15328 = n3438 & ~n15327 ;
  assign n15329 = n15328 ^ n9782 ^ 1'b0 ;
  assign n15330 = n4271 & ~n15329 ;
  assign n15331 = n15205 ^ n1473 ^ n950 ;
  assign n15332 = n11030 & n13578 ;
  assign n15333 = n15332 ^ n2172 ^ 1'b0 ;
  assign n15334 = n10098 ^ n7473 ^ 1'b0 ;
  assign n15335 = n6085 & ~n15334 ;
  assign n15336 = n4753 | n14976 ;
  assign n15337 = n8929 ^ n8040 ^ 1'b0 ;
  assign n15338 = n15336 & n15337 ;
  assign n15339 = ~n5293 & n11449 ;
  assign n15340 = n810 ^ n169 ^ 1'b0 ;
  assign n15341 = n5060 & ~n15340 ;
  assign n15342 = n15341 ^ n7008 ^ 1'b0 ;
  assign n15343 = n15342 ^ n5300 ^ 1'b0 ;
  assign n15344 = n15339 & n15343 ;
  assign n15345 = n1750 & n3059 ;
  assign n15346 = n11042 & n15345 ;
  assign n15347 = n15346 ^ n881 ^ 1'b0 ;
  assign n15348 = n15344 & ~n15347 ;
  assign n15349 = ( n391 & n5126 ) | ( n391 & ~n13110 ) | ( n5126 & ~n13110 ) ;
  assign n15350 = ( ~n2499 & n6553 ) | ( ~n2499 & n15349 ) | ( n6553 & n15349 ) ;
  assign n15351 = n5230 & n13863 ;
  assign n15352 = n15350 & n15351 ;
  assign n15353 = n1425 & ~n12178 ;
  assign n15354 = ~n5153 & n15353 ;
  assign n15355 = n4432 ^ n3434 ^ 1'b0 ;
  assign n15356 = n2508 & n7226 ;
  assign n15357 = n15356 ^ n6578 ^ n4257 ;
  assign n15358 = n1708 | n10488 ;
  assign n15359 = n15358 ^ n1573 ^ 1'b0 ;
  assign n15360 = ~n4495 & n15359 ;
  assign n15361 = n4542 & n15360 ;
  assign n15362 = n15361 ^ n2467 ^ 1'b0 ;
  assign n15363 = ~n597 & n4637 ;
  assign n15364 = ~n14158 & n15363 ;
  assign n15365 = n4704 & ~n14570 ;
  assign n15366 = ( ~n5954 & n15364 ) | ( ~n5954 & n15365 ) | ( n15364 & n15365 ) ;
  assign n15367 = n14750 ^ n13547 ^ 1'b0 ;
  assign n15368 = n12069 ^ n9406 ^ n6106 ;
  assign n15369 = n8737 ^ n8511 ^ 1'b0 ;
  assign n15370 = ~n194 & n12641 ;
  assign n15371 = ~n2121 & n9174 ;
  assign n15372 = n1135 ^ n248 ^ 1'b0 ;
  assign n15373 = n950 | n15372 ;
  assign n15374 = n8908 ^ n4271 ^ 1'b0 ;
  assign n15375 = n870 & ~n15374 ;
  assign n15376 = ~n15373 & n15375 ;
  assign n15377 = n15376 ^ n11591 ^ n4419 ;
  assign n15378 = n5076 & ~n15377 ;
  assign n15379 = n15378 ^ x107 ^ 1'b0 ;
  assign n15383 = n13360 | n14488 ;
  assign n15380 = ~n3327 & n7360 ;
  assign n15381 = n11875 ^ n8833 ^ n3679 ;
  assign n15382 = n15380 & ~n15381 ;
  assign n15384 = n15383 ^ n15382 ^ 1'b0 ;
  assign n15385 = n768 & n1648 ;
  assign n15386 = n13416 & n15385 ;
  assign n15388 = n2905 ^ n2248 ^ 1'b0 ;
  assign n15387 = n11524 ^ n2724 ^ n1913 ;
  assign n15389 = n15388 ^ n15387 ^ n12350 ;
  assign n15390 = ( ~n209 & n617 ) | ( ~n209 & n3597 ) | ( n617 & n3597 ) ;
  assign n15391 = ~n3595 & n15390 ;
  assign n15392 = n15391 ^ x13 ^ 1'b0 ;
  assign n15393 = ~n1483 & n15392 ;
  assign n15394 = n5955 ^ n5907 ^ 1'b0 ;
  assign n15395 = n5670 ^ n2557 ^ 1'b0 ;
  assign n15396 = x54 & n15395 ;
  assign n15397 = n5705 ^ n1665 ^ 1'b0 ;
  assign n15398 = ~n13480 & n15397 ;
  assign n15399 = ( ~n7758 & n15396 ) | ( ~n7758 & n15398 ) | ( n15396 & n15398 ) ;
  assign n15400 = n8611 & n14179 ;
  assign n15401 = n2873 & n15400 ;
  assign n15403 = n6770 & n8626 ;
  assign n15402 = n13281 ^ n9940 ^ 1'b0 ;
  assign n15404 = n15403 ^ n15402 ^ 1'b0 ;
  assign n15405 = n3284 | n13710 ;
  assign n15406 = n4253 & ~n11885 ;
  assign n15407 = n8953 & n15406 ;
  assign n15410 = n2763 & ~n11086 ;
  assign n15411 = n14058 ^ n402 ^ 1'b0 ;
  assign n15412 = n14106 & n15411 ;
  assign n15413 = ~n11268 & n15412 ;
  assign n15414 = n15410 & n15413 ;
  assign n15408 = ( n1654 & n11387 ) | ( n1654 & n11464 ) | ( n11387 & n11464 ) ;
  assign n15409 = n8341 | n15408 ;
  assign n15415 = n15414 ^ n15409 ^ 1'b0 ;
  assign n15420 = n917 & n6428 ;
  assign n15421 = n15420 ^ n5752 ^ n1491 ;
  assign n15416 = n3529 ^ n1317 ^ 1'b0 ;
  assign n15417 = ( ~n1729 & n8119 ) | ( ~n1729 & n15416 ) | ( n8119 & n15416 ) ;
  assign n15418 = n15417 ^ n9652 ^ n7918 ;
  assign n15419 = n15418 ^ n11779 ^ 1'b0 ;
  assign n15422 = n15421 ^ n15419 ^ n13306 ;
  assign n15423 = n810 | n1131 ;
  assign n15424 = n15423 ^ n11975 ^ 1'b0 ;
  assign n15425 = n7440 ^ n3578 ^ 1'b0 ;
  assign n15426 = n1124 & ~n15425 ;
  assign n15427 = n5977 | n9955 ;
  assign n15428 = n15427 ^ n7956 ^ 1'b0 ;
  assign n15431 = n9678 ^ n8366 ^ 1'b0 ;
  assign n15429 = n7502 ^ n3790 ^ 1'b0 ;
  assign n15430 = ~n12507 & n15429 ;
  assign n15432 = n15431 ^ n15430 ^ n8810 ;
  assign n15433 = n15432 ^ n11031 ^ n7144 ;
  assign n15434 = n15053 ^ n4748 ^ n1478 ;
  assign n15435 = n9734 ^ n2507 ^ 1'b0 ;
  assign n15436 = n12223 & ~n15435 ;
  assign n15437 = n4310 | n15436 ;
  assign n15440 = ( n4096 & n5241 ) | ( n4096 & ~n10050 ) | ( n5241 & ~n10050 ) ;
  assign n15441 = ( n7796 & n9607 ) | ( n7796 & ~n15440 ) | ( n9607 & ~n15440 ) ;
  assign n15438 = n4610 & n7021 ;
  assign n15439 = n15438 ^ n14001 ^ 1'b0 ;
  assign n15442 = n15441 ^ n15439 ^ n5821 ;
  assign n15443 = ( x100 & n7701 ) | ( x100 & n15213 ) | ( n7701 & n15213 ) ;
  assign n15444 = n13251 & n14585 ;
  assign n15445 = ~n4478 & n15444 ;
  assign n15446 = n15445 ^ n11181 ^ 1'b0 ;
  assign n15447 = n8697 ^ n1305 ^ 1'b0 ;
  assign n15448 = n438 | n15447 ;
  assign n15449 = ( n816 & n5111 ) | ( n816 & ~n7839 ) | ( n5111 & ~n7839 ) ;
  assign n15450 = n15449 ^ x63 ^ 1'b0 ;
  assign n15451 = x37 & n11500 ;
  assign n15452 = n15451 ^ n2326 ^ 1'b0 ;
  assign n15453 = n5165 | n15452 ;
  assign n15454 = n14855 & ~n15453 ;
  assign n15455 = x77 & ~n3390 ;
  assign n15456 = ~n1300 & n15455 ;
  assign n15457 = n15456 ^ n191 ^ 1'b0 ;
  assign n15458 = ~n1747 & n5669 ;
  assign n15459 = n1747 & n15458 ;
  assign n15460 = n1123 | n1299 ;
  assign n15461 = n1299 & ~n15460 ;
  assign n15462 = x39 & n15461 ;
  assign n15463 = n15459 | n15462 ;
  assign n15464 = n15457 & ~n15463 ;
  assign n15465 = n3800 | n9928 ;
  assign n15466 = n6129 & ~n11603 ;
  assign n15467 = ~n331 & n15466 ;
  assign n15468 = n2179 & ~n3538 ;
  assign n15469 = n1463 & ~n13205 ;
  assign n15470 = n7392 & n15469 ;
  assign n15471 = n1748 & n15470 ;
  assign n15472 = n15471 ^ n8418 ^ 1'b0 ;
  assign n15473 = n13853 ^ n11181 ^ x17 ;
  assign n15474 = n1860 & ~n3621 ;
  assign n15475 = n15474 ^ n1653 ^ 1'b0 ;
  assign n15476 = x44 & ~n13624 ;
  assign n15477 = ~n7627 & n15476 ;
  assign n15478 = ( n3856 & n10270 ) | ( n3856 & n11891 ) | ( n10270 & n11891 ) ;
  assign n15479 = ( n749 & n8552 ) | ( n749 & n15478 ) | ( n8552 & n15478 ) ;
  assign n15480 = ( n974 & n13258 ) | ( n974 & ~n13828 ) | ( n13258 & ~n13828 ) ;
  assign n15481 = n15480 ^ n6691 ^ 1'b0 ;
  assign n15482 = n14392 ^ n10211 ^ 1'b0 ;
  assign n15483 = n3241 & ~n15189 ;
  assign n15484 = ~n7765 & n15483 ;
  assign n15487 = n11143 ^ n5130 ^ n4095 ;
  assign n15485 = n5394 ^ n1433 ^ 1'b0 ;
  assign n15486 = n11360 & n15485 ;
  assign n15488 = n15487 ^ n15486 ^ 1'b0 ;
  assign n15491 = n10488 ^ n10087 ^ n7354 ;
  assign n15492 = n15491 ^ n6659 ^ n3126 ;
  assign n15493 = n15492 ^ n2625 ^ 1'b0 ;
  assign n15489 = n2034 & ~n6125 ;
  assign n15490 = n15489 ^ n13553 ^ 1'b0 ;
  assign n15494 = n15493 ^ n15490 ^ n13713 ;
  assign n15495 = n8380 ^ n5050 ^ 1'b0 ;
  assign n15496 = n2853 & ~n12725 ;
  assign n15497 = ( ~n6309 & n15495 ) | ( ~n6309 & n15496 ) | ( n15495 & n15496 ) ;
  assign n15498 = n5599 & ~n15497 ;
  assign n15499 = n5931 | n15498 ;
  assign n15500 = n4844 | n15499 ;
  assign n15503 = n11004 ^ n2275 ^ n1448 ;
  assign n15501 = n1183 ^ n288 ^ 1'b0 ;
  assign n15502 = ~n5641 & n15501 ;
  assign n15504 = n15503 ^ n15502 ^ 1'b0 ;
  assign n15505 = ~n2151 & n15504 ;
  assign n15506 = n4710 | n15505 ;
  assign n15507 = n15506 ^ n14711 ^ 1'b0 ;
  assign n15508 = n13552 ^ n186 ^ 1'b0 ;
  assign n15509 = n9703 ^ n3855 ^ 1'b0 ;
  assign n15510 = n2422 ^ n1171 ^ n1053 ;
  assign n15511 = n13869 ^ n2145 ^ n1538 ;
  assign n15512 = ~n1895 & n9136 ;
  assign n15513 = ~n9013 & n15512 ;
  assign n15514 = n9122 ^ n2499 ^ 1'b0 ;
  assign n15515 = n164 | n15514 ;
  assign n15516 = n5613 & ~n15515 ;
  assign n15517 = ( n2820 & ~n4156 ) | ( n2820 & n5013 ) | ( ~n4156 & n5013 ) ;
  assign n15518 = n9091 ^ n4269 ^ 1'b0 ;
  assign n15519 = n15517 & ~n15518 ;
  assign n15520 = ( n3517 & n7886 ) | ( n3517 & ~n15519 ) | ( n7886 & ~n15519 ) ;
  assign n15521 = n14760 ^ n14314 ^ 1'b0 ;
  assign n15522 = n9501 ^ n5558 ^ 1'b0 ;
  assign n15523 = n1143 | n6137 ;
  assign n15524 = n15523 ^ n14519 ^ 1'b0 ;
  assign n15525 = n15524 ^ n6282 ^ 1'b0 ;
  assign n15526 = n15522 & n15525 ;
  assign n15527 = n14591 ^ n12888 ^ n10653 ;
  assign n15528 = n14775 ^ n3534 ^ 1'b0 ;
  assign n15529 = n7077 ^ n4489 ^ x37 ;
  assign n15530 = n15529 ^ n7307 ^ 1'b0 ;
  assign n15531 = n6872 & n15530 ;
  assign n15532 = n8617 ^ n4003 ^ 1'b0 ;
  assign n15534 = n4392 ^ n1892 ^ 1'b0 ;
  assign n15533 = n4092 | n5328 ;
  assign n15535 = n15534 ^ n15533 ^ 1'b0 ;
  assign n15536 = ( ~n6208 & n6621 ) | ( ~n6208 & n8616 ) | ( n6621 & n8616 ) ;
  assign n15537 = n15536 ^ n7174 ^ 1'b0 ;
  assign n15538 = ~n15535 & n15537 ;
  assign n15539 = ( n3974 & n13752 ) | ( n3974 & n15538 ) | ( n13752 & n15538 ) ;
  assign n15540 = n7463 ^ n3317 ^ 1'b0 ;
  assign n15541 = ~n3012 & n15540 ;
  assign n15542 = n4462 & n15541 ;
  assign n15543 = n13128 & n15542 ;
  assign n15544 = ~n5609 & n5999 ;
  assign n15545 = n3790 & n15544 ;
  assign n15546 = n15545 ^ n13361 ^ n4699 ;
  assign n15547 = n928 | n5423 ;
  assign n15548 = n8112 | n15547 ;
  assign n15549 = n15548 ^ n11383 ^ 1'b0 ;
  assign n15550 = n13961 & n15549 ;
  assign n15551 = ~n15546 & n15550 ;
  assign n15552 = n15551 ^ n8945 ^ 1'b0 ;
  assign n15553 = n11727 ^ n8010 ^ n1796 ;
  assign n15554 = n12808 ^ n3748 ^ n2158 ;
  assign n15555 = n5777 | n9831 ;
  assign n15556 = n15555 ^ n13002 ^ n11352 ;
  assign n15557 = n11116 & ~n15135 ;
  assign n15558 = n3677 & n14620 ;
  assign n15559 = n15558 ^ n9366 ^ 1'b0 ;
  assign n15560 = ( n848 & n2224 ) | ( n848 & n7763 ) | ( n2224 & n7763 ) ;
  assign n15561 = ~n3991 & n5117 ;
  assign n15562 = ( n579 & n12953 ) | ( n579 & n15561 ) | ( n12953 & n15561 ) ;
  assign n15563 = n5352 ^ n3237 ^ 1'b0 ;
  assign n15564 = n10110 & ~n15563 ;
  assign n15565 = n15564 ^ n7990 ^ 1'b0 ;
  assign n15566 = n11165 | n15565 ;
  assign n15567 = ~n4126 & n4156 ;
  assign n15568 = n15566 & n15567 ;
  assign n15569 = n6889 | n10199 ;
  assign n15570 = n15569 ^ n1731 ^ 1'b0 ;
  assign n15571 = n10101 & ~n15037 ;
  assign n15572 = n15037 & n15571 ;
  assign n15573 = n9215 ^ n7448 ^ n3001 ;
  assign n15574 = n10423 ^ n6740 ^ n4720 ;
  assign n15575 = n10453 & n15574 ;
  assign n15576 = ~n10453 & n15575 ;
  assign n15577 = n6968 ^ n2981 ^ 1'b0 ;
  assign n15578 = ( n368 & n2640 ) | ( n368 & n13922 ) | ( n2640 & n13922 ) ;
  assign n15579 = n3248 ^ n3218 ^ 1'b0 ;
  assign n15580 = n9187 & ~n15579 ;
  assign n15581 = n9199 & n15580 ;
  assign n15582 = ~n7395 & n15581 ;
  assign n15583 = n327 & ~n2470 ;
  assign n15584 = n15583 ^ n8840 ^ 1'b0 ;
  assign n15585 = n15584 ^ n5755 ^ n2750 ;
  assign n15586 = ( ~n5297 & n15582 ) | ( ~n5297 & n15585 ) | ( n15582 & n15585 ) ;
  assign n15587 = ( n2285 & n12561 ) | ( n2285 & ~n14499 ) | ( n12561 & ~n14499 ) ;
  assign n15588 = ( n3828 & n6261 ) | ( n3828 & n15587 ) | ( n6261 & n15587 ) ;
  assign n15589 = n15588 ^ n8819 ^ n8527 ;
  assign n15590 = n7923 & ~n12600 ;
  assign n15591 = n6874 ^ n4906 ^ 1'b0 ;
  assign n15592 = n13605 | n15591 ;
  assign n15598 = n6730 ^ n6258 ^ 1'b0 ;
  assign n15593 = n8565 ^ n1802 ^ 1'b0 ;
  assign n15594 = n1116 & ~n15593 ;
  assign n15595 = n2492 & ~n5563 ;
  assign n15596 = ~n15594 & n15595 ;
  assign n15597 = n10512 | n15596 ;
  assign n15599 = n15598 ^ n15597 ^ 1'b0 ;
  assign n15600 = n13168 ^ n1725 ^ 1'b0 ;
  assign n15601 = ~n5024 & n15600 ;
  assign n15602 = n2212 & ~n9538 ;
  assign n15603 = n13484 | n15602 ;
  assign n15604 = n6623 & ~n7821 ;
  assign n15605 = ( n506 & ~n2947 ) | ( n506 & n5126 ) | ( ~n2947 & n5126 ) ;
  assign n15606 = n4975 ^ n3132 ^ 1'b0 ;
  assign n15607 = ~n15605 & n15606 ;
  assign n15608 = ( n2930 & n12266 ) | ( n2930 & n15607 ) | ( n12266 & n15607 ) ;
  assign n15610 = n4295 | n4409 ;
  assign n15611 = n15610 ^ n5621 ^ 1'b0 ;
  assign n15612 = n15611 ^ n1327 ^ 1'b0 ;
  assign n15613 = n6855 ^ n5352 ^ 1'b0 ;
  assign n15614 = n15612 & n15613 ;
  assign n15609 = n9042 & n14475 ;
  assign n15615 = n15614 ^ n15609 ^ 1'b0 ;
  assign n15616 = ( ~n1196 & n4694 ) | ( ~n1196 & n15615 ) | ( n4694 & n15615 ) ;
  assign n15617 = n1845 & ~n11024 ;
  assign n15618 = n12428 & ~n14655 ;
  assign n15619 = ~n10241 & n15618 ;
  assign n15621 = n12814 ^ n958 ^ 1'b0 ;
  assign n15622 = n9020 & n15621 ;
  assign n15620 = n10223 & ~n13978 ;
  assign n15623 = n15622 ^ n15620 ^ 1'b0 ;
  assign n15624 = n1797 | n7930 ;
  assign n15626 = ( n2261 & ~n4375 ) | ( n2261 & n6620 ) | ( ~n4375 & n6620 ) ;
  assign n15627 = n14641 & ~n15626 ;
  assign n15625 = n6332 ^ n6272 ^ n2869 ;
  assign n15628 = n15627 ^ n15625 ^ 1'b0 ;
  assign n15629 = n8680 ^ n5412 ^ 1'b0 ;
  assign n15630 = n5980 ^ n4405 ^ 1'b0 ;
  assign n15631 = n1383 | n15630 ;
  assign n15632 = ( ~n9214 & n15629 ) | ( ~n9214 & n15631 ) | ( n15629 & n15631 ) ;
  assign n15633 = n6229 & n15632 ;
  assign n15634 = ( ~n2306 & n4393 ) | ( ~n2306 & n6474 ) | ( n4393 & n6474 ) ;
  assign n15635 = n15193 ^ n6283 ^ 1'b0 ;
  assign n15636 = n8082 & ~n15635 ;
  assign n15637 = n14510 ^ n5954 ^ 1'b0 ;
  assign n15638 = ( n4243 & n15636 ) | ( n4243 & ~n15637 ) | ( n15636 & ~n15637 ) ;
  assign n15639 = n3140 ^ x46 ^ 1'b0 ;
  assign n15640 = n11496 & n15639 ;
  assign n15641 = n15640 ^ n8312 ^ 1'b0 ;
  assign n15642 = n2567 | n4343 ;
  assign n15643 = ~n8685 & n15642 ;
  assign n15644 = ~n15641 & n15643 ;
  assign n15645 = n11643 | n13490 ;
  assign n15646 = n2121 & ~n3700 ;
  assign n15647 = n6729 ^ n6419 ^ n2431 ;
  assign n15648 = n15647 ^ n972 ^ 1'b0 ;
  assign n15649 = ~n4096 & n15648 ;
  assign n15650 = n8762 | n12214 ;
  assign n15651 = n7312 & ~n15650 ;
  assign n15652 = ~n7402 & n11465 ;
  assign n15653 = n8984 & n10815 ;
  assign n15655 = n1704 | n2467 ;
  assign n15656 = ( n10110 & n10536 ) | ( n10110 & n15655 ) | ( n10536 & n15655 ) ;
  assign n15654 = ( n7980 & ~n11211 ) | ( n7980 & n14166 ) | ( ~n11211 & n14166 ) ;
  assign n15657 = n15656 ^ n15654 ^ n8994 ;
  assign n15661 = n15491 ^ n10755 ^ n9536 ;
  assign n15658 = ~n2746 & n2822 ;
  assign n15659 = n9866 & n15658 ;
  assign n15660 = n15659 ^ n7719 ^ n7700 ;
  assign n15662 = n15661 ^ n15660 ^ 1'b0 ;
  assign n15665 = n3015 & ~n3320 ;
  assign n15664 = ~n6345 & n13364 ;
  assign n15666 = n15665 ^ n15664 ^ 1'b0 ;
  assign n15663 = n4543 | n11409 ;
  assign n15667 = n15666 ^ n15663 ^ n15474 ;
  assign n15668 = n11268 ^ n5385 ^ 1'b0 ;
  assign n15669 = ~n3666 & n15668 ;
  assign n15670 = n5838 ^ n3088 ^ 1'b0 ;
  assign n15671 = n15669 & ~n15670 ;
  assign n15672 = n15318 ^ n801 ^ 1'b0 ;
  assign n15673 = n286 & n15672 ;
  assign n15674 = n15673 ^ n9499 ^ 1'b0 ;
  assign n15675 = n15674 ^ n3470 ^ 1'b0 ;
  assign n15676 = n7130 & n15675 ;
  assign n15677 = ~n10209 & n15676 ;
  assign n15678 = n15677 ^ n5851 ^ 1'b0 ;
  assign n15679 = ( ~n521 & n13382 ) | ( ~n521 & n15678 ) | ( n13382 & n15678 ) ;
  assign n15680 = n365 | n12071 ;
  assign n15686 = n10169 | n14342 ;
  assign n15687 = n4329 & n15686 ;
  assign n15681 = n7557 & n12961 ;
  assign n15682 = n4627 & n15681 ;
  assign n15683 = n14997 | n15682 ;
  assign n15684 = ~n13213 & n15683 ;
  assign n15685 = n4887 | n15684 ;
  assign n15688 = n15687 ^ n15685 ^ 1'b0 ;
  assign n15689 = ( n3503 & n4486 ) | ( n3503 & ~n5484 ) | ( n4486 & ~n5484 ) ;
  assign n15690 = ~n6638 & n15689 ;
  assign n15691 = n15690 ^ n15246 ^ 1'b0 ;
  assign n15692 = n11246 ^ n4904 ^ 1'b0 ;
  assign n15693 = n3961 & ~n6576 ;
  assign n15694 = ~n12338 & n15693 ;
  assign n15695 = n15694 ^ n2273 ^ 1'b0 ;
  assign n15696 = ( x32 & ~n1356 ) | ( x32 & n15695 ) | ( ~n1356 & n15695 ) ;
  assign n15697 = n9632 & n15696 ;
  assign n15698 = n12463 ^ n5890 ^ 1'b0 ;
  assign n15699 = n5197 ^ n1003 ^ 1'b0 ;
  assign n15700 = n15699 ^ n14286 ^ n163 ;
  assign n15701 = n6278 | n7671 ;
  assign n15702 = n8539 | n15701 ;
  assign n15703 = ~n3704 & n15702 ;
  assign n15704 = ( n3615 & ~n6422 ) | ( n3615 & n15703 ) | ( ~n6422 & n15703 ) ;
  assign n15705 = ( ~n987 & n5660 ) | ( ~n987 & n11875 ) | ( n5660 & n11875 ) ;
  assign n15706 = n6439 & n11823 ;
  assign n15707 = ~n15705 & n15706 ;
  assign n15708 = n9914 ^ n3845 ^ 1'b0 ;
  assign n15709 = ( n13290 & n15707 ) | ( n13290 & n15708 ) | ( n15707 & n15708 ) ;
  assign n15710 = ~x74 & n3651 ;
  assign n15711 = n15710 ^ n582 ^ 1'b0 ;
  assign n15712 = n12081 | n15711 ;
  assign n15713 = n2524 | n15712 ;
  assign n15714 = n15079 ^ n11741 ^ 1'b0 ;
  assign n15715 = n143 & ~n15714 ;
  assign n15716 = n1475 & n15153 ;
  assign n15717 = ( n2774 & n7177 ) | ( n2774 & ~n12297 ) | ( n7177 & ~n12297 ) ;
  assign n15718 = n15717 ^ n9370 ^ n4402 ;
  assign n15719 = n12951 & ~n15718 ;
  assign n15720 = ~n8504 & n15719 ;
  assign n15721 = ~n3616 & n7437 ;
  assign n15722 = n15721 ^ n2275 ^ 1'b0 ;
  assign n15723 = ~n1791 & n15707 ;
  assign n15724 = n2937 & n15723 ;
  assign n15725 = ( ~n4154 & n15722 ) | ( ~n4154 & n15724 ) | ( n15722 & n15724 ) ;
  assign n15726 = n15725 ^ n5695 ^ n3534 ;
  assign n15727 = n10429 ^ n5741 ^ 1'b0 ;
  assign n15728 = n8310 & ~n15727 ;
  assign n15729 = n6720 | n13296 ;
  assign n15730 = n12406 ^ n10384 ^ n7119 ;
  assign n15731 = n9126 | n10147 ;
  assign n15732 = n15731 ^ n14179 ^ 1'b0 ;
  assign n15733 = n1175 & n5499 ;
  assign n15734 = n14858 & n15733 ;
  assign n15735 = n6916 & ~n15734 ;
  assign n15736 = n661 & n15735 ;
  assign n15737 = ~n4748 & n4772 ;
  assign n15738 = n15737 ^ n1985 ^ 1'b0 ;
  assign n15739 = n3099 & ~n15738 ;
  assign n15740 = ~n6991 & n7017 ;
  assign n15741 = ~n15739 & n15740 ;
  assign n15742 = n15736 & n15741 ;
  assign n15743 = n7631 & ~n9429 ;
  assign n15744 = n5225 & ~n15743 ;
  assign n15745 = ~n3038 & n8373 ;
  assign n15746 = n3735 & ~n15745 ;
  assign n15747 = n3752 & n15746 ;
  assign n15748 = n15744 | n15747 ;
  assign n15749 = n11990 ^ n3164 ^ n2833 ;
  assign n15750 = n12062 ^ n11539 ^ n6318 ;
  assign n15751 = n8194 & n15750 ;
  assign n15754 = n14572 ^ x115 ^ 1'b0 ;
  assign n15755 = n11050 & ~n15754 ;
  assign n15752 = n4717 ^ n3319 ^ 1'b0 ;
  assign n15753 = n9755 | n15752 ;
  assign n15756 = n15755 ^ n15753 ^ 1'b0 ;
  assign n15757 = n11380 ^ n8221 ^ 1'b0 ;
  assign n15758 = n3323 & n13284 ;
  assign n15759 = n14827 ^ n4566 ^ 1'b0 ;
  assign n15760 = n15758 | n15759 ;
  assign n15761 = n1183 | n9455 ;
  assign n15762 = n3474 | n15761 ;
  assign n15763 = n4308 & n5895 ;
  assign n15764 = ~n15762 & n15763 ;
  assign n15765 = n7854 ^ n2419 ^ 1'b0 ;
  assign n15766 = n180 & n15765 ;
  assign n15768 = n7351 ^ n6115 ^ 1'b0 ;
  assign n15767 = ( n2472 & n4370 ) | ( n2472 & ~n10594 ) | ( n4370 & ~n10594 ) ;
  assign n15769 = n15768 ^ n15767 ^ 1'b0 ;
  assign n15770 = n5758 & n9763 ;
  assign n15771 = ~n15769 & n15770 ;
  assign n15772 = n15766 & ~n15771 ;
  assign n15773 = ~n3438 & n15772 ;
  assign n15774 = n10300 ^ n557 ^ 1'b0 ;
  assign n15775 = ~n3090 & n15774 ;
  assign n15776 = n4839 ^ n1141 ^ 1'b0 ;
  assign n15777 = ~n181 & n13334 ;
  assign n15778 = n8492 & n9617 ;
  assign n15779 = n8853 & ~n12453 ;
  assign n15780 = n15026 ^ n6796 ^ 1'b0 ;
  assign n15781 = n15780 ^ n10218 ^ 1'b0 ;
  assign n15782 = ( n7148 & n12403 ) | ( n7148 & n15781 ) | ( n12403 & n15781 ) ;
  assign n15789 = n12457 ^ n6857 ^ n6663 ;
  assign n15785 = n6282 ^ n3567 ^ 1'b0 ;
  assign n15786 = n9553 | n15785 ;
  assign n15787 = n3196 | n15786 ;
  assign n15788 = n15787 ^ n354 ^ 1'b0 ;
  assign n15783 = n7081 & n15469 ;
  assign n15784 = n15783 ^ n8897 ^ 1'b0 ;
  assign n15790 = n15789 ^ n15788 ^ n15784 ;
  assign n15791 = n4049 | n7447 ;
  assign n15792 = n11737 & ~n15791 ;
  assign n15793 = n5871 & n9598 ;
  assign n15794 = n229 & n15793 ;
  assign n15795 = ( n2377 & n5737 ) | ( n2377 & n15794 ) | ( n5737 & n15794 ) ;
  assign n15796 = n6110 & n6512 ;
  assign n15797 = ~n15795 & n15796 ;
  assign n15801 = n8290 ^ n3695 ^ n238 ;
  assign n15798 = ~n1853 & n11442 ;
  assign n15799 = n15798 ^ n14362 ^ 1'b0 ;
  assign n15800 = ~n6237 & n15799 ;
  assign n15802 = n15801 ^ n15800 ^ 1'b0 ;
  assign n15804 = n4240 ^ n3860 ^ 1'b0 ;
  assign n15803 = n1793 & n9930 ;
  assign n15805 = n15804 ^ n15803 ^ 1'b0 ;
  assign n15806 = n15549 & ~n15805 ;
  assign n15807 = n15806 ^ n1774 ^ 1'b0 ;
  assign n15808 = ( n582 & ~n8522 ) | ( n582 & n11936 ) | ( ~n8522 & n11936 ) ;
  assign n15809 = n2428 ^ n2049 ^ n730 ;
  assign n15810 = n1535 & ~n6940 ;
  assign n15811 = ~n11459 & n15810 ;
  assign n15812 = n15811 ^ n9562 ^ 1'b0 ;
  assign n15813 = n15809 & n15812 ;
  assign n15814 = n6647 | n10734 ;
  assign n15815 = n11643 & ~n15814 ;
  assign n15816 = n15813 | n15815 ;
  assign n15817 = n1499 & n3047 ;
  assign n15818 = n15817 ^ n4843 ^ 1'b0 ;
  assign n15819 = n12554 & n15818 ;
  assign n15820 = n14300 ^ n8847 ^ 1'b0 ;
  assign n15821 = n1823 & ~n15820 ;
  assign n15823 = n2172 & n12791 ;
  assign n15824 = ~n4722 & n15823 ;
  assign n15822 = n10847 | n15699 ;
  assign n15825 = n15824 ^ n15822 ^ 1'b0 ;
  assign n15826 = n4376 & ~n15825 ;
  assign n15828 = n4800 ^ n2107 ^ 1'b0 ;
  assign n15829 = ~n12367 & n15828 ;
  assign n15830 = n15829 ^ n10851 ^ n477 ;
  assign n15827 = n8369 ^ n1811 ^ 1'b0 ;
  assign n15831 = n15830 ^ n15827 ^ n5328 ;
  assign n15832 = ( n1722 & n10123 ) | ( n1722 & ~n11524 ) | ( n10123 & ~n11524 ) ;
  assign n15834 = n1699 & ~n5502 ;
  assign n15835 = n5412 & n15834 ;
  assign n15836 = n15835 ^ n14620 ^ n2445 ;
  assign n15833 = n4277 & n4625 ;
  assign n15837 = n15836 ^ n15833 ^ 1'b0 ;
  assign n15838 = ( n1586 & ~n9648 ) | ( n1586 & n15837 ) | ( ~n9648 & n15837 ) ;
  assign n15839 = n4011 & n10737 ;
  assign n15840 = ~n11278 & n15839 ;
  assign n15841 = n5116 ^ n2709 ^ n1485 ;
  assign n15842 = n13351 | n15841 ;
  assign n15843 = ~n15123 & n15842 ;
  assign n15844 = n5206 | n14908 ;
  assign n15845 = n8285 ^ n3375 ^ n270 ;
  assign n15846 = n9859 | n10189 ;
  assign n15847 = n15845 & ~n15846 ;
  assign n15848 = n11947 ^ n11014 ^ 1'b0 ;
  assign n15849 = n9089 & n15848 ;
  assign n15850 = n11900 ^ n8744 ^ 1'b0 ;
  assign n15851 = n8832 ^ n2723 ^ 1'b0 ;
  assign n15852 = n15851 ^ n4054 ^ 1'b0 ;
  assign n15853 = n2842 | n7160 ;
  assign n15854 = n15853 ^ n6227 ^ n1750 ;
  assign n15855 = n12707 | n15854 ;
  assign n15856 = n15855 ^ n4809 ^ 1'b0 ;
  assign n15857 = x35 & ~n15596 ;
  assign n15858 = ( n15852 & ~n15856 ) | ( n15852 & n15857 ) | ( ~n15856 & n15857 ) ;
  assign n15859 = n10680 ^ n1185 ^ 1'b0 ;
  assign n15866 = n2445 ^ n1642 ^ 1'b0 ;
  assign n15867 = ~n1928 & n15866 ;
  assign n15860 = n2635 & n4815 ;
  assign n15861 = n15860 ^ n6705 ^ 1'b0 ;
  assign n15862 = n11434 ^ n9553 ^ n3791 ;
  assign n15863 = ~n2590 & n15862 ;
  assign n15864 = ( ~n8953 & n14523 ) | ( ~n8953 & n15863 ) | ( n14523 & n15863 ) ;
  assign n15865 = ( n14289 & n15861 ) | ( n14289 & ~n15864 ) | ( n15861 & ~n15864 ) ;
  assign n15868 = n15867 ^ n15865 ^ x49 ;
  assign n15869 = n7410 ^ n5238 ^ n4394 ;
  assign n15870 = n2592 | n15869 ;
  assign n15871 = n15769 ^ n857 ^ 1'b0 ;
  assign n15872 = ( n4813 & n14506 ) | ( n4813 & ~n15871 ) | ( n14506 & ~n15871 ) ;
  assign n15873 = n6888 ^ n6126 ^ 1'b0 ;
  assign n15874 = n5855 | n15556 ;
  assign n15875 = n15874 ^ n6363 ^ 1'b0 ;
  assign n15876 = n7246 | n8156 ;
  assign n15877 = ~n11797 & n13457 ;
  assign n15878 = ( n6081 & ~n15876 ) | ( n6081 & n15877 ) | ( ~n15876 & n15877 ) ;
  assign n15879 = n2809 & ~n4781 ;
  assign n15880 = ( n3847 & ~n10280 ) | ( n3847 & n11368 ) | ( ~n10280 & n11368 ) ;
  assign n15881 = n15880 ^ n2869 ^ 1'b0 ;
  assign n15882 = n950 | n5264 ;
  assign n15883 = n15882 ^ n12693 ^ 1'b0 ;
  assign n15884 = ~n175 & n15883 ;
  assign n15885 = n1231 & n3614 ;
  assign n15886 = n15885 ^ n2494 ^ 1'b0 ;
  assign n15887 = n14305 ^ n10478 ^ 1'b0 ;
  assign n15888 = n15886 & n15887 ;
  assign n15889 = n360 | n15888 ;
  assign n15890 = n3704 ^ n2140 ^ 1'b0 ;
  assign n15891 = ~n3282 & n15890 ;
  assign n15892 = n8328 ^ n4052 ^ 1'b0 ;
  assign n15893 = ~n1729 & n15892 ;
  assign n15894 = n3286 ^ n1259 ^ 1'b0 ;
  assign n15895 = n3007 & n15894 ;
  assign n15896 = n15895 ^ n225 ^ 1'b0 ;
  assign n15897 = n4890 | n15896 ;
  assign n15898 = n15897 ^ x4 ^ 1'b0 ;
  assign n15899 = ( n13833 & ~n15893 ) | ( n13833 & n15898 ) | ( ~n15893 & n15898 ) ;
  assign n15900 = n10040 ^ n2687 ^ n2100 ;
  assign n15901 = n9432 ^ n8216 ^ x21 ;
  assign n15902 = ( n15899 & n15900 ) | ( n15899 & ~n15901 ) | ( n15900 & ~n15901 ) ;
  assign n15903 = ~n4239 & n10464 ;
  assign n15904 = n3358 ^ n2695 ^ 1'b0 ;
  assign n15905 = n6939 | n15904 ;
  assign n15906 = n2906 ^ n340 ^ 1'b0 ;
  assign n15907 = ~n15905 & n15906 ;
  assign n15908 = n15907 ^ n2202 ^ 1'b0 ;
  assign n15909 = n15903 & ~n15908 ;
  assign n15910 = n2434 & n15909 ;
  assign n15911 = n15910 ^ n14180 ^ 1'b0 ;
  assign n15912 = n8351 | n8785 ;
  assign n15913 = ~n8449 & n10433 ;
  assign n15914 = ~n11501 & n11834 ;
  assign n15915 = ~n12006 & n15914 ;
  assign n15916 = n5563 & n13497 ;
  assign n15917 = n15916 ^ n6832 ^ 1'b0 ;
  assign n15918 = ~n13707 & n15917 ;
  assign n15919 = n9639 ^ n2965 ^ 1'b0 ;
  assign n15920 = n8872 & ~n15919 ;
  assign n15921 = n5643 | n6763 ;
  assign n15922 = n1033 | n8019 ;
  assign n15923 = n7036 ^ n1173 ^ 1'b0 ;
  assign n15924 = n15923 ^ n14893 ^ 1'b0 ;
  assign n15925 = ~n8374 & n15924 ;
  assign n15926 = ~n11782 & n15925 ;
  assign n15927 = n15926 ^ n2748 ^ 1'b0 ;
  assign n15928 = n7873 ^ n6134 ^ 1'b0 ;
  assign n15929 = n15927 & ~n15928 ;
  assign n15930 = n13985 ^ n1793 ^ n404 ;
  assign n15931 = n15930 ^ n13112 ^ 1'b0 ;
  assign n15932 = ( ~n2695 & n5338 ) | ( ~n2695 & n9400 ) | ( n5338 & n9400 ) ;
  assign n15933 = ~n5117 & n5671 ;
  assign n15934 = n15933 ^ n5849 ^ 1'b0 ;
  assign n15935 = n5003 & ~n15934 ;
  assign n15936 = n15935 ^ n2260 ^ 1'b0 ;
  assign n15937 = ( n2299 & n6679 ) | ( n2299 & ~n15936 ) | ( n6679 & ~n15936 ) ;
  assign n15938 = n5037 & ~n12744 ;
  assign n15939 = ~n673 & n15938 ;
  assign n15940 = ~n11291 & n15939 ;
  assign n15941 = n9715 ^ n3006 ^ 1'b0 ;
  assign n15942 = n11916 & ~n15941 ;
  assign n15944 = ~n4824 & n8139 ;
  assign n15943 = n1246 & n2511 ;
  assign n15945 = n15944 ^ n15943 ^ 1'b0 ;
  assign n15946 = n15585 ^ n13302 ^ 1'b0 ;
  assign n15947 = n7607 | n15946 ;
  assign n15948 = ( n2638 & n6100 ) | ( n2638 & n13466 ) | ( n6100 & n13466 ) ;
  assign n15949 = n1351 & ~n11790 ;
  assign n15951 = n5223 ^ n3850 ^ n1959 ;
  assign n15950 = n913 & ~n10199 ;
  assign n15952 = n15951 ^ n15950 ^ 1'b0 ;
  assign n15954 = n1485 | n11079 ;
  assign n15955 = n746 & ~n15954 ;
  assign n15953 = n3659 & ~n11038 ;
  assign n15956 = n15955 ^ n15953 ^ 1'b0 ;
  assign n15957 = n15287 ^ n9809 ^ n1491 ;
  assign n15958 = ~n10009 & n15957 ;
  assign n15963 = ~n5561 & n14466 ;
  assign n15959 = n1184 ^ n1065 ^ n841 ;
  assign n15960 = n15959 ^ n3504 ^ 1'b0 ;
  assign n15961 = ~n6798 & n15960 ;
  assign n15962 = ~n14366 & n15961 ;
  assign n15964 = n15963 ^ n15962 ^ 1'b0 ;
  assign n15965 = n15189 ^ n4345 ^ 1'b0 ;
  assign n15966 = n15965 ^ n1502 ^ 1'b0 ;
  assign n15967 = ( ~n3349 & n6180 ) | ( ~n3349 & n15966 ) | ( n6180 & n15966 ) ;
  assign n15968 = n1751 & n1874 ;
  assign n15969 = n15968 ^ n322 ^ 1'b0 ;
  assign n15970 = n15969 ^ n13564 ^ n10333 ;
  assign n15971 = n14029 ^ n12467 ^ n4110 ;
  assign n15972 = n307 & ~n10234 ;
  assign n15973 = n1199 & ~n14838 ;
  assign n15974 = ~n14316 & n15973 ;
  assign n15975 = n3583 | n6256 ;
  assign n15976 = n15975 ^ n9766 ^ n4570 ;
  assign n15977 = n6778 & ~n15340 ;
  assign n15978 = n15977 ^ n4714 ^ 1'b0 ;
  assign n15979 = ~n5301 & n15978 ;
  assign n15980 = ~n2991 & n10146 ;
  assign n15981 = ( ~n9881 & n13567 ) | ( ~n9881 & n15980 ) | ( n13567 & n15980 ) ;
  assign n15982 = ~n4884 & n6057 ;
  assign n15983 = n15982 ^ n9593 ^ n8139 ;
  assign n15984 = n15983 ^ n9443 ^ 1'b0 ;
  assign n15985 = ~n15981 & n15984 ;
  assign n15986 = n11278 ^ n1832 ^ 1'b0 ;
  assign n15987 = n9348 & n15986 ;
  assign n15988 = n7514 & n8129 ;
  assign n15989 = n6652 & n15988 ;
  assign n15990 = ( n187 & n10958 ) | ( n187 & ~n15989 ) | ( n10958 & ~n15989 ) ;
  assign n15991 = n15990 ^ n6623 ^ 1'b0 ;
  assign n15992 = n8496 & ~n15991 ;
  assign n15993 = n15992 ^ n10024 ^ n4578 ;
  assign n15994 = n12609 ^ n7023 ^ 1'b0 ;
  assign n15995 = ( ~n3824 & n4654 ) | ( ~n3824 & n9925 ) | ( n4654 & n9925 ) ;
  assign n15996 = ( n10839 & ~n10985 ) | ( n10839 & n15995 ) | ( ~n10985 & n15995 ) ;
  assign n15997 = n15996 ^ n11797 ^ n1674 ;
  assign n15998 = n7795 ^ n1473 ^ 1'b0 ;
  assign n15999 = n1098 & ~n15998 ;
  assign n16000 = n10148 ^ n8786 ^ 1'b0 ;
  assign n16001 = ~n259 & n16000 ;
  assign n16002 = x103 & n16001 ;
  assign n16003 = n1739 & ~n12542 ;
  assign n16004 = n360 & n16003 ;
  assign n16005 = n9488 | n16004 ;
  assign n16006 = n16005 ^ n1200 ^ 1'b0 ;
  assign n16007 = n10234 ^ n3765 ^ 1'b0 ;
  assign n16008 = n4104 & n6854 ;
  assign n16009 = ( n7321 & n14151 ) | ( n7321 & ~n16008 ) | ( n14151 & ~n16008 ) ;
  assign n16010 = ~n9747 & n12118 ;
  assign n16011 = n14570 & n16010 ;
  assign n16012 = ( n5561 & n14347 ) | ( n5561 & ~n16011 ) | ( n14347 & ~n16011 ) ;
  assign n16013 = n8767 ^ n4091 ^ n2604 ;
  assign n16014 = n11321 | n14722 ;
  assign n16015 = n16014 ^ n3798 ^ 1'b0 ;
  assign n16016 = n7408 | n8374 ;
  assign n16017 = n6200 | n16016 ;
  assign n16018 = ~n11038 & n16017 ;
  assign n16019 = ~n4909 & n16018 ;
  assign n16020 = ~n1529 & n1637 ;
  assign n16021 = n16020 ^ n15969 ^ 1'b0 ;
  assign n16022 = n9002 ^ n6368 ^ 1'b0 ;
  assign n16023 = n16021 | n16022 ;
  assign n16024 = n3271 | n11115 ;
  assign n16025 = n16024 ^ n5317 ^ 1'b0 ;
  assign n16026 = n9292 & n16025 ;
  assign n16027 = ~n6601 & n16026 ;
  assign n16028 = n9001 & ~n12757 ;
  assign n16029 = n5158 ^ n1259 ^ 1'b0 ;
  assign n16030 = n4501 & n16029 ;
  assign n16031 = n16030 ^ n15745 ^ n2873 ;
  assign n16032 = n11960 | n16031 ;
  assign n16033 = n16028 & ~n16032 ;
  assign n16034 = n16033 ^ n15174 ^ n5384 ;
  assign n16038 = n15641 ^ n4966 ^ 1'b0 ;
  assign n16035 = n2740 & ~n3048 ;
  assign n16036 = ~n14628 & n16035 ;
  assign n16037 = n1848 & ~n16036 ;
  assign n16039 = n16038 ^ n16037 ^ 1'b0 ;
  assign n16040 = n15217 ^ n2082 ^ n1612 ;
  assign n16041 = ( ~n1587 & n2095 ) | ( ~n1587 & n4115 ) | ( n2095 & n4115 ) ;
  assign n16042 = ~n8952 & n16041 ;
  assign n16043 = ~n16040 & n16042 ;
  assign n16044 = ~n11564 & n16043 ;
  assign n16045 = n13755 ^ n12968 ^ n9675 ;
  assign n16046 = n8757 ^ n1674 ^ 1'b0 ;
  assign n16047 = n12617 & ~n16046 ;
  assign n16048 = n16047 ^ n16041 ^ 1'b0 ;
  assign n16049 = n16048 ^ n10834 ^ n6668 ;
  assign n16050 = ( ~n2445 & n6340 ) | ( ~n2445 & n7339 ) | ( n6340 & n7339 ) ;
  assign n16051 = ( n4939 & n5013 ) | ( n4939 & ~n11551 ) | ( n5013 & ~n11551 ) ;
  assign n16052 = n2377 & n12754 ;
  assign n16053 = n1519 & n16052 ;
  assign n16054 = n1600 | n16053 ;
  assign n16055 = n16051 & ~n16054 ;
  assign n16056 = n1049 | n7270 ;
  assign n16057 = n16056 ^ n2377 ^ 1'b0 ;
  assign n16058 = n14762 & ~n16057 ;
  assign n16060 = n816 | n1511 ;
  assign n16061 = n5224 & ~n16060 ;
  assign n16059 = n3317 & ~n9828 ;
  assign n16062 = n16061 ^ n16059 ^ 1'b0 ;
  assign n16063 = n12307 ^ n11562 ^ n6003 ;
  assign n16064 = n2645 & n8517 ;
  assign n16065 = ~n2383 & n14152 ;
  assign n16066 = n16065 ^ n1423 ^ 1'b0 ;
  assign n16067 = n3140 & ~n14560 ;
  assign n16068 = n16067 ^ n7986 ^ 1'b0 ;
  assign n16069 = n1107 ^ n802 ^ x98 ;
  assign n16070 = n16069 ^ n9073 ^ 1'b0 ;
  assign n16071 = n1732 & ~n15887 ;
  assign n16072 = ~n16070 & n16071 ;
  assign n16077 = ~n2624 & n4304 ;
  assign n16078 = n16077 ^ n1994 ^ 1'b0 ;
  assign n16074 = n6045 | n9393 ;
  assign n16073 = ( n2200 & n10304 ) | ( n2200 & n15016 ) | ( n10304 & n15016 ) ;
  assign n16075 = n16074 ^ n16073 ^ 1'b0 ;
  assign n16076 = n1260 | n16075 ;
  assign n16079 = n16078 ^ n16076 ^ n6536 ;
  assign n16080 = n16079 ^ n3837 ^ 1'b0 ;
  assign n16084 = n2161 | n2960 ;
  assign n16085 = n950 & ~n16084 ;
  assign n16081 = n1035 & n9710 ;
  assign n16082 = ~n6003 & n16081 ;
  assign n16083 = n16082 ^ n12628 ^ n2458 ;
  assign n16086 = n16085 ^ n16083 ^ n3051 ;
  assign n16087 = n10605 & n16086 ;
  assign n16088 = n16087 ^ n12419 ^ 1'b0 ;
  assign n16089 = n650 & n4722 ;
  assign n16090 = n16089 ^ n1304 ^ 1'b0 ;
  assign n16091 = n16090 ^ n10268 ^ 1'b0 ;
  assign n16093 = ( n652 & ~n7291 ) | ( n652 & n8253 ) | ( ~n7291 & n8253 ) ;
  assign n16094 = n16093 ^ n9094 ^ 1'b0 ;
  assign n16092 = ( ~n763 & n1876 ) | ( ~n763 & n5389 ) | ( n1876 & n5389 ) ;
  assign n16095 = n16094 ^ n16092 ^ n2195 ;
  assign n16096 = n13339 ^ n7877 ^ 1'b0 ;
  assign n16097 = ( n1794 & n11750 ) | ( n1794 & ~n16096 ) | ( n11750 & ~n16096 ) ;
  assign n16098 = n16097 ^ n7871 ^ n4571 ;
  assign n16099 = ~n331 & n8732 ;
  assign n16100 = n4468 & n16099 ;
  assign n16101 = n16100 ^ n934 ^ 1'b0 ;
  assign n16102 = n13332 & ~n16101 ;
  assign n16103 = ( n654 & n3695 ) | ( n654 & ~n11323 ) | ( n3695 & ~n11323 ) ;
  assign n16104 = n2731 & n6946 ;
  assign n16105 = n16104 ^ n7632 ^ n4206 ;
  assign n16106 = n1467 & n16105 ;
  assign n16107 = ~n16103 & n16106 ;
  assign n16108 = n8984 ^ n3880 ^ 1'b0 ;
  assign n16109 = n7375 & n16108 ;
  assign n16110 = n11201 | n15243 ;
  assign n16111 = n16109 | n16110 ;
  assign n16112 = ~n4882 & n7376 ;
  assign n16113 = n9435 & n16112 ;
  assign n16114 = n11038 ^ n11001 ^ n1295 ;
  assign n16115 = n3530 | n6053 ;
  assign n16116 = n16114 | n16115 ;
  assign n16117 = n15734 ^ n4188 ^ n1091 ;
  assign n16118 = n16117 ^ n12497 ^ 1'b0 ;
  assign n16119 = n16116 & n16118 ;
  assign n16120 = n4117 & n8923 ;
  assign n16121 = n16120 ^ n1756 ^ 1'b0 ;
  assign n16122 = n9536 & ~n16121 ;
  assign n16123 = n16122 ^ n6271 ^ 1'b0 ;
  assign n16125 = n10464 ^ n7573 ^ n1983 ;
  assign n16124 = n3447 | n4636 ;
  assign n16126 = n16125 ^ n16124 ^ 1'b0 ;
  assign n16127 = n16126 ^ n10688 ^ n2692 ;
  assign n16128 = n1406 ^ n740 ^ 1'b0 ;
  assign n16129 = n16127 & ~n16128 ;
  assign n16130 = n4978 ^ n2909 ^ 1'b0 ;
  assign n16131 = n16130 ^ n815 ^ n515 ;
  assign n16132 = n16131 ^ n3450 ^ 1'b0 ;
  assign n16133 = n3933 & ~n16132 ;
  assign n16134 = ~n7417 & n12255 ;
  assign n16135 = ~n8367 & n16134 ;
  assign n16136 = n469 & n16135 ;
  assign n16137 = n6679 & n16136 ;
  assign n16138 = ( ~n3756 & n5379 ) | ( ~n3756 & n7674 ) | ( n5379 & n7674 ) ;
  assign n16139 = n10110 ^ n4068 ^ n433 ;
  assign n16140 = n2570 & n16139 ;
  assign n16141 = ~n393 & n10647 ;
  assign n16142 = n9714 ^ n8147 ^ 1'b0 ;
  assign n16143 = ~n1281 & n5800 ;
  assign n16144 = ( ~n5318 & n6687 ) | ( ~n5318 & n12614 ) | ( n6687 & n12614 ) ;
  assign n16145 = n13786 ^ n6298 ^ 1'b0 ;
  assign n16146 = n16144 | n16145 ;
  assign n16147 = ( n3479 & n8319 ) | ( n3479 & n9945 ) | ( n8319 & n9945 ) ;
  assign n16148 = n9782 ^ n1430 ^ 1'b0 ;
  assign n16149 = n1862 & ~n12725 ;
  assign n16150 = n630 & ~n16149 ;
  assign n16151 = ( n10271 & n13334 ) | ( n10271 & n13553 ) | ( n13334 & n13553 ) ;
  assign n16152 = n16151 ^ n5107 ^ 1'b0 ;
  assign n16153 = ~n7324 & n16152 ;
  assign n16154 = n14215 ^ n13111 ^ n1914 ;
  assign n16155 = n16153 & ~n16154 ;
  assign n16156 = n607 | n10396 ;
  assign n16157 = n9788 | n16156 ;
  assign n16158 = n9441 ^ n7756 ^ 1'b0 ;
  assign n16159 = n16158 ^ n6182 ^ n3410 ;
  assign n16160 = ( n5348 & n6751 ) | ( n5348 & ~n16159 ) | ( n6751 & ~n16159 ) ;
  assign n16161 = ~n5780 & n15390 ;
  assign n16162 = ~n5230 & n16161 ;
  assign n16163 = n8363 & ~n14440 ;
  assign n16164 = n15869 ^ n3378 ^ 1'b0 ;
  assign n16165 = ~n14233 & n16164 ;
  assign n16166 = ~n8479 & n13883 ;
  assign n16167 = n8153 ^ n7289 ^ n3474 ;
  assign n16168 = n2156 & n16167 ;
  assign n16169 = n15149 ^ n10134 ^ 1'b0 ;
  assign n16170 = n7641 | n8901 ;
  assign n16174 = n4045 | n10752 ;
  assign n16175 = n16174 ^ n3859 ^ 1'b0 ;
  assign n16171 = n10315 ^ n1929 ^ 1'b0 ;
  assign n16172 = n7372 & ~n16171 ;
  assign n16173 = ~n644 & n16172 ;
  assign n16176 = n16175 ^ n16173 ^ n4148 ;
  assign n16177 = n1959 | n16176 ;
  assign n16181 = n3139 | n5356 ;
  assign n16178 = n6206 & ~n10757 ;
  assign n16179 = n9595 & n16178 ;
  assign n16180 = n16179 ^ n5460 ^ n4800 ;
  assign n16182 = n16181 ^ n16180 ^ x38 ;
  assign n16183 = n661 & n2527 ;
  assign n16188 = n4206 ^ n2105 ^ 1'b0 ;
  assign n16189 = n16188 ^ n3824 ^ 1'b0 ;
  assign n16184 = x22 & n9073 ;
  assign n16185 = ~n2577 & n16184 ;
  assign n16186 = n9283 | n16185 ;
  assign n16187 = n16186 ^ n5235 ^ 1'b0 ;
  assign n16190 = n16189 ^ n16187 ^ n6894 ;
  assign n16191 = n16183 | n16190 ;
  assign n16192 = ~n982 & n3777 ;
  assign n16196 = n9173 ^ n3392 ^ 1'b0 ;
  assign n16197 = x68 & ~n16196 ;
  assign n16193 = n6281 ^ n1276 ^ 1'b0 ;
  assign n16194 = n2456 & n16193 ;
  assign n16195 = n16194 ^ n9222 ^ 1'b0 ;
  assign n16198 = n16197 ^ n16195 ^ n12366 ;
  assign n16199 = n3777 ^ n370 ^ 1'b0 ;
  assign n16200 = n15520 ^ n10762 ^ 1'b0 ;
  assign n16201 = n6881 | n16200 ;
  assign n16202 = ~n1672 & n3785 ;
  assign n16203 = n16202 ^ n4870 ^ 1'b0 ;
  assign n16207 = ( n1150 & ~n3250 ) | ( n1150 & n5990 ) | ( ~n3250 & n5990 ) ;
  assign n16208 = n16207 ^ n11153 ^ n1895 ;
  assign n16204 = ~n4566 & n5026 ;
  assign n16205 = ~n10687 & n16204 ;
  assign n16206 = ~n1498 & n16205 ;
  assign n16209 = n16208 ^ n16206 ^ n378 ;
  assign n16210 = ~n5087 & n16209 ;
  assign n16211 = ( n1198 & n12403 ) | ( n1198 & ~n16210 ) | ( n12403 & ~n16210 ) ;
  assign n16212 = n1940 | n3463 ;
  assign n16213 = n16211 | n16212 ;
  assign n16214 = n4149 & n13418 ;
  assign n16215 = n9424 ^ n3832 ^ n2976 ;
  assign n16216 = n2233 | n6983 ;
  assign n16217 = n16216 ^ n7762 ^ 1'b0 ;
  assign n16222 = ( n3722 & n4052 ) | ( n3722 & n11187 ) | ( n4052 & n11187 ) ;
  assign n16221 = ( ~n140 & n2481 ) | ( ~n140 & n3923 ) | ( n2481 & n3923 ) ;
  assign n16218 = n14778 ^ n6216 ^ 1'b0 ;
  assign n16219 = n6121 | n16218 ;
  assign n16220 = ~n1228 & n16219 ;
  assign n16223 = n16222 ^ n16221 ^ n16220 ;
  assign n16224 = n5217 ^ n1358 ^ n1112 ;
  assign n16225 = n16224 ^ n5762 ^ 1'b0 ;
  assign n16226 = ( n9503 & n9598 ) | ( n9503 & ~n10982 ) | ( n9598 & ~n10982 ) ;
  assign n16227 = n5517 ^ n1777 ^ 1'b0 ;
  assign n16228 = ~n16226 & n16227 ;
  assign n16231 = n1335 | n3949 ;
  assign n16232 = n2888 | n16231 ;
  assign n16233 = n803 & ~n16232 ;
  assign n16229 = n7839 ^ n2256 ^ 1'b0 ;
  assign n16230 = ~n1552 & n16229 ;
  assign n16234 = n16233 ^ n16230 ^ 1'b0 ;
  assign n16235 = n4867 & ~n8900 ;
  assign n16236 = n10618 | n12451 ;
  assign n16237 = n16235 & ~n16236 ;
  assign n16238 = ~n4840 & n8441 ;
  assign n16239 = ~n4484 & n16238 ;
  assign n16240 = n3776 & n16239 ;
  assign n16241 = n146 | n2031 ;
  assign n16242 = ( n1915 & ~n9421 ) | ( n1915 & n16241 ) | ( ~n9421 & n16241 ) ;
  assign n16243 = n4242 & n10629 ;
  assign n16244 = ( n7304 & ~n16242 ) | ( n7304 & n16243 ) | ( ~n16242 & n16243 ) ;
  assign n16245 = ( n13743 & n16157 ) | ( n13743 & n16244 ) | ( n16157 & n16244 ) ;
  assign n16246 = n9709 ^ n1490 ^ 1'b0 ;
  assign n16247 = n16246 ^ n4451 ^ n2183 ;
  assign n16248 = ( n7648 & ~n10584 ) | ( n7648 & n16247 ) | ( ~n10584 & n16247 ) ;
  assign n16249 = n878 & ~n1458 ;
  assign n16250 = n8709 | n16249 ;
  assign n16251 = n9904 ^ n7592 ^ 1'b0 ;
  assign n16252 = n16251 ^ n8686 ^ 1'b0 ;
  assign n16253 = n16252 ^ n11915 ^ n10663 ;
  assign n16254 = n8489 & n11658 ;
  assign n16255 = n6776 ^ n1094 ^ 1'b0 ;
  assign n16256 = ( n2051 & n6104 ) | ( n2051 & n9920 ) | ( n6104 & n9920 ) ;
  assign n16257 = ( ~n219 & n8125 ) | ( ~n219 & n16256 ) | ( n8125 & n16256 ) ;
  assign n16259 = ~n2390 & n5147 ;
  assign n16260 = n16259 ^ n2016 ^ 1'b0 ;
  assign n16258 = ~n1502 & n2534 ;
  assign n16261 = n16260 ^ n16258 ^ 1'b0 ;
  assign n16262 = n6629 ^ n2897 ^ 1'b0 ;
  assign n16263 = n11525 | n16262 ;
  assign n16264 = n16263 ^ n11292 ^ n8969 ;
  assign n16265 = ( n3381 & n16261 ) | ( n3381 & ~n16264 ) | ( n16261 & ~n16264 ) ;
  assign n16266 = n6083 & ~n9611 ;
  assign n16267 = n2049 & ~n9683 ;
  assign n16268 = n16266 | n16267 ;
  assign n16269 = n7153 | n16268 ;
  assign n16270 = ~n15745 & n16217 ;
  assign n16271 = ~n1184 & n16270 ;
  assign n16272 = n2702 ^ n2186 ^ n1317 ;
  assign n16273 = n16272 ^ n10678 ^ 1'b0 ;
  assign n16274 = n16273 ^ x116 ^ 1'b0 ;
  assign n16275 = n7621 & ~n16274 ;
  assign n16276 = n13763 ^ n11128 ^ n10062 ;
  assign n16279 = ~n3613 & n5443 ;
  assign n16280 = n16279 ^ n13422 ^ 1'b0 ;
  assign n16277 = n15934 ^ n14427 ^ n2055 ;
  assign n16278 = n16277 ^ n16185 ^ n6544 ;
  assign n16281 = n16280 ^ n16278 ^ n14322 ;
  assign n16282 = n599 & ~n10276 ;
  assign n16283 = n6293 & n16282 ;
  assign n16284 = n10731 ^ n9579 ^ 1'b0 ;
  assign n16285 = n16284 ^ n6050 ^ 1'b0 ;
  assign n16287 = n258 & ~n1942 ;
  assign n16288 = n16287 ^ n5570 ^ 1'b0 ;
  assign n16286 = ( ~n11549 & n12137 ) | ( ~n11549 & n12357 ) | ( n12137 & n12357 ) ;
  assign n16289 = n16288 ^ n16286 ^ 1'b0 ;
  assign n16290 = n15003 ^ n8985 ^ 1'b0 ;
  assign n16291 = n6858 | n15522 ;
  assign n16292 = n3056 & ~n8056 ;
  assign n16293 = ~n4302 & n10681 ;
  assign n16294 = n6953 ^ n5493 ^ x61 ;
  assign n16295 = n16294 ^ n6411 ^ n1822 ;
  assign n16296 = n11764 ^ n3907 ^ 1'b0 ;
  assign n16297 = ( n576 & n4462 ) | ( n576 & n16296 ) | ( n4462 & n16296 ) ;
  assign n16298 = n2703 & ~n3682 ;
  assign n16299 = n708 & n16298 ;
  assign n16300 = ( ~n2552 & n15261 ) | ( ~n2552 & n16299 ) | ( n15261 & n16299 ) ;
  assign n16301 = ~n1840 & n2109 ;
  assign n16302 = ~n5461 & n16301 ;
  assign n16303 = n16302 ^ n13265 ^ n3284 ;
  assign n16304 = ( ~n2923 & n3961 ) | ( ~n2923 & n14517 ) | ( n3961 & n14517 ) ;
  assign n16305 = n15841 ^ n4378 ^ n2930 ;
  assign n16306 = n4473 & ~n16305 ;
  assign n16307 = n16306 ^ n15217 ^ 1'b0 ;
  assign n16308 = n16304 & n16307 ;
  assign n16309 = n357 & n16308 ;
  assign n16310 = n848 & ~n8867 ;
  assign n16311 = n16310 ^ n7295 ^ 1'b0 ;
  assign n16312 = ~n6978 & n13308 ;
  assign n16313 = n2867 & n8482 ;
  assign n16314 = ( n14293 & ~n16312 ) | ( n14293 & n16313 ) | ( ~n16312 & n16313 ) ;
  assign n16315 = n15328 ^ n12985 ^ 1'b0 ;
  assign n16316 = n16314 & n16315 ;
  assign n16317 = n11560 ^ n2584 ^ 1'b0 ;
  assign n16318 = n16317 ^ n9606 ^ 1'b0 ;
  assign n16319 = n14136 | n16318 ;
  assign n16320 = n6630 & ~n16319 ;
  assign n16321 = n10913 ^ n9871 ^ 1'b0 ;
  assign n16322 = n14654 & ~n16321 ;
  assign n16323 = n9959 & n16322 ;
  assign n16324 = n5111 & n16323 ;
  assign n16325 = n9955 | n14517 ;
  assign n16326 = n16325 ^ n10211 ^ 1'b0 ;
  assign n16327 = n6962 & n16326 ;
  assign n16328 = ~n5349 & n16327 ;
  assign n16329 = n16328 ^ n7723 ^ 1'b0 ;
  assign n16330 = ~n12343 & n16329 ;
  assign n16331 = n16330 ^ n1733 ^ n799 ;
  assign n16332 = ( ~n948 & n1691 ) | ( ~n948 & n2051 ) | ( n1691 & n2051 ) ;
  assign n16333 = n3583 ^ n950 ^ 1'b0 ;
  assign n16334 = n16333 ^ n9350 ^ 1'b0 ;
  assign n16335 = n9847 ^ n4566 ^ 1'b0 ;
  assign n16336 = n13771 & ~n16335 ;
  assign n16337 = n16336 ^ n12380 ^ n7131 ;
  assign n16338 = n10878 ^ n3554 ^ 1'b0 ;
  assign n16339 = ~n4065 & n6209 ;
  assign n16340 = n16339 ^ n5691 ^ 1'b0 ;
  assign n16341 = n8475 & n16340 ;
  assign n16342 = n16341 ^ n6475 ^ 1'b0 ;
  assign n16343 = n11562 | n16342 ;
  assign n16344 = n7237 ^ n2658 ^ n2273 ;
  assign n16345 = n16344 ^ n3749 ^ n260 ;
  assign n16346 = n16343 & ~n16345 ;
  assign n16347 = n8569 ^ n3716 ^ 1'b0 ;
  assign n16348 = n16286 & n16347 ;
  assign n16349 = ( ~n2318 & n6129 ) | ( ~n2318 & n16348 ) | ( n6129 & n16348 ) ;
  assign n16350 = n5771 ^ n3231 ^ n1521 ;
  assign n16351 = n16350 ^ n6999 ^ 1'b0 ;
  assign n16352 = ~n9587 & n16351 ;
  assign n16355 = n8708 & n9336 ;
  assign n16353 = n7293 & n9985 ;
  assign n16354 = ~n210 & n16353 ;
  assign n16356 = n16355 ^ n16354 ^ n5465 ;
  assign n16357 = n314 & ~n2391 ;
  assign n16358 = n2565 & n16357 ;
  assign n16359 = n2969 ^ n138 ^ 1'b0 ;
  assign n16360 = x97 & n16359 ;
  assign n16361 = ~n12383 & n16360 ;
  assign n16362 = n16358 & n16361 ;
  assign n16363 = n4717 ^ n307 ^ 1'b0 ;
  assign n16364 = n16362 | n16363 ;
  assign n16370 = ( n3721 & n10010 ) | ( n3721 & ~n12867 ) | ( n10010 & ~n12867 ) ;
  assign n16365 = n11950 ^ n10920 ^ 1'b0 ;
  assign n16366 = n13244 | n16365 ;
  assign n16367 = n9903 ^ n8395 ^ 1'b0 ;
  assign n16368 = n16366 | n16367 ;
  assign n16369 = n4088 | n16368 ;
  assign n16371 = n16370 ^ n16369 ^ 1'b0 ;
  assign n16384 = n7008 ^ n6281 ^ n2264 ;
  assign n16383 = ( n143 & n2296 ) | ( n143 & ~n7586 ) | ( n2296 & ~n7586 ) ;
  assign n16385 = n16384 ^ n16383 ^ n14205 ;
  assign n16378 = ( n3809 & ~n4401 ) | ( n3809 & n6575 ) | ( ~n4401 & n6575 ) ;
  assign n16379 = n4119 | n16378 ;
  assign n16377 = n15650 ^ n10295 ^ 1'b0 ;
  assign n16380 = n16379 ^ n16377 ^ n13110 ;
  assign n16373 = n2706 ^ n2489 ^ 1'b0 ;
  assign n16374 = n512 & ~n16373 ;
  assign n16372 = ~n5057 & n10986 ;
  assign n16375 = n16374 ^ n16372 ^ n10576 ;
  assign n16376 = n7268 | n16375 ;
  assign n16381 = n16380 ^ n16376 ^ 1'b0 ;
  assign n16382 = n325 | n16381 ;
  assign n16386 = n16385 ^ n16382 ^ 1'b0 ;
  assign n16387 = n14921 ^ n7737 ^ n7458 ;
  assign n16388 = n16387 ^ n1855 ^ 1'b0 ;
  assign n16389 = n5980 & ~n16388 ;
  assign n16390 = ~n160 & n6675 ;
  assign n16391 = n1669 & n16069 ;
  assign n16394 = n12302 ^ n1836 ^ 1'b0 ;
  assign n16395 = n4107 & n16394 ;
  assign n16392 = n1076 & ~n3357 ;
  assign n16393 = n16392 ^ n1358 ^ 1'b0 ;
  assign n16396 = n16395 ^ n16393 ^ n13291 ;
  assign n16397 = n16396 ^ n14494 ^ 1'b0 ;
  assign n16398 = n6794 ^ n281 ^ 1'b0 ;
  assign n16399 = ~n1502 & n4434 ;
  assign n16400 = n16399 ^ n9889 ^ 1'b0 ;
  assign n16401 = ( ~n8214 & n16398 ) | ( ~n8214 & n16400 ) | ( n16398 & n16400 ) ;
  assign n16402 = n16401 ^ n11917 ^ 1'b0 ;
  assign n16403 = ( n13914 & n14089 ) | ( n13914 & n16402 ) | ( n14089 & n16402 ) ;
  assign n16404 = n14930 ^ n3960 ^ 1'b0 ;
  assign n16405 = n6508 | n16404 ;
  assign n16406 = n7254 ^ n6306 ^ n5784 ;
  assign n16407 = n16405 | n16406 ;
  assign n16408 = ~n1440 & n13248 ;
  assign n16410 = n4413 & ~n5857 ;
  assign n16411 = n16410 ^ n5106 ^ 1'b0 ;
  assign n16409 = ~n440 & n9876 ;
  assign n16412 = n16411 ^ n16409 ^ 1'b0 ;
  assign n16413 = x78 & ~n16412 ;
  assign n16414 = n16408 & n16413 ;
  assign n16415 = n11140 ^ n8440 ^ 1'b0 ;
  assign n16416 = n5458 & ~n16415 ;
  assign n16417 = ( n2792 & n5461 ) | ( n2792 & ~n14678 ) | ( n5461 & ~n14678 ) ;
  assign n16418 = n8959 ^ n3289 ^ 1'b0 ;
  assign n16419 = n16418 ^ n8644 ^ n3316 ;
  assign n16420 = n16419 ^ n5635 ^ 1'b0 ;
  assign n16421 = n16417 & ~n16420 ;
  assign n16422 = n15896 ^ n10471 ^ n883 ;
  assign n16423 = n16422 ^ n13707 ^ 1'b0 ;
  assign n16424 = n7535 & n11315 ;
  assign n16425 = ( n5561 & ~n12900 ) | ( n5561 & n13034 ) | ( ~n12900 & n13034 ) ;
  assign n16426 = n13961 ^ n6381 ^ n5454 ;
  assign n16427 = n10323 ^ n8545 ^ 1'b0 ;
  assign n16428 = n10225 ^ n571 ^ 1'b0 ;
  assign n16429 = n7011 & ~n16428 ;
  assign n16430 = n1392 & n7130 ;
  assign n16431 = n6318 ^ n4242 ^ 1'b0 ;
  assign n16432 = n11070 & n16431 ;
  assign n16433 = ~n8036 & n14615 ;
  assign n16434 = n12410 ^ n493 ^ 1'b0 ;
  assign n16435 = ~n1123 & n16434 ;
  assign n16436 = n2957 | n16435 ;
  assign n16437 = n3136 ^ n2308 ^ 1'b0 ;
  assign n16438 = n9207 ^ n5613 ^ 1'b0 ;
  assign n16439 = n8139 & n16438 ;
  assign n16440 = n7196 & n13226 ;
  assign n16441 = ~n5290 & n10209 ;
  assign n16442 = n13991 ^ n6942 ^ 1'b0 ;
  assign n16445 = ~n1704 & n8044 ;
  assign n16443 = ( n1320 & ~n5759 ) | ( n1320 & n5792 ) | ( ~n5759 & n5792 ) ;
  assign n16444 = n3934 | n16443 ;
  assign n16446 = n16445 ^ n16444 ^ 1'b0 ;
  assign n16447 = n7023 | n16446 ;
  assign n16448 = n10537 | n16447 ;
  assign n16449 = ~n1324 & n1802 ;
  assign n16450 = ~x88 & n16449 ;
  assign n16451 = n16448 & ~n16450 ;
  assign n16452 = n6129 & n16451 ;
  assign n16456 = n6442 & n10699 ;
  assign n16457 = n16456 ^ n1068 ^ 1'b0 ;
  assign n16458 = ~n2499 & n16457 ;
  assign n16453 = n420 & n11581 ;
  assign n16454 = n16453 ^ n4301 ^ 1'b0 ;
  assign n16455 = n16454 ^ n3490 ^ 1'b0 ;
  assign n16459 = n16458 ^ n16455 ^ 1'b0 ;
  assign n16460 = n2380 | n16459 ;
  assign n16461 = n14471 ^ n2902 ^ 1'b0 ;
  assign n16462 = n9025 & ~n16461 ;
  assign n16463 = n16462 ^ n3772 ^ 1'b0 ;
  assign n16464 = n1865 | n4326 ;
  assign n16465 = ~n1086 & n16464 ;
  assign n16466 = ~x3 & n16465 ;
  assign n16467 = ( n1498 & ~n2961 ) | ( n1498 & n16466 ) | ( ~n2961 & n16466 ) ;
  assign n16468 = ~n510 & n736 ;
  assign n16469 = n16468 ^ n234 ^ 1'b0 ;
  assign n16478 = n1101 ^ n470 ^ 1'b0 ;
  assign n16479 = n4302 & n16478 ;
  assign n16480 = n7683 & n16479 ;
  assign n16470 = n12095 ^ n1949 ^ 1'b0 ;
  assign n16471 = n4699 ^ n2976 ^ 1'b0 ;
  assign n16472 = n16470 | n16471 ;
  assign n16473 = n2117 | n7064 ;
  assign n16474 = n807 & ~n16473 ;
  assign n16475 = n219 & ~n16474 ;
  assign n16476 = n16472 | n16475 ;
  assign n16477 = n10665 | n16476 ;
  assign n16481 = n16480 ^ n16477 ^ 1'b0 ;
  assign n16485 = n7768 ^ n447 ^ n264 ;
  assign n16482 = n9097 ^ n7373 ^ 1'b0 ;
  assign n16483 = n8550 & n15061 ;
  assign n16484 = n16482 & n16483 ;
  assign n16486 = n16485 ^ n16484 ^ 1'b0 ;
  assign n16487 = ~n6379 & n16486 ;
  assign n16490 = ( n1403 & n3068 ) | ( n1403 & n11116 ) | ( n3068 & n11116 ) ;
  assign n16491 = n853 | n16490 ;
  assign n16492 = n404 | n16491 ;
  assign n16488 = ( n3611 & ~n6533 ) | ( n3611 & n16374 ) | ( ~n6533 & n16374 ) ;
  assign n16489 = n16488 ^ n5154 ^ n1834 ;
  assign n16493 = n16492 ^ n16489 ^ n2606 ;
  assign n16494 = ~n1491 & n16493 ;
  assign n16495 = n804 & ~n7709 ;
  assign n16496 = ~n2272 & n4099 ;
  assign n16497 = n16496 ^ n4833 ^ 1'b0 ;
  assign n16498 = n1171 & ~n16497 ;
  assign n16499 = n3184 & ~n4596 ;
  assign n16500 = n16499 ^ n2801 ^ 1'b0 ;
  assign n16501 = ~n771 & n2527 ;
  assign n16502 = n11579 & n16501 ;
  assign n16503 = n7848 & n16502 ;
  assign n16504 = n16500 & n16503 ;
  assign n16505 = ( n2434 & n11612 ) | ( n2434 & ~n16504 ) | ( n11612 & ~n16504 ) ;
  assign n16506 = n11271 | n15959 ;
  assign n16507 = n9931 & ~n12185 ;
  assign n16508 = n16507 ^ n10998 ^ n9881 ;
  assign n16509 = n16508 ^ n802 ^ 1'b0 ;
  assign n16510 = n8688 & n16509 ;
  assign n16511 = ( n824 & ~n6193 ) | ( n824 & n13956 ) | ( ~n6193 & n13956 ) ;
  assign n16512 = n2588 & ~n12196 ;
  assign n16513 = n16512 ^ n15637 ^ 1'b0 ;
  assign n16514 = n2743 ^ n796 ^ 1'b0 ;
  assign n16515 = n1201 & n16514 ;
  assign n16516 = n2730 & ~n3864 ;
  assign n16517 = n16515 & n16516 ;
  assign n16518 = n4137 ^ n3620 ^ 1'b0 ;
  assign n16519 = n169 & n3688 ;
  assign n16520 = n16518 & n16519 ;
  assign n16521 = n2702 & n7180 ;
  assign n16522 = n16520 & n16521 ;
  assign n16523 = ~n5965 & n10549 ;
  assign n16524 = n16523 ^ n260 ^ 1'b0 ;
  assign n16525 = n2552 & n16524 ;
  assign n16526 = n16525 ^ n8903 ^ 1'b0 ;
  assign n16529 = n4343 ^ n1636 ^ 1'b0 ;
  assign n16530 = n16529 ^ n6137 ^ 1'b0 ;
  assign n16531 = n461 | n16530 ;
  assign n16528 = n3880 & n10566 ;
  assign n16532 = n16531 ^ n16528 ^ 1'b0 ;
  assign n16527 = ( n232 & ~n4511 ) | ( n232 & n5786 ) | ( ~n4511 & n5786 ) ;
  assign n16533 = n16532 ^ n16527 ^ n11923 ;
  assign n16534 = n11814 ^ n7750 ^ 1'b0 ;
  assign n16535 = n11946 ^ n5667 ^ n855 ;
  assign n16536 = n6356 & n16535 ;
  assign n16537 = n7059 & n16536 ;
  assign n16538 = ( n195 & n2061 ) | ( n195 & ~n9963 ) | ( n2061 & ~n9963 ) ;
  assign n16539 = n6605 ^ n2614 ^ 1'b0 ;
  assign n16540 = ( n8914 & ~n14587 ) | ( n8914 & n16539 ) | ( ~n14587 & n16539 ) ;
  assign n16541 = n4253 & n7107 ;
  assign n16542 = n9063 & ~n16541 ;
  assign n16543 = n16542 ^ n10030 ^ 1'b0 ;
  assign n16544 = n1709 | n16543 ;
  assign n16545 = ~n922 & n7908 ;
  assign n16546 = n16545 ^ n6432 ^ 1'b0 ;
  assign n16547 = n5304 & ~n13024 ;
  assign n16548 = n16547 ^ n138 ^ 1'b0 ;
  assign n16549 = ( n716 & ~n1186 ) | ( n716 & n16548 ) | ( ~n1186 & n16548 ) ;
  assign n16550 = ~n2040 & n3044 ;
  assign n16551 = n8438 ^ n1456 ^ 1'b0 ;
  assign n16552 = x40 & n13004 ;
  assign n16555 = n2931 & ~n6461 ;
  assign n16556 = n16555 ^ n2932 ^ 1'b0 ;
  assign n16553 = n11348 ^ n5293 ^ 1'b0 ;
  assign n16554 = n13867 | n16553 ;
  assign n16557 = n16556 ^ n16554 ^ 1'b0 ;
  assign n16558 = n4542 & n5842 ;
  assign n16559 = n7458 & n16558 ;
  assign n16560 = n1731 & n6148 ;
  assign n16561 = n16560 ^ n3431 ^ 1'b0 ;
  assign n16562 = n9903 ^ n7635 ^ n2401 ;
  assign n16563 = n4357 & ~n5138 ;
  assign n16564 = ~n6158 & n16563 ;
  assign n16565 = n16562 & n16564 ;
  assign n16566 = n1366 | n16565 ;
  assign n16567 = n7820 & ~n16566 ;
  assign n16568 = n11155 & n14100 ;
  assign n16569 = ~n10962 & n16568 ;
  assign n16570 = n11946 ^ n7618 ^ 1'b0 ;
  assign n16571 = n6834 & ~n8373 ;
  assign n16572 = ~n4190 & n9448 ;
  assign n16573 = n3413 & n16572 ;
  assign n16574 = n824 | n3340 ;
  assign n16575 = n7520 | n16574 ;
  assign n16576 = n15965 ^ n7200 ^ 1'b0 ;
  assign n16577 = n12768 | n16576 ;
  assign n16578 = n6752 & ~n16577 ;
  assign n16579 = n16578 ^ n6438 ^ 1'b0 ;
  assign n16580 = n8307 | n16579 ;
  assign n16581 = n16580 ^ n2193 ^ 1'b0 ;
  assign n16582 = n16581 ^ n12504 ^ 1'b0 ;
  assign n16583 = n5294 & ~n9781 ;
  assign n16584 = n16583 ^ n9744 ^ n2906 ;
  assign n16585 = n16584 ^ n4802 ^ 1'b0 ;
  assign n16586 = ( ~n5786 & n9850 ) | ( ~n5786 & n16175 ) | ( n9850 & n16175 ) ;
  assign n16587 = ~n2074 & n9831 ;
  assign n16588 = n16587 ^ n4591 ^ 1'b0 ;
  assign n16589 = n2599 & n4167 ;
  assign n16590 = n16589 ^ n7505 ^ 1'b0 ;
  assign n16591 = n6888 & ~n9603 ;
  assign n16592 = n16591 ^ n15626 ^ 1'b0 ;
  assign n16593 = ~n12882 & n16592 ;
  assign n16594 = n5164 & n16593 ;
  assign n16595 = n7130 | n8252 ;
  assign n16596 = n11100 & ~n16595 ;
  assign n16597 = n16594 & n16596 ;
  assign n16598 = n10807 ^ n10087 ^ 1'b0 ;
  assign n16599 = n2536 ^ n1200 ^ n389 ;
  assign n16600 = n2159 & n16599 ;
  assign n16601 = n4148 & n16600 ;
  assign n16602 = n11028 ^ n5784 ^ 1'b0 ;
  assign n16603 = ~n15410 & n16602 ;
  assign n16604 = n5689 ^ n2986 ^ 1'b0 ;
  assign n16605 = ~n16603 & n16604 ;
  assign n16606 = n3526 & ~n6349 ;
  assign n16607 = n12846 & n16606 ;
  assign n16609 = n3127 | n13505 ;
  assign n16610 = n16609 ^ n820 ^ 1'b0 ;
  assign n16608 = n3063 & ~n9177 ;
  assign n16611 = n16610 ^ n16608 ^ 1'b0 ;
  assign n16612 = ( n2285 & ~n5024 ) | ( n2285 & n16611 ) | ( ~n5024 & n16611 ) ;
  assign n16613 = n307 & n16612 ;
  assign n16614 = ~n13124 & n16613 ;
  assign n16615 = n3429 ^ n1450 ^ n380 ;
  assign n16616 = n3665 ^ n1340 ^ 1'b0 ;
  assign n16617 = ( n3787 & ~n10788 ) | ( n3787 & n16616 ) | ( ~n10788 & n16616 ) ;
  assign n16618 = ( n1770 & ~n6628 ) | ( n1770 & n16617 ) | ( ~n6628 & n16617 ) ;
  assign n16619 = ( n10751 & ~n13721 ) | ( n10751 & n16618 ) | ( ~n13721 & n16618 ) ;
  assign n16620 = n5274 & ~n13827 ;
  assign n16621 = n2138 & n9780 ;
  assign n16622 = n11089 ^ n10340 ^ 1'b0 ;
  assign n16623 = n16622 ^ n15168 ^ 1'b0 ;
  assign n16624 = x52 & ~n16623 ;
  assign n16625 = n8965 & n16624 ;
  assign n16626 = n16621 & n16625 ;
  assign n16627 = n1576 ^ n1078 ^ 1'b0 ;
  assign n16628 = n15061 & n16627 ;
  assign n16629 = n10189 ^ n9660 ^ n8955 ;
  assign n16630 = n586 & n1659 ;
  assign n16631 = ~n1612 & n6589 ;
  assign n16634 = n10609 ^ n4505 ^ n949 ;
  assign n16633 = n15762 & ~n16206 ;
  assign n16635 = n16634 ^ n16633 ^ 1'b0 ;
  assign n16632 = n1689 ^ n545 ^ 1'b0 ;
  assign n16636 = n16635 ^ n16632 ^ 1'b0 ;
  assign n16637 = n8033 ^ n4617 ^ 1'b0 ;
  assign n16638 = ~n4221 & n16637 ;
  assign n16639 = n16638 ^ n13505 ^ n11613 ;
  assign n16640 = ~n3803 & n3868 ;
  assign n16641 = n16640 ^ n1433 ^ 1'b0 ;
  assign n16642 = n16641 ^ n9869 ^ n6981 ;
  assign n16643 = n832 & n4343 ;
  assign n16644 = ( n4336 & n14605 ) | ( n4336 & n16643 ) | ( n14605 & n16643 ) ;
  assign n16645 = n16644 ^ n872 ^ 1'b0 ;
  assign n16646 = n5037 & ~n16645 ;
  assign n16647 = n2382 | n7058 ;
  assign n16648 = n10373 | n16647 ;
  assign n16649 = n2929 ^ n2648 ^ 1'b0 ;
  assign n16650 = n16649 ^ n10281 ^ n7023 ;
  assign n16651 = n16650 ^ n6191 ^ 1'b0 ;
  assign n16652 = n284 | n16651 ;
  assign n16653 = n6571 ^ n4797 ^ 1'b0 ;
  assign n16654 = n8032 ^ n2193 ^ 1'b0 ;
  assign n16655 = n16653 | n16654 ;
  assign n16656 = n16652 & n16655 ;
  assign n16657 = n16656 ^ n8196 ^ 1'b0 ;
  assign n16658 = n7769 ^ n3981 ^ 1'b0 ;
  assign n16659 = n1629 & ~n16658 ;
  assign n16660 = n4927 & n6476 ;
  assign n16661 = n16660 ^ n10489 ^ 1'b0 ;
  assign n16662 = ~n2869 & n14053 ;
  assign n16663 = n16662 ^ n10981 ^ 1'b0 ;
  assign n16664 = n13475 ^ n7987 ^ n2706 ;
  assign n16665 = n6986 ^ x20 ^ 1'b0 ;
  assign n16666 = n2171 & ~n16665 ;
  assign n16667 = n16666 ^ n10848 ^ 1'b0 ;
  assign n16668 = n16667 ^ n15520 ^ 1'b0 ;
  assign n16669 = n9625 ^ n8367 ^ 1'b0 ;
  assign n16670 = ( n3606 & ~n11617 ) | ( n3606 & n11633 ) | ( ~n11617 & n11633 ) ;
  assign n16671 = n14317 ^ n12336 ^ 1'b0 ;
  assign n16672 = n6127 | n16671 ;
  assign n16674 = n7568 & n13782 ;
  assign n16675 = n9153 ^ n5755 ^ 1'b0 ;
  assign n16676 = n16674 & ~n16675 ;
  assign n16673 = ( ~n3923 & n9439 ) | ( ~n3923 & n9872 ) | ( n9439 & n9872 ) ;
  assign n16677 = n16676 ^ n16673 ^ n10324 ;
  assign n16678 = n15028 ^ n12200 ^ 1'b0 ;
  assign n16679 = n16677 | n16678 ;
  assign n16680 = n5742 ^ n3114 ^ 1'b0 ;
  assign n16681 = ( n9868 & ~n12318 ) | ( n9868 & n16680 ) | ( ~n12318 & n16680 ) ;
  assign n16682 = n14183 ^ n1532 ^ 1'b0 ;
  assign n16683 = n3410 & n6005 ;
  assign n16684 = n11501 ^ n11368 ^ 1'b0 ;
  assign n16685 = ( n5284 & n16683 ) | ( n5284 & n16684 ) | ( n16683 & n16684 ) ;
  assign n16686 = n2874 ^ n849 ^ 1'b0 ;
  assign n16687 = n15992 & ~n16686 ;
  assign n16688 = ~n3553 & n11320 ;
  assign n16689 = n6713 | n9216 ;
  assign n16690 = n11128 ^ n4921 ^ 1'b0 ;
  assign n16691 = n16689 & n16690 ;
  assign n16692 = n11316 ^ n7981 ^ 1'b0 ;
  assign n16693 = n11327 & n16692 ;
  assign n16694 = n10429 & ~n16693 ;
  assign n16695 = n14957 ^ n6868 ^ 1'b0 ;
  assign n16696 = n7765 & n16695 ;
  assign n16697 = n11210 ^ n6453 ^ 1'b0 ;
  assign n16698 = ~n1354 & n16697 ;
  assign n16699 = ~n6636 & n9348 ;
  assign n16700 = n4149 & n16699 ;
  assign n16701 = n16700 ^ n9548 ^ n5351 ;
  assign n16702 = n824 & ~n3670 ;
  assign n16703 = n16702 ^ n12877 ^ n5127 ;
  assign n16704 = n16703 ^ n14452 ^ 1'b0 ;
  assign n16705 = ( x81 & n5049 ) | ( x81 & n6824 ) | ( n5049 & n6824 ) ;
  assign n16706 = n9556 ^ n9121 ^ 1'b0 ;
  assign n16707 = n1382 | n4645 ;
  assign n16708 = n16707 ^ n4274 ^ 1'b0 ;
  assign n16709 = ~n4981 & n11019 ;
  assign n16710 = n16708 & n16709 ;
  assign n16711 = n16710 ^ n755 ^ 1'b0 ;
  assign n16712 = ~n13268 & n16711 ;
  assign n16713 = n1867 & n16712 ;
  assign n16714 = n1808 & n16713 ;
  assign n16715 = n9197 & ~n14572 ;
  assign n16716 = n16715 ^ n10465 ^ 1'b0 ;
  assign n16717 = n4188 & n5461 ;
  assign n16718 = ( n8772 & n9145 ) | ( n8772 & n9182 ) | ( n9145 & n9182 ) ;
  assign n16720 = n318 & ~n4482 ;
  assign n16721 = n4621 & n16720 ;
  assign n16719 = n7221 | n11277 ;
  assign n16722 = n16721 ^ n16719 ^ 1'b0 ;
  assign n16723 = n16722 ^ n12353 ^ n802 ;
  assign n16728 = ~n8916 & n12573 ;
  assign n16726 = n13679 ^ n2912 ^ 1'b0 ;
  assign n16727 = n6200 & n16726 ;
  assign n16724 = n4519 & n7470 ;
  assign n16725 = n16724 ^ n14482 ^ 1'b0 ;
  assign n16729 = n16728 ^ n16727 ^ n16725 ;
  assign n16730 = n5821 & n14275 ;
  assign n16731 = n6926 & n16730 ;
  assign n16732 = n3318 ^ n3141 ^ 1'b0 ;
  assign n16733 = n13457 | n16732 ;
  assign n16734 = n5827 | n16733 ;
  assign n16735 = n16734 ^ n10988 ^ 1'b0 ;
  assign n16737 = ~n617 & n1856 ;
  assign n16738 = ~n5664 & n16737 ;
  assign n16736 = ~n2233 & n2586 ;
  assign n16739 = n16738 ^ n16736 ^ 1'b0 ;
  assign n16740 = n10564 ^ n7211 ^ n7066 ;
  assign n16741 = ( ~n11148 & n11457 ) | ( ~n11148 & n16740 ) | ( n11457 & n16740 ) ;
  assign n16742 = n9439 ^ n3123 ^ 1'b0 ;
  assign n16743 = n6874 & ~n16742 ;
  assign n16744 = n5999 & ~n16743 ;
  assign n16745 = n11647 ^ n2738 ^ 1'b0 ;
  assign n16746 = ~n6293 & n16745 ;
  assign n16747 = n16746 ^ n948 ^ 1'b0 ;
  assign n16748 = n12557 & ~n16747 ;
  assign n16749 = ~n3187 & n9897 ;
  assign n16750 = n16749 ^ n15851 ^ 1'b0 ;
  assign n16751 = n14401 ^ n10341 ^ 1'b0 ;
  assign n16752 = ~n7310 & n7566 ;
  assign n16753 = n16752 ^ n565 ^ 1'b0 ;
  assign n16754 = n16753 ^ n3453 ^ 1'b0 ;
  assign n16755 = ~n6232 & n16754 ;
  assign n16756 = n12827 & n16755 ;
  assign n16757 = n1856 ^ n251 ^ 1'b0 ;
  assign n16758 = n16757 ^ n15878 ^ n15745 ;
  assign n16759 = ~n7888 & n7918 ;
  assign n16760 = n5103 ^ n741 ^ 1'b0 ;
  assign n16761 = n1487 | n16760 ;
  assign n16762 = n15804 ^ n635 ^ 1'b0 ;
  assign n16763 = ~n3720 & n16762 ;
  assign n16764 = n7227 ^ n220 ^ 1'b0 ;
  assign n16765 = ( n16215 & n16763 ) | ( n16215 & n16764 ) | ( n16763 & n16764 ) ;
  assign n16766 = ~n3572 & n11155 ;
  assign n16767 = ~n9782 & n16766 ;
  assign n16768 = n2778 & n8974 ;
  assign n16769 = n4367 ^ n2076 ^ 1'b0 ;
  assign n16770 = n7692 ^ n1518 ^ 1'b0 ;
  assign n16771 = n6410 & n8033 ;
  assign n16772 = n2076 & n15944 ;
  assign n16773 = n13965 ^ n12786 ^ n12508 ;
  assign n16774 = n7103 ^ n1773 ^ 1'b0 ;
  assign n16775 = n7406 & n16774 ;
  assign n16776 = n14052 & ~n16490 ;
  assign n16777 = ~n16775 & n16776 ;
  assign n16778 = n867 & n16310 ;
  assign n16779 = n384 | n5238 ;
  assign n16780 = n2738 | n16779 ;
  assign n16781 = n9763 & n16780 ;
  assign n16782 = n1212 & n16781 ;
  assign n16783 = n6631 | n8445 ;
  assign n16784 = n16782 | n16783 ;
  assign n16785 = n16784 ^ n13536 ^ 1'b0 ;
  assign n16786 = n8891 ^ n2422 ^ 1'b0 ;
  assign n16787 = n6525 | n16786 ;
  assign n16788 = ( n1281 & n5587 ) | ( n1281 & ~n8271 ) | ( n5587 & ~n8271 ) ;
  assign n16789 = n207 & ~n3390 ;
  assign n16790 = n16789 ^ n497 ^ 1'b0 ;
  assign n16791 = n16740 ^ n7257 ^ 1'b0 ;
  assign n16792 = n16790 & ~n16791 ;
  assign n16793 = n16792 ^ n13332 ^ 1'b0 ;
  assign n16794 = n14661 ^ n6700 ^ n3728 ;
  assign n16795 = n7829 ^ n5715 ^ 1'b0 ;
  assign n16796 = n349 & n16795 ;
  assign n16797 = n12101 | n16796 ;
  assign n16798 = n138 & n14410 ;
  assign n16799 = n6838 & ~n13475 ;
  assign n16800 = n11666 & ~n12609 ;
  assign n16801 = n11685 & n16800 ;
  assign n16802 = n11738 ^ n7730 ^ 1'b0 ;
  assign n16803 = ~n16801 & n16802 ;
  assign n16804 = n16803 ^ n9778 ^ n2251 ;
  assign n16806 = n1689 & n6959 ;
  assign n16805 = n2487 & ~n10610 ;
  assign n16807 = n16806 ^ n16805 ^ 1'b0 ;
  assign n16808 = ~n1428 & n9538 ;
  assign n16809 = ~n3445 & n16808 ;
  assign n16810 = n16809 ^ n11079 ^ 1'b0 ;
  assign n16811 = n16807 & n16810 ;
  assign n16812 = n11697 ^ n1577 ^ 1'b0 ;
  assign n16813 = n2322 ^ n1490 ^ 1'b0 ;
  assign n16814 = n14595 ^ n6874 ^ n4664 ;
  assign n16815 = n16813 & ~n16814 ;
  assign n16816 = n16815 ^ n6152 ^ 1'b0 ;
  assign n16817 = n4387 & n6303 ;
  assign n16818 = n16817 ^ n7182 ^ 1'b0 ;
  assign n16819 = ( ~n3163 & n6768 ) | ( ~n3163 & n10049 ) | ( n6768 & n10049 ) ;
  assign n16820 = ~n12542 & n15927 ;
  assign n16821 = n1381 & n16820 ;
  assign n16822 = n1675 & n16821 ;
  assign n16823 = n1461 & n9384 ;
  assign n16824 = n7402 & n16823 ;
  assign n16825 = n16824 ^ n2402 ^ 1'b0 ;
  assign n16826 = ( n3307 & ~n14598 ) | ( n3307 & n16825 ) | ( ~n14598 & n16825 ) ;
  assign n16827 = n2591 | n7820 ;
  assign n16828 = n4245 & ~n8613 ;
  assign n16829 = n16828 ^ n15696 ^ 1'b0 ;
  assign n16830 = n7385 ^ n935 ^ 1'b0 ;
  assign n16831 = n12099 & n16830 ;
  assign n16832 = ( n3128 & ~n13973 ) | ( n3128 & n13997 ) | ( ~n13973 & n13997 ) ;
  assign n16833 = n16085 ^ n15305 ^ 1'b0 ;
  assign n16834 = n1579 ^ n1080 ^ 1'b0 ;
  assign n16835 = n4073 & ~n16834 ;
  assign n16836 = n749 & n2809 ;
  assign n16837 = n16836 ^ n4854 ^ 1'b0 ;
  assign n16838 = ( n10528 & ~n16835 ) | ( n10528 & n16837 ) | ( ~n16835 & n16837 ) ;
  assign n16839 = n9036 ^ n4104 ^ 1'b0 ;
  assign n16840 = n8257 | n16839 ;
  assign n16841 = ( n1162 & n12406 ) | ( n1162 & n16840 ) | ( n12406 & n16840 ) ;
  assign n16842 = n9277 ^ n7070 ^ 1'b0 ;
  assign n16843 = n6319 | n16842 ;
  assign n16844 = n3091 & ~n12870 ;
  assign n16845 = n16844 ^ n6110 ^ 1'b0 ;
  assign n16846 = n2604 ^ n173 ^ 1'b0 ;
  assign n16847 = n3247 & ~n16846 ;
  assign n16848 = n16847 ^ n10846 ^ 1'b0 ;
  assign n16849 = n9573 | n16848 ;
  assign n16850 = n16849 ^ n9548 ^ n9429 ;
  assign n16851 = n4553 ^ n3615 ^ n3002 ;
  assign n16852 = n7700 ^ n1719 ^ 1'b0 ;
  assign n16853 = ( n7276 & ~n16851 ) | ( n7276 & n16852 ) | ( ~n16851 & n16852 ) ;
  assign n16854 = n982 | n3257 ;
  assign n16855 = n16854 ^ n11731 ^ 1'b0 ;
  assign n16856 = ~n1454 & n6530 ;
  assign n16857 = n16856 ^ n575 ^ 1'b0 ;
  assign n16858 = n10690 ^ n5176 ^ 1'b0 ;
  assign n16859 = n14332 & ~n16858 ;
  assign n16860 = ~n9126 & n16859 ;
  assign n16861 = n16860 ^ n16502 ^ 1'b0 ;
  assign n16862 = n16861 ^ n10280 ^ n10112 ;
  assign n16863 = n6541 ^ n795 ^ 1'b0 ;
  assign n16864 = ~n2382 & n16863 ;
  assign n16865 = n1980 | n16864 ;
  assign n16866 = n11805 ^ n11377 ^ n2034 ;
  assign n16867 = n8508 ^ n3371 ^ 1'b0 ;
  assign n16868 = ~n7995 & n16867 ;
  assign n16869 = n16868 ^ n6646 ^ 1'b0 ;
  assign n16870 = n6924 ^ n5997 ^ 1'b0 ;
  assign n16871 = n1090 & n16870 ;
  assign n16872 = ( n3063 & n16869 ) | ( n3063 & ~n16871 ) | ( n16869 & ~n16871 ) ;
  assign n16873 = n14595 ^ n227 ^ 1'b0 ;
  assign n16874 = n16872 | n16873 ;
  assign n16875 = n3174 | n8627 ;
  assign n16879 = n8574 & n10559 ;
  assign n16880 = n16879 ^ n5694 ^ 1'b0 ;
  assign n16876 = n13889 ^ n353 ^ 1'b0 ;
  assign n16877 = n16876 ^ n5492 ^ 1'b0 ;
  assign n16878 = n16587 & ~n16877 ;
  assign n16881 = n16880 ^ n16878 ^ n12043 ;
  assign n16882 = n3037 ^ n2967 ^ 1'b0 ;
  assign n16883 = n1905 | n8482 ;
  assign n16884 = n16883 ^ n3506 ^ 1'b0 ;
  assign n16885 = n491 | n16265 ;
  assign n16886 = n16884 & ~n16885 ;
  assign n16887 = n14668 & ~n16610 ;
  assign n16888 = ~n14583 & n16887 ;
  assign n16889 = n7548 ^ n3513 ^ n1131 ;
  assign n16890 = ~n4593 & n6564 ;
  assign n16891 = n16890 ^ n13521 ^ n13137 ;
  assign n16892 = n1706 & n5352 ;
  assign n16893 = n16892 ^ n1532 ^ 1'b0 ;
  assign n16894 = n16893 ^ n10986 ^ n6327 ;
  assign n16895 = n4870 ^ n1257 ^ 1'b0 ;
  assign n16896 = n6906 & n13618 ;
  assign n16897 = n16895 & n16896 ;
  assign n16898 = n14119 ^ n9935 ^ 1'b0 ;
  assign n16899 = n2650 & ~n16898 ;
  assign n16900 = ( n1611 & n2053 ) | ( n1611 & n11414 ) | ( n2053 & n11414 ) ;
  assign n16901 = ( ~n1534 & n6905 ) | ( ~n1534 & n16900 ) | ( n6905 & n16900 ) ;
  assign n16902 = ~n3238 & n16901 ;
  assign n16903 = n3098 & ~n12948 ;
  assign n16904 = n7023 & ~n16903 ;
  assign n16905 = n5601 & ~n8121 ;
  assign n16906 = n7716 | n16905 ;
  assign n16907 = ( x123 & ~n1125 ) | ( x123 & n11667 ) | ( ~n1125 & n11667 ) ;
  assign n16908 = ( x123 & n6261 ) | ( x123 & n7505 ) | ( n6261 & n7505 ) ;
  assign n16909 = ( n2042 & ~n5754 ) | ( n2042 & n16908 ) | ( ~n5754 & n16908 ) ;
  assign n16910 = ~n16907 & n16909 ;
  assign n16911 = ( n8707 & ~n14803 ) | ( n8707 & n16910 ) | ( ~n14803 & n16910 ) ;
  assign n16912 = n16906 & n16911 ;
  assign n16913 = n2007 | n4878 ;
  assign n16914 = ~n201 & n16913 ;
  assign n16915 = n805 & n8283 ;
  assign n16916 = n16915 ^ n4581 ^ 1'b0 ;
  assign n16917 = ~n300 & n6539 ;
  assign n16918 = n16917 ^ n8188 ^ 1'b0 ;
  assign n16919 = n5357 ^ n2066 ^ 1'b0 ;
  assign n16920 = n16918 & n16919 ;
  assign n16921 = n10848 ^ n9705 ^ n4567 ;
  assign n16922 = n2236 & n16921 ;
  assign n16923 = n9945 ^ n201 ^ 1'b0 ;
  assign n16924 = ~n849 & n16923 ;
  assign n16925 = n16924 ^ n8566 ^ n4774 ;
  assign n16926 = n4709 & n8319 ;
  assign n16927 = ( ~n1678 & n16527 ) | ( ~n1678 & n16926 ) | ( n16527 & n16926 ) ;
  assign n16928 = n7360 ^ n4172 ^ 1'b0 ;
  assign n16929 = n16928 ^ n14169 ^ n13108 ;
  assign n16930 = n13795 & ~n16929 ;
  assign n16931 = n16930 ^ n13824 ^ 1'b0 ;
  assign n16932 = n1036 & ~n4901 ;
  assign n16933 = n16051 | n16932 ;
  assign n16934 = n16933 ^ n4621 ^ 1'b0 ;
  assign n16935 = n3962 & ~n11310 ;
  assign n16936 = n16935 ^ n12809 ^ n12071 ;
  assign n16937 = n12457 ^ n7844 ^ n560 ;
  assign n16938 = n16937 ^ n983 ^ 1'b0 ;
  assign n16939 = n2670 | n3323 ;
  assign n16940 = n11070 ^ n347 ^ 1'b0 ;
  assign n16941 = n4632 & ~n16940 ;
  assign n16942 = n14438 | n16941 ;
  assign n16943 = n16942 ^ n14452 ^ 1'b0 ;
  assign n16944 = n16939 | n16943 ;
  assign n16945 = n7225 & n8550 ;
  assign n16946 = n16944 & n16945 ;
  assign n16947 = ~n1096 & n3221 ;
  assign n16948 = n10768 & n16947 ;
  assign n16949 = n12048 ^ n1502 ^ 1'b0 ;
  assign n16950 = ~n16948 & n16949 ;
  assign n16951 = n11383 ^ n10864 ^ n8243 ;
  assign n16952 = ( n7083 & ~n10334 ) | ( n7083 & n10577 ) | ( ~n10334 & n10577 ) ;
  assign n16953 = n11307 ^ n8058 ^ 1'b0 ;
  assign n16954 = n11082 ^ n10575 ^ 1'b0 ;
  assign n16960 = n2483 & n6017 ;
  assign n16961 = ~n2875 & n16960 ;
  assign n16962 = n4521 | n16961 ;
  assign n16963 = n7219 | n12342 ;
  assign n16964 = n16962 | n16963 ;
  assign n16955 = n3355 ^ n3103 ^ 1'b0 ;
  assign n16956 = n6610 ^ n2315 ^ 1'b0 ;
  assign n16957 = ~n15133 & n16956 ;
  assign n16958 = n16957 ^ n8980 ^ n1731 ;
  assign n16959 = n16955 | n16958 ;
  assign n16965 = n16964 ^ n16959 ^ 1'b0 ;
  assign n16966 = n3974 & ~n12122 ;
  assign n16967 = ~n4402 & n16966 ;
  assign n16968 = n8217 & ~n16967 ;
  assign n16969 = n16968 ^ n14897 ^ 1'b0 ;
  assign n16970 = n589 ^ x15 ^ 1'b0 ;
  assign n16971 = n259 & n16970 ;
  assign n16972 = n16971 ^ n8112 ^ n186 ;
  assign n16973 = n16412 & ~n16972 ;
  assign n16974 = n7119 ^ n6711 ^ 1'b0 ;
  assign n16975 = n1343 & n16974 ;
  assign n16976 = n8432 & n16975 ;
  assign n16977 = n3517 & n16976 ;
  assign n16978 = ( n1094 & n7657 ) | ( n1094 & ~n16977 ) | ( n7657 & ~n16977 ) ;
  assign n16979 = n2364 ^ n2359 ^ 1'b0 ;
  assign n16980 = ~n1704 & n16979 ;
  assign n16981 = n761 | n16980 ;
  assign n16982 = ( n15327 & n15981 ) | ( n15327 & ~n16981 ) | ( n15981 & ~n16981 ) ;
  assign n16983 = n7956 ^ n4235 ^ 1'b0 ;
  assign n16984 = n3349 & n9988 ;
  assign n16985 = n11630 & n16984 ;
  assign n16986 = n16985 ^ n3650 ^ 1'b0 ;
  assign n16987 = n11164 & n16986 ;
  assign n16988 = n16472 ^ n9554 ^ 1'b0 ;
  assign n16989 = ~n8812 & n16988 ;
  assign n16990 = n4978 ^ n4070 ^ n2599 ;
  assign n16991 = n16990 ^ n3862 ^ n784 ;
  assign n16992 = ~n7130 & n16991 ;
  assign n16993 = n16992 ^ n2120 ^ 1'b0 ;
  assign n16994 = n1841 | n3083 ;
  assign n16995 = n4650 & ~n16994 ;
  assign n16996 = n9797 & ~n16995 ;
  assign n16997 = n16996 ^ n1878 ^ 1'b0 ;
  assign n16998 = ~n6851 & n16997 ;
  assign n16999 = n14922 | n16998 ;
  assign n17000 = n16999 ^ n3564 ^ 1'b0 ;
  assign n17001 = n9752 ^ n8184 ^ n3640 ;
  assign n17002 = ( n2905 & ~n4317 ) | ( n2905 & n5599 ) | ( ~n4317 & n5599 ) ;
  assign n17003 = n17002 ^ n16489 ^ n523 ;
  assign n17004 = n686 & n3438 ;
  assign n17005 = ~n445 & n5594 ;
  assign n17006 = n402 & n3802 ;
  assign n17007 = ~n3068 & n17006 ;
  assign n17008 = n14232 ^ n3689 ^ 1'b0 ;
  assign n17009 = n4757 | n17008 ;
  assign n17010 = n17009 ^ n10959 ^ 1'b0 ;
  assign n17011 = ~n17007 & n17010 ;
  assign n17012 = ~n3795 & n17011 ;
  assign n17013 = n17012 ^ n2270 ^ x52 ;
  assign n17014 = ~n1483 & n2982 ;
  assign n17015 = ( x102 & n9847 ) | ( x102 & ~n12024 ) | ( n9847 & ~n12024 ) ;
  assign n17016 = ( n4236 & n17014 ) | ( n4236 & ~n17015 ) | ( n17014 & ~n17015 ) ;
  assign n17017 = ( n3324 & n7520 ) | ( n3324 & ~n10646 ) | ( n7520 & ~n10646 ) ;
  assign n17018 = ( n201 & n3485 ) | ( n201 & ~n17017 ) | ( n3485 & ~n17017 ) ;
  assign n17019 = n1498 & ~n9793 ;
  assign n17020 = ~n6756 & n13984 ;
  assign n17021 = ( n12553 & n17019 ) | ( n12553 & n17020 ) | ( n17019 & n17020 ) ;
  assign n17022 = n12937 & n17021 ;
  assign n17023 = n17022 ^ n1932 ^ 1'b0 ;
  assign n17024 = n1723 & n8855 ;
  assign n17025 = n17024 ^ n2930 ^ 1'b0 ;
  assign n17026 = n6480 ^ n4529 ^ 1'b0 ;
  assign n17027 = n5559 ^ n1743 ^ n1632 ;
  assign n17028 = n17027 ^ n9392 ^ n2029 ;
  assign n17029 = n10952 ^ n3412 ^ n1923 ;
  assign n17030 = n3699 | n5806 ;
  assign n17031 = n13574 ^ n658 ^ 1'b0 ;
  assign n17032 = n6593 & n17031 ;
  assign n17035 = n10849 & ~n13584 ;
  assign n17033 = n1896 & ~n15270 ;
  assign n17034 = n10869 | n17033 ;
  assign n17036 = n17035 ^ n17034 ^ 1'b0 ;
  assign n17037 = ( n10264 & ~n12677 ) | ( n10264 & n13087 ) | ( ~n12677 & n13087 ) ;
  assign n17038 = n17037 ^ n2063 ^ 1'b0 ;
  assign n17039 = n15365 & n17038 ;
  assign n17040 = ( n12714 & ~n12918 ) | ( n12714 & n17039 ) | ( ~n12918 & n17039 ) ;
  assign n17041 = ~n4806 & n6590 ;
  assign n17042 = n8288 ^ n6733 ^ 1'b0 ;
  assign n17043 = ~n17041 & n17042 ;
  assign n17044 = ~n8126 & n11891 ;
  assign n17045 = ( n3525 & ~n17043 ) | ( n3525 & n17044 ) | ( ~n17043 & n17044 ) ;
  assign n17046 = ( ~n1728 & n6005 ) | ( ~n1728 & n17045 ) | ( n6005 & n17045 ) ;
  assign n17047 = n1489 ^ n858 ^ 1'b0 ;
  assign n17048 = n17047 ^ n15339 ^ 1'b0 ;
  assign n17049 = n17048 ^ n3514 ^ 1'b0 ;
  assign n17050 = n9406 & n17049 ;
  assign n17051 = n2236 | n13545 ;
  assign n17052 = n7629 ^ n7065 ^ 1'b0 ;
  assign n17053 = ~n11281 & n17052 ;
  assign n17054 = n4675 & n4901 ;
  assign n17055 = ~n7565 & n17054 ;
  assign n17056 = n17055 ^ n4303 ^ n401 ;
  assign n17057 = n9134 ^ n6003 ^ n4665 ;
  assign n17058 = n17056 & ~n17057 ;
  assign n17059 = ~n709 & n17058 ;
  assign n17061 = n4178 ^ n3406 ^ n2488 ;
  assign n17060 = ~n2342 & n6161 ;
  assign n17062 = n17061 ^ n17060 ^ 1'b0 ;
  assign n17063 = n11422 ^ n5272 ^ n4631 ;
  assign n17064 = n8473 ^ n7482 ^ 1'b0 ;
  assign n17065 = ~n11482 & n17064 ;
  assign n17066 = n8888 & n17065 ;
  assign n17067 = n17066 ^ n13635 ^ n6035 ;
  assign n17068 = ( ~n358 & n4610 ) | ( ~n358 & n13797 ) | ( n4610 & n13797 ) ;
  assign n17069 = n449 | n6676 ;
  assign n17070 = n15951 & ~n17069 ;
  assign n17071 = n11760 | n17070 ;
  assign n17072 = n8760 | n11879 ;
  assign n17073 = n316 & ~n2173 ;
  assign n17074 = n17073 ^ n2751 ^ 1'b0 ;
  assign n17075 = n7699 | n17074 ;
  assign n17076 = n17075 ^ n3912 ^ 1'b0 ;
  assign n17077 = ~n14853 & n17076 ;
  assign n17078 = n17072 & n17077 ;
  assign n17079 = n3755 | n6668 ;
  assign n17080 = n17079 ^ n9623 ^ 1'b0 ;
  assign n17081 = ~n6640 & n17080 ;
  assign n17082 = ( n8024 & ~n10164 ) | ( n8024 & n10180 ) | ( ~n10164 & n10180 ) ;
  assign n17083 = n1585 | n8255 ;
  assign n17084 = n17083 ^ n11471 ^ 1'b0 ;
  assign n17085 = ~n8041 & n17084 ;
  assign n17086 = n1990 & n17085 ;
  assign n17087 = n17086 ^ n15851 ^ n4061 ;
  assign n17088 = ( ~n7610 & n8830 ) | ( ~n7610 & n17087 ) | ( n8830 & n17087 ) ;
  assign n17089 = ( ~n2523 & n3241 ) | ( ~n2523 & n7327 ) | ( n3241 & n7327 ) ;
  assign n17090 = n17089 ^ n6166 ^ 1'b0 ;
  assign n17091 = n17090 ^ n13240 ^ 1'b0 ;
  assign n17092 = n10678 & ~n13426 ;
  assign n17093 = n7004 ^ n3474 ^ 1'b0 ;
  assign n17094 = n2688 & n17093 ;
  assign n17095 = ~n17092 & n17094 ;
  assign n17096 = n17091 & n17095 ;
  assign n17097 = n16061 ^ n3821 ^ 1'b0 ;
  assign n17098 = n14654 & n17097 ;
  assign n17099 = n13777 & ~n17077 ;
  assign n17100 = ( n1528 & n2624 ) | ( n1528 & ~n7821 ) | ( n2624 & ~n7821 ) ;
  assign n17101 = n17100 ^ n5826 ^ 1'b0 ;
  assign n17102 = n3410 ^ n817 ^ 1'b0 ;
  assign n17103 = n17101 & ~n17102 ;
  assign n17104 = n7937 ^ n6631 ^ 1'b0 ;
  assign n17105 = n17104 ^ n14895 ^ n3612 ;
  assign n17106 = ( n1517 & n1921 ) | ( n1517 & n11199 ) | ( n1921 & n11199 ) ;
  assign n17107 = n3193 & n4048 ;
  assign n17108 = n17107 ^ x78 ^ 1'b0 ;
  assign n17109 = n7816 ^ n882 ^ 1'b0 ;
  assign n17110 = n9156 | n17109 ;
  assign n17111 = ( n4148 & n12243 ) | ( n4148 & n16312 ) | ( n12243 & n16312 ) ;
  assign n17119 = n2796 & n4242 ;
  assign n17120 = n17119 ^ n7973 ^ 1'b0 ;
  assign n17121 = n17120 ^ n5094 ^ 1'b0 ;
  assign n17112 = n3515 & n6585 ;
  assign n17113 = n4779 & n17112 ;
  assign n17114 = n6345 ^ n5409 ^ 1'b0 ;
  assign n17115 = n14595 & ~n17114 ;
  assign n17116 = ~n17113 & n17115 ;
  assign n17117 = n17116 ^ n10485 ^ 1'b0 ;
  assign n17118 = x71 & n17117 ;
  assign n17122 = n17121 ^ n17118 ^ 1'b0 ;
  assign n17123 = n8225 ^ n3916 ^ 1'b0 ;
  assign n17127 = n1472 ^ n1390 ^ n440 ;
  assign n17124 = n6746 | n13532 ;
  assign n17125 = n1819 | n4271 ;
  assign n17126 = n17124 & n17125 ;
  assign n17128 = n17127 ^ n17126 ^ 1'b0 ;
  assign n17129 = ( n2462 & ~n11604 ) | ( n2462 & n17128 ) | ( ~n11604 & n17128 ) ;
  assign n17130 = n17129 ^ n4487 ^ n3790 ;
  assign n17131 = n17123 & n17130 ;
  assign n17132 = ~n4787 & n17131 ;
  assign n17133 = n14353 ^ n11733 ^ n4326 ;
  assign n17134 = n4863 & ~n15416 ;
  assign n17135 = n17134 ^ n12677 ^ 1'b0 ;
  assign n17136 = n15863 ^ n9656 ^ 1'b0 ;
  assign n17137 = n1709 & n17136 ;
  assign n17138 = n17137 ^ n7771 ^ n4716 ;
  assign n17139 = ~n1522 & n5137 ;
  assign n17141 = n9397 & n16425 ;
  assign n17142 = n16189 & n17141 ;
  assign n17140 = n1983 & ~n12756 ;
  assign n17143 = n17142 ^ n17140 ^ 1'b0 ;
  assign n17144 = n3866 ^ n2196 ^ 1'b0 ;
  assign n17145 = ~n14500 & n17144 ;
  assign n17146 = n8487 & n17145 ;
  assign n17147 = n16817 ^ n6103 ^ 1'b0 ;
  assign n17148 = n6172 | n17147 ;
  assign n17149 = n4090 | n17148 ;
  assign n17150 = n3366 ^ n1390 ^ 1'b0 ;
  assign n17151 = n17149 & n17150 ;
  assign n17157 = n1476 & ~n8573 ;
  assign n17154 = n7977 ^ n968 ^ 1'b0 ;
  assign n17152 = n727 ^ n458 ^ 1'b0 ;
  assign n17153 = n17152 ^ n6522 ^ 1'b0 ;
  assign n17155 = n17154 ^ n17153 ^ n972 ;
  assign n17156 = n2981 & ~n17155 ;
  assign n17158 = n17157 ^ n17156 ^ 1'b0 ;
  assign n17159 = n3910 & ~n7612 ;
  assign n17160 = n17159 ^ n2879 ^ 1'b0 ;
  assign n17161 = ~n3726 & n17160 ;
  assign n17162 = n9656 & n16379 ;
  assign n17163 = ( n1089 & ~n8513 ) | ( n1089 & n8933 ) | ( ~n8513 & n8933 ) ;
  assign n17164 = n8016 & ~n17163 ;
  assign n17165 = n16443 ^ n2563 ^ 1'b0 ;
  assign n17166 = n17165 ^ n452 ^ 1'b0 ;
  assign n17167 = n9113 & ~n17166 ;
  assign n17168 = n4267 & n17167 ;
  assign n17169 = n4154 & n8345 ;
  assign n17170 = n7376 & n7491 ;
  assign n17171 = n11944 ^ n6632 ^ n1309 ;
  assign n17172 = n17171 ^ n11056 ^ n6991 ;
  assign n17173 = ~n16948 & n17172 ;
  assign n17174 = n4805 & ~n15945 ;
  assign n17175 = n1121 & ~n5355 ;
  assign n17176 = n17175 ^ n2443 ^ 1'b0 ;
  assign n17177 = n17176 ^ n8489 ^ 1'b0 ;
  assign n17178 = n10431 | n17177 ;
  assign n17193 = n4271 ^ n4213 ^ n2638 ;
  assign n17179 = n16813 ^ n4141 ^ n1114 ;
  assign n17187 = n12297 ^ n1374 ^ 1'b0 ;
  assign n17188 = n4942 & ~n17187 ;
  assign n17189 = ~n9742 & n17188 ;
  assign n17190 = ~n713 & n17189 ;
  assign n17180 = ~n412 & n8325 ;
  assign n17181 = ~n3840 & n17180 ;
  assign n17182 = n6997 ^ n4921 ^ 1'b0 ;
  assign n17183 = n2969 | n17182 ;
  assign n17184 = n17181 | n17183 ;
  assign n17185 = n17184 ^ n5834 ^ 1'b0 ;
  assign n17186 = n735 & n17185 ;
  assign n17191 = n17190 ^ n17186 ^ 1'b0 ;
  assign n17192 = n17179 & n17191 ;
  assign n17194 = n17193 ^ n17192 ^ 1'b0 ;
  assign n17199 = ~n2909 & n11203 ;
  assign n17196 = n12742 ^ n4757 ^ n4382 ;
  assign n17195 = n1493 & n6560 ;
  assign n17197 = n17196 ^ n17195 ^ 1'b0 ;
  assign n17198 = n10101 & n17197 ;
  assign n17200 = n17199 ^ n17198 ^ 1'b0 ;
  assign n17201 = n17200 ^ n13476 ^ n992 ;
  assign n17202 = ~n347 & n8551 ;
  assign n17203 = n6517 & ~n9237 ;
  assign n17204 = n8700 ^ n8200 ^ 1'b0 ;
  assign n17205 = ~n7110 & n17204 ;
  assign n17206 = n13347 & n17205 ;
  assign n17207 = n2999 & n17206 ;
  assign n17208 = n17203 | n17207 ;
  assign n17210 = ( n2552 & ~n4009 ) | ( n2552 & n5367 ) | ( ~n4009 & n5367 ) ;
  assign n17209 = ~n10821 & n15966 ;
  assign n17211 = n17210 ^ n17209 ^ n13946 ;
  assign n17212 = n13738 & ~n17211 ;
  assign n17214 = n3734 | n9914 ;
  assign n17215 = n17214 ^ n4601 ^ 1'b0 ;
  assign n17213 = n8994 & ~n14768 ;
  assign n17216 = n17215 ^ n17213 ^ 1'b0 ;
  assign n17217 = n15989 ^ n252 ^ 1'b0 ;
  assign n17218 = n12825 ^ n8382 ^ n626 ;
  assign n17219 = n8801 ^ n7071 ^ 1'b0 ;
  assign n17220 = n9880 & n17219 ;
  assign n17221 = ~n4211 & n17220 ;
  assign n17222 = n17221 ^ n12689 ^ 1'b0 ;
  assign n17223 = ( ~n551 & n1828 ) | ( ~n551 & n2898 ) | ( n1828 & n2898 ) ;
  assign n17224 = n17223 ^ n572 ^ 1'b0 ;
  assign n17225 = n1643 | n17224 ;
  assign n17226 = n1132 | n17225 ;
  assign n17227 = n9680 & ~n11625 ;
  assign n17228 = n17227 ^ n13099 ^ 1'b0 ;
  assign n17229 = ( n10960 & n11310 ) | ( n10960 & ~n17228 ) | ( n11310 & ~n17228 ) ;
  assign n17230 = n2863 | n12614 ;
  assign n17231 = n17230 ^ n7438 ^ 1'b0 ;
  assign n17232 = n4822 ^ x17 ^ 1'b0 ;
  assign n17233 = n17231 & n17232 ;
  assign n17234 = n8205 | n9585 ;
  assign n17235 = n3147 ^ n393 ^ 1'b0 ;
  assign n17236 = n9178 | n17235 ;
  assign n17237 = n17236 ^ n1086 ^ 1'b0 ;
  assign n17238 = ~n2400 & n17237 ;
  assign n17239 = n17238 ^ n7225 ^ n2554 ;
  assign n17240 = ( n2246 & n3015 ) | ( n2246 & ~n7060 ) | ( n3015 & ~n7060 ) ;
  assign n17241 = ~n5887 & n17240 ;
  assign n17242 = n4498 | n5007 ;
  assign n17243 = n10559 ^ n8741 ^ n6439 ;
  assign n17244 = ( ~n16880 & n17242 ) | ( ~n16880 & n17243 ) | ( n17242 & n17243 ) ;
  assign n17245 = n2213 & n17244 ;
  assign n17246 = n9164 & n17245 ;
  assign n17250 = ( n7662 & n10720 ) | ( n7662 & n14247 ) | ( n10720 & n14247 ) ;
  assign n17251 = n1815 | n17250 ;
  assign n17252 = n15536 | n17251 ;
  assign n17247 = ~n9843 & n16980 ;
  assign n17248 = n7383 & n17247 ;
  assign n17249 = n4658 & ~n17248 ;
  assign n17253 = n17252 ^ n17249 ^ 1'b0 ;
  assign n17254 = n8529 ^ n7004 ^ 1'b0 ;
  assign n17255 = n165 | n17254 ;
  assign n17256 = n2064 & ~n12235 ;
  assign n17257 = n17255 & n17256 ;
  assign n17258 = n13707 | n17257 ;
  assign n17259 = n10257 & n17258 ;
  assign n17260 = n7023 ^ n1110 ^ n975 ;
  assign n17261 = n4697 | n17260 ;
  assign n17262 = n14316 | n17261 ;
  assign n17263 = n13724 ^ n8576 ^ 1'b0 ;
  assign n17265 = ~n194 & n11694 ;
  assign n17264 = n9652 ^ n7923 ^ 1'b0 ;
  assign n17266 = n17265 ^ n17264 ^ 1'b0 ;
  assign n17267 = n6889 & n16448 ;
  assign n17268 = n15044 ^ n10328 ^ 1'b0 ;
  assign n17269 = n6877 & ~n17268 ;
  assign n17270 = ~n11304 & n13816 ;
  assign n17271 = ( n3318 & n17269 ) | ( n3318 & n17270 ) | ( n17269 & n17270 ) ;
  assign n17272 = n5465 ^ n3042 ^ 1'b0 ;
  assign n17273 = n3581 & ~n17272 ;
  assign n17274 = n168 & n17273 ;
  assign n17275 = n17274 ^ n7717 ^ 1'b0 ;
  assign n17276 = ~n8585 & n17275 ;
  assign n17277 = n17276 ^ n5402 ^ 1'b0 ;
  assign n17278 = n2098 & ~n11134 ;
  assign n17279 = n9697 & n17278 ;
  assign n17280 = n17277 & n17279 ;
  assign n17282 = ~n6878 & n15755 ;
  assign n17281 = ~n1418 & n11802 ;
  assign n17283 = n17282 ^ n17281 ^ 1'b0 ;
  assign n17284 = n5543 & ~n17283 ;
  assign n17285 = n17284 ^ n13582 ^ 1'b0 ;
  assign n17286 = ~n181 & n2924 ;
  assign n17287 = n17286 ^ n1651 ^ 1'b0 ;
  assign n17288 = ( ~n5328 & n6746 ) | ( ~n5328 & n17287 ) | ( n6746 & n17287 ) ;
  assign n17289 = ( n1794 & n1929 ) | ( n1794 & ~n17288 ) | ( n1929 & ~n17288 ) ;
  assign n17290 = ( n320 & n2834 ) | ( n320 & ~n8406 ) | ( n2834 & ~n8406 ) ;
  assign n17291 = n9046 & ~n9864 ;
  assign n17292 = n17290 & n17291 ;
  assign n17293 = n3485 & n4337 ;
  assign n17294 = ~n16395 & n17293 ;
  assign n17295 = n17292 & ~n17294 ;
  assign n17296 = x92 & n3540 ;
  assign n17297 = n5851 | n10290 ;
  assign n17298 = n4128 | n8522 ;
  assign n17299 = n17298 ^ n16595 ^ 1'b0 ;
  assign n17300 = n6064 & n10857 ;
  assign n17301 = n14012 & n17300 ;
  assign n17302 = ~n210 & n4188 ;
  assign n17303 = ~n13361 & n17302 ;
  assign n17304 = n5726 ^ n1318 ^ 1'b0 ;
  assign n17305 = n7295 & ~n8727 ;
  assign n17306 = n10398 & n17305 ;
  assign n17307 = n16720 & n17306 ;
  assign n17308 = n3719 ^ n2799 ^ 1'b0 ;
  assign n17309 = n3375 & ~n6671 ;
  assign n17310 = n16358 & n17309 ;
  assign n17311 = n8631 & ~n17310 ;
  assign n17312 = n14221 ^ n8065 ^ 1'b0 ;
  assign n17313 = n2738 & ~n17312 ;
  assign n17314 = n5384 ^ n3449 ^ 1'b0 ;
  assign n17315 = n12361 & n17314 ;
  assign n17316 = n17313 & ~n17315 ;
  assign n17317 = n17316 ^ n1160 ^ 1'b0 ;
  assign n17318 = ( n6226 & n11352 ) | ( n6226 & n17317 ) | ( n11352 & n17317 ) ;
  assign n17319 = n17318 ^ n2087 ^ 1'b0 ;
  assign n17320 = n13646 | n17319 ;
  assign n17321 = ( n17308 & ~n17311 ) | ( n17308 & n17320 ) | ( ~n17311 & n17320 ) ;
  assign n17322 = n14087 & ~n17321 ;
  assign n17323 = n17307 & n17322 ;
  assign n17324 = n5385 ^ n2002 ^ 1'b0 ;
  assign n17325 = n10734 | n16850 ;
  assign n17326 = n17324 | n17325 ;
  assign n17330 = n7182 ^ n3654 ^ n3564 ;
  assign n17331 = ( n4881 & ~n13796 ) | ( n4881 & n17330 ) | ( ~n13796 & n17330 ) ;
  assign n17328 = ~n5199 & n10753 ;
  assign n17327 = n10888 & n16634 ;
  assign n17329 = n17328 ^ n17327 ^ 1'b0 ;
  assign n17332 = n17331 ^ n17329 ^ 1'b0 ;
  assign n17333 = n10656 ^ n2524 ^ 1'b0 ;
  assign n17334 = n11555 ^ n3413 ^ 1'b0 ;
  assign n17335 = n17333 | n17334 ;
  assign n17336 = n17335 ^ n5501 ^ 1'b0 ;
  assign n17337 = n17332 & ~n17336 ;
  assign n17338 = n4207 & ~n11084 ;
  assign n17339 = n3613 & n17338 ;
  assign n17340 = n1798 ^ n391 ^ 1'b0 ;
  assign n17341 = ( n2048 & n17339 ) | ( n2048 & n17340 ) | ( n17339 & n17340 ) ;
  assign n17342 = ( n8426 & n13368 ) | ( n8426 & n17341 ) | ( n13368 & n17341 ) ;
  assign n17343 = ( ~n1782 & n2972 ) | ( ~n1782 & n16103 ) | ( n2972 & n16103 ) ;
  assign n17344 = n17342 | n17343 ;
  assign n17345 = n13868 | n17344 ;
  assign n17346 = n9324 | n16876 ;
  assign n17347 = ( n4867 & ~n5864 ) | ( n4867 & n17346 ) | ( ~n5864 & n17346 ) ;
  assign n17348 = ~n793 & n12786 ;
  assign n17349 = ( n1139 & n3597 ) | ( n1139 & ~n3678 ) | ( n3597 & ~n3678 ) ;
  assign n17350 = n17348 | n17349 ;
  assign n17351 = ( n12852 & n15229 ) | ( n12852 & n17350 ) | ( n15229 & n17350 ) ;
  assign n17352 = n16564 ^ n11259 ^ 1'b0 ;
  assign n17353 = n1362 & ~n2976 ;
  assign n17354 = n3923 & ~n5678 ;
  assign n17355 = ~n3923 & n17354 ;
  assign n17356 = n1969 | n8746 ;
  assign n17357 = n8746 & ~n17356 ;
  assign n17358 = n859 | n1973 ;
  assign n17359 = n17357 & ~n17358 ;
  assign n17360 = n17355 | n17359 ;
  assign n17361 = n17355 & ~n17360 ;
  assign n17362 = n10411 | n17361 ;
  assign n17363 = n10411 & ~n17362 ;
  assign n17364 = n148 & ~n1014 ;
  assign n17365 = ~n148 & n17364 ;
  assign n17366 = ~n2680 & n17365 ;
  assign n17367 = n3173 | n3831 ;
  assign n17368 = n17366 & ~n17367 ;
  assign n17369 = ~n660 & n17368 ;
  assign n17370 = n5419 & n17369 ;
  assign n17371 = ~n5419 & n17370 ;
  assign n17372 = n3278 ^ n2243 ^ 1'b0 ;
  assign n17373 = n17371 | n17372 ;
  assign n17374 = n17363 | n17373 ;
  assign n17375 = n17353 | n17374 ;
  assign n17376 = n17375 ^ n11247 ^ 1'b0 ;
  assign n17377 = n5347 & n13426 ;
  assign n17379 = n13961 ^ n2666 ^ 1'b0 ;
  assign n17380 = ~n9260 & n17379 ;
  assign n17381 = n17380 ^ n5406 ^ 1'b0 ;
  assign n17378 = n2018 & ~n8146 ;
  assign n17382 = n17381 ^ n17378 ^ 1'b0 ;
  assign n17383 = ~n3244 & n11645 ;
  assign n17384 = n17383 ^ n15442 ^ 1'b0 ;
  assign n17386 = n14058 ^ n6297 ^ 1'b0 ;
  assign n17387 = n7534 & ~n17386 ;
  assign n17385 = n7469 | n9078 ;
  assign n17388 = n17387 ^ n17385 ^ 1'b0 ;
  assign n17389 = ( n1532 & n1997 ) | ( n1532 & ~n9044 ) | ( n1997 & ~n9044 ) ;
  assign n17390 = n2625 & n10080 ;
  assign n17391 = n17390 ^ n8156 ^ 1'b0 ;
  assign n17392 = ( n14812 & ~n17389 ) | ( n14812 & n17391 ) | ( ~n17389 & n17391 ) ;
  assign n17393 = n9171 ^ n8791 ^ n142 ;
  assign n17394 = n16023 ^ n7035 ^ 1'b0 ;
  assign n17395 = ( n2753 & n6140 ) | ( n2753 & n9970 ) | ( n6140 & n9970 ) ;
  assign n17396 = n17395 ^ n8033 ^ 1'b0 ;
  assign n17398 = n3788 ^ n2041 ^ n1408 ;
  assign n17397 = ~n3722 & n11443 ;
  assign n17399 = n17398 ^ n17397 ^ 1'b0 ;
  assign n17400 = ( ~n447 & n1096 ) | ( ~n447 & n5568 ) | ( n1096 & n5568 ) ;
  assign n17401 = n17400 ^ n11697 ^ 1'b0 ;
  assign n17402 = n17399 & n17401 ;
  assign n17404 = n11266 ^ n9092 ^ n8201 ;
  assign n17403 = n2416 & n17053 ;
  assign n17405 = n17404 ^ n17403 ^ 1'b0 ;
  assign n17409 = n1186 & n3505 ;
  assign n17410 = n17409 ^ n1238 ^ 1'b0 ;
  assign n17406 = n12552 ^ n1808 ^ 1'b0 ;
  assign n17407 = n2740 & ~n17406 ;
  assign n17408 = n990 | n17407 ;
  assign n17411 = n17410 ^ n17408 ^ n4756 ;
  assign n17412 = n13880 ^ n6772 ^ n3739 ;
  assign n17413 = ~n1233 & n17412 ;
  assign n17414 = ~n3218 & n17413 ;
  assign n17415 = n9345 | n17414 ;
  assign n17416 = n17415 ^ n8217 ^ 1'b0 ;
  assign n17417 = n4199 | n15863 ;
  assign n17418 = n13314 & ~n17417 ;
  assign n17419 = n998 & n6875 ;
  assign n17420 = n17419 ^ n5040 ^ 1'b0 ;
  assign n17421 = n8335 & ~n17420 ;
  assign n17422 = ~n7870 & n17421 ;
  assign n17423 = n17422 ^ n15440 ^ 1'b0 ;
  assign n17424 = n5397 ^ n2728 ^ 1'b0 ;
  assign n17425 = n14768 | n17424 ;
  assign n17426 = n10909 & ~n17425 ;
  assign n17427 = ( n923 & n6237 ) | ( n923 & n6388 ) | ( n6237 & n6388 ) ;
  assign n17428 = n4155 & ~n5831 ;
  assign n17429 = ( ~n4239 & n17427 ) | ( ~n4239 & n17428 ) | ( n17427 & n17428 ) ;
  assign n17430 = ( n4422 & n7085 ) | ( n4422 & ~n13268 ) | ( n7085 & ~n13268 ) ;
  assign n17431 = n17430 ^ n16187 ^ n15111 ;
  assign n17432 = n6271 ^ n1177 ^ x81 ;
  assign n17433 = n17432 ^ n1906 ^ 1'b0 ;
  assign n17434 = n3407 & n17433 ;
  assign n17438 = n1564 & n9894 ;
  assign n17435 = n9921 | n9970 ;
  assign n17436 = n7398 | n17435 ;
  assign n17437 = n712 & n17436 ;
  assign n17439 = n17438 ^ n17437 ^ 1'b0 ;
  assign n17440 = n16261 ^ n8955 ^ n5997 ;
  assign n17441 = n4971 & ~n17440 ;
  assign n17442 = n17441 ^ n4328 ^ 1'b0 ;
  assign n17443 = n3316 ^ n2278 ^ n2041 ;
  assign n17444 = ~n3469 & n5599 ;
  assign n17445 = n7657 & n17444 ;
  assign n17446 = n8209 ^ n3222 ^ n3102 ;
  assign n17448 = ~n3851 & n6439 ;
  assign n17449 = n17448 ^ n4442 ^ 1'b0 ;
  assign n17450 = n2262 | n17449 ;
  assign n17447 = n2501 & n3988 ;
  assign n17451 = n17450 ^ n17447 ^ 1'b0 ;
  assign n17452 = n17451 ^ n6851 ^ n4414 ;
  assign n17453 = ( ~n17445 & n17446 ) | ( ~n17445 & n17452 ) | ( n17446 & n17452 ) ;
  assign n17454 = n12783 ^ n5237 ^ 1'b0 ;
  assign n17455 = n9630 | n17454 ;
  assign n17456 = ~n441 & n5224 ;
  assign n17457 = n12940 & ~n17456 ;
  assign n17458 = n1214 & n17457 ;
  assign n17459 = n8692 ^ n2607 ^ 1'b0 ;
  assign n17460 = n1723 & n17459 ;
  assign n17461 = ~n6789 & n10168 ;
  assign n17462 = ~n17460 & n17461 ;
  assign n17463 = ( n1894 & n12004 ) | ( n1894 & n17462 ) | ( n12004 & n17462 ) ;
  assign n17464 = ~n293 & n7307 ;
  assign n17465 = n10369 ^ n7246 ^ 1'b0 ;
  assign n17466 = n14208 & n17465 ;
  assign n17467 = ~n9591 & n11422 ;
  assign n17468 = n17467 ^ n9260 ^ 1'b0 ;
  assign n17469 = n17468 ^ n13530 ^ 1'b0 ;
  assign n17470 = n2215 & ~n15291 ;
  assign n17471 = ~n17469 & n17470 ;
  assign n17474 = n4422 & ~n4861 ;
  assign n17473 = n14737 ^ n1347 ^ 1'b0 ;
  assign n17472 = n7234 ^ n1928 ^ n540 ;
  assign n17475 = n17474 ^ n17473 ^ n17472 ;
  assign n17476 = n5219 ^ n2366 ^ 1'b0 ;
  assign n17477 = n17476 ^ n10335 ^ 1'b0 ;
  assign n17478 = n11557 ^ n8033 ^ n4627 ;
  assign n17479 = n17478 ^ n9279 ^ 1'b0 ;
  assign n17480 = ~n4719 & n17479 ;
  assign n17481 = n1713 | n8573 ;
  assign n17482 = n17481 ^ n701 ^ 1'b0 ;
  assign n17483 = n7192 & ~n12209 ;
  assign n17484 = n5986 | n17483 ;
  assign n17485 = n17484 ^ n2077 ^ 1'b0 ;
  assign n17486 = n2575 & ~n17485 ;
  assign n17487 = ~n17482 & n17486 ;
  assign n17488 = ~n17480 & n17487 ;
  assign n17489 = n15402 ^ n3342 ^ n2651 ;
  assign n17490 = n17489 ^ n11255 ^ 1'b0 ;
  assign n17491 = ~n13378 & n17490 ;
  assign n17492 = n7011 | n11536 ;
  assign n17493 = n5873 & ~n17492 ;
  assign n17494 = n8695 ^ n7006 ^ 1'b0 ;
  assign n17495 = ~n11128 & n17494 ;
  assign n17499 = n12361 ^ n4360 ^ 1'b0 ;
  assign n17500 = n4300 | n17499 ;
  assign n17496 = n1280 | n6996 ;
  assign n17497 = x92 | n17496 ;
  assign n17498 = n17497 ^ n9401 ^ n594 ;
  assign n17501 = n17500 ^ n17498 ^ n7803 ;
  assign n17502 = n17501 ^ n2582 ^ 1'b0 ;
  assign n17503 = n17495 & n17502 ;
  assign n17506 = n693 & n7213 ;
  assign n17505 = n6085 & n10699 ;
  assign n17507 = n17506 ^ n17505 ^ 1'b0 ;
  assign n17504 = n15817 ^ n14781 ^ 1'b0 ;
  assign n17508 = n17507 ^ n17504 ^ n9924 ;
  assign n17509 = ~n2741 & n9655 ;
  assign n17510 = n3787 & n17509 ;
  assign n17511 = n17510 ^ n16935 ^ n15777 ;
  assign n17512 = n6846 & n7962 ;
  assign n17513 = ( ~n2388 & n3019 ) | ( ~n2388 & n5225 ) | ( n3019 & n5225 ) ;
  assign n17520 = ( n1469 & n1645 ) | ( n1469 & n3728 ) | ( n1645 & n3728 ) ;
  assign n17514 = n14336 ^ n10956 ^ n8029 ;
  assign n17517 = n12442 ^ n3693 ^ 1'b0 ;
  assign n17515 = n4488 ^ n2878 ^ n972 ;
  assign n17516 = n2471 & n17515 ;
  assign n17518 = n17517 ^ n17516 ^ 1'b0 ;
  assign n17519 = n17514 & ~n17518 ;
  assign n17521 = n17520 ^ n17519 ^ 1'b0 ;
  assign n17522 = n4991 ^ n1626 ^ x7 ;
  assign n17523 = ( ~n3122 & n14543 ) | ( ~n3122 & n17522 ) | ( n14543 & n17522 ) ;
  assign n17524 = ( n3412 & n14113 ) | ( n3412 & n17523 ) | ( n14113 & n17523 ) ;
  assign n17525 = ~n15943 & n17524 ;
  assign n17526 = ~n6111 & n11808 ;
  assign n17527 = n2595 | n9392 ;
  assign n17528 = n16851 & ~n17527 ;
  assign n17529 = ( ~n3330 & n8218 ) | ( ~n3330 & n12277 ) | ( n8218 & n12277 ) ;
  assign n17530 = n10154 ^ n4889 ^ n302 ;
  assign n17531 = n15256 & ~n17530 ;
  assign n17532 = ~n1080 & n5514 ;
  assign n17533 = n17532 ^ n5526 ^ 1'b0 ;
  assign n17534 = n11776 ^ n8736 ^ 1'b0 ;
  assign n17535 = n17533 | n17534 ;
  assign n17536 = n12801 ^ n1230 ^ n381 ;
  assign n17537 = ( n4802 & ~n6756 ) | ( n4802 & n16274 ) | ( ~n6756 & n16274 ) ;
  assign n17538 = n2365 & n6539 ;
  assign n17539 = n17538 ^ n1351 ^ 1'b0 ;
  assign n17540 = n5159 & n5241 ;
  assign n17541 = n17540 ^ n2779 ^ 1'b0 ;
  assign n17542 = n17541 ^ n8299 ^ 1'b0 ;
  assign n17543 = ~n17539 & n17542 ;
  assign n17544 = n16500 ^ n360 ^ 1'b0 ;
  assign n17545 = n17544 ^ n11315 ^ n2273 ;
  assign n17546 = ( n9121 & n10080 ) | ( n9121 & n15431 ) | ( n10080 & n15431 ) ;
  assign n17547 = n8777 ^ n7408 ^ n641 ;
  assign n17548 = n6442 & ~n17547 ;
  assign n17549 = n7021 ^ n6808 ^ 1'b0 ;
  assign n17550 = ( n3648 & n3650 ) | ( n3648 & n5841 ) | ( n3650 & n5841 ) ;
  assign n17551 = n17550 ^ x114 ^ 1'b0 ;
  assign n17552 = n593 | n17551 ;
  assign n17553 = n14471 & ~n14620 ;
  assign n17554 = ( n3540 & ~n17552 ) | ( n3540 & n17553 ) | ( ~n17552 & n17553 ) ;
  assign n17555 = ( n7665 & n9158 ) | ( n7665 & ~n14736 ) | ( n9158 & ~n14736 ) ;
  assign n17556 = n17555 ^ n6017 ^ 1'b0 ;
  assign n17557 = n4950 & ~n17556 ;
  assign n17558 = n17557 ^ n2082 ^ n2030 ;
  assign n17560 = n2408 & ~n9439 ;
  assign n17561 = n3142 & ~n6818 ;
  assign n17562 = n17561 ^ n1389 ^ 1'b0 ;
  assign n17563 = ~n17560 & n17562 ;
  assign n17564 = ~n12514 & n17563 ;
  assign n17559 = n3968 & ~n6909 ;
  assign n17565 = n17564 ^ n17559 ^ 1'b0 ;
  assign n17566 = n8276 & n9969 ;
  assign n17567 = ~n13922 & n17566 ;
  assign n17568 = ~n3389 & n7844 ;
  assign n17569 = n17568 ^ n12621 ^ 1'b0 ;
  assign n17570 = n17569 ^ n10106 ^ 1'b0 ;
  assign n17571 = n12834 ^ n9135 ^ 1'b0 ;
  assign n17572 = n10011 & n17571 ;
  assign n17576 = n6195 | n8460 ;
  assign n17573 = n11743 ^ n3393 ^ n517 ;
  assign n17574 = n8316 & n17573 ;
  assign n17575 = ~n5895 & n17574 ;
  assign n17577 = n17576 ^ n17575 ^ n10731 ;
  assign n17578 = n11632 ^ n5453 ^ 1'b0 ;
  assign n17579 = n7356 ^ n1928 ^ 1'b0 ;
  assign n17580 = n162 & n17579 ;
  assign n17581 = n6769 & n17580 ;
  assign n17582 = n4616 & n10791 ;
  assign n17583 = n3935 & ~n12841 ;
  assign n17584 = n16076 & n17583 ;
  assign n17585 = n3905 ^ n3326 ^ 1'b0 ;
  assign n17586 = ( ~x31 & n6043 ) | ( ~x31 & n6775 ) | ( n6043 & n6775 ) ;
  assign n17587 = n17586 ^ n8129 ^ n2248 ;
  assign n17588 = n17587 ^ n10692 ^ n1955 ;
  assign n17589 = ( n12183 & ~n15431 ) | ( n12183 & n16847 ) | ( ~n15431 & n16847 ) ;
  assign n17590 = n7497 ^ n5700 ^ 1'b0 ;
  assign n17591 = n4088 ^ n2592 ^ n327 ;
  assign n17592 = x64 & ~n17591 ;
  assign n17593 = ~n12303 & n17592 ;
  assign n17594 = ~n3123 & n17593 ;
  assign n17595 = n17594 ^ n7784 ^ 1'b0 ;
  assign n17596 = n11514 ^ n9906 ^ 1'b0 ;
  assign n17597 = n12516 & n17596 ;
  assign n17598 = n16149 ^ n4483 ^ n2756 ;
  assign n17599 = n398 & ~n8100 ;
  assign n17600 = n725 | n8348 ;
  assign n17601 = n11915 | n17600 ;
  assign n17602 = n2182 & ~n16997 ;
  assign n17603 = ( ~n1463 & n17601 ) | ( ~n1463 & n17602 ) | ( n17601 & n17602 ) ;
  assign n17604 = ( n17598 & ~n17599 ) | ( n17598 & n17603 ) | ( ~n17599 & n17603 ) ;
  assign n17606 = n1700 & ~n3441 ;
  assign n17607 = n8677 & n17606 ;
  assign n17605 = n9901 & n14705 ;
  assign n17608 = n17607 ^ n17605 ^ 1'b0 ;
  assign n17609 = n2595 | n4704 ;
  assign n17610 = n17609 ^ n6326 ^ 1'b0 ;
  assign n17611 = n10925 & ~n17610 ;
  assign n17612 = n1715 & n17611 ;
  assign n17618 = n10922 ^ n4052 ^ 1'b0 ;
  assign n17619 = ~n2285 & n17618 ;
  assign n17613 = n4994 | n9176 ;
  assign n17614 = n17613 ^ n3621 ^ 1'b0 ;
  assign n17615 = n7183 ^ n6988 ^ 1'b0 ;
  assign n17616 = ~n17614 & n17615 ;
  assign n17617 = ~n1867 & n17616 ;
  assign n17620 = n17619 ^ n17617 ^ 1'b0 ;
  assign n17621 = n2846 & ~n7077 ;
  assign n17622 = n17046 & n17621 ;
  assign n17623 = n16529 ^ n4052 ^ 1'b0 ;
  assign n17624 = n13362 ^ n1528 ^ 1'b0 ;
  assign n17625 = n17623 & ~n17624 ;
  assign n17626 = ( n3466 & n3541 ) | ( n3466 & n3785 ) | ( n3541 & n3785 ) ;
  assign n17627 = ~n6635 & n17626 ;
  assign n17628 = n4286 & n5440 ;
  assign n17629 = ( n8599 & n17627 ) | ( n8599 & n17628 ) | ( n17627 & n17628 ) ;
  assign n17630 = n6717 & ~n8643 ;
  assign n17631 = ( n775 & n2269 ) | ( n775 & ~n2493 ) | ( n2269 & ~n2493 ) ;
  assign n17632 = n11643 & n17631 ;
  assign n17633 = n11107 ^ n5195 ^ 1'b0 ;
  assign n17634 = ~n17632 & n17633 ;
  assign n17635 = ~n6747 & n15236 ;
  assign n17636 = n9791 ^ n459 ^ 1'b0 ;
  assign n17637 = n1330 ^ n1320 ^ 1'b0 ;
  assign n17638 = n17636 & ~n17637 ;
  assign n17639 = n1687 | n3900 ;
  assign n17640 = n5183 & ~n17639 ;
  assign n17641 = ~n4667 & n13451 ;
  assign n17642 = n10867 & n17641 ;
  assign n17643 = ~n7978 & n17642 ;
  assign n17644 = n9302 & ~n17643 ;
  assign n17645 = n3317 | n7527 ;
  assign n17646 = n12302 ^ n4956 ^ 1'b0 ;
  assign n17647 = n10048 & ~n17646 ;
  assign n17648 = n4543 & n17647 ;
  assign n17649 = n4785 & n7311 ;
  assign n17650 = n17649 ^ n9215 ^ 1'b0 ;
  assign n17651 = ~n2296 & n5323 ;
  assign n17652 = n17651 ^ n5208 ^ 1'b0 ;
  assign n17653 = n17652 ^ n6758 ^ n2822 ;
  assign n17654 = ( n1907 & n5263 ) | ( n1907 & ~n17653 ) | ( n5263 & ~n17653 ) ;
  assign n17655 = n1537 & n3910 ;
  assign n17656 = n17655 ^ n1129 ^ 1'b0 ;
  assign n17657 = n17656 ^ n10335 ^ 1'b0 ;
  assign n17658 = n12234 ^ n1818 ^ 1'b0 ;
  assign n17659 = n17658 ^ n9314 ^ n982 ;
  assign n17660 = n3568 & n16957 ;
  assign n17661 = n17660 ^ n788 ^ 1'b0 ;
  assign n17662 = ~n7753 & n10036 ;
  assign n17663 = n2823 ^ n2768 ^ 1'b0 ;
  assign n17664 = n2650 & n17663 ;
  assign n17665 = x63 & ~n17664 ;
  assign n17666 = ( ~n1150 & n2159 ) | ( ~n1150 & n16299 ) | ( n2159 & n16299 ) ;
  assign n17667 = n12052 ^ n5357 ^ n2870 ;
  assign n17668 = n14421 & n17667 ;
  assign n17669 = ~n17666 & n17668 ;
  assign n17670 = n8346 & ~n12289 ;
  assign n17671 = n17670 ^ n16786 ^ 1'b0 ;
  assign n17672 = ~n12632 & n17146 ;
  assign n17673 = n15549 ^ n14135 ^ n11339 ;
  assign n17674 = n6938 & n15236 ;
  assign n17675 = ~n12144 & n17674 ;
  assign n17676 = n15809 ^ n10335 ^ 1'b0 ;
  assign n17677 = n2443 & ~n17676 ;
  assign n17678 = n4614 & n15093 ;
  assign n17679 = n12681 ^ n11118 ^ n10652 ;
  assign n17680 = n11147 ^ n6949 ^ 1'b0 ;
  assign n17681 = n3025 | n17680 ;
  assign n17682 = n17681 ^ n4550 ^ 1'b0 ;
  assign n17683 = n12781 ^ n1033 ^ 1'b0 ;
  assign n17684 = n7296 ^ n4312 ^ 1'b0 ;
  assign n17685 = n9177 | n17684 ;
  assign n17686 = ( n8478 & n12521 ) | ( n8478 & ~n17685 ) | ( n12521 & ~n17685 ) ;
  assign n17687 = n2268 | n17686 ;
  assign n17688 = n302 & n6605 ;
  assign n17689 = ( ~n1475 & n5236 ) | ( ~n1475 & n7287 ) | ( n5236 & n7287 ) ;
  assign n17690 = n5537 & ~n17689 ;
  assign n17691 = n17690 ^ n14553 ^ n550 ;
  assign n17692 = n5258 & ~n11027 ;
  assign n17693 = n7333 ^ n4393 ^ n2524 ;
  assign n17694 = ( ~n8217 & n17692 ) | ( ~n8217 & n17693 ) | ( n17692 & n17693 ) ;
  assign n17695 = ~n6852 & n17694 ;
  assign n17696 = n17695 ^ n219 ^ 1'b0 ;
  assign n17700 = n4618 ^ n1818 ^ n1076 ;
  assign n17697 = n3022 & ~n14395 ;
  assign n17698 = n17697 ^ n284 ^ 1'b0 ;
  assign n17699 = ( n1825 & n5698 ) | ( n1825 & n17698 ) | ( n5698 & n17698 ) ;
  assign n17701 = n17700 ^ n17699 ^ 1'b0 ;
  assign n17703 = n8052 & n8467 ;
  assign n17704 = ~n10030 & n17703 ;
  assign n17705 = n17704 ^ n6412 ^ 1'b0 ;
  assign n17702 = n1441 & n16668 ;
  assign n17706 = n17705 ^ n17702 ^ 1'b0 ;
  assign n17707 = n4295 & ~n9168 ;
  assign n17708 = ( ~n3245 & n10340 ) | ( ~n3245 & n11769 ) | ( n10340 & n11769 ) ;
  assign n17709 = n3372 | n17708 ;
  assign n17710 = n9125 ^ n2090 ^ 1'b0 ;
  assign n17711 = n17709 & ~n17710 ;
  assign n17712 = n3962 & n14757 ;
  assign n17713 = ~n14189 & n17712 ;
  assign n17714 = n17713 ^ n10495 ^ 1'b0 ;
  assign n17715 = n1173 & ~n17714 ;
  assign n17716 = n8033 ^ n2497 ^ 1'b0 ;
  assign n17717 = n2748 | n17716 ;
  assign n17718 = n11315 & ~n17717 ;
  assign n17719 = n10611 & n17718 ;
  assign n17720 = n17719 ^ n12697 ^ 1'b0 ;
  assign n17721 = n10912 & n17720 ;
  assign n17722 = n3392 & n7479 ;
  assign n17723 = n17722 ^ n12949 ^ n11161 ;
  assign n17724 = ~n8065 & n16304 ;
  assign n17725 = ( n1354 & ~n1552 ) | ( n1354 & n15229 ) | ( ~n1552 & n15229 ) ;
  assign n17726 = n634 & n4660 ;
  assign n17727 = ~n3428 & n17726 ;
  assign n17728 = n2303 & n4574 ;
  assign n17729 = n17727 & n17728 ;
  assign n17730 = n1394 & n9784 ;
  assign n17731 = ~n9744 & n17730 ;
  assign n17732 = n11465 ^ n2236 ^ n1721 ;
  assign n17733 = n1515 | n7897 ;
  assign n17734 = n17733 ^ n12554 ^ 1'b0 ;
  assign n17735 = n8609 ^ n3441 ^ 1'b0 ;
  assign n17736 = n17734 & ~n17735 ;
  assign n17737 = n17736 ^ n9961 ^ n5832 ;
  assign n17738 = x77 & ~n16895 ;
  assign n17739 = n14773 & n17738 ;
  assign n17740 = n5076 & n9052 ;
  assign n17741 = n17740 ^ n773 ^ 1'b0 ;
  assign n17742 = ( ~n7466 & n17739 ) | ( ~n7466 & n17741 ) | ( n17739 & n17741 ) ;
  assign n17743 = ( n7121 & n7458 ) | ( n7121 & ~n17742 ) | ( n7458 & ~n17742 ) ;
  assign n17744 = ( ~n4623 & n9472 ) | ( ~n4623 & n10204 ) | ( n9472 & n10204 ) ;
  assign n17745 = n6714 ^ n4559 ^ 1'b0 ;
  assign n17746 = n9383 | n17745 ;
  assign n17747 = n17746 ^ n6984 ^ 1'b0 ;
  assign n17748 = n15561 | n17747 ;
  assign n17749 = ( n4050 & ~n5614 ) | ( n4050 & n13868 ) | ( ~n5614 & n13868 ) ;
  assign n17750 = n6305 & ~n17749 ;
  assign n17751 = n6758 & n17750 ;
  assign n17752 = n1465 & n14149 ;
  assign n17754 = n14201 ^ n3877 ^ n2622 ;
  assign n17755 = ~n1510 & n17754 ;
  assign n17753 = n5597 & ~n10789 ;
  assign n17756 = n17755 ^ n17753 ^ 1'b0 ;
  assign n17757 = ~n378 & n4733 ;
  assign n17758 = n12255 & ~n17757 ;
  assign n17759 = ~n6715 & n17758 ;
  assign n17760 = x15 & n9406 ;
  assign n17761 = n6832 & n17760 ;
  assign n17762 = n17759 | n17761 ;
  assign n17763 = n17380 | n17762 ;
  assign n17764 = n7734 ^ n1738 ^ 1'b0 ;
  assign n17765 = n6255 | n17764 ;
  assign n17766 = n1374 & n1588 ;
  assign n17767 = n5967 & n6822 ;
  assign n17768 = n1246 ^ n942 ^ 1'b0 ;
  assign n17769 = n17767 | n17768 ;
  assign n17770 = ~n3423 & n6921 ;
  assign n17771 = n17769 & n17770 ;
  assign n17772 = n17771 ^ n17704 ^ 1'b0 ;
  assign n17773 = n16088 ^ n1173 ^ 1'b0 ;
  assign n17774 = ~n13083 & n17773 ;
  assign n17775 = ~n1789 & n9748 ;
  assign n17776 = n17775 ^ n1212 ^ 1'b0 ;
  assign n17777 = n13846 & n17776 ;
  assign n17778 = n6058 & n13466 ;
  assign n17779 = n9648 | n17778 ;
  assign n17780 = n17779 ^ n1728 ^ 1'b0 ;
  assign n17781 = n2469 & n6265 ;
  assign n17782 = ( n4616 & ~n4982 ) | ( n4616 & n17781 ) | ( ~n4982 & n17781 ) ;
  assign n17783 = ( n1728 & n13621 ) | ( n1728 & ~n16824 ) | ( n13621 & ~n16824 ) ;
  assign n17784 = ( n1602 & n2104 ) | ( n1602 & n9575 ) | ( n2104 & n9575 ) ;
  assign n17785 = n3191 | n17784 ;
  assign n17786 = n17785 ^ x103 ^ 1'b0 ;
  assign n17787 = x106 & ~n292 ;
  assign n17788 = n5050 & ~n6220 ;
  assign n17789 = n17788 ^ n1593 ^ 1'b0 ;
  assign n17790 = n8430 | n17789 ;
  assign n17792 = n6356 ^ n5286 ^ 1'b0 ;
  assign n17791 = n1850 & ~n17205 ;
  assign n17793 = n17792 ^ n17791 ^ n7287 ;
  assign n17794 = n16539 | n17793 ;
  assign n17795 = ( ~n17787 & n17790 ) | ( ~n17787 & n17794 ) | ( n17790 & n17794 ) ;
  assign n17796 = ( n4792 & ~n7658 ) | ( n4792 & n8712 ) | ( ~n7658 & n8712 ) ;
  assign n17797 = n3817 & n17796 ;
  assign n17798 = n6319 | n9554 ;
  assign n17799 = n17798 ^ n14011 ^ 1'b0 ;
  assign n17800 = ~n8839 & n17799 ;
  assign n17801 = n6552 | n8113 ;
  assign n17802 = n17801 ^ n279 ^ 1'b0 ;
  assign n17803 = n1779 ^ n1629 ^ n1162 ;
  assign n17804 = n17803 ^ n9310 ^ 1'b0 ;
  assign n17805 = ~n6098 & n17804 ;
  assign n17806 = ~n4174 & n7780 ;
  assign n17807 = n17806 ^ n9688 ^ 1'b0 ;
  assign n17808 = n17311 | n17807 ;
  assign n17809 = n17805 | n17808 ;
  assign n17810 = ~n5092 & n13120 ;
  assign n17811 = ( n5284 & n5844 ) | ( n5284 & n7487 ) | ( n5844 & n7487 ) ;
  assign n17812 = n17811 ^ n3847 ^ 1'b0 ;
  assign n17813 = n5228 & ~n13040 ;
  assign n17814 = n17813 ^ n15644 ^ 1'b0 ;
  assign n17815 = n1314 | n8243 ;
  assign n17817 = n1157 & n7323 ;
  assign n17818 = n17817 ^ n16021 ^ 1'b0 ;
  assign n17816 = ~n1538 & n5322 ;
  assign n17819 = n17818 ^ n17816 ^ n10776 ;
  assign n17820 = n17819 ^ n697 ^ 1'b0 ;
  assign n17821 = ~n17815 & n17820 ;
  assign n17824 = n2247 & n10693 ;
  assign n17822 = ( n4914 & ~n6433 ) | ( n4914 & n8663 ) | ( ~n6433 & n8663 ) ;
  assign n17823 = n17822 ^ n12343 ^ 1'b0 ;
  assign n17825 = n17824 ^ n17823 ^ 1'b0 ;
  assign n17826 = n518 & n684 ;
  assign n17827 = ~n17792 & n17826 ;
  assign n17828 = ( n8874 & n13677 ) | ( n8874 & n17827 ) | ( n13677 & n17827 ) ;
  assign n17829 = n10713 ^ n593 ^ 1'b0 ;
  assign n17830 = n11651 & ~n17829 ;
  assign n17831 = n12112 & ~n17830 ;
  assign n17832 = n4809 ^ n2251 ^ n2193 ;
  assign n17833 = n11964 & n17832 ;
  assign n17834 = ~n7763 & n17833 ;
  assign n17835 = n13568 ^ n4485 ^ 1'b0 ;
  assign n17836 = n8009 ^ n5328 ^ n1126 ;
  assign n17837 = n17836 ^ n12713 ^ n2184 ;
  assign n17838 = n2242 & ~n17837 ;
  assign n17839 = n17838 ^ n11860 ^ 1'b0 ;
  assign n17840 = ~n14585 & n16612 ;
  assign n17841 = n1739 & n16622 ;
  assign n17842 = ~n2404 & n17841 ;
  assign n17843 = x2 | n12311 ;
  assign n17844 = ~n2999 & n17843 ;
  assign n17845 = n6640 | n17811 ;
  assign n17846 = n10255 | n17845 ;
  assign n17847 = n14106 & ~n15144 ;
  assign n17848 = n17847 ^ n11897 ^ 1'b0 ;
  assign n17849 = ~n1965 & n16011 ;
  assign n17851 = ( n2609 & n6126 ) | ( n2609 & n10271 ) | ( n6126 & n10271 ) ;
  assign n17852 = n17851 ^ n7697 ^ n5952 ;
  assign n17850 = n523 | n8378 ;
  assign n17853 = n17852 ^ n17850 ^ n6874 ;
  assign n17854 = n6428 | n8949 ;
  assign n17855 = n5623 | n17854 ;
  assign n17856 = n9921 ^ n6620 ^ 1'b0 ;
  assign n17857 = n13349 ^ n970 ^ 1'b0 ;
  assign n17858 = n5899 & ~n17857 ;
  assign n17859 = ~n6329 & n11862 ;
  assign n17860 = n17859 ^ n5824 ^ 1'b0 ;
  assign n17861 = ( ~n148 & n3660 ) | ( ~n148 & n6550 ) | ( n3660 & n6550 ) ;
  assign n17862 = n17861 ^ n11699 ^ 1'b0 ;
  assign n17863 = n12467 | n17862 ;
  assign n17864 = n3942 & ~n17863 ;
  assign n17865 = n17864 ^ n17278 ^ 1'b0 ;
  assign n17866 = ~n3850 & n8601 ;
  assign n17867 = n1491 & n17866 ;
  assign n17868 = n10643 ^ n8936 ^ n5110 ;
  assign n17871 = n812 | n6317 ;
  assign n17872 = n17871 ^ n3915 ^ 1'b0 ;
  assign n17873 = n17872 ^ n3079 ^ 1'b0 ;
  assign n17869 = n9456 ^ n2182 ^ 1'b0 ;
  assign n17870 = ( n2919 & n5929 ) | ( n2919 & n17869 ) | ( n5929 & n17869 ) ;
  assign n17874 = n17873 ^ n17870 ^ 1'b0 ;
  assign n17875 = ( n4160 & n4252 ) | ( n4160 & ~n9247 ) | ( n4252 & ~n9247 ) ;
  assign n17876 = n2586 & ~n14368 ;
  assign n17877 = n17876 ^ n2573 ^ 1'b0 ;
  assign n17878 = n2796 & n17877 ;
  assign n17879 = n17875 & ~n17878 ;
  assign n17880 = ~n5357 & n17879 ;
  assign n17881 = n1622 | n15965 ;
  assign n17882 = n152 & ~n17881 ;
  assign n17883 = n12870 ^ n8487 ^ 1'b0 ;
  assign n17884 = ~n17882 & n17883 ;
  assign n17885 = ( x87 & ~n14891 ) | ( x87 & n17875 ) | ( ~n14891 & n17875 ) ;
  assign n17886 = n3146 | n5389 ;
  assign n17887 = n3974 | n17886 ;
  assign n17888 = n3581 & ~n17887 ;
  assign n17889 = ( n1450 & ~n4959 ) | ( n1450 & n17888 ) | ( ~n4959 & n17888 ) ;
  assign n17890 = ~n2907 & n3040 ;
  assign n17891 = ( n8545 & n15809 ) | ( n8545 & ~n17890 ) | ( n15809 & ~n17890 ) ;
  assign n17892 = n17891 ^ n12537 ^ 1'b0 ;
  assign n17893 = n201 | n17892 ;
  assign n17894 = ( n1402 & n6924 ) | ( n1402 & n16480 ) | ( n6924 & n16480 ) ;
  assign n17895 = n16004 ^ n3852 ^ 1'b0 ;
  assign n17896 = n17894 & n17895 ;
  assign n17897 = ~n17893 & n17896 ;
  assign n17898 = ~n14559 & n17897 ;
  assign n17899 = ~x47 & n11368 ;
  assign n17900 = n3999 ^ n2599 ^ n986 ;
  assign n17901 = ( n2310 & n11763 ) | ( n2310 & n17900 ) | ( n11763 & n17900 ) ;
  assign n17902 = n17901 ^ n1532 ^ 1'b0 ;
  assign n17903 = n12785 & n14008 ;
  assign n17904 = n1185 & n17903 ;
  assign n17905 = n17904 ^ n12328 ^ n8028 ;
  assign n17906 = n13433 ^ n12316 ^ n3926 ;
  assign n17907 = n13478 ^ n12768 ^ n710 ;
  assign n17908 = n11868 & n12497 ;
  assign n17909 = ( n10681 & ~n12412 ) | ( n10681 & n17908 ) | ( ~n12412 & n17908 ) ;
  assign n17910 = n11256 & n17909 ;
  assign n17911 = ~n1485 & n17039 ;
  assign n17912 = n17911 ^ n15989 ^ 1'b0 ;
  assign n17913 = n10646 & n13477 ;
  assign n17914 = n8353 & n17913 ;
  assign n17915 = n13097 ^ n5955 ^ 1'b0 ;
  assign n17916 = n17915 ^ n2502 ^ n950 ;
  assign n17917 = n15622 ^ n7308 ^ n2064 ;
  assign n17918 = ( n5076 & n7059 ) | ( n5076 & n8859 ) | ( n7059 & n8859 ) ;
  assign n17919 = n17918 ^ n456 ^ 1'b0 ;
  assign n17920 = n5753 ^ n5394 ^ 1'b0 ;
  assign n17921 = n17920 ^ n7725 ^ n6675 ;
  assign n17922 = n6166 | n12626 ;
  assign n17923 = n17922 ^ n6724 ^ 1'b0 ;
  assign n17924 = n17554 ^ n14538 ^ n6855 ;
  assign n17925 = ( n798 & n5374 ) | ( n798 & ~n7349 ) | ( n5374 & ~n7349 ) ;
  assign n17926 = n7760 ^ n793 ^ 1'b0 ;
  assign n17927 = n17926 ^ n8598 ^ 1'b0 ;
  assign n17928 = ~n4399 & n17927 ;
  assign n17929 = n758 | n8864 ;
  assign n17930 = n17929 ^ n12905 ^ 1'b0 ;
  assign n17931 = ~n9135 & n17811 ;
  assign n17932 = n12635 ^ n3002 ^ 1'b0 ;
  assign n17933 = n2018 & ~n17932 ;
  assign n17936 = ~n7140 & n11306 ;
  assign n17934 = n5616 & ~n9223 ;
  assign n17935 = n11879 & n17934 ;
  assign n17937 = n17936 ^ n17935 ^ n3060 ;
  assign n17938 = ( n4331 & ~n6515 ) | ( n4331 & n12024 ) | ( ~n6515 & n12024 ) ;
  assign n17942 = n2877 | n3376 ;
  assign n17943 = n7364 | n17942 ;
  assign n17944 = n2563 ^ n1419 ^ 1'b0 ;
  assign n17945 = n17943 & n17944 ;
  assign n17939 = n1985 ^ n292 ^ 1'b0 ;
  assign n17940 = n17939 ^ n7411 ^ 1'b0 ;
  assign n17941 = n1231 & n17940 ;
  assign n17946 = n17945 ^ n17941 ^ n1135 ;
  assign n17947 = n9228 ^ n2806 ^ 1'b0 ;
  assign n17948 = ( n17938 & n17946 ) | ( n17938 & ~n17947 ) | ( n17946 & ~n17947 ) ;
  assign n17949 = n2526 & ~n15224 ;
  assign n17950 = n17949 ^ n14780 ^ n14042 ;
  assign n17951 = n9212 ^ n4419 ^ 1'b0 ;
  assign n17952 = ~n12437 & n12626 ;
  assign n17953 = n2653 | n17952 ;
  assign n17954 = n14112 & n17953 ;
  assign n17955 = ~n1716 & n17954 ;
  assign n17956 = n17955 ^ n1907 ^ 1'b0 ;
  assign n17957 = ( n2706 & ~n6022 ) | ( n2706 & n15229 ) | ( ~n6022 & n15229 ) ;
  assign n17958 = ~n4048 & n17957 ;
  assign n17959 = n1287 & n17958 ;
  assign n17960 = n4059 | n15356 ;
  assign n17961 = n17960 ^ n7283 ^ 1'b0 ;
  assign n17962 = ~n17959 & n17961 ;
  assign n17963 = n6747 | n10308 ;
  assign n17964 = n893 & ~n3469 ;
  assign n17965 = n17964 ^ n3158 ^ 1'b0 ;
  assign n17966 = n17965 ^ n1995 ^ 1'b0 ;
  assign n17967 = ( n129 & n3869 ) | ( n129 & n16926 ) | ( n3869 & n16926 ) ;
  assign n17968 = n8196 & ~n17967 ;
  assign n17969 = n17449 & n17968 ;
  assign n17970 = n11655 | n17969 ;
  assign n17971 = n16674 | n17970 ;
  assign n17972 = ( n4170 & n13514 ) | ( n4170 & n16466 ) | ( n13514 & n16466 ) ;
  assign n17973 = n17972 ^ n694 ^ 1'b0 ;
  assign n17974 = n17971 & ~n17973 ;
  assign n17975 = n14759 ^ n5596 ^ 1'b0 ;
  assign n17976 = ~n12757 & n17975 ;
  assign n17977 = n13473 ^ n11430 ^ n4016 ;
  assign n17978 = n8199 & ~n17977 ;
  assign n17979 = n3376 & ~n5445 ;
  assign n17980 = n3995 | n16757 ;
  assign n17981 = n958 | n17980 ;
  assign n17982 = n17981 ^ n3976 ^ 1'b0 ;
  assign n17983 = n17982 ^ n12188 ^ n3022 ;
  assign n17987 = n7603 ^ x30 ^ 1'b0 ;
  assign n17988 = n17900 & ~n17987 ;
  assign n17984 = ~n260 & n1199 ;
  assign n17985 = n15321 ^ n5347 ^ n4182 ;
  assign n17986 = ( n11842 & n17984 ) | ( n11842 & n17985 ) | ( n17984 & n17985 ) ;
  assign n17989 = n17988 ^ n17986 ^ 1'b0 ;
  assign n17990 = n9573 ^ n701 ^ 1'b0 ;
  assign n17991 = n10756 & n17990 ;
  assign n17992 = ~n2662 & n17991 ;
  assign n17993 = n381 & ~n17992 ;
  assign n17994 = ~n10280 & n17993 ;
  assign n17995 = ~n1663 & n13713 ;
  assign n17996 = n6812 & ~n17995 ;
  assign n17997 = n17996 ^ n8730 ^ 1'b0 ;
  assign n17998 = ~n4166 & n11806 ;
  assign n17999 = n9169 ^ n6245 ^ 1'b0 ;
  assign n18000 = n6743 ^ n1858 ^ 1'b0 ;
  assign n18001 = n17999 | n18000 ;
  assign n18002 = ( n6903 & n8004 ) | ( n6903 & n10214 ) | ( n8004 & n10214 ) ;
  assign n18003 = ~n13584 & n18002 ;
  assign n18004 = n18003 ^ n13291 ^ 1'b0 ;
  assign n18005 = n8856 & ~n18004 ;
  assign n18006 = n5364 & n18005 ;
  assign n18007 = n18006 ^ n12316 ^ n10824 ;
  assign n18008 = n10537 | n16884 ;
  assign n18009 = n18008 ^ n3507 ^ n1895 ;
  assign n18019 = ( n2731 & n6778 ) | ( n2731 & n8100 ) | ( n6778 & n8100 ) ;
  assign n18020 = n18019 ^ n9303 ^ n6700 ;
  assign n18021 = ( n4115 & n11198 ) | ( n4115 & ~n18020 ) | ( n11198 & ~n18020 ) ;
  assign n18015 = x80 & ~n10066 ;
  assign n18010 = n6616 ^ n6388 ^ 1'b0 ;
  assign n18011 = n2419 | n18010 ;
  assign n18012 = ~n514 & n18011 ;
  assign n18013 = n8466 & n14620 ;
  assign n18014 = ~n18012 & n18013 ;
  assign n18016 = n18015 ^ n18014 ^ 1'b0 ;
  assign n18017 = n5725 & n18016 ;
  assign n18018 = n18017 ^ n3252 ^ 1'b0 ;
  assign n18022 = n18021 ^ n18018 ^ 1'b0 ;
  assign n18023 = n4176 & n18022 ;
  assign n18024 = n3863 ^ n2942 ^ 1'b0 ;
  assign n18025 = n6838 & n17924 ;
  assign n18026 = n14037 & n18025 ;
  assign n18027 = n18024 & ~n18026 ;
  assign n18028 = n9603 & n18027 ;
  assign n18029 = n13873 ^ n650 ^ 1'b0 ;
  assign n18030 = n16267 ^ n13742 ^ 1'b0 ;
  assign n18031 = ~n16185 & n16599 ;
  assign n18032 = n17412 | n18031 ;
  assign n18033 = n9775 ^ n7518 ^ 1'b0 ;
  assign n18034 = n18033 ^ n13060 ^ n787 ;
  assign n18036 = ~n11046 & n12621 ;
  assign n18037 = ~x47 & n18036 ;
  assign n18038 = ( n1768 & n9099 ) | ( n1768 & ~n18037 ) | ( n9099 & ~n18037 ) ;
  assign n18035 = ~n2737 & n5966 ;
  assign n18039 = n18038 ^ n18035 ^ 1'b0 ;
  assign n18040 = n6275 & n12782 ;
  assign n18041 = n1677 & ~n2752 ;
  assign n18042 = n18041 ^ n8348 ^ n4957 ;
  assign n18043 = n18040 & n18042 ;
  assign n18044 = n18043 ^ n16262 ^ 1'b0 ;
  assign n18045 = n3337 | n18044 ;
  assign n18046 = ~n5332 & n16207 ;
  assign n18047 = n5880 & n8788 ;
  assign n18048 = n14907 & n18047 ;
  assign n18049 = n5874 & ~n8728 ;
  assign n18050 = n10903 ^ n5931 ^ n2420 ;
  assign n18051 = n3563 & ~n16790 ;
  assign n18052 = n7005 & ~n18051 ;
  assign n18053 = n2459 & n18052 ;
  assign n18054 = ( n13959 & ~n18050 ) | ( n13959 & n18053 ) | ( ~n18050 & n18053 ) ;
  assign n18055 = n4104 & ~n18054 ;
  assign n18056 = n18049 & n18055 ;
  assign n18057 = n2774 & n4862 ;
  assign n18058 = n1373 & n7212 ;
  assign n18059 = ( ~n3172 & n18057 ) | ( ~n3172 & n18058 ) | ( n18057 & n18058 ) ;
  assign n18060 = ~n7408 & n9683 ;
  assign n18061 = n18060 ^ n4326 ^ n1691 ;
  assign n18062 = ( n3168 & n4037 ) | ( n3168 & n16489 ) | ( n4037 & n16489 ) ;
  assign n18064 = n1739 ^ n1539 ^ 1'b0 ;
  assign n18065 = ~x78 & n8431 ;
  assign n18066 = n6374 & ~n12523 ;
  assign n18067 = n18065 & n18066 ;
  assign n18068 = ( n2874 & n18064 ) | ( n2874 & n18067 ) | ( n18064 & n18067 ) ;
  assign n18063 = n7682 | n11158 ;
  assign n18069 = n18068 ^ n18063 ^ 1'b0 ;
  assign n18070 = ~n12519 & n14466 ;
  assign n18071 = n13436 ^ n2365 ^ 1'b0 ;
  assign n18072 = n1200 & n1893 ;
  assign n18073 = ( n10343 & n13127 ) | ( n10343 & n18072 ) | ( n13127 & n18072 ) ;
  assign n18074 = ( ~n313 & n786 ) | ( ~n313 & n3423 ) | ( n786 & n3423 ) ;
  assign n18075 = n18074 ^ n14279 ^ 1'b0 ;
  assign n18076 = n15056 ^ n2553 ^ 1'b0 ;
  assign n18077 = n6591 & ~n15396 ;
  assign n18078 = ~n855 & n18077 ;
  assign n18079 = n18078 ^ n6408 ^ 1'b0 ;
  assign n18080 = n5285 & n18079 ;
  assign n18081 = n18080 ^ n17337 ^ 1'b0 ;
  assign n18082 = n10086 & ~n17182 ;
  assign n18083 = n18082 ^ n14474 ^ 1'b0 ;
  assign n18084 = n4424 ^ n1743 ^ 1'b0 ;
  assign n18085 = n18084 ^ n4753 ^ 1'b0 ;
  assign n18086 = n1498 & ~n18085 ;
  assign n18087 = n18086 ^ n15007 ^ 1'b0 ;
  assign n18088 = n3714 & ~n18087 ;
  assign n18089 = n18088 ^ n10214 ^ 1'b0 ;
  assign n18090 = n6505 | n9393 ;
  assign n18091 = n18090 ^ n12185 ^ n3574 ;
  assign n18092 = n6527 ^ n2138 ^ 1'b0 ;
  assign n18093 = n18091 & ~n18092 ;
  assign n18097 = n7494 | n16539 ;
  assign n18098 = n18097 ^ n9820 ^ 1'b0 ;
  assign n18094 = ( ~n3651 & n5499 ) | ( ~n3651 & n13059 ) | ( n5499 & n13059 ) ;
  assign n18095 = n5794 | n18094 ;
  assign n18096 = n18095 ^ n12043 ^ 1'b0 ;
  assign n18099 = n18098 ^ n18096 ^ n6929 ;
  assign n18100 = ( n7036 & n7158 ) | ( n7036 & ~n10737 ) | ( n7158 & ~n10737 ) ;
  assign n18101 = n16948 | n18100 ;
  assign n18102 = n12306 & n17480 ;
  assign n18103 = n18102 ^ n17282 ^ 1'b0 ;
  assign n18104 = n1221 | n16445 ;
  assign n18105 = ( ~n1546 & n3806 ) | ( ~n1546 & n8718 ) | ( n3806 & n8718 ) ;
  assign n18106 = n11813 ^ n8350 ^ 1'b0 ;
  assign n18107 = n6163 | n14416 ;
  assign n18108 = ~n4043 & n18107 ;
  assign n18109 = ( n4921 & n13094 ) | ( n4921 & n18108 ) | ( n13094 & n18108 ) ;
  assign n18110 = n17432 ^ n139 ^ 1'b0 ;
  assign n18111 = n8223 & ~n18110 ;
  assign n18112 = n4111 & n18111 ;
  assign n18113 = n726 & n18112 ;
  assign n18114 = n18113 ^ n7360 ^ 1'b0 ;
  assign n18115 = ( n341 & n4058 ) | ( n341 & n4722 ) | ( n4058 & n4722 ) ;
  assign n18116 = n18115 ^ n5527 ^ 1'b0 ;
  assign n18117 = n5954 & ~n16650 ;
  assign n18118 = n2200 & n4197 ;
  assign n18119 = n9137 ^ n8064 ^ 1'b0 ;
  assign n18120 = ~n18118 & n18119 ;
  assign n18121 = n14424 & n18120 ;
  assign n18122 = n6571 ^ n5721 ^ 1'b0 ;
  assign n18123 = n9412 | n18122 ;
  assign n18124 = n14934 ^ n8958 ^ 1'b0 ;
  assign n18125 = n18124 ^ n14105 ^ 1'b0 ;
  assign n18126 = n18125 ^ n10822 ^ n2592 ;
  assign n18128 = n14571 & ~n17324 ;
  assign n18127 = n3776 & n7546 ;
  assign n18129 = n18128 ^ n18127 ^ n13615 ;
  assign n18130 = n14055 ^ n3679 ^ 1'b0 ;
  assign n18131 = n12235 ^ n7351 ^ 1'b0 ;
  assign n18132 = n1160 & n18131 ;
  assign n18133 = n7438 ^ n2531 ^ 1'b0 ;
  assign n18134 = n697 & ~n7110 ;
  assign n18135 = n18134 ^ n2111 ^ 1'b0 ;
  assign n18136 = n18135 ^ n7632 ^ 1'b0 ;
  assign n18137 = n15262 ^ n6164 ^ x60 ;
  assign n18138 = n14413 ^ n10394 ^ n7310 ;
  assign n18139 = n18138 ^ n16048 ^ n726 ;
  assign n18140 = n2079 & n17231 ;
  assign n18141 = ~n3621 & n4580 ;
  assign n18142 = n18141 ^ n12704 ^ 1'b0 ;
  assign n18143 = n9868 ^ n7669 ^ 1'b0 ;
  assign n18144 = n13851 ^ n9150 ^ x118 ;
  assign n18145 = n1441 ^ n429 ^ 1'b0 ;
  assign n18146 = ~n6942 & n18145 ;
  assign n18147 = ~n11576 & n18146 ;
  assign n18148 = n18147 ^ n9059 ^ 1'b0 ;
  assign n18149 = ( n134 & n2397 ) | ( n134 & ~n3525 ) | ( n2397 & ~n3525 ) ;
  assign n18150 = n18149 ^ n7116 ^ n3323 ;
  assign n18151 = n15027 ^ n4863 ^ n3831 ;
  assign n18152 = n7900 & ~n18151 ;
  assign n18153 = n6665 & n11694 ;
  assign n18154 = n15144 ^ n1316 ^ 1'b0 ;
  assign n18155 = ~n18153 & n18154 ;
  assign n18156 = ~n4118 & n7699 ;
  assign n18157 = n15686 & n18156 ;
  assign n18158 = x100 & n18157 ;
  assign n18159 = ~n1352 & n17108 ;
  assign n18160 = n18159 ^ n6955 ^ 1'b0 ;
  assign n18161 = n13073 ^ n12146 ^ 1'b0 ;
  assign n18162 = n4900 & n12686 ;
  assign n18163 = n1761 & n18162 ;
  assign n18164 = n12545 | n18163 ;
  assign n18165 = n18161 | n18164 ;
  assign n18166 = ~n1992 & n2593 ;
  assign n18167 = ~n4726 & n8092 ;
  assign n18168 = ( n4864 & n18166 ) | ( n4864 & n18167 ) | ( n18166 & n18167 ) ;
  assign n18169 = n10800 ^ n8573 ^ n5988 ;
  assign n18170 = n3925 | n11292 ;
  assign n18171 = n6685 | n18170 ;
  assign n18172 = n7624 & ~n12246 ;
  assign n18173 = n18172 ^ x38 ^ 1'b0 ;
  assign n18174 = n2172 & n12885 ;
  assign n18177 = n14086 ^ n13112 ^ 1'b0 ;
  assign n18175 = n9066 ^ n1867 ^ 1'b0 ;
  assign n18176 = n10908 & ~n18175 ;
  assign n18178 = n18177 ^ n18176 ^ n2072 ;
  assign n18179 = n5937 | n12585 ;
  assign n18180 = ~n6041 & n10284 ;
  assign n18181 = ~n15992 & n18180 ;
  assign n18182 = n5417 ^ n3096 ^ 1'b0 ;
  assign n18183 = ( n3063 & n11725 ) | ( n3063 & n13771 ) | ( n11725 & n13771 ) ;
  assign n18184 = n8721 ^ n7938 ^ n7864 ;
  assign n18185 = n18184 ^ n13436 ^ 1'b0 ;
  assign n18186 = n13594 & ~n18185 ;
  assign n18187 = n15016 ^ n11538 ^ n3083 ;
  assign n18188 = n4483 & n18187 ;
  assign n18189 = ~n10992 & n18188 ;
  assign n18190 = ( n2687 & ~n8761 ) | ( n2687 & n10769 ) | ( ~n8761 & n10769 ) ;
  assign n18191 = ( n6586 & n8767 ) | ( n6586 & ~n16131 ) | ( n8767 & ~n16131 ) ;
  assign n18192 = n17380 ^ n4797 ^ 1'b0 ;
  assign n18193 = n3783 & n18192 ;
  assign n18197 = n9441 & n12012 ;
  assign n18198 = n5793 ^ n3787 ^ 1'b0 ;
  assign n18199 = ( n2182 & n18197 ) | ( n2182 & ~n18198 ) | ( n18197 & ~n18198 ) ;
  assign n18196 = ~n3954 & n13060 ;
  assign n18194 = n7440 | n12326 ;
  assign n18195 = n6203 | n18194 ;
  assign n18200 = n18199 ^ n18196 ^ n18195 ;
  assign n18201 = n2237 | n10323 ;
  assign n18202 = n18201 ^ n9000 ^ n6136 ;
  assign n18203 = ~n13361 & n18202 ;
  assign n18204 = n1532 | n18203 ;
  assign n18205 = n18204 ^ n3174 ^ 1'b0 ;
  assign n18206 = n1878 ^ n1419 ^ 1'b0 ;
  assign n18207 = ( n6254 & n6610 ) | ( n6254 & n18206 ) | ( n6610 & n18206 ) ;
  assign n18208 = n18207 ^ n12685 ^ n6316 ;
  assign n18209 = ~n10225 & n18208 ;
  assign n18210 = n18209 ^ n4414 ^ 1'b0 ;
  assign n18211 = n17007 ^ n2665 ^ n1899 ;
  assign n18220 = ~n8648 & n16929 ;
  assign n18217 = ~n4986 & n6070 ;
  assign n18218 = ~n5878 & n18217 ;
  assign n18219 = ( ~n212 & n6228 ) | ( ~n212 & n18218 ) | ( n6228 & n18218 ) ;
  assign n18212 = n3999 ^ n2547 ^ 1'b0 ;
  assign n18213 = ( n3677 & ~n14667 ) | ( n3677 & n18212 ) | ( ~n14667 & n18212 ) ;
  assign n18214 = ~n6313 & n18213 ;
  assign n18215 = ~n10605 & n18214 ;
  assign n18216 = ( n13466 & ~n17523 ) | ( n13466 & n18215 ) | ( ~n17523 & n18215 ) ;
  assign n18221 = n18220 ^ n18219 ^ n18216 ;
  assign n18222 = ~n18211 & n18221 ;
  assign n18223 = n18222 ^ n8313 ^ 1'b0 ;
  assign n18224 = n17811 ^ n5659 ^ 1'b0 ;
  assign n18225 = n17445 | n18224 ;
  assign n18226 = ( n2174 & n3187 ) | ( n2174 & n10843 ) | ( n3187 & n10843 ) ;
  assign n18227 = n1167 | n9480 ;
  assign n18228 = n18227 ^ n3928 ^ n637 ;
  assign n18229 = n8565 | n18228 ;
  assign n18230 = n18229 ^ n9894 ^ 1'b0 ;
  assign n18231 = ~n573 & n18230 ;
  assign n18232 = ~n5043 & n18231 ;
  assign n18233 = n145 & n4523 ;
  assign n18234 = n4841 ^ n2000 ^ 1'b0 ;
  assign n18235 = ~n5104 & n18234 ;
  assign n18236 = ~n18233 & n18235 ;
  assign n18237 = ~n1639 & n18236 ;
  assign n18238 = ~n477 & n18237 ;
  assign n18239 = ( n4922 & ~n13244 ) | ( n4922 & n18238 ) | ( ~n13244 & n18238 ) ;
  assign n18240 = ~n1621 & n3277 ;
  assign n18241 = x53 & ~n18240 ;
  assign n18242 = n18241 ^ n11256 ^ 1'b0 ;
  assign n18243 = ( n3469 & n14210 ) | ( n3469 & n18242 ) | ( n14210 & n18242 ) ;
  assign n18244 = n6498 & ~n14403 ;
  assign n18245 = n18244 ^ n11821 ^ 1'b0 ;
  assign n18246 = ( ~n6084 & n6121 ) | ( ~n6084 & n10698 ) | ( n6121 & n10698 ) ;
  assign n18247 = n13497 & n18246 ;
  assign n18248 = ~n18245 & n18247 ;
  assign n18250 = n15529 ^ n9445 ^ n6872 ;
  assign n18249 = n8973 & n11406 ;
  assign n18251 = n18250 ^ n18249 ^ n17949 ;
  assign n18252 = n15168 ^ n1862 ^ n862 ;
  assign n18253 = n4601 ^ n2095 ^ n874 ;
  assign n18254 = n18253 ^ n11982 ^ 1'b0 ;
  assign n18255 = n3513 & n11594 ;
  assign n18256 = n1565 & n8682 ;
  assign n18257 = ~n17035 & n18256 ;
  assign n18258 = ~n4367 & n9924 ;
  assign n18259 = n9199 ^ n1758 ^ 1'b0 ;
  assign n18260 = n2450 & ~n18259 ;
  assign n18261 = n18260 ^ n11751 ^ n10611 ;
  assign n18262 = n5929 & ~n6939 ;
  assign n18263 = n10387 ^ n8837 ^ 1'b0 ;
  assign n18264 = n15060 & n18263 ;
  assign n18265 = ( n10068 & n18262 ) | ( n10068 & n18264 ) | ( n18262 & n18264 ) ;
  assign n18266 = n3386 & ~n15542 ;
  assign n18267 = ( ~n740 & n9284 ) | ( ~n740 & n9894 ) | ( n9284 & n9894 ) ;
  assign n18268 = n212 & n18253 ;
  assign n18269 = n18268 ^ n7398 ^ 1'b0 ;
  assign n18270 = n18269 ^ n334 ^ 1'b0 ;
  assign n18271 = n3362 & ~n17020 ;
  assign n18272 = n6243 & n18271 ;
  assign n18273 = ( n1061 & n2568 ) | ( n1061 & n5726 ) | ( n2568 & n5726 ) ;
  assign n18274 = n10315 | n18273 ;
  assign n18275 = n286 | n18274 ;
  assign n18276 = n5584 & n5783 ;
  assign n18277 = ~n844 & n1690 ;
  assign n18278 = n18277 ^ n7966 ^ 1'b0 ;
  assign n18279 = n6852 | n8332 ;
  assign n18280 = n9505 ^ n5089 ^ 1'b0 ;
  assign n18281 = n3824 & n18280 ;
  assign n18282 = n12494 ^ n8017 ^ 1'b0 ;
  assign n18283 = n2546 & n18282 ;
  assign n18284 = n15725 ^ n8140 ^ 1'b0 ;
  assign n18285 = ( n6333 & n18283 ) | ( n6333 & n18284 ) | ( n18283 & n18284 ) ;
  assign n18286 = ( n5475 & ~n6333 ) | ( n5475 & n8711 ) | ( ~n6333 & n8711 ) ;
  assign n18287 = n18286 ^ n17741 ^ n15496 ;
  assign n18288 = n15777 ^ n8232 ^ n5037 ;
  assign n18289 = n1152 | n3395 ;
  assign n18290 = n18289 ^ n8783 ^ n7045 ;
  assign n18291 = ~n2863 & n18290 ;
  assign n18292 = n13469 ^ n2177 ^ 1'b0 ;
  assign n18293 = ~n18291 & n18292 ;
  assign n18294 = n419 & n9857 ;
  assign n18295 = n18294 ^ n9441 ^ 1'b0 ;
  assign n18296 = ( n2395 & n9345 ) | ( n2395 & n18295 ) | ( n9345 & n18295 ) ;
  assign n18297 = n12452 & n18296 ;
  assign n18298 = ( n3546 & n6299 ) | ( n3546 & n7727 ) | ( n6299 & n7727 ) ;
  assign n18299 = ( n9221 & n9837 ) | ( n9221 & ~n18298 ) | ( n9837 & ~n18298 ) ;
  assign n18300 = n2280 & ~n15000 ;
  assign n18301 = n18300 ^ n2875 ^ 1'b0 ;
  assign n18302 = n14172 & ~n17177 ;
  assign n18303 = n4181 & n18302 ;
  assign n18304 = n3525 ^ n2641 ^ 1'b0 ;
  assign n18305 = n4338 & ~n18304 ;
  assign n18306 = n9199 & ~n18305 ;
  assign n18307 = n6962 & n12264 ;
  assign n18308 = n12087 & ~n14788 ;
  assign n18309 = ( n9233 & ~n18307 ) | ( n9233 & n18308 ) | ( ~n18307 & n18308 ) ;
  assign n18310 = n6433 ^ n4173 ^ n4156 ;
  assign n18311 = n18310 ^ n10116 ^ 1'b0 ;
  assign n18312 = n7769 ^ n1740 ^ n1683 ;
  assign n18313 = n18312 ^ n8523 ^ 1'b0 ;
  assign n18314 = n9203 & ~n18313 ;
  assign n18315 = n8818 & ~n9920 ;
  assign n18316 = ~n11916 & n18315 ;
  assign n18317 = ~n4051 & n5419 ;
  assign n18318 = n6281 & n18317 ;
  assign n18319 = n4885 | n14201 ;
  assign n18320 = n4184 | n6826 ;
  assign n18321 = ~n4723 & n7038 ;
  assign n18322 = n18321 ^ n15547 ^ n3252 ;
  assign n18323 = n18322 ^ n14195 ^ 1'b0 ;
  assign n18324 = n15689 & n18323 ;
  assign n18325 = ~n18320 & n18324 ;
  assign n18326 = n18325 ^ n12618 ^ 1'b0 ;
  assign n18327 = n3011 & ~n7914 ;
  assign n18328 = ~n2099 & n9096 ;
  assign n18329 = n8839 & ~n18328 ;
  assign n18330 = n11813 & ~n18329 ;
  assign n18331 = n14370 ^ n9068 ^ n7197 ;
  assign n18332 = ( n2415 & n10057 ) | ( n2415 & ~n18331 ) | ( n10057 & ~n18331 ) ;
  assign n18333 = n13699 ^ n5683 ^ 1'b0 ;
  assign n18334 = n18333 ^ n3035 ^ 1'b0 ;
  assign n18335 = n10002 ^ n6376 ^ 1'b0 ;
  assign n18336 = n1031 & n15619 ;
  assign n18337 = n8249 | n10698 ;
  assign n18338 = n9291 & ~n18337 ;
  assign n18339 = n18338 ^ n15845 ^ 1'b0 ;
  assign n18340 = ( n8294 & n9524 ) | ( n8294 & n18339 ) | ( n9524 & n18339 ) ;
  assign n18341 = n6446 ^ n736 ^ 1'b0 ;
  assign n18342 = n15805 ^ n12882 ^ 1'b0 ;
  assign n18343 = n18341 & n18342 ;
  assign n18344 = n18343 ^ n8286 ^ n679 ;
  assign n18345 = ( n1736 & n9533 ) | ( n1736 & n17179 ) | ( n9533 & n17179 ) ;
  assign n18346 = n3027 | n18345 ;
  assign n18347 = n18346 ^ n13446 ^ 1'b0 ;
  assign n18348 = ~n4774 & n5960 ;
  assign n18349 = n14294 ^ n12866 ^ 1'b0 ;
  assign n18350 = n927 | n18349 ;
  assign n18351 = n4803 ^ n2242 ^ 1'b0 ;
  assign n18352 = ~n7166 & n18351 ;
  assign n18353 = n7672 | n10680 ;
  assign n18354 = n18353 ^ n974 ^ 1'b0 ;
  assign n18355 = n12361 | n18354 ;
  assign n18356 = n15001 ^ n6737 ^ n5043 ;
  assign n18357 = n11967 & ~n13869 ;
  assign n18358 = n2048 & n7966 ;
  assign n18359 = n6138 & n18358 ;
  assign n18360 = ~n4994 & n18359 ;
  assign n18361 = n15642 ^ n4837 ^ 1'b0 ;
  assign n18362 = ~n2046 & n3059 ;
  assign n18363 = ( n1431 & n6603 ) | ( n1431 & ~n12513 ) | ( n6603 & ~n12513 ) ;
  assign n18364 = ( n6028 & n15159 ) | ( n6028 & n18363 ) | ( n15159 & n18363 ) ;
  assign n18365 = ( ~n18361 & n18362 ) | ( ~n18361 & n18364 ) | ( n18362 & n18364 ) ;
  assign n18366 = n4806 ^ n3337 ^ 1'b0 ;
  assign n18367 = n11460 & ~n18366 ;
  assign n18368 = ~n9728 & n18367 ;
  assign n18369 = ~n3695 & n18368 ;
  assign n18370 = n18369 ^ n3136 ^ 1'b0 ;
  assign n18371 = n15599 ^ n12858 ^ 1'b0 ;
  assign n18372 = n18370 & n18371 ;
  assign n18373 = n10757 ^ n9755 ^ 1'b0 ;
  assign n18374 = n14135 ^ n8072 ^ 1'b0 ;
  assign n18375 = n4867 | n18374 ;
  assign n18376 = n850 & ~n3400 ;
  assign n18377 = n2961 & n9013 ;
  assign n18378 = n9709 | n18377 ;
  assign n18379 = n18378 ^ n616 ^ 1'b0 ;
  assign n18380 = ~n11349 & n18379 ;
  assign n18381 = n18376 & ~n18380 ;
  assign n18382 = ( n7934 & ~n16412 ) | ( n7934 & n18381 ) | ( ~n16412 & n18381 ) ;
  assign n18383 = n10170 ^ n2602 ^ 1'b0 ;
  assign n18384 = n18383 ^ n7184 ^ 1'b0 ;
  assign n18385 = n12421 & n18384 ;
  assign n18386 = n10018 ^ n4646 ^ 1'b0 ;
  assign n18387 = n13380 & n18386 ;
  assign n18388 = n4426 ^ n390 ^ 1'b0 ;
  assign n18389 = n950 ^ n795 ^ 1'b0 ;
  assign n18390 = n8442 & n11909 ;
  assign n18391 = n1065 | n18390 ;
  assign n18392 = n18389 | n18391 ;
  assign n18393 = n10961 | n16490 ;
  assign n18394 = n10446 ^ n2158 ^ 1'b0 ;
  assign n18395 = n6732 | n12092 ;
  assign n18396 = n16738 & ~n18395 ;
  assign n18397 = n5879 & ~n13913 ;
  assign n18398 = n11007 ^ n7938 ^ n7701 ;
  assign n18399 = n18398 ^ n13819 ^ n3807 ;
  assign n18400 = ~n906 & n3042 ;
  assign n18401 = n2637 | n18400 ;
  assign n18402 = ~n6669 & n9566 ;
  assign n18403 = n18402 ^ n3749 ^ 1'b0 ;
  assign n18404 = n18403 ^ n2340 ^ 1'b0 ;
  assign n18405 = n10873 & ~n18404 ;
  assign n18406 = n2801 | n18405 ;
  assign n18407 = n2831 ^ n1937 ^ 1'b0 ;
  assign n18408 = n1996 & n8395 ;
  assign n18409 = n4951 | n18408 ;
  assign n18410 = n2051 | n5385 ;
  assign n18411 = n18410 ^ n8960 ^ 1'b0 ;
  assign n18412 = n1175 | n12818 ;
  assign n18413 = n18412 ^ n13700 ^ 1'b0 ;
  assign n18414 = n6255 | n8138 ;
  assign n18415 = n9482 & ~n18414 ;
  assign n18416 = n4090 & n7953 ;
  assign n18417 = ~n1444 & n18416 ;
  assign n18418 = n13691 ^ n4909 ^ 1'b0 ;
  assign n18419 = n17353 ^ n10299 ^ n4593 ;
  assign n18420 = n9202 & n15674 ;
  assign n18421 = ( n13502 & n18419 ) | ( n13502 & n18420 ) | ( n18419 & n18420 ) ;
  assign n18422 = ~n1430 & n13460 ;
  assign n18423 = ( n593 & n8688 ) | ( n593 & ~n12559 ) | ( n8688 & ~n12559 ) ;
  assign n18424 = n18423 ^ n7021 ^ n1297 ;
  assign n18425 = n18422 & ~n18424 ;
  assign n18426 = n3699 | n4491 ;
  assign n18427 = n9678 & ~n18426 ;
  assign n18428 = n2573 | n18427 ;
  assign n18429 = n1782 | n18428 ;
  assign n18430 = ( ~n2413 & n7417 ) | ( ~n2413 & n18429 ) | ( n7417 & n18429 ) ;
  assign n18431 = ( ~n4662 & n18425 ) | ( ~n4662 & n18430 ) | ( n18425 & n18430 ) ;
  assign n18432 = ( n211 & n3300 ) | ( n211 & ~n8487 ) | ( n3300 & ~n8487 ) ;
  assign n18433 = n1682 | n12168 ;
  assign n18434 = n18432 | n18433 ;
  assign n18435 = n18434 ^ n7632 ^ 1'b0 ;
  assign n18436 = n4333 | n6872 ;
  assign n18437 = n4657 | n10398 ;
  assign n18438 = n18436 & n18437 ;
  assign n18439 = n18438 ^ n7258 ^ 1'b0 ;
  assign n18440 = n13673 ^ n6919 ^ n4603 ;
  assign n18441 = ( n2868 & ~n15365 ) | ( n2868 & n17120 ) | ( ~n15365 & n17120 ) ;
  assign n18442 = n16131 | n17544 ;
  assign n18443 = n6996 | n13054 ;
  assign n18444 = n6206 | n18443 ;
  assign n18445 = n6092 ^ n3610 ^ n3442 ;
  assign n18446 = n18444 | n18445 ;
  assign n18447 = n1280 & n8395 ;
  assign n18448 = n9546 | n13423 ;
  assign n18449 = n18448 ^ n14934 ^ 1'b0 ;
  assign n18450 = n969 & ~n8793 ;
  assign n18451 = n17394 & ~n18450 ;
  assign n18452 = n5278 & n16274 ;
  assign n18453 = n18452 ^ n3240 ^ 1'b0 ;
  assign n18454 = n1569 & n18453 ;
  assign n18455 = n9240 & n10474 ;
  assign n18456 = n18455 ^ n7511 ^ 1'b0 ;
  assign n18457 = n13767 ^ n4110 ^ n3474 ;
  assign n18458 = n18457 ^ n620 ^ 1'b0 ;
  assign n18459 = n2992 & n18458 ;
  assign n18460 = n9174 & ~n15739 ;
  assign n18461 = ~n9649 & n18460 ;
  assign n18462 = ~n2180 & n4572 ;
  assign n18463 = n18461 & n18462 ;
  assign n18464 = n10164 ^ n242 ^ 1'b0 ;
  assign n18465 = n5641 | n13627 ;
  assign n18466 = n5641 & ~n18465 ;
  assign n18467 = n18466 ^ n8376 ^ n4800 ;
  assign n18468 = ~n9199 & n15699 ;
  assign n18469 = n8311 ^ n6928 ^ n1441 ;
  assign n18470 = ~n3858 & n6994 ;
  assign n18471 = n18469 & n18470 ;
  assign n18473 = n2200 | n3752 ;
  assign n18474 = n18473 ^ n4805 ^ 1'b0 ;
  assign n18475 = n18474 ^ n16362 ^ 1'b0 ;
  assign n18472 = n1114 & n1450 ;
  assign n18476 = n18475 ^ n18472 ^ 1'b0 ;
  assign n18477 = n6118 & n18394 ;
  assign n18478 = n11770 & n18477 ;
  assign n18479 = ( ~n3456 & n3869 ) | ( ~n3456 & n5425 ) | ( n3869 & n5425 ) ;
  assign n18480 = n249 & n4854 ;
  assign n18481 = ~n4707 & n18480 ;
  assign n18482 = n18479 & ~n18481 ;
  assign n18483 = n17269 & n17661 ;
  assign n18484 = n6828 ^ n421 ^ 1'b0 ;
  assign n18485 = n18484 ^ n5654 ^ 1'b0 ;
  assign n18486 = n5176 | n18485 ;
  assign n18487 = n11127 | n17142 ;
  assign n18488 = n2919 | n18487 ;
  assign n18489 = n15505 ^ n2207 ^ 1'b0 ;
  assign n18490 = n15012 | n18489 ;
  assign n18491 = n811 & ~n15092 ;
  assign n18492 = ~n1522 & n18491 ;
  assign n18493 = ( n8644 & ~n9812 ) | ( n8644 & n18492 ) | ( ~n9812 & n18492 ) ;
  assign n18494 = n18493 ^ n13525 ^ 1'b0 ;
  assign n18495 = n18490 | n18494 ;
  assign n18496 = n13750 ^ n11161 ^ n9372 ;
  assign n18497 = ~n8551 & n18048 ;
  assign n18498 = n712 & ~n15752 ;
  assign n18499 = n11045 ^ n7193 ^ n1710 ;
  assign n18500 = ~n10790 & n18099 ;
  assign n18501 = ~n10941 & n18500 ;
  assign n18502 = ~n11384 & n14316 ;
  assign n18503 = n18502 ^ n1678 ^ 1'b0 ;
  assign n18504 = n701 & n18503 ;
  assign n18506 = n3615 & n6810 ;
  assign n18507 = n18506 ^ n3751 ^ 1'b0 ;
  assign n18505 = n3108 | n7128 ;
  assign n18508 = n18507 ^ n18505 ^ 1'b0 ;
  assign n18512 = n1545 & ~n13412 ;
  assign n18509 = n670 & n1493 ;
  assign n18510 = ~n8525 & n18509 ;
  assign n18511 = n18510 ^ n3930 ^ 1'b0 ;
  assign n18513 = n18512 ^ n18511 ^ n6247 ;
  assign n18514 = n18513 ^ n14085 ^ 1'b0 ;
  assign n18515 = ( n3945 & n8565 ) | ( n3945 & ~n18419 ) | ( n8565 & ~n18419 ) ;
  assign n18516 = ( n3042 & n4414 ) | ( n3042 & ~n14176 ) | ( n4414 & ~n14176 ) ;
  assign n18517 = n15496 ^ n14201 ^ n734 ;
  assign n18520 = n7214 & ~n9323 ;
  assign n18521 = n1712 & n18520 ;
  assign n18518 = n15396 ^ n6537 ^ n5469 ;
  assign n18519 = ( n8922 & n12428 ) | ( n8922 & ~n18518 ) | ( n12428 & ~n18518 ) ;
  assign n18522 = n18521 ^ n18519 ^ 1'b0 ;
  assign n18524 = n5329 & n6226 ;
  assign n18523 = n10072 & ~n18481 ;
  assign n18525 = n18524 ^ n18523 ^ 1'b0 ;
  assign n18526 = n490 & n2077 ;
  assign n18527 = ( n494 & n8762 ) | ( n494 & ~n18526 ) | ( n8762 & ~n18526 ) ;
  assign n18528 = n18527 ^ n13226 ^ n5933 ;
  assign n18529 = ~n2502 & n6681 ;
  assign n18530 = n11923 ^ n8014 ^ n5526 ;
  assign n18531 = n18530 ^ n17048 ^ n2113 ;
  assign n18532 = n11336 & ~n18531 ;
  assign n18533 = n16091 & n18532 ;
  assign n18534 = n838 & ~n8565 ;
  assign n18535 = n2122 & ~n13724 ;
  assign n18536 = n18535 ^ n3722 ^ 1'b0 ;
  assign n18537 = ( ~n5613 & n18534 ) | ( ~n5613 & n18536 ) | ( n18534 & n18536 ) ;
  assign n18541 = n4580 ^ n1664 ^ 1'b0 ;
  assign n18542 = n14387 | n18541 ;
  assign n18538 = n10223 ^ n8869 ^ n4294 ;
  assign n18539 = n9155 | n18538 ;
  assign n18540 = n18539 ^ n11549 ^ 1'b0 ;
  assign n18543 = n18542 ^ n18540 ^ 1'b0 ;
  assign n18544 = n1760 | n2635 ;
  assign n18545 = n18544 ^ n7760 ^ n1150 ;
  assign n18546 = n3780 ^ n3699 ^ n2888 ;
  assign n18547 = n18546 ^ n11908 ^ n5784 ;
  assign n18548 = n14392 ^ n3316 ^ 1'b0 ;
  assign n18549 = ~n8150 & n18548 ;
  assign n18550 = n18549 ^ n1390 ^ 1'b0 ;
  assign n18551 = n12372 ^ n1619 ^ 1'b0 ;
  assign n18552 = n7481 | n18551 ;
  assign n18553 = n3070 | n18552 ;
  assign n18554 = n17830 ^ n12283 ^ 1'b0 ;
  assign n18555 = n13881 ^ n10848 ^ n4792 ;
  assign n18556 = ~n1614 & n13141 ;
  assign n18557 = n9064 ^ n1571 ^ 1'b0 ;
  assign n18558 = n15877 ^ n7888 ^ 1'b0 ;
  assign n18559 = n5876 ^ n5737 ^ 1'b0 ;
  assign n18560 = n1014 | n18559 ;
  assign n18561 = ~n14095 & n18560 ;
  assign n18562 = n18561 ^ n10340 ^ n4292 ;
  assign n18563 = n10760 & n16817 ;
  assign n18564 = n18563 ^ n6764 ^ 1'b0 ;
  assign n18565 = n2771 ^ n951 ^ 1'b0 ;
  assign n18566 = n2758 | n18565 ;
  assign n18567 = n169 & n18566 ;
  assign n18568 = ~n1139 & n14097 ;
  assign n18569 = n13541 & n18568 ;
  assign n18570 = n17730 ^ n599 ^ 1'b0 ;
  assign n18571 = n18569 | n18570 ;
  assign n18572 = ~n1890 & n6047 ;
  assign n18573 = n7564 & ~n13339 ;
  assign n18574 = n18573 ^ n2250 ^ 1'b0 ;
  assign n18575 = ( n5116 & n8759 ) | ( n5116 & n8839 ) | ( n8759 & n8839 ) ;
  assign n18576 = ( n4407 & n6820 ) | ( n4407 & n18575 ) | ( n6820 & n18575 ) ;
  assign n18577 = n18576 ^ n13793 ^ n1205 ;
  assign n18578 = n13690 ^ n4712 ^ n2117 ;
  assign n18579 = ~n229 & n4756 ;
  assign n18580 = ~n11442 & n18579 ;
  assign n18581 = n8276 & n18580 ;
  assign n18582 = n18206 & ~n18581 ;
  assign n18583 = n14595 ^ n566 ^ 1'b0 ;
  assign n18584 = n18583 ^ n4507 ^ n368 ;
  assign n18585 = n4717 & ~n11731 ;
  assign n18586 = n18585 ^ n857 ^ 1'b0 ;
  assign n18587 = n1307 | n18586 ;
  assign n18588 = ~n3027 & n5011 ;
  assign n18589 = ( ~n8229 & n13366 ) | ( ~n8229 & n18588 ) | ( n13366 & n18588 ) ;
  assign n18590 = n10005 ^ n5789 ^ 1'b0 ;
  assign n18591 = n12931 ^ n4964 ^ 1'b0 ;
  assign n18592 = n12771 ^ n5368 ^ 1'b0 ;
  assign n18593 = ( n1761 & ~n13085 ) | ( n1761 & n18592 ) | ( ~n13085 & n18592 ) ;
  assign n18594 = n13712 | n16814 ;
  assign n18595 = n18593 & ~n18594 ;
  assign n18596 = n13620 ^ n3388 ^ 1'b0 ;
  assign n18597 = n2085 & n2769 ;
  assign n18598 = n18597 ^ n14571 ^ 1'b0 ;
  assign n18599 = n18598 ^ n11160 ^ n2368 ;
  assign n18600 = n5904 & n11857 ;
  assign n18601 = n18600 ^ n13163 ^ n1940 ;
  assign n18602 = ~n6701 & n12171 ;
  assign n18603 = n15206 | n18602 ;
  assign n18604 = n8991 ^ n7973 ^ n6715 ;
  assign n18605 = ~n1230 & n18604 ;
  assign n18606 = n13014 & n18605 ;
  assign n18607 = n9786 ^ n523 ^ 1'b0 ;
  assign n18608 = ( n1472 & n9445 ) | ( n1472 & n18604 ) | ( n9445 & n18604 ) ;
  assign n18609 = n4618 | n18608 ;
  assign n18610 = ~n5746 & n12124 ;
  assign n18611 = ~n1410 & n2684 ;
  assign n18612 = n18611 ^ n2428 ^ 1'b0 ;
  assign n18613 = ( ~n3677 & n4863 ) | ( ~n3677 & n18612 ) | ( n4863 & n18612 ) ;
  assign n18614 = n18613 ^ n872 ^ 1'b0 ;
  assign n18615 = n3827 ^ n1747 ^ n665 ;
  assign n18616 = n10460 ^ n10335 ^ 1'b0 ;
  assign n18617 = n1478 & ~n7391 ;
  assign n18618 = ~n8143 & n11826 ;
  assign n18619 = ( n965 & ~n11219 ) | ( n965 & n18618 ) | ( ~n11219 & n18618 ) ;
  assign n18620 = ~n4061 & n18619 ;
  assign n18621 = n18620 ^ n10400 ^ 1'b0 ;
  assign n18623 = n9184 ^ n7236 ^ n4261 ;
  assign n18624 = ~x28 & n18623 ;
  assign n18622 = ~n6779 & n9345 ;
  assign n18625 = n18624 ^ n18622 ^ n17771 ;
  assign n18626 = n18625 ^ n2104 ^ 1'b0 ;
  assign n18627 = n18626 ^ n7361 ^ 1'b0 ;
  assign n18628 = n2231 | n3771 ;
  assign n18629 = n18628 ^ n13087 ^ n3323 ;
  assign n18630 = n3672 & ~n6986 ;
  assign n18631 = n15019 ^ n12749 ^ 1'b0 ;
  assign n18632 = ( n8787 & n10343 ) | ( n8787 & ~n15308 ) | ( n10343 & ~n15308 ) ;
  assign n18633 = ( n2497 & ~n4341 ) | ( n2497 & n9949 ) | ( ~n4341 & n9949 ) ;
  assign n18634 = n7176 & ~n8012 ;
  assign n18635 = ( ~n15496 & n18633 ) | ( ~n15496 & n18634 ) | ( n18633 & n18634 ) ;
  assign n18636 = n2889 ^ n1043 ^ 1'b0 ;
  assign n18637 = ~n4653 & n13336 ;
  assign n18638 = n18637 ^ n17380 ^ 1'b0 ;
  assign n18639 = n6513 | n16874 ;
  assign n18640 = n17128 | n18639 ;
  assign n18641 = ~n1133 & n4501 ;
  assign n18642 = ~x84 & n18641 ;
  assign n18643 = n1745 & n1892 ;
  assign n18644 = n18643 ^ n10885 ^ 1'b0 ;
  assign n18645 = n18644 ^ n17914 ^ 1'b0 ;
  assign n18646 = ~n3649 & n15857 ;
  assign n18647 = n6641 ^ n5228 ^ n4462 ;
  assign n18648 = n12948 & ~n16220 ;
  assign n18649 = n18648 ^ n5552 ^ 1'b0 ;
  assign n18650 = n18649 ^ n18167 ^ 1'b0 ;
  assign n18651 = n3252 & ~n18650 ;
  assign n18652 = n18651 ^ n17257 ^ n1123 ;
  assign n18653 = n5033 & ~n17183 ;
  assign n18654 = ~n16227 & n18653 ;
  assign n18655 = n14768 ^ n9844 ^ n3173 ;
  assign n18659 = ( n6764 & n7573 ) | ( n6764 & n8742 ) | ( n7573 & n8742 ) ;
  assign n18656 = n13410 ^ n3519 ^ 1'b0 ;
  assign n18657 = ~n14858 & n18656 ;
  assign n18658 = n18657 ^ n6166 ^ 1'b0 ;
  assign n18660 = n18659 ^ n18658 ^ 1'b0 ;
  assign n18661 = n18655 | n18660 ;
  assign n18662 = n1900 | n4142 ;
  assign n18663 = ~n2217 & n13886 ;
  assign n18664 = n18662 & n18663 ;
  assign n18665 = n9632 ^ n6991 ^ n3384 ;
  assign n18666 = n15614 ^ n6199 ^ 1'b0 ;
  assign n18667 = n11071 ^ n5223 ^ 1'b0 ;
  assign n18668 = n13389 & n18667 ;
  assign n18669 = n6269 & ~n9412 ;
  assign n18670 = ~n11329 & n15819 ;
  assign n18671 = ~n1921 & n18670 ;
  assign n18672 = n3659 | n8412 ;
  assign n18673 = n5657 | n16053 ;
  assign n18674 = n18673 ^ n5653 ^ 1'b0 ;
  assign n18676 = n14461 ^ n11148 ^ n3012 ;
  assign n18677 = n3056 & n18676 ;
  assign n18675 = x122 & ~n10209 ;
  assign n18678 = n18677 ^ n18675 ^ 1'b0 ;
  assign n18679 = ~n5098 & n11352 ;
  assign n18680 = ~n4519 & n18679 ;
  assign n18681 = n15026 & ~n18680 ;
  assign n18682 = n474 & ~n4925 ;
  assign n18683 = n2855 & ~n6321 ;
  assign n18684 = n5537 & n18683 ;
  assign n18685 = ( n2549 & ~n4013 ) | ( n2549 & n18684 ) | ( ~n4013 & n18684 ) ;
  assign n18686 = n6136 ^ n3260 ^ 1'b0 ;
  assign n18687 = n15028 ^ n3693 ^ 1'b0 ;
  assign n18688 = ( ~n4102 & n12191 ) | ( ~n4102 & n17700 ) | ( n12191 & n17700 ) ;
  assign n18689 = n18688 ^ n2315 ^ n1447 ;
  assign n18690 = n18689 ^ n4102 ^ 1'b0 ;
  assign n18691 = ~n1768 & n5038 ;
  assign n18692 = ~n13142 & n18691 ;
  assign n18693 = ~n2768 & n18692 ;
  assign n18694 = n6148 ^ n4417 ^ 1'b0 ;
  assign n18695 = ~n8785 & n18694 ;
  assign n18696 = n2566 & n12647 ;
  assign n18697 = n8437 ^ n7910 ^ 1'b0 ;
  assign n18698 = n453 & ~n18697 ;
  assign n18699 = n4566 | n18698 ;
  assign n18700 = n18699 ^ n3224 ^ 1'b0 ;
  assign n18701 = n10142 & ~n18700 ;
  assign n18702 = n8668 ^ n3147 ^ n808 ;
  assign n18704 = n15977 ^ n9087 ^ n6214 ;
  assign n18703 = n7861 & n9858 ;
  assign n18705 = n18704 ^ n18703 ^ 1'b0 ;
  assign n18706 = n18702 | n18705 ;
  assign n18707 = n11095 ^ n3482 ^ 1'b0 ;
  assign n18708 = n18707 ^ n748 ^ 1'b0 ;
  assign n18709 = n17700 ^ n15566 ^ n10014 ;
  assign n18710 = ( n9190 & ~n18322 ) | ( n9190 & n18709 ) | ( ~n18322 & n18709 ) ;
  assign n18711 = n5539 & ~n7691 ;
  assign n18712 = n18711 ^ n15883 ^ 1'b0 ;
  assign n18713 = n4815 & n11596 ;
  assign n18714 = n18713 ^ n3168 ^ 1'b0 ;
  assign n18715 = n1458 & ~n11868 ;
  assign n18716 = n4199 ^ n2819 ^ 1'b0 ;
  assign n18717 = n17269 & ~n18716 ;
  assign n18720 = n12677 | n14744 ;
  assign n18718 = n201 & n10591 ;
  assign n18719 = n18718 ^ n11834 ^ n7561 ;
  assign n18721 = n18720 ^ n18719 ^ 1'b0 ;
  assign n18722 = ~n4593 & n5031 ;
  assign n18723 = n7627 & ~n14051 ;
  assign n18724 = n18723 ^ n9794 ^ 1'b0 ;
  assign n18725 = n7099 ^ n5987 ^ n5689 ;
  assign n18726 = ~n14737 & n15013 ;
  assign n18727 = n18725 & n18726 ;
  assign n18734 = n8488 ^ n5698 ^ 1'b0 ;
  assign n18735 = n16868 & ~n18734 ;
  assign n18728 = ~n1123 & n4167 ;
  assign n18729 = n18728 ^ n639 ^ 1'b0 ;
  assign n18730 = n298 & ~n18729 ;
  assign n18731 = n5483 ^ n1449 ^ n866 ;
  assign n18732 = n18731 ^ n14208 ^ 1'b0 ;
  assign n18733 = n18730 & n18732 ;
  assign n18736 = n18735 ^ n18733 ^ 1'b0 ;
  assign n18737 = ( n191 & n423 ) | ( n191 & n609 ) | ( n423 & n609 ) ;
  assign n18738 = n18737 ^ n12052 ^ n2626 ;
  assign n18739 = n11233 & n12161 ;
  assign n18740 = ~n7658 & n7817 ;
  assign n18741 = n15081 & n18740 ;
  assign n18742 = n18741 ^ n4271 ^ 1'b0 ;
  assign n18743 = n18739 & ~n18742 ;
  assign n18744 = n18743 ^ n2552 ^ 1'b0 ;
  assign n18746 = n7689 ^ n1373 ^ 1'b0 ;
  assign n18745 = n5882 | n8290 ;
  assign n18747 = n18746 ^ n18745 ^ 1'b0 ;
  assign n18748 = n5630 | n17236 ;
  assign n18749 = n18748 ^ n8031 ^ 1'b0 ;
  assign n18750 = n7594 ^ n6846 ^ 1'b0 ;
  assign n18752 = ( n859 & n2462 ) | ( n859 & ~n4230 ) | ( n2462 & ~n4230 ) ;
  assign n18753 = n2721 & ~n18752 ;
  assign n18751 = n11707 ^ n11402 ^ n7813 ;
  assign n18754 = n18753 ^ n18751 ^ n2350 ;
  assign n18755 = ~n5425 & n7020 ;
  assign n18756 = n6696 & n18755 ;
  assign n18757 = n18756 ^ n219 ^ 1'b0 ;
  assign n18758 = n14184 ^ n8341 ^ n2134 ;
  assign n18759 = n4294 & n18758 ;
  assign n18760 = n18759 ^ n9941 ^ 1'b0 ;
  assign n18761 = n14045 ^ n7665 ^ 1'b0 ;
  assign n18762 = n14189 ^ n9426 ^ n3191 ;
  assign n18763 = n5895 & ~n18762 ;
  assign n18764 = n3413 & n18763 ;
  assign n18765 = n985 & ~n14858 ;
  assign n18766 = n16600 ^ n13334 ^ n1712 ;
  assign n18767 = ~n14657 & n18766 ;
  assign n18768 = n2976 & n18767 ;
  assign n18769 = n6255 ^ n3792 ^ 1'b0 ;
  assign n18770 = n5116 & n18769 ;
  assign n18771 = n14877 ^ n12062 ^ n2341 ;
  assign n18772 = n18771 ^ n4126 ^ n3704 ;
  assign n18773 = ( n3180 & n18770 ) | ( n3180 & ~n18772 ) | ( n18770 & ~n18772 ) ;
  assign n18774 = n2591 | n16794 ;
  assign n18775 = n18774 ^ n15248 ^ 1'b0 ;
  assign n18776 = n9144 ^ n2296 ^ 1'b0 ;
  assign n18777 = n14503 & n18776 ;
  assign n18778 = n18777 ^ n9058 ^ 1'b0 ;
  assign n18782 = n8709 & n12937 ;
  assign n18783 = n1137 & n18782 ;
  assign n18784 = n18783 ^ n820 ^ 1'b0 ;
  assign n18779 = n10822 ^ n3673 ^ 1'b0 ;
  assign n18780 = n7648 & ~n18779 ;
  assign n18781 = ~n14437 & n18780 ;
  assign n18785 = n18784 ^ n18781 ^ n4147 ;
  assign n18786 = n6605 ^ n6390 ^ 1'b0 ;
  assign n18787 = n5198 | n18786 ;
  assign n18788 = n5225 & n18787 ;
  assign n18789 = n15323 & n18788 ;
  assign n18790 = ~n9547 & n13922 ;
  assign n18791 = n7587 & n17882 ;
  assign n18792 = n7266 & n10827 ;
  assign n18793 = n8429 | n8921 ;
  assign n18794 = n7082 ^ n3303 ^ 1'b0 ;
  assign n18795 = ~n7947 & n18794 ;
  assign n18796 = ~n14418 & n18795 ;
  assign n18797 = n1167 & ~n2121 ;
  assign n18798 = n3530 & n18797 ;
  assign n18799 = n18196 | n18798 ;
  assign n18800 = ( n2458 & n9477 ) | ( n2458 & n9738 ) | ( n9477 & n9738 ) ;
  assign n18801 = ( ~n6934 & n9862 ) | ( ~n6934 & n13929 ) | ( n9862 & n13929 ) ;
  assign n18802 = n8826 ^ n477 ^ 1'b0 ;
  assign n18803 = n6818 & n18802 ;
  assign n18804 = n4709 | n17352 ;
  assign n18806 = ~n4124 & n10558 ;
  assign n18805 = ~n2217 & n17957 ;
  assign n18807 = n18806 ^ n18805 ^ 1'b0 ;
  assign n18808 = n9712 ^ n9242 ^ 1'b0 ;
  assign n18809 = n5759 ^ n4757 ^ 1'b0 ;
  assign n18810 = ~n10224 & n18809 ;
  assign n18811 = n18810 ^ n13406 ^ 1'b0 ;
  assign n18812 = ~n1184 & n18811 ;
  assign n18813 = ( n4233 & n4893 ) | ( n4233 & n16831 ) | ( n4893 & n16831 ) ;
  assign n18814 = n3887 ^ n3065 ^ 1'b0 ;
  assign n18815 = n18814 ^ n15819 ^ n10033 ;
  assign n18816 = n713 ^ n416 ^ 1'b0 ;
  assign n18817 = n9531 | n18816 ;
  assign n18818 = n8773 ^ n6254 ^ n3159 ;
  assign n18819 = n3254 & n17522 ;
  assign n18820 = n18819 ^ n13087 ^ 1'b0 ;
  assign n18821 = n18818 & n18820 ;
  assign n18822 = n1047 & ~n15780 ;
  assign n18823 = n18822 ^ n9390 ^ 1'b0 ;
  assign n18824 = n11101 & ~n17105 ;
  assign n18825 = n18824 ^ n9054 ^ 1'b0 ;
  assign n18827 = n5367 & ~n6186 ;
  assign n18826 = n652 | n868 ;
  assign n18828 = n18827 ^ n18826 ^ 1'b0 ;
  assign n18830 = n14922 ^ n13519 ^ n5406 ;
  assign n18829 = n1803 | n4601 ;
  assign n18831 = n18830 ^ n18829 ^ n4372 ;
  assign n18833 = n5552 ^ n1915 ^ 1'b0 ;
  assign n18832 = n945 | n4875 ;
  assign n18834 = n18833 ^ n18832 ^ 1'b0 ;
  assign n18835 = n1921 ^ n763 ^ 1'b0 ;
  assign n18836 = n6573 ^ n1336 ^ 1'b0 ;
  assign n18838 = n13700 ^ x59 ^ 1'b0 ;
  assign n18837 = n5812 ^ n3224 ^ 1'b0 ;
  assign n18839 = n18838 ^ n18837 ^ n10262 ;
  assign n18840 = n4433 | n15755 ;
  assign n18841 = n18840 ^ n8042 ^ 1'b0 ;
  assign n18842 = n4463 | n18841 ;
  assign n18843 = n11781 | n18842 ;
  assign n18844 = n1674 | n4926 ;
  assign n18845 = n18844 ^ n1124 ^ 1'b0 ;
  assign n18846 = n18845 ^ n5770 ^ n4356 ;
  assign n18847 = n7133 | n9820 ;
  assign n18848 = n18846 & ~n18847 ;
  assign n18849 = x2 | n5475 ;
  assign n18850 = ( n1748 & n2939 ) | ( n1748 & ~n16130 ) | ( n2939 & ~n16130 ) ;
  assign n18851 = n13830 | n18850 ;
  assign n18852 = n12858 & ~n16311 ;
  assign n18853 = n15534 ^ n3272 ^ 1'b0 ;
  assign n18854 = ( n2215 & ~n2395 ) | ( n2215 & n9857 ) | ( ~n2395 & n9857 ) ;
  assign n18855 = n18854 ^ n5257 ^ 1'b0 ;
  assign n18856 = n5438 ^ n1718 ^ n997 ;
  assign n18857 = n5382 & ~n18856 ;
  assign n18858 = n478 & ~n17115 ;
  assign n18859 = n14765 ^ n12771 ^ 1'b0 ;
  assign n18860 = ~n7658 & n8532 ;
  assign n18861 = n18860 ^ n12662 ^ 1'b0 ;
  assign n18862 = n18861 ^ n7832 ^ 1'b0 ;
  assign n18863 = n3651 & n18862 ;
  assign n18864 = n801 | n5348 ;
  assign n18865 = n3522 & ~n18864 ;
  assign n18866 = n18767 & n18865 ;
  assign n18867 = ( n4714 & n13475 ) | ( n4714 & ~n18866 ) | ( n13475 & ~n18866 ) ;
  assign n18868 = n4908 | n8231 ;
  assign n18869 = n2513 & ~n18868 ;
  assign n18870 = n18869 ^ n11989 ^ n2242 ;
  assign n18871 = n12496 ^ n6293 ^ 1'b0 ;
  assign n18872 = n16876 & ~n18871 ;
  assign n18873 = n18872 ^ n5370 ^ 1'b0 ;
  assign n18874 = n8538 ^ n3765 ^ 1'b0 ;
  assign n18875 = ~n1958 & n5948 ;
  assign n18876 = n6730 & n18875 ;
  assign n18877 = n18876 ^ n3920 ^ 1'b0 ;
  assign n18878 = n6585 & ~n18877 ;
  assign n18879 = n9409 ^ n9023 ^ 1'b0 ;
  assign n18880 = n18878 & n18879 ;
  assign n18881 = x47 | n6041 ;
  assign n18882 = n18881 ^ n9467 ^ 1'b0 ;
  assign n18883 = ( n1069 & n17533 ) | ( n1069 & n18882 ) | ( n17533 & n18882 ) ;
  assign n18884 = n3010 | n8562 ;
  assign n18885 = n11958 | n18884 ;
  assign n18886 = n15501 ^ n7481 ^ 1'b0 ;
  assign n18887 = ~n751 & n18886 ;
  assign n18888 = n18887 ^ n1988 ^ 1'b0 ;
  assign n18889 = n10210 ^ n8007 ^ n3132 ;
  assign n18890 = n5706 & n18889 ;
  assign n18891 = n18890 ^ n6537 ^ 1'b0 ;
  assign n18892 = n3159 & ~n10931 ;
  assign n18893 = ~n18891 & n18892 ;
  assign n18894 = n18893 ^ n15209 ^ 1'b0 ;
  assign n18895 = ~n4593 & n18894 ;
  assign n18896 = n10581 & ~n11281 ;
  assign n18897 = n5190 & ~n10024 ;
  assign n18898 = n18897 ^ n4926 ^ 1'b0 ;
  assign n18899 = n7482 & n8078 ;
  assign n18900 = n18899 ^ n2904 ^ 1'b0 ;
  assign n18901 = n18898 & n18900 ;
  assign n18902 = n18901 ^ n2657 ^ 1'b0 ;
  assign n18903 = n13881 ^ n13587 ^ 1'b0 ;
  assign n18904 = n18903 ^ n17945 ^ n916 ;
  assign n18905 = n8503 ^ n1371 ^ 1'b0 ;
  assign n18906 = n456 | n18905 ;
  assign n18907 = n18906 ^ n5284 ^ 1'b0 ;
  assign n18909 = n15133 ^ n11199 ^ n1805 ;
  assign n18908 = n3484 & ~n5885 ;
  assign n18910 = n18909 ^ n18908 ^ 1'b0 ;
  assign n18911 = n1822 & ~n6363 ;
  assign n18912 = ~n2510 & n18911 ;
  assign n18913 = n18903 ^ n6638 ^ 1'b0 ;
  assign n18914 = ~n18912 & n18913 ;
  assign n18915 = n4181 | n11071 ;
  assign n18916 = n18914 | n18915 ;
  assign n18917 = n9770 ^ n6003 ^ 1'b0 ;
  assign n18918 = n8308 ^ n1252 ^ 1'b0 ;
  assign n18919 = x52 & ~n584 ;
  assign n18920 = ( ~n3386 & n8527 ) | ( ~n3386 & n18919 ) | ( n8527 & n18919 ) ;
  assign n18921 = n4432 & ~n18920 ;
  assign n18922 = n17057 ^ n5535 ^ n3238 ;
  assign n18923 = n3159 & ~n9608 ;
  assign n18924 = n9688 ^ n3710 ^ 1'b0 ;
  assign n18925 = n18924 ^ n6361 ^ 1'b0 ;
  assign n18926 = n15869 ^ n5286 ^ 1'b0 ;
  assign n18927 = n13222 | n18926 ;
  assign n18928 = n18925 & ~n18927 ;
  assign n18929 = n18928 ^ n5901 ^ 1'b0 ;
  assign n18930 = n9526 ^ n2890 ^ 1'b0 ;
  assign n18931 = n16685 & n18930 ;
  assign n18932 = n7076 ^ n1576 ^ 1'b0 ;
  assign n18933 = n3512 ^ n2499 ^ 1'b0 ;
  assign n18934 = n18932 | n18933 ;
  assign n18935 = n6135 | n9947 ;
  assign n18936 = n14705 & ~n18935 ;
  assign n18937 = n8190 ^ n3225 ^ 1'b0 ;
  assign n18938 = n11195 & ~n18937 ;
  assign n18939 = ~n12550 & n18938 ;
  assign n18940 = n17982 ^ n6822 ^ n2730 ;
  assign n18944 = n2655 ^ x69 ^ 1'b0 ;
  assign n18945 = n1414 | n18944 ;
  assign n18941 = n7295 ^ n2597 ^ 1'b0 ;
  assign n18942 = n7122 | n18941 ;
  assign n18943 = n8225 | n18942 ;
  assign n18946 = n18945 ^ n18943 ^ 1'b0 ;
  assign n18947 = n4042 & n16712 ;
  assign n18948 = n2954 & ~n7641 ;
  assign n18949 = n18948 ^ n6647 ^ n3240 ;
  assign n18950 = n4431 ^ n1201 ^ 1'b0 ;
  assign n18951 = n18949 & ~n18950 ;
  assign n18952 = n3805 & ~n9538 ;
  assign n18953 = n8123 & ~n18952 ;
  assign n18954 = n18953 ^ n1819 ^ 1'b0 ;
  assign n18955 = n4149 ^ n1721 ^ n1276 ;
  assign n18956 = n3837 & ~n12968 ;
  assign n18957 = ( n1205 & n14012 ) | ( n1205 & ~n18956 ) | ( n14012 & ~n18956 ) ;
  assign n18958 = ( n4482 & ~n4581 ) | ( n4482 & n7775 ) | ( ~n4581 & n7775 ) ;
  assign n18959 = ( n2382 & n10352 ) | ( n2382 & n18958 ) | ( n10352 & n18958 ) ;
  assign n18960 = n6138 ^ n2077 ^ 1'b0 ;
  assign n18961 = n6239 ^ n5935 ^ 1'b0 ;
  assign n18962 = n4704 ^ n1914 ^ 1'b0 ;
  assign n18963 = n18962 ^ n6956 ^ 1'b0 ;
  assign n18964 = n18963 ^ n10914 ^ n4709 ;
  assign n18965 = ( n4681 & n15158 ) | ( n4681 & ~n18964 ) | ( n15158 & ~n18964 ) ;
  assign n18966 = n18961 | n18965 ;
  assign n18968 = n2500 & n5068 ;
  assign n18969 = n18968 ^ n4074 ^ 1'b0 ;
  assign n18967 = n2967 | n16922 ;
  assign n18970 = n18969 ^ n18967 ^ 1'b0 ;
  assign n18971 = n9645 ^ n7537 ^ n2595 ;
  assign n18972 = ~n1704 & n3757 ;
  assign n18973 = n18972 ^ n5694 ^ 1'b0 ;
  assign n18974 = n4882 | n18973 ;
  assign n18975 = n1162 | n2854 ;
  assign n18976 = n15456 ^ n719 ^ n191 ;
  assign n18977 = n18975 | n18976 ;
  assign n18978 = n14064 ^ n13973 ^ 1'b0 ;
  assign n18979 = n10747 | n18978 ;
  assign n18980 = n523 & n3077 ;
  assign n18981 = ~n3134 & n9926 ;
  assign n18982 = n18981 ^ n6515 ^ 1'b0 ;
  assign n18983 = x52 & n3957 ;
  assign n18984 = n1441 & n4321 ;
  assign n18985 = n727 & n18984 ;
  assign n18986 = n18985 ^ n5402 ^ 1'b0 ;
  assign n18987 = n18983 & ~n18986 ;
  assign n18988 = ( n4314 & ~n6007 ) | ( n4314 & n18987 ) | ( ~n6007 & n18987 ) ;
  assign n18989 = n3365 ^ x105 ^ 1'b0 ;
  assign n18990 = n737 & ~n18989 ;
  assign n18991 = n15944 & n18990 ;
  assign n18992 = n18991 ^ n8815 ^ 1'b0 ;
  assign n18993 = x127 & ~n18992 ;
  assign n18994 = n9113 ^ n8130 ^ n5784 ;
  assign n18995 = ( ~n12644 & n18993 ) | ( ~n12644 & n18994 ) | ( n18993 & n18994 ) ;
  assign n18996 = n7595 | n11063 ;
  assign n18997 = n6988 & n10708 ;
  assign n18998 = n18997 ^ n11283 ^ 1'b0 ;
  assign n18999 = n949 & ~n4967 ;
  assign n19000 = n18999 ^ n5355 ^ 1'b0 ;
  assign n19001 = n8853 ^ n8019 ^ n5044 ;
  assign n19002 = ( n12083 & ~n19000 ) | ( n12083 & n19001 ) | ( ~n19000 & n19001 ) ;
  assign n19003 = ~n1805 & n14191 ;
  assign n19004 = n3315 ^ n499 ^ 1'b0 ;
  assign n19005 = n9358 ^ n8299 ^ 1'b0 ;
  assign n19006 = n16981 & ~n18057 ;
  assign n19007 = n19006 ^ n3776 ^ n2484 ;
  assign n19008 = n5525 & n19007 ;
  assign n19009 = ~n19005 & n19008 ;
  assign n19010 = n2004 & n12805 ;
  assign n19011 = n19010 ^ n13933 ^ 1'b0 ;
  assign n19012 = ~n1942 & n2651 ;
  assign n19013 = n19012 ^ n2140 ^ 1'b0 ;
  assign n19014 = n19013 ^ n11430 ^ 1'b0 ;
  assign n19015 = ( n13088 & n15101 ) | ( n13088 & n19014 ) | ( n15101 & n19014 ) ;
  assign n19016 = n14778 ^ n3264 ^ 1'b0 ;
  assign n19018 = ( ~n3811 & n4921 ) | ( ~n3811 & n14189 ) | ( n4921 & n14189 ) ;
  assign n19017 = n8819 ^ n4942 ^ n2328 ;
  assign n19019 = n19018 ^ n19017 ^ 1'b0 ;
  assign n19020 = n12508 ^ n4523 ^ 1'b0 ;
  assign n19021 = ~n1469 & n4833 ;
  assign n19022 = n19021 ^ n18838 ^ n12341 ;
  assign n19023 = n7203 & ~n19022 ;
  assign n19024 = n3856 ^ n2352 ^ 1'b0 ;
  assign n19025 = n19024 ^ n6013 ^ 1'b0 ;
  assign n19026 = x77 & n19025 ;
  assign n19027 = n4889 & n9599 ;
  assign n19028 = n7977 | n8482 ;
  assign n19029 = n1331 & ~n19028 ;
  assign n19030 = n11235 ^ n7581 ^ n3257 ;
  assign n19031 = ( ~n19013 & n19029 ) | ( ~n19013 & n19030 ) | ( n19029 & n19030 ) ;
  assign n19032 = ( x81 & n343 ) | ( x81 & n19031 ) | ( n343 & n19031 ) ;
  assign n19033 = n7518 & ~n19032 ;
  assign n19034 = n5630 | n9714 ;
  assign n19035 = n19034 ^ n18361 ^ 1'b0 ;
  assign n19036 = n795 | n990 ;
  assign n19037 = n4580 ^ n2641 ^ 1'b0 ;
  assign n19038 = n3391 & ~n19037 ;
  assign n19039 = ( n3673 & n7984 ) | ( n3673 & ~n9859 ) | ( n7984 & ~n9859 ) ;
  assign n19040 = n19039 ^ n3634 ^ 1'b0 ;
  assign n19041 = ~n2475 & n19040 ;
  assign n19042 = n17151 ^ n14667 ^ n10217 ;
  assign n19043 = n16104 ^ n6324 ^ n3030 ;
  assign n19044 = n967 | n1373 ;
  assign n19046 = ~n6876 & n12171 ;
  assign n19047 = n3838 & n19046 ;
  assign n19045 = n8129 & ~n15556 ;
  assign n19048 = n19047 ^ n19045 ^ 1'b0 ;
  assign n19049 = n3537 | n6126 ;
  assign n19050 = n19049 ^ n6524 ^ 1'b0 ;
  assign n19051 = n6283 ^ n3964 ^ 1'b0 ;
  assign n19052 = n5005 | n19051 ;
  assign n19053 = ~n6659 & n9215 ;
  assign n19054 = n19053 ^ n8225 ^ n5228 ;
  assign n19055 = n19052 | n19054 ;
  assign n19061 = ~n2371 & n6283 ;
  assign n19057 = n7518 ^ n1393 ^ 1'b0 ;
  assign n19056 = n1236 & ~n4085 ;
  assign n19058 = n19057 ^ n19056 ^ 1'b0 ;
  assign n19059 = n19058 ^ n4489 ^ 1'b0 ;
  assign n19060 = n3202 | n19059 ;
  assign n19062 = n19061 ^ n19060 ^ 1'b0 ;
  assign n19063 = n13743 | n19062 ;
  assign n19064 = n19063 ^ n17656 ^ 1'b0 ;
  assign n19065 = n17708 ^ n6640 ^ n1791 ;
  assign n19066 = n12750 ^ n5423 ^ n2823 ;
  assign n19067 = n2750 ^ n2739 ^ n1709 ;
  assign n19068 = n4043 | n19067 ;
  assign n19069 = n1619 & ~n19068 ;
  assign n19070 = ~n1345 & n4512 ;
  assign n19071 = n6889 & n19070 ;
  assign n19072 = n19071 ^ n10875 ^ 1'b0 ;
  assign n19073 = n13248 & n13432 ;
  assign n19074 = n19073 ^ n3975 ^ 1'b0 ;
  assign n19075 = ~n551 & n7888 ;
  assign n19076 = n2416 ^ n1524 ^ 1'b0 ;
  assign n19077 = n2358 & n19076 ;
  assign n19078 = ~n1251 & n19077 ;
  assign n19079 = n19078 ^ n11421 ^ n7119 ;
  assign n19080 = n6935 | n19079 ;
  assign n19081 = x22 & ~n10601 ;
  assign n19082 = n19081 ^ n8756 ^ 1'b0 ;
  assign n19083 = n857 ^ n467 ^ 1'b0 ;
  assign n19084 = ~n3638 & n19083 ;
  assign n19085 = x77 & n19084 ;
  assign n19086 = n19085 ^ n15467 ^ 1'b0 ;
  assign n19087 = n19086 ^ n9705 ^ n4107 ;
  assign n19088 = ~n905 & n14410 ;
  assign n19089 = n13362 ^ n2597 ^ 1'b0 ;
  assign n19090 = n4607 & n19089 ;
  assign n19091 = n15116 & n19090 ;
  assign n19092 = n19091 ^ n14844 ^ n2282 ;
  assign n19093 = n1351 & ~n9000 ;
  assign n19094 = ~n2678 & n19093 ;
  assign n19095 = n16783 ^ n4897 ^ 1'b0 ;
  assign n19096 = n1046 | n19095 ;
  assign n19097 = n2868 & ~n4238 ;
  assign n19098 = n19097 ^ n16595 ^ 1'b0 ;
  assign n19099 = n2141 ^ x74 ^ 1'b0 ;
  assign n19100 = n4197 & n19099 ;
  assign n19101 = n6668 & ~n10567 ;
  assign n19102 = ~n2774 & n19101 ;
  assign n19103 = ( ~n9190 & n13819 ) | ( ~n9190 & n19102 ) | ( n13819 & n19102 ) ;
  assign n19104 = ~n19100 & n19103 ;
  assign n19105 = ( ~n7266 & n10305 ) | ( ~n7266 & n15403 ) | ( n10305 & n15403 ) ;
  assign n19106 = n5368 & n15944 ;
  assign n19107 = n19106 ^ n10865 ^ 1'b0 ;
  assign n19108 = ~n5493 & n19107 ;
  assign n19109 = ~n11824 & n19108 ;
  assign n19114 = n3091 | n12163 ;
  assign n19110 = n8037 & n9229 ;
  assign n19111 = n19110 ^ n8711 ^ 1'b0 ;
  assign n19112 = ( ~n7707 & n15708 ) | ( ~n7707 & n16288 ) | ( n15708 & n16288 ) ;
  assign n19113 = n19111 & n19112 ;
  assign n19115 = n19114 ^ n19113 ^ 1'b0 ;
  assign n19116 = n14282 & ~n14294 ;
  assign n19117 = n5370 | n15140 ;
  assign n19118 = n10045 | n19117 ;
  assign n19119 = n19118 ^ n4296 ^ 1'b0 ;
  assign n19120 = n17225 | n19119 ;
  assign n19121 = n6676 | n8616 ;
  assign n19122 = n17144 ^ n2854 ^ 1'b0 ;
  assign n19123 = n18361 ^ n15789 ^ 1'b0 ;
  assign n19124 = ( ~n1794 & n2454 ) | ( ~n1794 & n3881 ) | ( n2454 & n3881 ) ;
  assign n19125 = n19124 ^ n7293 ^ n5703 ;
  assign n19126 = n15768 ^ n4316 ^ 1'b0 ;
  assign n19128 = n138 & n9407 ;
  assign n19129 = n19128 ^ n6718 ^ 1'b0 ;
  assign n19127 = n822 | n1129 ;
  assign n19130 = n19129 ^ n19127 ^ 1'b0 ;
  assign n19131 = n3317 ^ n740 ^ 1'b0 ;
  assign n19132 = n15584 & ~n19131 ;
  assign n19133 = n5001 & n19132 ;
  assign n19134 = ( n12351 & n18456 ) | ( n12351 & ~n19133 ) | ( n18456 & ~n19133 ) ;
  assign n19135 = ( n3850 & n4676 ) | ( n3850 & n13401 ) | ( n4676 & n13401 ) ;
  assign n19136 = n8204 & ~n19135 ;
  assign n19137 = n8759 ^ n6641 ^ 1'b0 ;
  assign n19138 = ( ~n6226 & n19136 ) | ( ~n6226 & n19137 ) | ( n19136 & n19137 ) ;
  assign n19139 = ( ~n6884 & n14510 ) | ( ~n6884 & n16935 ) | ( n14510 & n16935 ) ;
  assign n19140 = ~n2261 & n10974 ;
  assign n19141 = n15863 & n19140 ;
  assign n19143 = n9131 ^ n7226 ^ 1'b0 ;
  assign n19144 = ( n2498 & n15734 ) | ( n2498 & n19143 ) | ( n15734 & n19143 ) ;
  assign n19142 = n12875 ^ n3240 ^ 1'b0 ;
  assign n19145 = n19144 ^ n19142 ^ 1'b0 ;
  assign n19146 = n19141 | n19145 ;
  assign n19147 = n16529 ^ n8334 ^ 1'b0 ;
  assign n19148 = ~n19146 & n19147 ;
  assign n19149 = n19148 ^ n8023 ^ 1'b0 ;
  assign n19150 = n4186 ^ n820 ^ 1'b0 ;
  assign n19151 = n8667 & n19150 ;
  assign n19152 = n8513 ^ n2913 ^ n992 ;
  assign n19153 = n19152 ^ n10218 ^ n6991 ;
  assign n19154 = n19151 & n19153 ;
  assign n19155 = n19154 ^ n862 ^ 1'b0 ;
  assign n19156 = ~n3679 & n18267 ;
  assign n19157 = n19156 ^ n12307 ^ 1'b0 ;
  assign n19158 = n14630 & n15250 ;
  assign n19159 = n19158 ^ n9992 ^ 1'b0 ;
  assign n19160 = n10545 ^ n4588 ^ 1'b0 ;
  assign n19164 = n2748 | n10558 ;
  assign n19162 = ~n3373 & n7160 ;
  assign n19161 = n13345 ^ n1362 ^ 1'b0 ;
  assign n19163 = n19162 ^ n19161 ^ n10503 ;
  assign n19165 = n19164 ^ n19163 ^ n10031 ;
  assign n19166 = n18764 ^ n2546 ^ 1'b0 ;
  assign n19167 = n17016 ^ n1502 ^ 1'b0 ;
  assign n19168 = n5317 & ~n19167 ;
  assign n19169 = n2399 & n16105 ;
  assign n19170 = ~n18283 & n19169 ;
  assign n19171 = n2390 | n8445 ;
  assign n19172 = n2705 | n19171 ;
  assign n19173 = n19172 ^ n8746 ^ n2384 ;
  assign n19174 = n2418 & n3677 ;
  assign n19175 = ~n19173 & n19174 ;
  assign n19176 = n13865 ^ n9556 ^ 1'b0 ;
  assign n19177 = n6075 & n19176 ;
  assign n19178 = n19177 ^ n11126 ^ 1'b0 ;
  assign n19179 = ( n1440 & n9869 ) | ( n1440 & n15584 ) | ( n9869 & n15584 ) ;
  assign n19180 = n1000 & ~n9771 ;
  assign n19181 = n19180 ^ n9692 ^ 1'b0 ;
  assign n19182 = n8961 | n19181 ;
  assign n19183 = n6057 ^ n3615 ^ 1'b0 ;
  assign n19185 = ~n3694 & n14815 ;
  assign n19184 = n3095 ^ n1345 ^ 1'b0 ;
  assign n19186 = n19185 ^ n19184 ^ n4271 ;
  assign n19187 = n4104 ^ x123 ^ x92 ;
  assign n19188 = n19187 ^ n462 ^ 1'b0 ;
  assign n19189 = n7385 | n19188 ;
  assign n19190 = n18569 ^ n491 ^ 1'b0 ;
  assign n19191 = n1617 & n19190 ;
  assign n19192 = n5552 ^ n3482 ^ 1'b0 ;
  assign n19193 = n15238 & n19192 ;
  assign n19194 = n19193 ^ n10362 ^ 1'b0 ;
  assign n19195 = n13146 | n19194 ;
  assign n19196 = n13614 ^ n11004 ^ n1445 ;
  assign n19197 = n14410 & ~n19196 ;
  assign n19198 = n14247 & n19197 ;
  assign n19199 = n19198 ^ n6430 ^ 1'b0 ;
  assign n19203 = n11763 ^ n3856 ^ 1'b0 ;
  assign n19204 = n5570 | n19203 ;
  assign n19200 = n8524 ^ n949 ^ 1'b0 ;
  assign n19201 = n19200 ^ n18662 ^ 1'b0 ;
  assign n19202 = n5901 & n19201 ;
  assign n19205 = n19204 ^ n19202 ^ 1'b0 ;
  assign n19206 = n1656 & ~n19205 ;
  assign n19207 = ~n15659 & n17067 ;
  assign n19208 = ~n433 & n19207 ;
  assign n19209 = n12124 & n17243 ;
  assign n19210 = n19209 ^ n10656 ^ 1'b0 ;
  assign n19211 = n11221 ^ n8342 ^ n5525 ;
  assign n19212 = n10168 & ~n19211 ;
  assign n19213 = n19212 ^ n14119 ^ n5817 ;
  assign n19214 = n271 & ~n1034 ;
  assign n19215 = n1436 & ~n7301 ;
  assign n19216 = n19215 ^ n14215 ^ n12251 ;
  assign n19217 = ( ~n1314 & n7047 ) | ( ~n1314 & n15314 ) | ( n7047 & n15314 ) ;
  assign n19218 = ~n827 & n1943 ;
  assign n19219 = n1805 & n7706 ;
  assign n19220 = n19219 ^ n2397 ^ 1'b0 ;
  assign n19221 = n6536 ^ n3412 ^ 1'b0 ;
  assign n19222 = n12729 & ~n15625 ;
  assign n19223 = n19221 & n19222 ;
  assign n19224 = ( ~n7066 & n13841 ) | ( ~n7066 & n17863 ) | ( n13841 & n17863 ) ;
  assign n19225 = ( ~n7798 & n9126 ) | ( ~n7798 & n19224 ) | ( n9126 & n19224 ) ;
  assign n19226 = n6196 | n8826 ;
  assign n19227 = n19226 ^ n15373 ^ n9101 ;
  assign n19228 = n8482 ^ n3421 ^ n611 ;
  assign n19229 = ( n11469 & ~n19227 ) | ( n11469 & n19228 ) | ( ~n19227 & n19228 ) ;
  assign n19230 = n784 | n7292 ;
  assign n19231 = ( ~n4038 & n4834 ) | ( ~n4038 & n7976 ) | ( n4834 & n7976 ) ;
  assign n19232 = n7355 | n10088 ;
  assign n19233 = n19231 | n19232 ;
  assign n19234 = ~n2304 & n7518 ;
  assign n19235 = n4164 & ~n12116 ;
  assign n19236 = ~n19234 & n19235 ;
  assign n19237 = n11562 ^ n5583 ^ n4120 ;
  assign n19238 = n10980 ^ n4699 ^ 1'b0 ;
  assign n19239 = n19238 ^ n4523 ^ n3037 ;
  assign n19240 = n13512 ^ n6810 ^ 1'b0 ;
  assign n19241 = ~n5421 & n19240 ;
  assign n19242 = n1325 | n12470 ;
  assign n19243 = n19242 ^ n219 ^ 1'b0 ;
  assign n19244 = n6598 ^ n3320 ^ 1'b0 ;
  assign n19245 = ~n19243 & n19244 ;
  assign n19246 = ~n1214 & n2197 ;
  assign n19247 = ~n5166 & n19246 ;
  assign n19248 = n7085 & ~n19247 ;
  assign n19249 = n19248 ^ n15824 ^ 1'b0 ;
  assign n19250 = n491 & n8065 ;
  assign n19251 = ( ~n781 & n2828 ) | ( ~n781 & n16556 ) | ( n2828 & n16556 ) ;
  assign n19252 = n19251 ^ n17926 ^ n4778 ;
  assign n19253 = n10164 | n14531 ;
  assign n19254 = n19253 ^ n13582 ^ 1'b0 ;
  assign n19255 = n4246 | n19254 ;
  assign n19256 = n16948 ^ n5201 ^ n4524 ;
  assign n19257 = n7927 & ~n19256 ;
  assign n19258 = n16806 & n19257 ;
  assign n19259 = ( n5252 & n9403 ) | ( n5252 & ~n10840 ) | ( n9403 & ~n10840 ) ;
  assign n19260 = ( n3606 & ~n14820 ) | ( n3606 & n19259 ) | ( ~n14820 & n19259 ) ;
  assign n19261 = ~n19258 & n19260 ;
  assign n19262 = n7391 | n8431 ;
  assign n19263 = n10882 ^ n6962 ^ 1'b0 ;
  assign n19264 = n19262 & n19263 ;
  assign n19265 = n12048 ^ n7545 ^ 1'b0 ;
  assign n19266 = n13796 & n19265 ;
  assign n19267 = n19266 ^ n16908 ^ 1'b0 ;
  assign n19268 = n4221 ^ n905 ^ 1'b0 ;
  assign n19269 = n13821 & ~n19268 ;
  assign n19270 = ( n6055 & ~n9246 ) | ( n6055 & n12046 ) | ( ~n9246 & n12046 ) ;
  assign n19271 = n13477 ^ n5753 ^ 1'b0 ;
  assign n19272 = n17130 | n19271 ;
  assign n19273 = n3626 ^ n2312 ^ 1'b0 ;
  assign n19274 = n2462 | n11249 ;
  assign n19275 = n6814 | n19115 ;
  assign n19276 = n19275 ^ n9699 ^ 1'b0 ;
  assign n19277 = n1354 & n6519 ;
  assign n19278 = n15667 ^ n379 ^ 1'b0 ;
  assign n19279 = n5919 | n19278 ;
  assign n19280 = n18281 ^ n2724 ^ 1'b0 ;
  assign n19281 = ( x110 & n8160 ) | ( x110 & ~n19280 ) | ( n8160 & ~n19280 ) ;
  assign n19282 = n9803 ^ n7554 ^ n6950 ;
  assign n19283 = n10700 | n17653 ;
  assign n19284 = n6057 ^ n3743 ^ 1'b0 ;
  assign n19285 = ~n9729 & n19284 ;
  assign n19286 = ( n7765 & ~n8918 ) | ( n7765 & n14011 ) | ( ~n8918 & n14011 ) ;
  assign n19287 = n1575 & n19286 ;
  assign n19288 = ~n15718 & n19287 ;
  assign n19289 = n3756 & ~n9220 ;
  assign n19290 = ~n1440 & n19289 ;
  assign n19291 = ( n706 & n6428 ) | ( n706 & ~n12813 ) | ( n6428 & ~n12813 ) ;
  assign n19292 = n19291 ^ n11549 ^ n920 ;
  assign n19293 = n1093 & ~n9672 ;
  assign n19294 = n19293 ^ n616 ^ 1'b0 ;
  assign n19295 = n13322 | n19294 ;
  assign n19296 = ~n1603 & n9642 ;
  assign n19297 = n19296 ^ n6126 ^ 1'b0 ;
  assign n19303 = ( n2478 & n7962 ) | ( n2478 & ~n10800 ) | ( n7962 & ~n10800 ) ;
  assign n19304 = n3554 | n19303 ;
  assign n19305 = n19304 ^ n2054 ^ 1'b0 ;
  assign n19301 = n3706 & n3969 ;
  assign n19302 = n19301 ^ n8084 ^ 1'b0 ;
  assign n19306 = n19305 ^ n19302 ^ n2036 ;
  assign n19298 = n1215 | n3638 ;
  assign n19299 = ( x126 & n10640 ) | ( x126 & ~n19298 ) | ( n10640 & ~n19298 ) ;
  assign n19300 = n4091 & n19299 ;
  assign n19307 = n19306 ^ n19300 ^ n18563 ;
  assign n19308 = n12046 ^ n908 ^ 1'b0 ;
  assign n19309 = n11964 & n19308 ;
  assign n19310 = n19309 ^ n2557 ^ 1'b0 ;
  assign n19311 = ~n2299 & n5526 ;
  assign n19312 = n1011 & n19311 ;
  assign n19313 = n12584 & ~n19312 ;
  assign n19314 = n6108 ^ n2530 ^ 1'b0 ;
  assign n19315 = n19313 & ~n19314 ;
  assign n19316 = n19315 ^ n1935 ^ 1'b0 ;
  assign n19318 = n7286 ^ n2512 ^ 1'b0 ;
  assign n19319 = n397 | n19318 ;
  assign n19320 = n4954 | n19319 ;
  assign n19321 = n3728 & ~n19320 ;
  assign n19322 = ( n2679 & n4429 ) | ( n2679 & n19321 ) | ( n4429 & n19321 ) ;
  assign n19317 = n16131 ^ n3911 ^ 1'b0 ;
  assign n19323 = n19322 ^ n19317 ^ 1'b0 ;
  assign n19324 = n6240 ^ n4403 ^ 1'b0 ;
  assign n19325 = n19324 ^ n10287 ^ n5460 ;
  assign n19326 = n14648 ^ n295 ^ 1'b0 ;
  assign n19327 = n19326 ^ n2680 ^ n1485 ;
  assign n19328 = n2542 & ~n4964 ;
  assign n19329 = ~n9462 & n19328 ;
  assign n19330 = n9291 & ~n13627 ;
  assign n19331 = n19330 ^ n770 ^ 1'b0 ;
  assign n19332 = ( ~n15270 & n19329 ) | ( ~n15270 & n19331 ) | ( n19329 & n19331 ) ;
  assign n19333 = n3778 & ~n7717 ;
  assign n19334 = n19333 ^ n18546 ^ 1'b0 ;
  assign n19335 = n4810 & ~n7725 ;
  assign n19336 = n19335 ^ n7695 ^ 1'b0 ;
  assign n19337 = n2201 & ~n8232 ;
  assign n19338 = n19336 & n19337 ;
  assign n19339 = n4005 & n19018 ;
  assign n19340 = ~n12199 & n19339 ;
  assign n19341 = n8353 | n18258 ;
  assign n19342 = ~n9945 & n19305 ;
  assign n19343 = n12153 & n19342 ;
  assign n19344 = n19343 ^ n12508 ^ 1'b0 ;
  assign n19345 = n6087 & ~n19344 ;
  assign n19346 = n19345 ^ x24 ^ 1'b0 ;
  assign n19347 = n18622 & ~n19346 ;
  assign n19348 = n15750 ^ n3228 ^ 1'b0 ;
  assign n19349 = n16139 ^ n13595 ^ 1'b0 ;
  assign n19350 = ( n16293 & n19348 ) | ( n16293 & ~n19349 ) | ( n19348 & ~n19349 ) ;
  assign n19351 = n5977 ^ x105 ^ 1'b0 ;
  assign n19352 = n16612 ^ n4720 ^ 1'b0 ;
  assign n19354 = ( n597 & n10049 ) | ( n597 & ~n11213 ) | ( n10049 & ~n11213 ) ;
  assign n19353 = n12373 & n13629 ;
  assign n19355 = n19354 ^ n19353 ^ 1'b0 ;
  assign n19356 = n182 | n901 ;
  assign n19357 = n19356 ^ n4028 ^ 1'b0 ;
  assign n19358 = ~n2664 & n12366 ;
  assign n19359 = n13119 ^ n6995 ^ 1'b0 ;
  assign n19360 = n15835 ^ n8854 ^ n3821 ;
  assign n19361 = ( ~n3503 & n14326 ) | ( ~n3503 & n19360 ) | ( n14326 & n19360 ) ;
  assign n19362 = n9665 ^ n6852 ^ 1'b0 ;
  assign n19363 = n1073 & n19362 ;
  assign n19364 = n5234 ^ n3318 ^ 1'b0 ;
  assign n19365 = ~n19314 & n19364 ;
  assign n19366 = n3284 & ~n6934 ;
  assign n19367 = n2389 & ~n19366 ;
  assign n19368 = n7998 & ~n18050 ;
  assign n19370 = n11682 ^ n10264 ^ 1'b0 ;
  assign n19371 = n7937 & n19370 ;
  assign n19369 = n1314 | n11079 ;
  assign n19372 = n19371 ^ n19369 ^ 1'b0 ;
  assign n19373 = n19372 ^ n16766 ^ 1'b0 ;
  assign n19374 = n19368 & n19373 ;
  assign n19376 = n5584 ^ n3173 ^ 1'b0 ;
  assign n19375 = n6408 ^ n5080 ^ 1'b0 ;
  assign n19377 = n19376 ^ n19375 ^ n9407 ;
  assign n19378 = ( n6530 & n12908 ) | ( n6530 & n19377 ) | ( n12908 & n19377 ) ;
  assign n19379 = n5226 ^ n3217 ^ 1'b0 ;
  assign n19380 = n946 | n19379 ;
  assign n19381 = n13085 & n17165 ;
  assign n19382 = n19381 ^ n1741 ^ 1'b0 ;
  assign n19383 = ( n142 & n19380 ) | ( n142 & n19382 ) | ( n19380 & n19382 ) ;
  assign n19384 = n10980 ^ n5313 ^ 1'b0 ;
  assign n19385 = n7513 & ~n13705 ;
  assign n19386 = n19385 ^ n5537 ^ n1743 ;
  assign n19387 = n2573 & n8103 ;
  assign n19388 = ~n2224 & n17223 ;
  assign n19389 = ~n6239 & n19388 ;
  assign n19390 = n1499 | n19389 ;
  assign n19391 = n3858 | n19390 ;
  assign n19392 = n19387 & ~n19391 ;
  assign n19393 = n5504 | n19392 ;
  assign n19394 = n3362 | n15734 ;
  assign n19395 = n4263 & n19394 ;
  assign n19396 = n2499 | n19395 ;
  assign n19397 = n13614 ^ n6766 ^ 1'b0 ;
  assign n19419 = n7293 & ~n7570 ;
  assign n19420 = n7570 & n19419 ;
  assign n19416 = n4217 & n13997 ;
  assign n19417 = ~n13997 & n19416 ;
  assign n19418 = n19417 ^ n9969 ^ 1'b0 ;
  assign n19398 = n6271 & ~n14612 ;
  assign n19399 = n14612 & n19398 ;
  assign n19400 = n19399 ^ n16817 ^ 1'b0 ;
  assign n19401 = n2792 | n19400 ;
  assign n19402 = n19401 ^ n10878 ^ 1'b0 ;
  assign n19412 = n2133 | n18932 ;
  assign n19413 = n2133 & ~n19412 ;
  assign n19404 = ~n270 & n5451 ;
  assign n19405 = ~n968 & n19404 ;
  assign n19406 = ( x19 & ~n7752 ) | ( x19 & n12744 ) | ( ~n7752 & n12744 ) ;
  assign n19407 = n4193 & n19406 ;
  assign n19408 = n19407 ^ n15040 ^ 1'b0 ;
  assign n19409 = n19405 | n19408 ;
  assign n19410 = n19409 ^ n1139 ^ 1'b0 ;
  assign n19403 = n15207 ^ n7319 ^ 1'b0 ;
  assign n19411 = n19410 ^ n19403 ^ 1'b0 ;
  assign n19414 = n19413 ^ n19411 ^ 1'b0 ;
  assign n19415 = n19402 & ~n19414 ;
  assign n19421 = n19420 ^ n19418 ^ n19415 ;
  assign n19422 = n19421 ^ n6527 ^ 1'b0 ;
  assign n19423 = n19397 & n19422 ;
  assign n19424 = n13771 ^ n5719 ^ 1'b0 ;
  assign n19425 = ~n3277 & n15782 ;
  assign n19426 = n19425 ^ n8901 ^ 1'b0 ;
  assign n19432 = n10536 ^ n1114 ^ 1'b0 ;
  assign n19433 = n5686 & n19432 ;
  assign n19430 = ( n620 & n1438 ) | ( n620 & n5130 ) | ( n1438 & n5130 ) ;
  assign n19429 = ~n4631 & n6718 ;
  assign n19431 = n19430 ^ n19429 ^ 1'b0 ;
  assign n19434 = n19433 ^ n19431 ^ n2767 ;
  assign n19427 = n11232 ^ n2296 ^ 1'b0 ;
  assign n19428 = ~n17552 & n19427 ;
  assign n19435 = n19434 ^ n19428 ^ 1'b0 ;
  assign n19436 = ( n10960 & ~n11183 ) | ( n10960 & n17736 ) | ( ~n11183 & n17736 ) ;
  assign n19437 = n19436 ^ n18370 ^ n17436 ;
  assign n19438 = n19437 ^ n12734 ^ n10024 ;
  assign n19439 = n7314 & ~n12568 ;
  assign n19440 = n19439 ^ n5060 ^ n2260 ;
  assign n19441 = ~n2932 & n5583 ;
  assign n19442 = n19441 ^ n3813 ^ 1'b0 ;
  assign n19443 = n15498 ^ n4257 ^ 1'b0 ;
  assign n19444 = n2519 & n15465 ;
  assign n19445 = ~n5826 & n19256 ;
  assign n19446 = n19445 ^ n12545 ^ 1'b0 ;
  assign n19447 = n11221 & n19446 ;
  assign n19449 = n1564 & n19077 ;
  assign n19448 = n8332 | n17626 ;
  assign n19450 = n19449 ^ n19448 ^ 1'b0 ;
  assign n19451 = ( n3250 & n13739 ) | ( n3250 & ~n19450 ) | ( n13739 & ~n19450 ) ;
  assign n19452 = n1788 ^ n1714 ^ 1'b0 ;
  assign n19453 = n8311 | n19452 ;
  assign n19454 = n19451 & ~n19453 ;
  assign n19455 = ~n19447 & n19454 ;
  assign n19456 = n6348 & ~n6456 ;
  assign n19457 = ~n11568 & n19456 ;
  assign n19458 = n2321 & n19457 ;
  assign n19459 = n19458 ^ n11053 ^ 1'b0 ;
  assign n19460 = n19459 ^ n5168 ^ 1'b0 ;
  assign n19461 = n7435 | n19460 ;
  assign n19462 = n19461 ^ n12485 ^ n11215 ;
  assign n19463 = n15430 ^ n4669 ^ n1150 ;
  assign n19464 = n12307 & n16646 ;
  assign n19465 = ~n2148 & n5701 ;
  assign n19466 = n5032 | n8467 ;
  assign n19467 = ( n798 & ~n1304 ) | ( n798 & n19466 ) | ( ~n1304 & n19466 ) ;
  assign n19468 = n19467 ^ n2661 ^ 1'b0 ;
  assign n19469 = n19468 ^ x126 ^ 1'b0 ;
  assign n19470 = n19465 | n19469 ;
  assign n19471 = n7721 & n8614 ;
  assign n19472 = n19471 ^ n9228 ^ 1'b0 ;
  assign n19473 = n18752 ^ n5935 ^ n5533 ;
  assign n19474 = n15204 ^ n1871 ^ 1'b0 ;
  assign n19475 = ~n9539 & n19474 ;
  assign n19476 = n19475 ^ n7681 ^ 1'b0 ;
  assign n19477 = n4859 | n12946 ;
  assign n19478 = n19476 & ~n19477 ;
  assign n19479 = n11788 ^ n181 ^ 1'b0 ;
  assign n19480 = n9640 | n19479 ;
  assign n19481 = ( ~n19473 & n19478 ) | ( ~n19473 & n19480 ) | ( n19478 & n19480 ) ;
  assign n19482 = ~n3787 & n14601 ;
  assign n19483 = n19482 ^ n7895 ^ 1'b0 ;
  assign n19484 = n19483 ^ n13771 ^ n4277 ;
  assign n19485 = n18345 ^ n11049 ^ 1'b0 ;
  assign n19486 = n138 & n9628 ;
  assign n19487 = n1356 & n6110 ;
  assign n19493 = ~n5092 & n11457 ;
  assign n19494 = n6968 & n19493 ;
  assign n19488 = n8763 ^ n848 ^ 1'b0 ;
  assign n19489 = n1524 | n19488 ;
  assign n19490 = ~n5417 & n19489 ;
  assign n19491 = ( n5428 & n11645 ) | ( n5428 & ~n19490 ) | ( n11645 & ~n19490 ) ;
  assign n19492 = n2408 & n19491 ;
  assign n19495 = n19494 ^ n19492 ^ 1'b0 ;
  assign n19496 = n3421 & n5873 ;
  assign n19497 = ~n11743 & n19496 ;
  assign n19499 = n8712 & ~n12427 ;
  assign n19500 = n19499 ^ n7672 ^ 1'b0 ;
  assign n19498 = ~n5117 & n11839 ;
  assign n19501 = n19500 ^ n19498 ^ 1'b0 ;
  assign n19502 = n11181 ^ n773 ^ 1'b0 ;
  assign n19503 = n18074 & n19502 ;
  assign n19504 = ( n2333 & n6269 ) | ( n2333 & n19007 ) | ( n6269 & n19007 ) ;
  assign n19505 = n7807 ^ n1542 ^ 1'b0 ;
  assign n19509 = n6908 & ~n15981 ;
  assign n19510 = n4170 & n11719 ;
  assign n19511 = ~n19509 & n19510 ;
  assign n19506 = n1587 & ~n1918 ;
  assign n19507 = n1814 & ~n19506 ;
  assign n19508 = n7824 & n19507 ;
  assign n19512 = n19511 ^ n19508 ^ 1'b0 ;
  assign n19513 = ( n870 & n3894 ) | ( n870 & ~n6702 ) | ( n3894 & ~n6702 ) ;
  assign n19514 = n19513 ^ n8298 ^ x43 ;
  assign n19515 = n7401 & ~n14113 ;
  assign n19516 = n19515 ^ n11718 ^ 1'b0 ;
  assign n19517 = ( ~n11833 & n19514 ) | ( ~n11833 & n19516 ) | ( n19514 & n19516 ) ;
  assign n19518 = ~n1632 & n16398 ;
  assign n19519 = n16273 ^ n11534 ^ 1'b0 ;
  assign n19520 = n3974 & ~n8637 ;
  assign n19521 = n19520 ^ n3291 ^ n2870 ;
  assign n19522 = n19077 ^ n3252 ^ n860 ;
  assign n19523 = ( n2770 & ~n16284 ) | ( n2770 & n19522 ) | ( ~n16284 & n19522 ) ;
  assign n19524 = n16728 ^ n7191 ^ 1'b0 ;
  assign n19525 = n19524 ^ n4714 ^ 1'b0 ;
  assign n19526 = n9258 | n19525 ;
  assign n19527 = n776 & ~n4216 ;
  assign n19528 = ~n9715 & n18861 ;
  assign n19529 = n6625 ^ n4633 ^ 1'b0 ;
  assign n19530 = ~n19528 & n19529 ;
  assign n19531 = n3056 & n6342 ;
  assign n19532 = n19531 ^ x25 ^ 1'b0 ;
  assign n19533 = n8848 & n19532 ;
  assign n19536 = n4331 & n18549 ;
  assign n19537 = n19536 ^ n12398 ^ 1'b0 ;
  assign n19534 = ~n8043 & n18437 ;
  assign n19535 = n19534 ^ n173 ^ 1'b0 ;
  assign n19538 = n19537 ^ n19535 ^ 1'b0 ;
  assign n19539 = n3470 ^ n953 ^ 1'b0 ;
  assign n19540 = n3678 | n11723 ;
  assign n19541 = n13276 | n19540 ;
  assign n19542 = ( n19001 & ~n19539 ) | ( n19001 & n19541 ) | ( ~n19539 & n19541 ) ;
  assign n19546 = n5291 | n14201 ;
  assign n19547 = n2304 | n19546 ;
  assign n19543 = ~n6696 & n8532 ;
  assign n19544 = ~n3212 & n19543 ;
  assign n19545 = n19544 ^ n16085 ^ 1'b0 ;
  assign n19548 = n19547 ^ n19545 ^ n18124 ;
  assign n19549 = n16768 ^ n341 ^ 1'b0 ;
  assign n19550 = ( x83 & n1212 ) | ( x83 & n4871 ) | ( n1212 & n4871 ) ;
  assign n19551 = n8543 & ~n19550 ;
  assign n19552 = n143 & ~n1914 ;
  assign n19553 = n8953 & n19552 ;
  assign n19554 = n10548 ^ n845 ^ 1'b0 ;
  assign n19555 = n19553 | n19554 ;
  assign n19556 = ( n4424 & ~n8491 ) | ( n4424 & n19555 ) | ( ~n8491 & n19555 ) ;
  assign n19557 = n6339 & n16243 ;
  assign n19558 = n4781 | n13052 ;
  assign n19559 = n1184 | n19558 ;
  assign n19560 = n6948 | n8072 ;
  assign n19561 = n8924 | n19560 ;
  assign n19562 = n19561 ^ n12962 ^ 1'b0 ;
  assign n19563 = n5958 | n8970 ;
  assign n19564 = n5543 ^ n1224 ^ 1'b0 ;
  assign n19565 = n4216 | n19564 ;
  assign n19566 = n290 & ~n19565 ;
  assign n19567 = n19566 ^ n17483 ^ 1'b0 ;
  assign n19568 = n19563 & n19567 ;
  assign n19569 = n13853 ^ n3522 ^ 1'b0 ;
  assign n19570 = n13771 & n19569 ;
  assign n19571 = n4473 & n12176 ;
  assign n19572 = n19571 ^ n4797 ^ 1'b0 ;
  assign n19573 = n6530 & ~n12706 ;
  assign n19574 = n19572 & n19573 ;
  assign n19576 = n9869 | n12311 ;
  assign n19577 = n3732 | n19576 ;
  assign n19575 = n853 & n6632 ;
  assign n19578 = n19577 ^ n19575 ^ 1'b0 ;
  assign n19579 = ( n8817 & n13234 ) | ( n8817 & n18798 ) | ( n13234 & n18798 ) ;
  assign n19580 = n14770 ^ n1417 ^ 1'b0 ;
  assign n19581 = n807 | n6060 ;
  assign n19582 = n5048 & ~n6636 ;
  assign n19583 = ~n6497 & n19582 ;
  assign n19584 = n771 | n7986 ;
  assign n19585 = n19584 ^ n5663 ^ 1'b0 ;
  assign n19586 = n19585 ^ n8365 ^ 1'b0 ;
  assign n19587 = n3589 ^ n2417 ^ n888 ;
  assign n19588 = n4605 & ~n19587 ;
  assign n19589 = n11103 & n19588 ;
  assign n19590 = ( n2428 & n5206 ) | ( n2428 & ~n14620 ) | ( n5206 & ~n14620 ) ;
  assign n19594 = n6445 ^ n548 ^ 1'b0 ;
  assign n19595 = n4384 | n19594 ;
  assign n19591 = ~n1381 & n12612 ;
  assign n19592 = n19591 ^ n9439 ^ 1'b0 ;
  assign n19593 = n16935 | n19592 ;
  assign n19596 = n19595 ^ n19593 ^ 1'b0 ;
  assign n19597 = ( ~n16249 & n17960 ) | ( ~n16249 & n19596 ) | ( n17960 & n19596 ) ;
  assign n19598 = n12982 ^ n3700 ^ 1'b0 ;
  assign n19599 = n7400 | n19598 ;
  assign n19600 = n19599 ^ n2954 ^ 1'b0 ;
  assign n19601 = n654 & ~n12193 ;
  assign n19602 = n10322 ^ n10071 ^ n8823 ;
  assign n19603 = n19602 ^ n4768 ^ 1'b0 ;
  assign n19604 = ~n19601 & n19603 ;
  assign n19605 = n496 & n4885 ;
  assign n19606 = ~n270 & n19605 ;
  assign n19607 = ( n4131 & n8824 ) | ( n4131 & n11278 ) | ( n8824 & n11278 ) ;
  assign n19608 = n1770 | n19607 ;
  assign n19609 = n14173 | n19608 ;
  assign n19610 = n14622 | n19609 ;
  assign n19611 = n4829 ^ n997 ^ 1'b0 ;
  assign n19612 = n5416 & n19611 ;
  assign n19613 = n2355 | n19612 ;
  assign n19614 = n3926 | n13650 ;
  assign n19615 = n1947 | n19614 ;
  assign n19616 = n19615 ^ n5268 ^ 1'b0 ;
  assign n19617 = ( n2982 & n5939 ) | ( n2982 & ~n8325 ) | ( n5939 & ~n8325 ) ;
  assign n19618 = n19617 ^ n8441 ^ 1'b0 ;
  assign n19619 = n5588 & n7587 ;
  assign n19620 = ~n19618 & n19619 ;
  assign n19621 = n19620 ^ n14630 ^ 1'b0 ;
  assign n19626 = ~n9001 & n18283 ;
  assign n19624 = n6594 & n9806 ;
  assign n19622 = n1854 & n5384 ;
  assign n19623 = n10106 & n19622 ;
  assign n19625 = n19624 ^ n19623 ^ n932 ;
  assign n19627 = n19626 ^ n19625 ^ 1'b0 ;
  assign n19628 = n19627 ^ n4554 ^ 1'b0 ;
  assign n19629 = n16757 & ~n18196 ;
  assign n19630 = n19005 ^ n14105 ^ 1'b0 ;
  assign n19631 = n8359 ^ n7291 ^ 1'b0 ;
  assign n19632 = ~n6216 & n19631 ;
  assign n19633 = n9402 & n10526 ;
  assign n19634 = n19633 ^ n2891 ^ 1'b0 ;
  assign n19635 = n19634 ^ n7337 ^ 1'b0 ;
  assign n19636 = ( ~n3728 & n8472 ) | ( ~n3728 & n11123 ) | ( n8472 & n11123 ) ;
  assign n19637 = ( n1575 & n3420 ) | ( n1575 & ~n19636 ) | ( n3420 & ~n19636 ) ;
  assign n19638 = ( n982 & n19635 ) | ( n982 & ~n19637 ) | ( n19635 & ~n19637 ) ;
  assign n19639 = n5338 ^ n3537 ^ n1135 ;
  assign n19640 = ( n12898 & n14083 ) | ( n12898 & n15893 ) | ( n14083 & n15893 ) ;
  assign n19641 = n8099 ^ n7568 ^ n1297 ;
  assign n19642 = n9699 | n19641 ;
  assign n19643 = n19642 ^ n9904 ^ 1'b0 ;
  assign n19644 = n12724 ^ n8916 ^ 1'b0 ;
  assign n19645 = n972 | n4011 ;
  assign n19646 = n4095 | n19645 ;
  assign n19647 = n19646 ^ n17076 ^ 1'b0 ;
  assign n19648 = n10699 & n19647 ;
  assign n19649 = ( n10458 & n19644 ) | ( n10458 & ~n19648 ) | ( n19644 & ~n19648 ) ;
  assign n19650 = n5558 | n6788 ;
  assign n19651 = n19650 ^ n3512 ^ 1'b0 ;
  assign n19655 = n6811 & ~n18783 ;
  assign n19656 = n19655 ^ n2246 ^ 1'b0 ;
  assign n19652 = n6651 | n8631 ;
  assign n19653 = n5385 & ~n19652 ;
  assign n19654 = n19653 ^ n4277 ^ n3817 ;
  assign n19657 = n19656 ^ n19654 ^ 1'b0 ;
  assign n19658 = ( n408 & n1423 ) | ( n408 & n6825 ) | ( n1423 & n6825 ) ;
  assign n19659 = ( n3552 & ~n6628 ) | ( n3552 & n7504 ) | ( ~n6628 & n7504 ) ;
  assign n19660 = ~n2648 & n5380 ;
  assign n19661 = ~n14941 & n19660 ;
  assign n19662 = n4273 | n8780 ;
  assign n19663 = n8673 & ~n19662 ;
  assign n19664 = n194 & ~n19663 ;
  assign n19665 = n12882 & n19664 ;
  assign n19666 = x75 & n19665 ;
  assign n19667 = n1268 & ~n1940 ;
  assign n19668 = n9420 & n19667 ;
  assign n19669 = n2141 & ~n14556 ;
  assign n19670 = n19669 ^ n3790 ^ 1'b0 ;
  assign n19671 = ~n19668 & n19670 ;
  assign n19672 = n18846 & n19671 ;
  assign n19673 = n9077 & ~n13708 ;
  assign n19674 = n19673 ^ n7431 ^ 1'b0 ;
  assign n19675 = n9960 ^ n7789 ^ n2993 ;
  assign n19676 = n19675 ^ n16033 ^ n855 ;
  assign n19677 = n16007 ^ n15878 ^ n10527 ;
  assign n19678 = n3988 ^ n1794 ^ 1'b0 ;
  assign n19679 = n3718 & n19678 ;
  assign n19680 = ~n10044 & n14601 ;
  assign n19681 = ( n15740 & n19679 ) | ( n15740 & ~n19680 ) | ( n19679 & ~n19680 ) ;
  assign n19682 = ( n5512 & ~n7197 ) | ( n5512 & n11432 ) | ( ~n7197 & n11432 ) ;
  assign n19683 = n13746 ^ n2148 ^ 1'b0 ;
  assign n19684 = ~n19682 & n19683 ;
  assign n19685 = n2379 & n4461 ;
  assign n19686 = ~n16474 & n19685 ;
  assign n19687 = n12714 ^ n9603 ^ x80 ;
  assign n19688 = ~n19686 & n19687 ;
  assign n19689 = n4001 | n16009 ;
  assign n19690 = n15412 | n19689 ;
  assign n19691 = n11418 ^ n7740 ^ 1'b0 ;
  assign n19692 = ~n4504 & n19691 ;
  assign n19694 = n613 | n2702 ;
  assign n19695 = n8033 | n18238 ;
  assign n19696 = n6185 | n19695 ;
  assign n19697 = ~n5630 & n19696 ;
  assign n19698 = ~n19694 & n19697 ;
  assign n19699 = n19698 ^ n11296 ^ n6219 ;
  assign n19693 = n3809 & n6972 ;
  assign n19700 = n19699 ^ n19693 ^ 1'b0 ;
  assign n19701 = n18125 ^ n9533 ^ n136 ;
  assign n19702 = n15574 ^ n7207 ^ 1'b0 ;
  assign n19703 = n2481 & n2706 ;
  assign n19704 = n19702 & n19703 ;
  assign n19705 = n19704 ^ n7803 ^ n6271 ;
  assign n19706 = n6152 | n7663 ;
  assign n19707 = n6103 & ~n19706 ;
  assign n19708 = n3371 & n9204 ;
  assign n19709 = n2734 & n19708 ;
  assign n19710 = n18551 & n19709 ;
  assign n19711 = n2388 & n8707 ;
  assign n19712 = n13426 & n19711 ;
  assign n19713 = n6271 ^ n1094 ^ 1'b0 ;
  assign n19714 = ( n350 & n8807 ) | ( n350 & n10554 ) | ( n8807 & n10554 ) ;
  assign n19715 = ~n1147 & n6984 ;
  assign n19716 = n19715 ^ n1327 ^ 1'b0 ;
  assign n19717 = n5955 & n19716 ;
  assign n19718 = n19717 ^ n3915 ^ 1'b0 ;
  assign n19719 = n351 | n3459 ;
  assign n19720 = n17576 ^ n15501 ^ n10873 ;
  assign n19721 = n19356 ^ n10890 ^ n3150 ;
  assign n19722 = ( ~n19719 & n19720 ) | ( ~n19719 & n19721 ) | ( n19720 & n19721 ) ;
  assign n19723 = n5465 ^ n1829 ^ 1'b0 ;
  assign n19724 = n19723 ^ n14166 ^ 1'b0 ;
  assign n19725 = n18719 & n19724 ;
  assign n19726 = n13864 & n15907 ;
  assign n19727 = ~n3182 & n19726 ;
  assign n19728 = n11376 & ~n19727 ;
  assign n19729 = n15963 ^ n13188 ^ n6285 ;
  assign n19730 = ( n12150 & n13754 ) | ( n12150 & n14878 ) | ( n13754 & n14878 ) ;
  assign n19731 = n206 & ~n4213 ;
  assign n19732 = ~n5322 & n19731 ;
  assign n19733 = n5929 | n6059 ;
  assign n19734 = n808 | n7433 ;
  assign n19735 = ( n10651 & n16650 ) | ( n10651 & n19734 ) | ( n16650 & n19734 ) ;
  assign n19736 = ( n1049 & ~n16564 ) | ( n1049 & n19735 ) | ( ~n16564 & n19735 ) ;
  assign n19737 = ( n3231 & ~n14994 ) | ( n3231 & n16111 ) | ( ~n14994 & n16111 ) ;
  assign n19738 = n1441 & n6010 ;
  assign n19739 = ~n6997 & n19738 ;
  assign n19740 = ~n2549 & n5768 ;
  assign n19741 = n19739 & n19740 ;
  assign n19742 = n12488 ^ n6040 ^ 1'b0 ;
  assign n19743 = n17037 & ~n19742 ;
  assign n19744 = n5551 ^ n2956 ^ 1'b0 ;
  assign n19745 = n17063 ^ n5132 ^ 1'b0 ;
  assign n19746 = n10464 & n19745 ;
  assign n19747 = x34 & n11609 ;
  assign n19748 = n9332 & ~n19747 ;
  assign n19749 = n8139 ^ n1230 ^ 1'b0 ;
  assign n19750 = n17803 & ~n19749 ;
  assign n19751 = n9393 ^ n5417 ^ n3931 ;
  assign n19752 = n18312 ^ n625 ^ 1'b0 ;
  assign n19753 = ~n7219 & n19752 ;
  assign n19755 = n3428 ^ n2601 ^ 1'b0 ;
  assign n19756 = n18836 ^ n8538 ^ 1'b0 ;
  assign n19757 = n19755 & ~n19756 ;
  assign n19754 = n2371 | n9039 ;
  assign n19758 = n19757 ^ n19754 ^ 1'b0 ;
  assign n19759 = n8236 ^ n951 ^ n820 ;
  assign n19760 = x85 & n19759 ;
  assign n19761 = n16953 & ~n19760 ;
  assign n19762 = n7301 & n19761 ;
  assign n19763 = n7861 ^ n2211 ^ 1'b0 ;
  assign n19764 = ~n19762 & n19763 ;
  assign n19766 = n4329 ^ n3356 ^ 1'b0 ;
  assign n19767 = n293 & n19766 ;
  assign n19765 = n9844 ^ n7308 ^ 1'b0 ;
  assign n19768 = n19767 ^ n19765 ^ n11851 ;
  assign n19769 = n16314 ^ n16256 ^ n12673 ;
  assign n19770 = n7862 ^ n1515 ^ 1'b0 ;
  assign n19771 = n7648 & ~n19770 ;
  assign n19772 = n19771 ^ n16583 ^ 1'b0 ;
  assign n19773 = n10374 ^ n4789 ^ 1'b0 ;
  assign n19774 = n8103 & n19773 ;
  assign n19775 = n9976 | n19774 ;
  assign n19776 = n18424 ^ n3600 ^ 1'b0 ;
  assign n19777 = n19775 & ~n19776 ;
  assign n19778 = n13186 ^ n8374 ^ 1'b0 ;
  assign n19779 = n19778 ^ n5746 ^ 1'b0 ;
  assign n19780 = n12867 & ~n19779 ;
  assign n19781 = n9648 | n14744 ;
  assign n19782 = n3975 & ~n19781 ;
  assign n19783 = n19782 ^ n7081 ^ n4548 ;
  assign n19784 = n1205 | n19783 ;
  assign n19785 = n5317 ^ n932 ^ 1'b0 ;
  assign n19786 = ~n11455 & n16417 ;
  assign n19787 = n19786 ^ n1733 ^ 1'b0 ;
  assign n19788 = n4758 | n19787 ;
  assign n19789 = n5345 & n7769 ;
  assign n19790 = n2489 & ~n19789 ;
  assign n19791 = ( n10299 & ~n12336 ) | ( n10299 & n19790 ) | ( ~n12336 & n19790 ) ;
  assign n19792 = n3676 ^ n3142 ^ 1'b0 ;
  assign n19793 = n19792 ^ n8935 ^ 1'b0 ;
  assign n19796 = ( x113 & n1634 ) | ( x113 & n10465 ) | ( n1634 & n10465 ) ;
  assign n19794 = n15983 ^ n14205 ^ 1'b0 ;
  assign n19795 = n7695 & ~n19794 ;
  assign n19797 = n19796 ^ n19795 ^ n15841 ;
  assign n19798 = n17803 ^ n5857 ^ 1'b0 ;
  assign n19799 = n1714 & ~n19798 ;
  assign n19800 = ~n2761 & n9183 ;
  assign n19801 = n2087 & n19800 ;
  assign n19802 = n1748 | n19801 ;
  assign n19803 = n2145 & ~n19802 ;
  assign n19804 = n16911 ^ n9614 ^ 1'b0 ;
  assign n19806 = n7013 ^ n2748 ^ 1'b0 ;
  assign n19807 = n3667 | n19806 ;
  assign n19805 = n9182 & ~n16674 ;
  assign n19808 = n19807 ^ n19805 ^ 1'b0 ;
  assign n19809 = n771 ^ n320 ^ 1'b0 ;
  assign n19810 = n13224 | n18712 ;
  assign n19811 = n5894 | n19810 ;
  assign n19813 = n9139 ^ n7504 ^ n1734 ;
  assign n19812 = n4664 | n7469 ;
  assign n19814 = n19813 ^ n19812 ^ 1'b0 ;
  assign n19815 = ~n2972 & n5836 ;
  assign n19816 = ~n19814 & n19815 ;
  assign n19817 = n19816 ^ n6207 ^ 1'b0 ;
  assign n19818 = n7718 ^ n3980 ^ n2773 ;
  assign n19821 = n3238 | n6533 ;
  assign n19819 = n11158 ^ n6255 ^ 1'b0 ;
  assign n19820 = n5175 | n19819 ;
  assign n19822 = n19821 ^ n19820 ^ n1899 ;
  assign n19826 = n14876 ^ n298 ^ 1'b0 ;
  assign n19827 = n5187 & n19826 ;
  assign n19824 = n2200 & n3981 ;
  assign n19825 = n19824 ^ n14840 ^ 1'b0 ;
  assign n19823 = n5358 & n6289 ;
  assign n19828 = n19827 ^ n19825 ^ n19823 ;
  assign n19829 = n5002 | n11435 ;
  assign n19831 = n14711 & ~n16577 ;
  assign n19830 = n2828 & ~n18741 ;
  assign n19832 = n19831 ^ n19830 ^ 1'b0 ;
  assign n19833 = n5214 & ~n14826 ;
  assign n19834 = n19833 ^ n7685 ^ 1'b0 ;
  assign n19835 = n12718 & ~n19834 ;
  assign n19836 = n8285 & n19835 ;
  assign n19837 = n6571 & n7740 ;
  assign n19838 = n8657 ^ n7277 ^ 1'b0 ;
  assign n19839 = n9097 & n19838 ;
  assign n19840 = ~n19837 & n19839 ;
  assign n19841 = n15340 ^ n11420 ^ n5162 ;
  assign n19842 = n3194 & ~n4789 ;
  assign n19843 = n19842 ^ n404 ^ 1'b0 ;
  assign n19844 = n19843 ^ n13438 ^ 1'b0 ;
  assign n19845 = ( ~n800 & n8768 ) | ( ~n800 & n19844 ) | ( n8768 & n19844 ) ;
  assign n19846 = n7482 & n8793 ;
  assign n19847 = n15596 & n19846 ;
  assign n19848 = ( n4038 & n12264 ) | ( n4038 & n19847 ) | ( n12264 & n19847 ) ;
  assign n19852 = n16496 ^ n10257 ^ n7817 ;
  assign n19849 = n3171 & n18735 ;
  assign n19850 = n9173 & n19849 ;
  assign n19851 = n17449 | n19850 ;
  assign n19853 = n19852 ^ n19851 ^ 1'b0 ;
  assign n19854 = n2100 ^ n201 ^ 1'b0 ;
  assign n19855 = n19853 & n19854 ;
  assign n19856 = ( n5929 & ~n18572 ) | ( n5929 & n19855 ) | ( ~n18572 & n19855 ) ;
  assign n19857 = n16085 ^ n8609 ^ n327 ;
  assign n19858 = ~n7545 & n7908 ;
  assign n19859 = ( n4971 & n5374 ) | ( n4971 & ~n19858 ) | ( n5374 & ~n19858 ) ;
  assign n19860 = ( n1355 & n5233 ) | ( n1355 & n11954 ) | ( n5233 & n11954 ) ;
  assign n19861 = ( n7005 & n10309 ) | ( n7005 & ~n19860 ) | ( n10309 & ~n19860 ) ;
  assign n19862 = ~n5945 & n19861 ;
  assign n19863 = ~n2946 & n14293 ;
  assign n19864 = n19863 ^ n14288 ^ 1'b0 ;
  assign n19865 = ( n13041 & n16272 ) | ( n13041 & ~n19864 ) | ( n16272 & ~n19864 ) ;
  assign n19866 = ~n2687 & n13534 ;
  assign n19867 = n6032 & n19866 ;
  assign n19868 = n17440 | n19867 ;
  assign n19869 = n19868 ^ n2204 ^ 1'b0 ;
  assign n19870 = ~n7672 & n18948 ;
  assign n19871 = ~n5177 & n19870 ;
  assign n19872 = n4743 & n6798 ;
  assign n19873 = x5 & ~n272 ;
  assign n19874 = n3760 | n16543 ;
  assign n19875 = n18238 & ~n19874 ;
  assign n19876 = n11187 | n19875 ;
  assign n19877 = n19876 ^ n16564 ^ 1'b0 ;
  assign n19878 = n2347 & ~n10602 ;
  assign n19879 = n19878 ^ n6855 ^ 1'b0 ;
  assign n19880 = n7356 ^ n5960 ^ n3267 ;
  assign n19881 = n19880 ^ n9660 ^ 1'b0 ;
  assign n19882 = n5506 | n19881 ;
  assign n19883 = n1733 & ~n19882 ;
  assign n19884 = n19883 ^ n13052 ^ 1'b0 ;
  assign n19885 = n17074 ^ n12191 ^ 1'b0 ;
  assign n19886 = n625 & ~n15736 ;
  assign n19887 = ~n3642 & n19886 ;
  assign n19888 = ( n599 & ~n3330 ) | ( n599 & n19887 ) | ( ~n3330 & n19887 ) ;
  assign n19889 = n9078 & n19888 ;
  assign n19890 = n19885 & n19889 ;
  assign n19891 = n9778 ^ n1329 ^ 1'b0 ;
  assign n19892 = n10831 | n19891 ;
  assign n19893 = n1685 | n19892 ;
  assign n19894 = n13813 ^ n7196 ^ 1'b0 ;
  assign n19895 = n14261 ^ n7370 ^ 1'b0 ;
  assign n19896 = x65 & n5784 ;
  assign n19897 = n19896 ^ n1352 ^ 1'b0 ;
  assign n19898 = x56 & ~n16512 ;
  assign n19899 = ~n9482 & n17385 ;
  assign n19900 = n15269 ^ n1605 ^ 1'b0 ;
  assign n19901 = n822 | n19900 ;
  assign n19902 = n19211 ^ n15621 ^ 1'b0 ;
  assign n19904 = n5488 ^ n1445 ^ 1'b0 ;
  assign n19905 = n9943 & n19904 ;
  assign n19906 = n19905 ^ n10259 ^ n8493 ;
  assign n19907 = n19906 ^ n5379 ^ n4724 ;
  assign n19903 = n3826 | n4917 ;
  assign n19908 = n19907 ^ n19903 ^ n10898 ;
  assign n19909 = n14682 & ~n19908 ;
  assign n19910 = ( n17891 & n19615 ) | ( n17891 & ~n19909 ) | ( n19615 & ~n19909 ) ;
  assign n19911 = n9935 ^ n9405 ^ n1264 ;
  assign n19912 = n12036 & ~n19911 ;
  assign n19913 = n19912 ^ n2843 ^ 1'b0 ;
  assign n19914 = n18912 ^ n4593 ^ 1'b0 ;
  assign n19915 = n15123 & ~n19914 ;
  assign n19916 = n19915 ^ n540 ^ 1'b0 ;
  assign n19917 = n3096 | n12803 ;
  assign n19918 = n2795 | n19917 ;
  assign n19919 = n10049 & ~n19918 ;
  assign n19920 = ~n398 & n874 ;
  assign n19921 = n398 & n19920 ;
  assign n19922 = n19921 ^ n10554 ^ n7758 ;
  assign n19923 = n3538 ^ n2149 ^ 1'b0 ;
  assign n19924 = n11496 & ~n19923 ;
  assign n19926 = n4712 & n14595 ;
  assign n19925 = n3552 | n5765 ;
  assign n19927 = n19926 ^ n19925 ^ 1'b0 ;
  assign n19928 = n6744 & n19927 ;
  assign n19929 = n5673 & n8382 ;
  assign n19930 = n19929 ^ n7486 ^ 1'b0 ;
  assign n19931 = ~n5540 & n19930 ;
  assign n19932 = ~n6380 & n19931 ;
  assign n19933 = ~n13961 & n19932 ;
  assign n19934 = n19933 ^ n11211 ^ 1'b0 ;
  assign n19935 = ~n17875 & n19934 ;
  assign n19936 = n19935 ^ n17700 ^ 1'b0 ;
  assign n19938 = n9600 & ~n16078 ;
  assign n19939 = n19938 ^ n5181 ^ 1'b0 ;
  assign n19937 = n8263 ^ n4592 ^ 1'b0 ;
  assign n19940 = n19939 ^ n19937 ^ n19208 ;
  assign n19941 = n18658 ^ n9533 ^ 1'b0 ;
  assign n19943 = n1815 ^ n781 ^ 1'b0 ;
  assign n19942 = n6996 ^ n5442 ^ 1'b0 ;
  assign n19944 = n19943 ^ n19942 ^ n2082 ;
  assign n19945 = ( n4292 & ~n17278 ) | ( n4292 & n19944 ) | ( ~n17278 & n19944 ) ;
  assign n19946 = ( n6017 & n7176 ) | ( n6017 & n8791 ) | ( n7176 & n8791 ) ;
  assign n19947 = n19946 ^ n10072 ^ n3341 ;
  assign n19948 = ~n14964 & n19947 ;
  assign n19949 = ~n6998 & n8024 ;
  assign n19950 = n19949 ^ n13682 ^ 1'b0 ;
  assign n19954 = n1062 & ~n9509 ;
  assign n19951 = n9755 ^ n5533 ^ 1'b0 ;
  assign n19952 = n11357 | n19951 ;
  assign n19953 = n11022 & ~n19952 ;
  assign n19955 = n19954 ^ n19953 ^ 1'b0 ;
  assign n19956 = ( ~n2226 & n3323 ) | ( ~n2226 & n7359 ) | ( n3323 & n7359 ) ;
  assign n19957 = ~n19702 & n19939 ;
  assign n19958 = n6818 | n8657 ;
  assign n19959 = n6118 | n14436 ;
  assign n19960 = ( n13586 & ~n19958 ) | ( n13586 & n19959 ) | ( ~n19958 & n19959 ) ;
  assign n19961 = n10918 ^ n9073 ^ 1'b0 ;
  assign n19962 = ~n7501 & n19961 ;
  assign n19963 = ~n4938 & n17623 ;
  assign n19964 = ~n9881 & n19963 ;
  assign n19965 = n514 | n19754 ;
  assign n19966 = n8310 ^ n3403 ^ 1'b0 ;
  assign n19967 = ( n16418 & n17233 ) | ( n16418 & n19966 ) | ( n17233 & n19966 ) ;
  assign n19968 = ~n1956 & n19967 ;
  assign n19969 = ~n4290 & n12857 ;
  assign n19970 = ( n3978 & n14762 ) | ( n3978 & n19969 ) | ( n14762 & n19969 ) ;
  assign n19971 = n17893 ^ n3629 ^ 1'b0 ;
  assign n19972 = n19970 & n19971 ;
  assign n19973 = n6306 & ~n7099 ;
  assign n19974 = n5012 ^ n1462 ^ 1'b0 ;
  assign n19975 = ~n19973 & n19974 ;
  assign n19976 = n4160 & ~n13006 ;
  assign n19977 = n266 & ~n19976 ;
  assign n19978 = n5072 | n6059 ;
  assign n19979 = n236 & n686 ;
  assign n19980 = ~n19978 & n19979 ;
  assign n19981 = n15221 ^ n5537 ^ 1'b0 ;
  assign n19982 = n9359 & n19981 ;
  assign n19983 = ( ~n5965 & n19980 ) | ( ~n5965 & n19982 ) | ( n19980 & n19982 ) ;
  assign n19984 = n1205 | n17051 ;
  assign n19985 = n13413 ^ n4700 ^ 1'b0 ;
  assign n19986 = n12016 & ~n19985 ;
  assign n19987 = n9955 | n19361 ;
  assign n19988 = n14601 | n19987 ;
  assign n19989 = n10618 | n14854 ;
  assign n19990 = n19989 ^ n5387 ^ 1'b0 ;
  assign n19994 = n3925 | n6758 ;
  assign n19995 = n3925 & ~n19994 ;
  assign n19996 = n4712 | n19995 ;
  assign n19997 = n19995 & ~n19996 ;
  assign n19998 = n2626 & n7200 ;
  assign n19999 = ~n7200 & n19998 ;
  assign n20000 = n19999 ^ n568 ^ 1'b0 ;
  assign n20001 = ~n568 & n20000 ;
  assign n20002 = ~n5502 & n20001 ;
  assign n20003 = n5502 & n20002 ;
  assign n20004 = n353 | n20003 ;
  assign n20005 = n19997 & ~n20004 ;
  assign n19991 = x41 & n148 ;
  assign n19992 = ~x41 & n19991 ;
  assign n19993 = n18333 | n19992 ;
  assign n20006 = n20005 ^ n19993 ^ n819 ;
  assign n20007 = n2770 & n5241 ;
  assign n20008 = n20007 ^ n12827 ^ 1'b0 ;
  assign n20009 = n7314 ^ x111 ^ 1'b0 ;
  assign n20010 = n9109 & n16307 ;
  assign n20011 = n20010 ^ n16070 ^ 1'b0 ;
  assign n20012 = n20009 | n20011 ;
  assign n20013 = ~n3393 & n5331 ;
  assign n20014 = n784 | n9892 ;
  assign n20015 = n20014 ^ x73 ^ 1'b0 ;
  assign n20016 = n7073 & ~n16231 ;
  assign n20017 = n20016 ^ n7479 ^ 1'b0 ;
  assign n20018 = n16266 | n20017 ;
  assign n20019 = n3005 & ~n6513 ;
  assign n20020 = n19172 ^ n11460 ^ n11376 ;
  assign n20024 = ( n3802 & n6214 ) | ( n3802 & n6664 ) | ( n6214 & n6664 ) ;
  assign n20022 = n5002 & ~n13927 ;
  assign n20023 = n17057 & n20022 ;
  assign n20021 = n138 | n17784 ;
  assign n20025 = n20024 ^ n20023 ^ n20021 ;
  assign n20026 = n7331 & ~n7506 ;
  assign n20027 = n1996 & n11101 ;
  assign n20028 = n20027 ^ n2445 ^ 1'b0 ;
  assign n20029 = n5057 | n14166 ;
  assign n20030 = x63 | n20029 ;
  assign n20031 = n6675 ^ n4661 ^ n3942 ;
  assign n20032 = n10605 ^ n5045 ^ 1'b0 ;
  assign n20033 = n20031 & ~n20032 ;
  assign n20034 = ( n2930 & n5049 ) | ( n2930 & ~n6750 ) | ( n5049 & ~n6750 ) ;
  assign n20035 = n8644 ^ n2593 ^ 1'b0 ;
  assign n20036 = ~n20034 & n20035 ;
  assign n20037 = n8880 ^ n1845 ^ 1'b0 ;
  assign n20038 = n8005 & n20037 ;
  assign n20039 = n20038 ^ n13542 ^ n797 ;
  assign n20040 = n20039 ^ n17102 ^ n15637 ;
  assign n20041 = ( n1554 & ~n3949 ) | ( n1554 & n11313 ) | ( ~n3949 & n11313 ) ;
  assign n20042 = ~n6567 & n12813 ;
  assign n20043 = n9369 ^ n1369 ^ 1'b0 ;
  assign n20044 = n18215 | n20043 ;
  assign n20045 = n20044 ^ n10050 ^ n9820 ;
  assign n20046 = n20045 ^ n19144 ^ 1'b0 ;
  assign n20047 = n2592 | n4211 ;
  assign n20048 = n20047 ^ n6185 ^ n3541 ;
  assign n20049 = ~n9302 & n20048 ;
  assign n20050 = ( n5125 & n7798 ) | ( n5125 & n9892 ) | ( n7798 & n9892 ) ;
  assign n20051 = n3862 ^ n3222 ^ 1'b0 ;
  assign n20052 = ~n9467 & n20051 ;
  assign n20053 = n19343 | n20052 ;
  assign n20054 = n10080 | n19480 ;
  assign n20055 = n20054 ^ n13650 ^ 1'b0 ;
  assign n20056 = n14001 | n20055 ;
  assign n20057 = ( n173 & n5314 ) | ( n173 & n14714 ) | ( n5314 & n14714 ) ;
  assign n20058 = n6471 & ~n20057 ;
  assign n20059 = n15036 ^ n6428 ^ n3533 ;
  assign n20060 = n986 | n20059 ;
  assign n20061 = ~n6249 & n13827 ;
  assign n20062 = n2937 | n10243 ;
  assign n20063 = n20062 ^ n14210 ^ n6867 ;
  assign n20064 = ( x49 & n3274 ) | ( x49 & n16474 ) | ( n3274 & n16474 ) ;
  assign n20065 = n20064 ^ n8204 ^ n1856 ;
  assign n20066 = n3745 ^ n3664 ^ 1'b0 ;
  assign n20067 = n15554 ^ n8127 ^ 1'b0 ;
  assign n20068 = ~n4844 & n20067 ;
  assign n20069 = n14323 ^ n13846 ^ 1'b0 ;
  assign n20070 = ( n1691 & n5172 ) | ( n1691 & ~n17552 ) | ( n5172 & ~n17552 ) ;
  assign n20071 = n17191 & ~n20070 ;
  assign n20072 = n17859 ^ n13983 ^ 1'b0 ;
  assign n20073 = n19760 | n20072 ;
  assign n20074 = ~n3717 & n13155 ;
  assign n20075 = n13499 & ~n19524 ;
  assign n20076 = ~n3772 & n10420 ;
  assign n20077 = ~n2402 & n20076 ;
  assign n20078 = n18781 ^ n8138 ^ 1'b0 ;
  assign n20080 = n2124 & n10210 ;
  assign n20079 = n13528 & ~n13856 ;
  assign n20081 = n20080 ^ n20079 ^ 1'b0 ;
  assign n20082 = ~n2942 & n3923 ;
  assign n20083 = n20082 ^ n15535 ^ n7852 ;
  assign n20084 = ( n15390 & ~n20081 ) | ( n15390 & n20083 ) | ( ~n20081 & n20083 ) ;
  assign n20085 = ( ~n16828 & n17196 ) | ( ~n16828 & n20084 ) | ( n17196 & n20084 ) ;
  assign n20086 = ~n561 & n6530 ;
  assign n20087 = n17717 | n20086 ;
  assign n20088 = n13819 ^ n4095 ^ 1'b0 ;
  assign n20089 = ~n4749 & n20088 ;
  assign n20090 = n10703 ^ n154 ^ 1'b0 ;
  assign n20091 = n225 & n11555 ;
  assign n20092 = ~n19567 & n20091 ;
  assign n20097 = n1320 & n7479 ;
  assign n20096 = n157 | n13844 ;
  assign n20098 = n20097 ^ n20096 ^ 1'b0 ;
  assign n20099 = n12333 | n20098 ;
  assign n20100 = n20099 ^ n14127 ^ 1'b0 ;
  assign n20093 = n9163 ^ n5988 ^ 1'b0 ;
  assign n20094 = n20093 ^ n5522 ^ n1146 ;
  assign n20095 = ( n5612 & n11458 ) | ( n5612 & n20094 ) | ( n11458 & n20094 ) ;
  assign n20101 = n20100 ^ n20095 ^ 1'b0 ;
  assign n20104 = ( n1414 & n4054 ) | ( n1414 & ~n6297 ) | ( n4054 & ~n6297 ) ;
  assign n20102 = n6793 & n13620 ;
  assign n20103 = ( n146 & n9883 ) | ( n146 & ~n20102 ) | ( n9883 & ~n20102 ) ;
  assign n20105 = n20104 ^ n20103 ^ n1490 ;
  assign n20106 = n2974 | n20105 ;
  assign n20107 = n20106 ^ n17980 ^ 1'b0 ;
  assign n20109 = n12289 ^ n10918 ^ 1'b0 ;
  assign n20108 = n4904 & n7624 ;
  assign n20110 = n20109 ^ n20108 ^ 1'b0 ;
  assign n20111 = n4978 ^ x117 ^ 1'b0 ;
  assign n20112 = n3005 & n20111 ;
  assign n20113 = ~n12183 & n20112 ;
  assign n20114 = n20113 ^ n2504 ^ 1'b0 ;
  assign n20115 = n20114 ^ n11853 ^ 1'b0 ;
  assign n20117 = n1856 & ~n2619 ;
  assign n20118 = n20117 ^ n7056 ^ 1'b0 ;
  assign n20119 = n20118 ^ n1143 ^ 1'b0 ;
  assign n20116 = ~n5233 & n9271 ;
  assign n20120 = n20119 ^ n20116 ^ 1'b0 ;
  assign n20121 = ~n1075 & n1881 ;
  assign n20122 = n5748 ^ n2824 ^ 1'b0 ;
  assign n20123 = ~n929 & n6030 ;
  assign n20124 = n6035 ^ n2113 ^ 1'b0 ;
  assign n20125 = n20123 & ~n20124 ;
  assign n20126 = ~n1680 & n5568 ;
  assign n20127 = ~n2401 & n9764 ;
  assign n20128 = n14620 ^ n10709 ^ 1'b0 ;
  assign n20129 = ~n6974 & n20128 ;
  assign n20130 = n1039 & ~n10232 ;
  assign n20131 = n20130 ^ n1118 ^ 1'b0 ;
  assign n20132 = n11531 ^ n7370 ^ n259 ;
  assign n20133 = n10036 ^ n4926 ^ n4359 ;
  assign n20134 = n319 & ~n6661 ;
  assign n20139 = n11541 ^ n5159 ^ 1'b0 ;
  assign n20137 = n5341 ^ n1042 ^ 1'b0 ;
  assign n20135 = n805 & ~n880 ;
  assign n20136 = n20135 ^ n2849 ^ 1'b0 ;
  assign n20138 = n20137 ^ n20136 ^ n15768 ;
  assign n20140 = n20139 ^ n20138 ^ 1'b0 ;
  assign n20141 = x69 & n20140 ;
  assign n20142 = n16502 & n20141 ;
  assign n20143 = n2952 & n14994 ;
  assign n20144 = ( n617 & n6079 ) | ( n617 & ~n16840 ) | ( n6079 & ~n16840 ) ;
  assign n20145 = ~n1657 & n11100 ;
  assign n20146 = n3848 | n5252 ;
  assign n20147 = n229 & ~n20146 ;
  assign n20148 = n653 & ~n6372 ;
  assign n20149 = n20148 ^ n11207 ^ 1'b0 ;
  assign n20150 = n16455 ^ n12160 ^ 1'b0 ;
  assign n20151 = n10806 & ~n11787 ;
  assign n20152 = n20151 ^ n19029 ^ 1'b0 ;
  assign n20153 = n20152 ^ n2334 ^ 1'b0 ;
  assign n20154 = n4295 ^ n270 ^ 1'b0 ;
  assign n20155 = n1806 | n12248 ;
  assign n20156 = n2554 | n20155 ;
  assign n20157 = n11471 ^ n10527 ^ n8325 ;
  assign n20158 = n4694 ^ n3507 ^ 1'b0 ;
  assign n20159 = ( n398 & n10784 ) | ( n398 & ~n20158 ) | ( n10784 & ~n20158 ) ;
  assign n20160 = ( n1331 & n3141 ) | ( n1331 & ~n5131 ) | ( n3141 & ~n5131 ) ;
  assign n20161 = n2372 ^ n644 ^ 1'b0 ;
  assign n20162 = n17666 ^ n1064 ^ 1'b0 ;
  assign n20163 = ( n14820 & n20161 ) | ( n14820 & n20162 ) | ( n20161 & n20162 ) ;
  assign n20164 = n14697 ^ n9963 ^ 1'b0 ;
  assign n20165 = n4927 & n20164 ;
  assign n20166 = n401 & n9432 ;
  assign n20167 = n1644 & ~n4978 ;
  assign n20168 = n768 | n20167 ;
  assign n20169 = n10644 ^ n5945 ^ 1'b0 ;
  assign n20170 = ~n20168 & n20169 ;
  assign n20171 = n20170 ^ n16656 ^ 1'b0 ;
  assign n20172 = ( n2846 & ~n3493 ) | ( n2846 & n4216 ) | ( ~n3493 & n4216 ) ;
  assign n20173 = ~n1276 & n5671 ;
  assign n20174 = ~n20172 & n20173 ;
  assign n20175 = n14514 ^ n3968 ^ n1770 ;
  assign n20176 = ~n12207 & n20175 ;
  assign n20177 = n13568 & n20176 ;
  assign n20178 = n7469 & ~n20177 ;
  assign n20179 = n20178 ^ n17041 ^ n16144 ;
  assign n20180 = n5009 ^ n2553 ^ 1'b0 ;
  assign n20181 = n9133 ^ n6750 ^ 1'b0 ;
  assign n20182 = n5557 | n20181 ;
  assign n20183 = n1689 & n5539 ;
  assign n20184 = ~n10222 & n20183 ;
  assign n20185 = ( n15755 & n20182 ) | ( n15755 & ~n20184 ) | ( n20182 & ~n20184 ) ;
  assign n20186 = n20180 & n20185 ;
  assign n20187 = n16230 ^ n9790 ^ 1'b0 ;
  assign n20188 = ~n3122 & n20187 ;
  assign n20189 = n8860 ^ n1485 ^ 1'b0 ;
  assign n20191 = ~n10180 & n11946 ;
  assign n20190 = n3357 | n8265 ;
  assign n20192 = n20191 ^ n20190 ^ 1'b0 ;
  assign n20193 = n20192 ^ n5655 ^ 1'b0 ;
  assign n20194 = ~n20189 & n20193 ;
  assign n20196 = n3576 | n5231 ;
  assign n20197 = n2573 & ~n20196 ;
  assign n20198 = ( n6264 & ~n17441 ) | ( n6264 & n20197 ) | ( ~n17441 & n20197 ) ;
  assign n20195 = n9064 | n10646 ;
  assign n20199 = n20198 ^ n20195 ^ 1'b0 ;
  assign n20200 = n16728 ^ n8949 ^ n7758 ;
  assign n20201 = n20200 ^ n6915 ^ n5798 ;
  assign n20202 = ~n5196 & n20201 ;
  assign n20203 = n10114 & n20202 ;
  assign n20204 = n2903 | n20191 ;
  assign n20205 = n1774 & ~n20204 ;
  assign n20206 = n10331 & ~n20205 ;
  assign n20207 = n8909 & n20206 ;
  assign n20208 = ( n7396 & n7499 ) | ( n7396 & ~n11170 ) | ( n7499 & ~n11170 ) ;
  assign n20209 = n20208 ^ n13519 ^ n5937 ;
  assign n20210 = n20209 ^ n1326 ^ 1'b0 ;
  assign n20211 = ~n18090 & n20210 ;
  assign n20212 = n20211 ^ n15781 ^ 1'b0 ;
  assign n20213 = ~n7153 & n17992 ;
  assign n20214 = n10480 ^ n4927 ^ 1'b0 ;
  assign n20215 = ~n17427 & n20214 ;
  assign n20218 = n5828 | n12333 ;
  assign n20219 = n20218 ^ n10155 ^ 1'b0 ;
  assign n20216 = n16030 ^ n5360 ^ 1'b0 ;
  assign n20217 = n20216 ^ n9844 ^ n8318 ;
  assign n20220 = n20219 ^ n20217 ^ 1'b0 ;
  assign n20221 = n206 & ~n11430 ;
  assign n20222 = ~n19827 & n20221 ;
  assign n20223 = n3146 ^ n877 ^ 1'b0 ;
  assign n20224 = n12168 | n20223 ;
  assign n20225 = n20224 ^ n2817 ^ 1'b0 ;
  assign n20226 = n9383 | n10676 ;
  assign n20227 = ( n13715 & n19529 ) | ( n13715 & n20226 ) | ( n19529 & n20226 ) ;
  assign n20229 = ( n2231 & ~n2573 ) | ( n2231 & n19539 ) | ( ~n2573 & n19539 ) ;
  assign n20228 = n3856 & ~n5421 ;
  assign n20230 = n20229 ^ n20228 ^ n5206 ;
  assign n20231 = n9147 ^ n618 ^ 1'b0 ;
  assign n20232 = n20231 ^ n13553 ^ 1'b0 ;
  assign n20233 = n20230 | n20232 ;
  assign n20234 = n20233 ^ n2976 ^ 1'b0 ;
  assign n20237 = n1175 | n8677 ;
  assign n20235 = ( ~n2688 & n2865 ) | ( ~n2688 & n6640 ) | ( n2865 & n6640 ) ;
  assign n20236 = ( ~n3987 & n6098 ) | ( ~n3987 & n20235 ) | ( n6098 & n20235 ) ;
  assign n20238 = n20237 ^ n20236 ^ n8299 ;
  assign n20239 = ( n2532 & ~n10015 ) | ( n2532 & n18269 ) | ( ~n10015 & n18269 ) ;
  assign n20240 = n20239 ^ n7196 ^ n6571 ;
  assign n20241 = n10313 ^ n3956 ^ 1'b0 ;
  assign n20242 = n20240 | n20241 ;
  assign n20243 = n5147 & n6264 ;
  assign n20244 = n2985 & n20243 ;
  assign n20245 = ~n10008 & n15395 ;
  assign n20246 = n7551 & n7986 ;
  assign n20247 = ( x80 & n10883 ) | ( x80 & ~n20246 ) | ( n10883 & ~n20246 ) ;
  assign n20248 = n16468 & n20247 ;
  assign n20249 = n4372 | n18308 ;
  assign n20250 = n16372 & ~n20249 ;
  assign n20251 = n11875 ^ n5967 ^ n4706 ;
  assign n20252 = ~n9126 & n20251 ;
  assign n20253 = n2565 | n5575 ;
  assign n20254 = n20252 & ~n20253 ;
  assign n20255 = n12452 ^ n9509 ^ 1'b0 ;
  assign n20256 = n8732 & n20255 ;
  assign n20257 = ( ~n1781 & n12186 ) | ( ~n1781 & n20256 ) | ( n12186 & n20256 ) ;
  assign n20259 = n14312 ^ n7486 ^ 1'b0 ;
  assign n20260 = n918 & ~n20259 ;
  assign n20258 = n3981 & ~n14334 ;
  assign n20261 = n20260 ^ n20258 ^ 1'b0 ;
  assign n20262 = ~n7553 & n15093 ;
  assign n20263 = ~n19677 & n20262 ;
  assign n20264 = n3433 | n5053 ;
  assign n20265 = n7038 | n20264 ;
  assign n20266 = n7316 ^ n5169 ^ n1491 ;
  assign n20267 = n5380 & n18340 ;
  assign n20268 = n3525 & n20267 ;
  assign n20269 = n20268 ^ n4332 ^ 1'b0 ;
  assign n20270 = n11900 | n16935 ;
  assign n20271 = n20270 ^ n12363 ^ 1'b0 ;
  assign n20272 = n9588 ^ n7865 ^ 1'b0 ;
  assign n20273 = ~n20271 & n20272 ;
  assign n20274 = n6550 & n16524 ;
  assign n20275 = n20274 ^ n9734 ^ 1'b0 ;
  assign n20276 = ~n6178 & n20275 ;
  assign n20277 = ~n11376 & n20276 ;
  assign n20278 = n8609 ^ n2148 ^ 1'b0 ;
  assign n20279 = ~n2616 & n20278 ;
  assign n20280 = ( n5100 & ~n5458 ) | ( n5100 & n6675 ) | ( ~n5458 & n6675 ) ;
  assign n20281 = ( n4199 & n20279 ) | ( n4199 & n20280 ) | ( n20279 & n20280 ) ;
  assign n20282 = n8614 & n16643 ;
  assign n20283 = n20282 ^ n9841 ^ n4336 ;
  assign n20284 = n1442 & n2044 ;
  assign n20285 = ~n12858 & n20284 ;
  assign n20286 = ( n4397 & n5477 ) | ( n4397 & n20285 ) | ( n5477 & n20285 ) ;
  assign n20287 = ( ~n2211 & n4658 ) | ( ~n2211 & n12635 ) | ( n4658 & n12635 ) ;
  assign n20288 = ~n3534 & n15540 ;
  assign n20289 = n11887 & n20288 ;
  assign n20290 = ( n4296 & ~n9573 ) | ( n4296 & n9946 ) | ( ~n9573 & n9946 ) ;
  assign n20291 = n3923 & ~n16829 ;
  assign n20292 = ~n20290 & n20291 ;
  assign n20293 = n15321 ^ n10250 ^ n9384 ;
  assign n20294 = ~n1781 & n3816 ;
  assign n20295 = ~n20293 & n20294 ;
  assign n20296 = ~n5278 & n13467 ;
  assign n20297 = n20296 ^ n7427 ^ 1'b0 ;
  assign n20298 = n20297 ^ n12314 ^ 1'b0 ;
  assign n20299 = n18861 ^ n9158 ^ 1'b0 ;
  assign n20300 = ~n7448 & n20299 ;
  assign n20301 = n19185 ^ n4623 ^ n4505 ;
  assign n20302 = n10624 | n20301 ;
  assign n20303 = n20300 | n20302 ;
  assign n20304 = ( ~x123 & n12219 ) | ( ~x123 & n20303 ) | ( n12219 & n20303 ) ;
  assign n20307 = n5956 ^ x72 ^ 1'b0 ;
  assign n20308 = n11095 | n20307 ;
  assign n20305 = n2743 ^ n2581 ^ 1'b0 ;
  assign n20306 = ( ~n7925 & n17074 ) | ( ~n7925 & n20305 ) | ( n17074 & n20305 ) ;
  assign n20309 = n20308 ^ n20306 ^ n7931 ;
  assign n20310 = ( n7803 & n8599 ) | ( n7803 & ~n13125 ) | ( n8599 & ~n13125 ) ;
  assign n20311 = n3012 | n20310 ;
  assign n20312 = n20311 ^ n10474 ^ 1'b0 ;
  assign n20313 = ( n1375 & ~n18403 ) | ( n1375 & n19258 ) | ( ~n18403 & n19258 ) ;
  assign n20314 = n15356 ^ n11651 ^ 1'b0 ;
  assign n20315 = n20313 & ~n20314 ;
  assign n20316 = n5523 | n16541 ;
  assign n20317 = n5483 ^ n1708 ^ 1'b0 ;
  assign n20320 = n915 & ~n3521 ;
  assign n20318 = n17110 ^ n2946 ^ 1'b0 ;
  assign n20319 = n10660 & ~n20318 ;
  assign n20321 = n20320 ^ n20319 ^ x24 ;
  assign n20322 = n18178 ^ n7094 ^ 1'b0 ;
  assign n20323 = ( n5329 & n11989 ) | ( n5329 & n16682 ) | ( n11989 & n16682 ) ;
  assign n20324 = n20323 ^ n5484 ^ n4820 ;
  assign n20325 = n10155 ^ n5568 ^ 1'b0 ;
  assign n20326 = n18369 & ~n20325 ;
  assign n20327 = n15493 ^ n7892 ^ 1'b0 ;
  assign n20328 = n11940 & ~n18772 ;
  assign n20329 = n10625 ^ n753 ^ 1'b0 ;
  assign n20330 = x2 & n1569 ;
  assign n20331 = n20330 ^ n838 ^ 1'b0 ;
  assign n20332 = ( n15242 & n20329 ) | ( n15242 & n20331 ) | ( n20329 & n20331 ) ;
  assign n20335 = ( n2581 & n2947 ) | ( n2581 & ~n4273 ) | ( n2947 & ~n4273 ) ;
  assign n20336 = n20335 ^ n16185 ^ n3417 ;
  assign n20333 = ( n3108 & n4407 ) | ( n3108 & ~n20007 ) | ( n4407 & ~n20007 ) ;
  assign n20334 = n20333 ^ n12901 ^ n9751 ;
  assign n20337 = n20336 ^ n20334 ^ 1'b0 ;
  assign n20338 = n16344 ^ n9384 ^ n2189 ;
  assign n20339 = n1404 | n13603 ;
  assign n20340 = n20339 ^ n3873 ^ 1'b0 ;
  assign n20341 = n12024 ^ n7413 ^ x114 ;
  assign n20342 = ( n20338 & n20340 ) | ( n20338 & n20341 ) | ( n20340 & n20341 ) ;
  assign n20343 = n4636 & n7420 ;
  assign n20344 = n8282 & ~n20343 ;
  assign n20345 = n3138 | n7442 ;
  assign n20346 = n10859 & n20345 ;
  assign n20347 = n20346 ^ n17011 ^ 1'b0 ;
  assign n20348 = ( n6003 & ~n11321 ) | ( n6003 & n13872 ) | ( ~n11321 & n13872 ) ;
  assign n20349 = ~n1678 & n2945 ;
  assign n20352 = ( x7 & ~n324 ) | ( x7 & n4246 ) | ( ~n324 & n4246 ) ;
  assign n20350 = n2044 & n2269 ;
  assign n20351 = ~n5899 & n20350 ;
  assign n20353 = n20352 ^ n20351 ^ 1'b0 ;
  assign n20354 = n9107 | n20353 ;
  assign n20355 = n11028 ^ n10218 ^ 1'b0 ;
  assign n20356 = n17727 ^ n4329 ^ n1511 ;
  assign n20357 = n9314 & ~n20356 ;
  assign n20358 = ( n3436 & n6055 ) | ( n3436 & ~n6346 ) | ( n6055 & ~n6346 ) ;
  assign n20362 = ( n8200 & ~n8994 ) | ( n8200 & n11944 ) | ( ~n8994 & n11944 ) ;
  assign n20363 = n8516 ^ n5269 ^ 1'b0 ;
  assign n20364 = n3079 | n20363 ;
  assign n20365 = n20362 & ~n20364 ;
  assign n20366 = n20365 ^ n10644 ^ 1'b0 ;
  assign n20367 = ~n8850 & n20366 ;
  assign n20368 = n5387 & n20367 ;
  assign n20359 = ~n16892 & n17851 ;
  assign n20360 = n20359 ^ n2058 ^ 1'b0 ;
  assign n20361 = n4512 & n20360 ;
  assign n20369 = n20368 ^ n20361 ^ 1'b0 ;
  assign n20370 = n16861 ^ n7317 ^ 1'b0 ;
  assign n20372 = n6273 ^ n1491 ^ 1'b0 ;
  assign n20373 = n3887 | n20372 ;
  assign n20371 = ~n1524 & n6203 ;
  assign n20374 = n20373 ^ n20371 ^ 1'b0 ;
  assign n20375 = ( ~n2611 & n3695 ) | ( ~n2611 & n6849 ) | ( n3695 & n6849 ) ;
  assign n20376 = n1338 | n7543 ;
  assign n20377 = n20375 & ~n20376 ;
  assign n20378 = ~n1272 & n19529 ;
  assign n20379 = n679 & ~n19457 ;
  assign n20380 = x29 & n2130 ;
  assign n20381 = n10500 & n20380 ;
  assign n20382 = n20381 ^ n2616 ^ 1'b0 ;
  assign n20383 = n1173 & n20382 ;
  assign n20384 = n20383 ^ n3341 ^ 1'b0 ;
  assign n20385 = n508 ^ x58 ^ 1'b0 ;
  assign n20386 = n818 & n6003 ;
  assign n20387 = n20385 & n20386 ;
  assign n20388 = ~n2390 & n7338 ;
  assign n20389 = ~n5154 & n20388 ;
  assign n20390 = ~n14053 & n20389 ;
  assign n20391 = n10086 ^ n8037 ^ 1'b0 ;
  assign n20392 = n11891 | n17007 ;
  assign n20393 = n20392 ^ n11136 ^ n2828 ;
  assign n20394 = ( ~n2165 & n9711 ) | ( ~n2165 & n20393 ) | ( n9711 & n20393 ) ;
  assign n20395 = ( n5689 & n6164 ) | ( n5689 & n18980 ) | ( n6164 & n18980 ) ;
  assign n20396 = n2779 & n14872 ;
  assign n20397 = n808 & n20396 ;
  assign n20398 = n5352 & ~n8033 ;
  assign n20399 = ~n2406 & n20398 ;
  assign n20400 = ( n5565 & n20397 ) | ( n5565 & ~n20399 ) | ( n20397 & ~n20399 ) ;
  assign n20401 = n804 | n14136 ;
  assign n20402 = ~n3399 & n4900 ;
  assign n20403 = n20402 ^ n913 ^ 1'b0 ;
  assign n20404 = n932 | n12217 ;
  assign n20405 = n14992 ^ n7785 ^ 1'b0 ;
  assign n20406 = n20404 & n20405 ;
  assign n20407 = n3638 | n14064 ;
  assign n20408 = n3119 & ~n11954 ;
  assign n20409 = n8130 & n11099 ;
  assign n20410 = ~n947 & n20409 ;
  assign n20411 = n9532 | n20410 ;
  assign n20412 = n12781 & ~n12936 ;
  assign n20413 = n20412 ^ n13442 ^ 1'b0 ;
  assign n20414 = n20413 ^ n8585 ^ n4674 ;
  assign n20415 = n7404 ^ x6 ^ 1'b0 ;
  assign n20416 = n12284 ^ n2792 ^ n1195 ;
  assign n20417 = n3027 | n20416 ;
  assign n20418 = n20415 | n20417 ;
  assign n20419 = n13974 ^ n4942 ^ n4235 ;
  assign n20420 = ~n5888 & n8835 ;
  assign n20421 = n20419 & n20420 ;
  assign n20422 = n20421 ^ n7663 ^ 1'b0 ;
  assign n20423 = ( n946 & n5522 ) | ( n946 & ~n9132 ) | ( n5522 & ~n9132 ) ;
  assign n20424 = n12336 ^ n8194 ^ n1163 ;
  assign n20425 = n16636 & ~n20424 ;
  assign n20426 = n20423 & n20425 ;
  assign n20427 = ( n1972 & n3709 ) | ( n1972 & ~n12950 ) | ( n3709 & ~n12950 ) ;
  assign n20428 = ( n322 & n5883 ) | ( n322 & ~n20427 ) | ( n5883 & ~n20427 ) ;
  assign n20429 = n12014 & n16766 ;
  assign n20430 = x113 | n1839 ;
  assign n20431 = n5997 ^ n2653 ^ x87 ;
  assign n20432 = n19474 ^ n4385 ^ 1'b0 ;
  assign n20433 = n20431 & n20432 ;
  assign n20434 = n607 | n2338 ;
  assign n20435 = n20434 ^ x126 ^ 1'b0 ;
  assign n20436 = ( n4945 & n15980 ) | ( n4945 & ~n20435 ) | ( n15980 & ~n20435 ) ;
  assign n20437 = n686 & n12317 ;
  assign n20438 = n3327 & n15612 ;
  assign n20439 = ~n831 & n7075 ;
  assign n20440 = n5333 & n8217 ;
  assign n20441 = ~n10757 & n20440 ;
  assign n20442 = n20439 | n20441 ;
  assign n20445 = n13594 ^ n8390 ^ 1'b0 ;
  assign n20446 = n7528 & n20445 ;
  assign n20443 = n5402 ^ n3938 ^ n2126 ;
  assign n20444 = ( ~n8712 & n9940 ) | ( ~n8712 & n20443 ) | ( n9940 & n20443 ) ;
  assign n20447 = n20446 ^ n20444 ^ n8169 ;
  assign n20454 = ~n4896 & n6378 ;
  assign n20450 = n9967 ^ n9216 ^ n5954 ;
  assign n20451 = n13892 & n20450 ;
  assign n20452 = n14702 & n20451 ;
  assign n20448 = n10970 ^ n8255 ^ 1'b0 ;
  assign n20449 = n9644 | n20448 ;
  assign n20453 = n20452 ^ n20449 ^ 1'b0 ;
  assign n20455 = n20454 ^ n20453 ^ 1'b0 ;
  assign n20456 = n20455 ^ x4 ^ 1'b0 ;
  assign n20457 = n8342 & n9973 ;
  assign n20458 = ( ~n11409 & n13422 ) | ( ~n11409 & n20457 ) | ( n13422 & n20457 ) ;
  assign n20459 = n20458 ^ n9647 ^ n6778 ;
  assign n20460 = n10172 & ~n20351 ;
  assign n20461 = n20460 ^ n10762 ^ 1'b0 ;
  assign n20462 = n6560 ^ n1532 ^ 1'b0 ;
  assign n20463 = n5926 & ~n20462 ;
  assign n20464 = n4264 & n20463 ;
  assign n20465 = n5607 & ~n18644 ;
  assign n20466 = ~n8901 & n20465 ;
  assign n20467 = n3589 & n14594 ;
  assign n20468 = n5868 ^ n3789 ^ n1791 ;
  assign n20469 = n2304 & ~n20468 ;
  assign n20470 = n20469 ^ n6068 ^ 1'b0 ;
  assign n20471 = n20467 & n20470 ;
  assign n20472 = x61 & ~n4227 ;
  assign n20473 = n1271 & n20472 ;
  assign n20474 = n20471 | n20473 ;
  assign n20475 = ( n1603 & n11063 ) | ( n1603 & n20474 ) | ( n11063 & n20474 ) ;
  assign n20476 = n2944 ^ n2823 ^ 1'b0 ;
  assign n20477 = ( n7687 & n14364 ) | ( n7687 & n20476 ) | ( n14364 & n20476 ) ;
  assign n20478 = n6420 & n12367 ;
  assign n20479 = ( ~n319 & n4142 ) | ( ~n319 & n17287 ) | ( n4142 & n17287 ) ;
  assign n20484 = n1777 | n12628 ;
  assign n20485 = n12628 & ~n20484 ;
  assign n20486 = n5517 | n20485 ;
  assign n20480 = n148 | n2540 ;
  assign n20481 = n2540 & ~n20480 ;
  assign n20482 = n15319 & ~n20481 ;
  assign n20483 = n1222 & ~n20482 ;
  assign n20487 = n20486 ^ n20483 ^ 1'b0 ;
  assign n20488 = n9778 & ~n20487 ;
  assign n20489 = n13087 ^ n11851 ^ 1'b0 ;
  assign n20490 = n1383 & n20489 ;
  assign n20491 = n11215 & n20490 ;
  assign n20492 = n3763 | n12588 ;
  assign n20493 = n15546 | n20492 ;
  assign n20494 = n15112 ^ n353 ^ 1'b0 ;
  assign n20495 = n13663 & ~n14957 ;
  assign n20496 = n13953 & ~n20495 ;
  assign n20497 = ( n1312 & n4341 ) | ( n1312 & ~n9005 ) | ( n4341 & ~n9005 ) ;
  assign n20498 = n11088 & ~n20497 ;
  assign n20499 = ~n8528 & n20498 ;
  assign n20502 = n7052 ^ x71 ^ 1'b0 ;
  assign n20503 = ~n19143 & n20502 ;
  assign n20500 = n451 | n4253 ;
  assign n20501 = n3589 & ~n20500 ;
  assign n20504 = n20503 ^ n20501 ^ n11499 ;
  assign n20505 = n10014 ^ n6114 ^ n5349 ;
  assign n20506 = n6001 & ~n19624 ;
  assign n20507 = ~n16371 & n20506 ;
  assign n20508 = n2976 ^ n1276 ^ n1036 ;
  assign n20509 = n11927 & ~n20508 ;
  assign n20510 = n1170 ^ n950 ^ 1'b0 ;
  assign n20511 = ( ~n3255 & n5525 ) | ( ~n3255 & n20510 ) | ( n5525 & n20510 ) ;
  assign n20512 = n20511 ^ n11879 ^ 1'b0 ;
  assign n20513 = n4632 & ~n20512 ;
  assign n20514 = n8058 & ~n10423 ;
  assign n20515 = ~n20513 & n20514 ;
  assign n20516 = ( n7246 & n20509 ) | ( n7246 & n20515 ) | ( n20509 & n20515 ) ;
  assign n20517 = n8507 | n20516 ;
  assign n20518 = n6971 ^ n2506 ^ 1'b0 ;
  assign n20519 = n19394 & n20518 ;
  assign n20520 = n11645 ^ n7938 ^ 1'b0 ;
  assign n20521 = n19680 & n20520 ;
  assign n20522 = n925 | n16073 ;
  assign n20523 = n798 & ~n20522 ;
  assign n20524 = n18390 | n20523 ;
  assign n20525 = n4574 ^ n1839 ^ x77 ;
  assign n20526 = n9359 & n20525 ;
  assign n20527 = ( n962 & ~n14234 ) | ( n962 & n20526 ) | ( ~n14234 & n20526 ) ;
  assign n20528 = ( n8695 & n11370 ) | ( n8695 & ~n20527 ) | ( n11370 & ~n20527 ) ;
  assign n20529 = n19057 ^ n9501 ^ 1'b0 ;
  assign n20530 = n1880 | n6340 ;
  assign n20531 = ~n499 & n20530 ;
  assign n20536 = n4139 | n16294 ;
  assign n20537 = n12803 & ~n20536 ;
  assign n20532 = n4029 & n10296 ;
  assign n20533 = n438 & n20532 ;
  assign n20534 = n20533 ^ n13045 ^ 1'b0 ;
  assign n20535 = n13088 | n20534 ;
  assign n20538 = n20537 ^ n20535 ^ 1'b0 ;
  assign n20539 = n7076 ^ n145 ^ 1'b0 ;
  assign n20540 = n9113 & n20539 ;
  assign n20541 = n18193 ^ n6632 ^ n5364 ;
  assign n20542 = ~n10598 & n20541 ;
  assign n20543 = ~n20540 & n20542 ;
  assign n20545 = ( n2158 & n7598 ) | ( n2158 & ~n8623 ) | ( n7598 & ~n8623 ) ;
  assign n20546 = n20545 ^ n5177 ^ 1'b0 ;
  assign n20544 = ( n4103 & n6163 ) | ( n4103 & ~n11954 ) | ( n6163 & ~n11954 ) ;
  assign n20547 = n20546 ^ n20544 ^ n16857 ;
  assign n20548 = ( n4699 & n12336 ) | ( n4699 & ~n13446 ) | ( n12336 & ~n13446 ) ;
  assign n20549 = ~n3414 & n9969 ;
  assign n20550 = n20548 | n20549 ;
  assign n20551 = n16926 ^ n6256 ^ n3658 ;
  assign n20552 = ~n12563 & n20551 ;
  assign n20553 = n13928 & ~n16733 ;
  assign n20554 = n20552 & n20553 ;
  assign n20555 = n6765 ^ n4211 ^ 1'b0 ;
  assign n20556 = n4426 | n15626 ;
  assign n20557 = n20555 & ~n20556 ;
  assign n20558 = n5965 & ~n20393 ;
  assign n20559 = n20558 ^ n13889 ^ n12507 ;
  assign n20560 = n20080 ^ n725 ^ 1'b0 ;
  assign n20561 = n5278 & n20560 ;
  assign n20562 = n2215 | n17089 ;
  assign n20563 = x39 & ~n9469 ;
  assign n20564 = n20563 ^ n20415 ^ 1'b0 ;
  assign n20565 = n20564 ^ n7168 ^ 1'b0 ;
  assign n20566 = ~n18361 & n20565 ;
  assign n20567 = n11879 ^ n10653 ^ 1'b0 ;
  assign n20568 = ~n7530 & n20567 ;
  assign n20569 = n1881 & ~n11454 ;
  assign n20570 = ~n8744 & n20569 ;
  assign n20571 = n20570 ^ n8916 ^ 1'b0 ;
  assign n20572 = ~n9234 & n20571 ;
  assign n20573 = n20572 ^ n5320 ^ n1640 ;
  assign n20574 = n20568 & n20573 ;
  assign n20575 = ~n13696 & n17308 ;
  assign n20576 = n3845 | n20575 ;
  assign n20577 = n8823 & ~n20576 ;
  assign n20578 = n6772 & ~n20577 ;
  assign n20579 = n3756 & n20578 ;
  assign n20580 = ~n10421 & n12282 ;
  assign n20581 = n11711 ^ n2496 ^ 1'b0 ;
  assign n20582 = n18837 & ~n20581 ;
  assign n20583 = n1441 & n16401 ;
  assign n20584 = ~n20582 & n20583 ;
  assign n20585 = n18019 ^ n13789 ^ 1'b0 ;
  assign n20586 = n20585 ^ n9523 ^ n2419 ;
  assign n20587 = ~n800 & n8382 ;
  assign n20588 = n4146 & n20587 ;
  assign n20589 = n20588 ^ n2331 ^ n1575 ;
  assign n20590 = n18703 ^ n16832 ^ n13422 ;
  assign n20591 = n7790 & ~n12852 ;
  assign n20592 = ~n525 & n18963 ;
  assign n20593 = n20592 ^ n8487 ^ 1'b0 ;
  assign n20594 = n6007 ^ n1389 ^ 1'b0 ;
  assign n20595 = ~n20593 & n20594 ;
  assign n20596 = n14326 ^ n9879 ^ 1'b0 ;
  assign n20597 = n20595 & n20596 ;
  assign n20598 = n2909 ^ n935 ^ 1'b0 ;
  assign n20599 = n14782 & ~n20598 ;
  assign n20600 = n10849 & n20599 ;
  assign n20601 = n8980 ^ n6404 ^ 1'b0 ;
  assign n20602 = n11432 ^ n2930 ^ 1'b0 ;
  assign n20603 = ~n7256 & n20602 ;
  assign n20604 = n19085 & n20603 ;
  assign n20605 = n20604 ^ n15678 ^ 1'b0 ;
  assign n20606 = n8231 ^ n2120 ^ 1'b0 ;
  assign n20607 = n10241 & n20606 ;
  assign n20610 = n5654 ^ n4971 ^ 1'b0 ;
  assign n20611 = n13351 & ~n20610 ;
  assign n20612 = ( n1660 & n6661 ) | ( n1660 & n20611 ) | ( n6661 & n20611 ) ;
  assign n20608 = ~n7241 & n20201 ;
  assign n20609 = n20608 ^ n9099 ^ 1'b0 ;
  assign n20613 = n20612 ^ n20609 ^ 1'b0 ;
  assign n20614 = ( n974 & ~n4216 ) | ( n974 & n9358 ) | ( ~n4216 & n9358 ) ;
  assign n20615 = ~n20613 & n20614 ;
  assign n20616 = n2898 | n7027 ;
  assign n20617 = n15133 & n20616 ;
  assign n20618 = ( ~n9625 & n11440 ) | ( ~n9625 & n19514 ) | ( n11440 & n19514 ) ;
  assign n20619 = n1960 | n20618 ;
  assign n20620 = n16992 ^ n12516 ^ n9242 ;
  assign n20621 = n20620 ^ n7557 ^ 1'b0 ;
  assign n20622 = n14598 ^ n7514 ^ n4459 ;
  assign n20623 = n7984 ^ n1101 ^ 1'b0 ;
  assign n20624 = n20623 ^ n8590 ^ n413 ;
  assign n20625 = n2609 & ~n6550 ;
  assign n20626 = n20625 ^ n15499 ^ 1'b0 ;
  assign n20627 = ~n4863 & n18457 ;
  assign n20628 = n3240 & ~n14994 ;
  assign n20629 = n20628 ^ n15436 ^ n12118 ;
  assign n20630 = n8799 ^ n6803 ^ n1008 ;
  assign n20631 = n5242 ^ n969 ^ 1'b0 ;
  assign n20632 = ~n15176 & n20631 ;
  assign n20633 = n6249 & ~n7047 ;
  assign n20634 = n20633 ^ n5537 ^ 1'b0 ;
  assign n20635 = n15966 ^ n3278 ^ 1'b0 ;
  assign n20636 = n3239 | n12250 ;
  assign n20637 = n20636 ^ n11207 ^ 1'b0 ;
  assign n20638 = ~n2278 & n12593 ;
  assign n20641 = n13112 ^ n8484 ^ 1'b0 ;
  assign n20639 = n16219 ^ n15321 ^ 1'b0 ;
  assign n20640 = n20639 ^ n11947 ^ n7226 ;
  assign n20642 = n20641 ^ n20640 ^ 1'b0 ;
  assign n20645 = n7612 ^ n6308 ^ 1'b0 ;
  assign n20646 = n11177 & n20645 ;
  assign n20643 = n14697 & ~n19430 ;
  assign n20644 = ( ~n9704 & n12414 ) | ( ~n9704 & n20643 ) | ( n12414 & n20643 ) ;
  assign n20647 = n20646 ^ n20644 ^ 1'b0 ;
  assign n20648 = n12959 | n20647 ;
  assign n20649 = n7270 & n10072 ;
  assign n20650 = n20649 ^ n18733 ^ 1'b0 ;
  assign n20651 = n20650 ^ n286 ^ 1'b0 ;
  assign n20652 = n14357 | n20651 ;
  assign n20653 = n11620 ^ n7502 ^ 1'b0 ;
  assign n20654 = ~n10220 & n20653 ;
  assign n20655 = n1326 & n3830 ;
  assign n20656 = n20655 ^ n11527 ^ n8392 ;
  assign n20657 = n14669 & n20656 ;
  assign n20658 = n13052 ^ n4507 ^ n1025 ;
  assign n20659 = ( n3821 & n17730 ) | ( n3821 & ~n19864 ) | ( n17730 & ~n19864 ) ;
  assign n20660 = n4708 & n16157 ;
  assign n20665 = n16224 ^ n16222 ^ 1'b0 ;
  assign n20661 = n522 & ~n992 ;
  assign n20662 = n10119 & n16393 ;
  assign n20663 = ~n18990 & n20662 ;
  assign n20664 = n20661 & ~n20663 ;
  assign n20666 = n20665 ^ n20664 ^ 1'b0 ;
  assign n20667 = n3729 ^ n2404 ^ 1'b0 ;
  assign n20668 = n20667 ^ n3121 ^ 1'b0 ;
  assign n20670 = n6497 ^ n190 ^ 1'b0 ;
  assign n20671 = n14201 & ~n20670 ;
  assign n20669 = n12414 ^ n11767 ^ n6901 ;
  assign n20672 = n20671 ^ n20669 ^ 1'b0 ;
  assign n20673 = n20668 & n20672 ;
  assign n20674 = n7393 ^ n2939 ^ n1113 ;
  assign n20675 = n8156 | n12714 ;
  assign n20676 = ( ~n9535 & n20674 ) | ( ~n9535 & n20675 ) | ( n20674 & n20675 ) ;
  assign n20677 = n2760 & n20676 ;
  assign n20678 = n15896 & n20677 ;
  assign n20679 = ( ~n629 & n8644 ) | ( ~n629 & n14311 ) | ( n8644 & n14311 ) ;
  assign n20682 = n140 & ~n4201 ;
  assign n20683 = n893 & n20682 ;
  assign n20680 = ~n3622 & n4154 ;
  assign n20681 = n20680 ^ n7091 ^ 1'b0 ;
  assign n20684 = n20683 ^ n20681 ^ n9260 ;
  assign n20685 = n4073 ^ n313 ^ 1'b0 ;
  assign n20686 = n4538 | n13961 ;
  assign n20687 = n13075 & ~n13342 ;
  assign n20688 = n13083 ^ n3488 ^ 1'b0 ;
  assign n20689 = n2813 & n20688 ;
  assign n20690 = n11095 & n11688 ;
  assign n20692 = n1481 | n4792 ;
  assign n20693 = n20692 ^ n9775 ^ 1'b0 ;
  assign n20691 = n13133 ^ n11565 ^ 1'b0 ;
  assign n20694 = n20693 ^ n20691 ^ 1'b0 ;
  assign n20695 = n20690 | n20694 ;
  assign n20696 = n2297 & ~n14300 ;
  assign n20697 = ~n5773 & n20696 ;
  assign n20698 = n17523 ^ n5539 ^ n4664 ;
  assign n20699 = ( n603 & ~n4057 ) | ( n603 & n4346 ) | ( ~n4057 & n4346 ) ;
  assign n20700 = n20699 ^ n11676 ^ n11489 ;
  assign n20701 = ( n18479 & n20698 ) | ( n18479 & n20700 ) | ( n20698 & n20700 ) ;
  assign n20702 = n9862 ^ n9806 ^ n2344 ;
  assign n20703 = n9880 & ~n20702 ;
  assign n20704 = n20703 ^ n8383 ^ 1'b0 ;
  assign n20705 = ( ~n11459 & n11915 ) | ( ~n11459 & n20704 ) | ( n11915 & n20704 ) ;
  assign n20706 = ( n6698 & n8179 ) | ( n6698 & ~n17685 ) | ( n8179 & ~n17685 ) ;
  assign n20707 = n18419 & n20706 ;
  assign n20708 = ~n4197 & n17347 ;
  assign n20709 = ( n3844 & n4852 ) | ( n3844 & n10605 ) | ( n4852 & n10605 ) ;
  assign n20711 = n16085 ^ n4652 ^ 1'b0 ;
  assign n20710 = n4934 ^ n3083 ^ 1'b0 ;
  assign n20712 = n20711 ^ n20710 ^ n17901 ;
  assign n20713 = n12020 & n20712 ;
  assign n20714 = n296 | n17341 ;
  assign n20715 = n20714 ^ n16375 ^ 1'b0 ;
  assign n20716 = n12098 ^ n7406 ^ 1'b0 ;
  assign n20722 = n16224 ^ n187 ^ 1'b0 ;
  assign n20723 = n657 & n2687 ;
  assign n20724 = ~n20722 & n20723 ;
  assign n20720 = n1435 ^ n1318 ^ 1'b0 ;
  assign n20721 = n20720 ^ n12029 ^ 1'b0 ;
  assign n20717 = n5621 ^ n4078 ^ 1'b0 ;
  assign n20718 = n2143 & ~n20717 ;
  assign n20719 = n20718 ^ n2991 ^ 1'b0 ;
  assign n20725 = n20724 ^ n20721 ^ n20719 ;
  assign n20726 = n6289 ^ n4706 ^ 1'b0 ;
  assign n20727 = n5673 & ~n7219 ;
  assign n20728 = n20727 ^ n4051 ^ 1'b0 ;
  assign n20729 = n2957 & ~n3964 ;
  assign n20730 = ( n5639 & ~n15437 ) | ( n5639 & n20729 ) | ( ~n15437 & n20729 ) ;
  assign n20731 = ~n7869 & n10125 ;
  assign n20732 = n20731 ^ n9084 ^ 1'b0 ;
  assign n20733 = n18880 ^ n15420 ^ 1'b0 ;
  assign n20734 = n20732 & ~n20733 ;
  assign n20735 = n391 | n13584 ;
  assign n20736 = n20735 ^ n6281 ^ 1'b0 ;
  assign n20737 = x120 & n13061 ;
  assign n20738 = n20737 ^ n475 ^ 1'b0 ;
  assign n20739 = ( n15769 & n19702 ) | ( n15769 & ~n20738 ) | ( n19702 & ~n20738 ) ;
  assign n20740 = n3300 & ~n20739 ;
  assign n20741 = n20740 ^ n7916 ^ 1'b0 ;
  assign n20742 = n8050 ^ n5007 ^ 1'b0 ;
  assign n20743 = n2105 | n20742 ;
  assign n20744 = ( n2897 & ~n8184 ) | ( n2897 & n15710 ) | ( ~n8184 & n15710 ) ;
  assign n20745 = ~n8809 & n10446 ;
  assign n20746 = n411 & ~n20745 ;
  assign n20747 = n20746 ^ n2534 ^ 1'b0 ;
  assign n20748 = ( n4665 & n5227 ) | ( n4665 & n15684 ) | ( n5227 & n15684 ) ;
  assign n20749 = n6974 ^ n4483 ^ 1'b0 ;
  assign n20750 = n9034 | n18945 ;
  assign n20751 = n20749 & ~n20750 ;
  assign n20752 = n6110 ^ n2034 ^ n1069 ;
  assign n20753 = n20752 ^ n15614 ^ 1'b0 ;
  assign n20754 = n19820 | n20753 ;
  assign n20755 = n20754 ^ n16384 ^ 1'b0 ;
  assign n20756 = n19347 ^ n13615 ^ n10462 ;
  assign n20757 = ( ~n2595 & n5882 ) | ( ~n2595 & n11854 ) | ( n5882 & n11854 ) ;
  assign n20758 = n15388 ^ n3414 ^ 1'b0 ;
  assign n20759 = ~n2551 & n15893 ;
  assign n20760 = ~n20758 & n20759 ;
  assign n20761 = n20760 ^ n1175 ^ 1'b0 ;
  assign n20762 = n20757 | n20761 ;
  assign n20763 = n20762 ^ n9670 ^ 1'b0 ;
  assign n20764 = n886 | n5776 ;
  assign n20765 = n20764 ^ x100 ^ 1'b0 ;
  assign n20767 = n14858 ^ n3343 ^ 1'b0 ;
  assign n20766 = n14101 & ~n14631 ;
  assign n20768 = n20767 ^ n20766 ^ 1'b0 ;
  assign n20769 = ~n13566 & n20768 ;
  assign n20770 = ~n20427 & n20769 ;
  assign n20771 = n13795 ^ n345 ^ 1'b0 ;
  assign n20772 = n1159 & ~n1748 ;
  assign n20773 = n1146 ^ n374 ^ 1'b0 ;
  assign n20774 = n1181 & n20773 ;
  assign n20775 = n6818 ^ n1066 ^ 1'b0 ;
  assign n20776 = ( n20772 & n20774 ) | ( n20772 & n20775 ) | ( n20774 & n20775 ) ;
  assign n20777 = n12861 ^ n8759 ^ 1'b0 ;
  assign n20778 = n6239 ^ n5274 ^ n3582 ;
  assign n20779 = n20777 | n20778 ;
  assign n20780 = ( n1470 & n10407 ) | ( n1470 & ~n12306 ) | ( n10407 & ~n12306 ) ;
  assign n20781 = n15299 ^ n5355 ^ 1'b0 ;
  assign n20782 = ~n7166 & n20781 ;
  assign n20783 = n20782 ^ n11689 ^ n9434 ;
  assign n20784 = n10706 & n12277 ;
  assign n20785 = n4753 ^ n2366 ^ 1'b0 ;
  assign n20786 = n3012 | n20785 ;
  assign n20787 = ( ~x103 & n4357 ) | ( ~x103 & n9211 ) | ( n4357 & n9211 ) ;
  assign n20788 = n20787 ^ n1427 ^ n1126 ;
  assign n20789 = n584 | n20788 ;
  assign n20790 = n8129 & ~n20789 ;
  assign n20791 = n16002 & ~n16317 ;
  assign n20792 = n20791 ^ n18043 ^ 1'b0 ;
  assign n20793 = n13546 ^ n1351 ^ 1'b0 ;
  assign n20794 = n5802 & n20793 ;
  assign n20795 = n2976 ^ n2138 ^ 1'b0 ;
  assign n20796 = ~n10423 & n20795 ;
  assign n20797 = ( n11097 & n11412 ) | ( n11097 & ~n20796 ) | ( n11412 & ~n20796 ) ;
  assign n20798 = ( n1132 & n8380 ) | ( n1132 & n8890 ) | ( n8380 & n8890 ) ;
  assign n20799 = ~n18269 & n20798 ;
  assign n20800 = ( n540 & n16242 ) | ( n540 & ~n20799 ) | ( n16242 & ~n20799 ) ;
  assign n20801 = n10692 & ~n12095 ;
  assign n20802 = n20801 ^ n8332 ^ 1'b0 ;
  assign n20803 = n4216 & n10049 ;
  assign n20804 = n20803 ^ n2515 ^ 1'b0 ;
  assign n20805 = n6969 ^ n6571 ^ 1'b0 ;
  assign n20806 = n9712 & n20805 ;
  assign n20807 = n1537 & ~n3925 ;
  assign n20808 = n9571 & n20807 ;
  assign n20809 = n10234 | n10687 ;
  assign n20810 = ~n1199 & n5530 ;
  assign n20811 = ( ~n16665 & n20809 ) | ( ~n16665 & n20810 ) | ( n20809 & n20810 ) ;
  assign n20812 = n3832 | n13752 ;
  assign n20813 = n5418 ^ n4084 ^ 1'b0 ;
  assign n20814 = n3524 & n20813 ;
  assign n20815 = n12062 ^ n4121 ^ n1306 ;
  assign n20816 = ~n20814 & n20815 ;
  assign n20817 = n20724 & n20816 ;
  assign n20818 = n2008 & ~n17171 ;
  assign n20819 = n20818 ^ n7744 ^ 1'b0 ;
  assign n20820 = ( n3873 & n9599 ) | ( n3873 & n20819 ) | ( n9599 & n20819 ) ;
  assign n20821 = n1515 & ~n20820 ;
  assign n20822 = n20821 ^ n18233 ^ 1'b0 ;
  assign n20823 = ~n3776 & n6157 ;
  assign n20824 = ~n9349 & n20823 ;
  assign n20825 = n5793 & ~n20824 ;
  assign n20826 = ( ~n8272 & n13754 ) | ( ~n8272 & n14967 ) | ( n13754 & n14967 ) ;
  assign n20827 = ( ~n1216 & n3522 ) | ( ~n1216 & n20826 ) | ( n3522 & n20826 ) ;
  assign n20828 = n5050 | n8571 ;
  assign n20829 = n20827 | n20828 ;
  assign n20830 = n19844 ^ n13545 ^ 1'b0 ;
  assign n20831 = n3076 & ~n16211 ;
  assign n20832 = n20831 ^ n14667 ^ 1'b0 ;
  assign n20833 = ( n820 & n7829 ) | ( n820 & n11500 ) | ( n7829 & n11500 ) ;
  assign n20834 = n20833 ^ n726 ^ 1'b0 ;
  assign n20835 = n3658 | n20834 ;
  assign n20836 = ~n1354 & n3393 ;
  assign n20837 = n2449 & n8271 ;
  assign n20838 = n20836 & n20837 ;
  assign n20839 = n7226 & ~n20838 ;
  assign n20840 = n20839 ^ n221 ^ 1'b0 ;
  assign n20841 = n413 & ~n20840 ;
  assign n20844 = n14288 ^ n8702 ^ n4407 ;
  assign n20842 = ( n557 & ~n1314 ) | ( n557 & n15836 ) | ( ~n1314 & n15836 ) ;
  assign n20843 = n18514 & ~n20842 ;
  assign n20845 = n20844 ^ n20843 ^ 1'b0 ;
  assign n20846 = n12542 ^ n8709 ^ 1'b0 ;
  assign n20847 = n14754 & ~n20846 ;
  assign n20848 = n20847 ^ n4897 ^ 1'b0 ;
  assign n20849 = n3482 | n15835 ;
  assign n20850 = n194 | n20849 ;
  assign n20851 = n4447 & ~n20850 ;
  assign n20852 = n8863 ^ n3241 ^ n1345 ;
  assign n20853 = ( ~n6556 & n20851 ) | ( ~n6556 & n20852 ) | ( n20851 & n20852 ) ;
  assign n20854 = n6570 & n14158 ;
  assign n20855 = n20854 ^ n6702 ^ n1273 ;
  assign n20856 = ~n17994 & n18429 ;
  assign n20857 = ~n18128 & n20856 ;
  assign n20858 = ( n8108 & n8585 ) | ( n8108 & ~n16632 ) | ( n8585 & ~n16632 ) ;
  assign n20859 = n20858 ^ n10432 ^ 1'b0 ;
  assign n20860 = ~n1905 & n2815 ;
  assign n20861 = ( n4295 & n6513 ) | ( n4295 & n20860 ) | ( n6513 & n20860 ) ;
  assign n20862 = n6895 & ~n12467 ;
  assign n20863 = n7535 & ~n20862 ;
  assign n20864 = n20861 & n20863 ;
  assign n20868 = n6053 | n12672 ;
  assign n20869 = n14016 | n20868 ;
  assign n20865 = n6438 ^ n3820 ^ n3265 ;
  assign n20866 = n13438 & ~n20865 ;
  assign n20867 = n14973 & n20866 ;
  assign n20870 = n20869 ^ n20867 ^ 1'b0 ;
  assign n20871 = n9772 ^ n8988 ^ 1'b0 ;
  assign n20872 = ~n14855 & n20871 ;
  assign n20873 = n3228 ^ n2884 ^ n2717 ;
  assign n20874 = n14166 | n20873 ;
  assign n20875 = n20874 ^ n15629 ^ n11155 ;
  assign n20876 = n15898 ^ n11719 ^ n7490 ;
  assign n20877 = n6723 | n9418 ;
  assign n20878 = n11410 & n19187 ;
  assign n20879 = n20877 & n20878 ;
  assign n20880 = n20879 ^ n2400 ^ 1'b0 ;
  assign n20881 = ~n7432 & n13673 ;
  assign n20882 = n20881 ^ n6880 ^ 1'b0 ;
  assign n20886 = n2781 & ~n7977 ;
  assign n20884 = n3215 | n17061 ;
  assign n20883 = n11979 ^ n10592 ^ 1'b0 ;
  assign n20885 = n20884 ^ n20883 ^ n13767 ;
  assign n20887 = n20886 ^ n20885 ^ n5322 ;
  assign n20888 = n11730 & n20887 ;
  assign n20889 = n10756 ^ n4592 ^ 1'b0 ;
  assign n20890 = ~n1269 & n20889 ;
  assign n20891 = n20890 ^ n8212 ^ n7284 ;
  assign n20892 = n3684 | n20891 ;
  assign n20893 = n6733 | n6749 ;
  assign n20894 = n6632 & ~n8151 ;
  assign n20895 = n12825 | n20894 ;
  assign n20896 = n3541 | n9925 ;
  assign n20897 = n20896 ^ n1388 ^ 1'b0 ;
  assign n20898 = n20422 ^ n915 ^ 1'b0 ;
  assign n20899 = n1104 & n8199 ;
  assign n20900 = n20899 ^ n18530 ^ 1'b0 ;
  assign n20901 = ( n2306 & ~n2913 ) | ( n2306 & n5281 ) | ( ~n2913 & n5281 ) ;
  assign n20902 = ( n1908 & ~n5046 ) | ( n1908 & n18976 ) | ( ~n5046 & n18976 ) ;
  assign n20903 = n14341 ^ n12590 ^ n319 ;
  assign n20904 = n1311 ^ n474 ^ 1'b0 ;
  assign n20905 = n20904 ^ n12405 ^ 1'b0 ;
  assign n20906 = n3820 ^ n2265 ^ 1'b0 ;
  assign n20907 = n2186 ^ n1647 ^ 1'b0 ;
  assign n20908 = n20907 ^ n3323 ^ 1'b0 ;
  assign n20909 = n6731 ^ n5430 ^ 1'b0 ;
  assign n20910 = n20909 ^ n20103 ^ n6994 ;
  assign n20911 = ~n843 & n1690 ;
  assign n20912 = n20911 ^ n4495 ^ 1'b0 ;
  assign n20913 = n20912 ^ n9448 ^ n3964 ;
  assign n20914 = n14920 | n20913 ;
  assign n20915 = n20914 ^ n11129 ^ 1'b0 ;
  assign n20916 = ( n1725 & n7697 ) | ( n1725 & n20915 ) | ( n7697 & n20915 ) ;
  assign n20917 = n13868 ^ n3707 ^ 1'b0 ;
  assign n20918 = n7649 ^ n6367 ^ n2650 ;
  assign n20919 = n20918 ^ n13138 ^ n2601 ;
  assign n20920 = n13937 ^ n8608 ^ 1'b0 ;
  assign n20921 = n20919 & ~n20920 ;
  assign n20922 = x30 | n1253 ;
  assign n20923 = ~n2224 & n2293 ;
  assign n20924 = n20923 ^ n19627 ^ 1'b0 ;
  assign n20925 = n13750 ^ n9131 ^ 1'b0 ;
  assign n20926 = ~n18943 & n19831 ;
  assign n20927 = ~n15135 & n20926 ;
  assign n20928 = n14404 ^ n10674 ^ n4132 ;
  assign n20929 = n9583 & ~n19047 ;
  assign n20930 = n9259 ^ n1476 ^ 1'b0 ;
  assign n20931 = ~n16531 & n20930 ;
  assign n20932 = n20707 ^ n9664 ^ n4495 ;
  assign n20933 = ( n3242 & ~n4454 ) | ( n3242 & n7036 ) | ( ~n4454 & n7036 ) ;
  assign n20934 = n16452 ^ n13160 ^ 1'b0 ;
  assign n20935 = ~n12744 & n20934 ;
  assign n20936 = n10173 & n10978 ;
  assign n20937 = n20936 ^ n15504 ^ 1'b0 ;
  assign n20938 = ~n17994 & n20937 ;
  assign n20939 = n4656 ^ n4274 ^ n401 ;
  assign n20940 = n20939 ^ n15150 ^ n9655 ;
  assign n20941 = n20938 & n20940 ;
  assign n20942 = n1145 & ~n12203 ;
  assign n20943 = n10752 | n20942 ;
  assign n20944 = n1141 & ~n20943 ;
  assign n20945 = n20944 ^ n9682 ^ n7383 ;
  assign n20946 = n2763 | n5308 ;
  assign n20947 = n20946 ^ n16462 ^ 1'b0 ;
  assign n20948 = n1342 ^ n1124 ^ 1'b0 ;
  assign n20949 = n14078 & ~n20948 ;
  assign n20950 = n20949 ^ n3303 ^ 1'b0 ;
  assign n20951 = n4756 & ~n20950 ;
  assign n20952 = n9903 & ~n17794 ;
  assign n20956 = n4714 ^ n1996 ^ 1'b0 ;
  assign n20957 = ~n10031 & n20956 ;
  assign n20953 = n9367 ^ n719 ^ 1'b0 ;
  assign n20954 = ~n9427 & n20953 ;
  assign n20955 = ~n2074 & n20954 ;
  assign n20958 = n20957 ^ n20955 ^ 1'b0 ;
  assign n20959 = ( n12242 & ~n15222 ) | ( n12242 & n20958 ) | ( ~n15222 & n20958 ) ;
  assign n20960 = n8686 ^ n6649 ^ n5274 ;
  assign n20961 = n12897 ^ n7105 ^ 1'b0 ;
  assign n20962 = n4554 | n20961 ;
  assign n20963 = ( n3954 & n7706 ) | ( n3954 & ~n20962 ) | ( n7706 & ~n20962 ) ;
  assign n20964 = n16401 ^ n12881 ^ n3718 ;
  assign n20965 = ~n6884 & n19926 ;
  assign n20966 = n20965 ^ n2089 ^ 1'b0 ;
  assign n20967 = n20966 ^ x9 ^ 1'b0 ;
  assign n20968 = n8861 ^ n1631 ^ 1'b0 ;
  assign n20969 = n2265 | n20968 ;
  assign n20970 = n9190 & ~n20969 ;
  assign n20971 = n20970 ^ n6186 ^ 1'b0 ;
  assign n20972 = n17123 & n20971 ;
  assign n20973 = n3016 ^ n2448 ^ 1'b0 ;
  assign n20974 = n1713 | n20973 ;
  assign n20975 = n17449 & n19934 ;
  assign n20976 = n9619 ^ n5306 ^ 1'b0 ;
  assign n20977 = ~n5467 & n20976 ;
  assign n20978 = n4805 & n20977 ;
  assign n20980 = ~n2196 & n8839 ;
  assign n20981 = n20980 ^ x98 ^ 1'b0 ;
  assign n20982 = n11440 & ~n20981 ;
  assign n20979 = n16405 ^ n12537 ^ n6237 ;
  assign n20983 = n20982 ^ n20979 ^ n2658 ;
  assign n20984 = n18766 ^ n11651 ^ 1'b0 ;
  assign n20985 = n1146 | n7984 ;
  assign n20986 = n20985 ^ n2931 ^ 1'b0 ;
  assign n20987 = n15794 ^ n11743 ^ n7481 ;
  assign n20988 = n20986 | n20987 ;
  assign n20989 = n5643 | n7156 ;
  assign n20990 = n12350 & ~n20989 ;
  assign n20991 = n20990 ^ n9020 ^ 1'b0 ;
  assign n20992 = n7930 ^ n4043 ^ 1'b0 ;
  assign n20993 = ~n20991 & n20992 ;
  assign n20994 = n17900 ^ n17055 ^ 1'b0 ;
  assign n20995 = n9595 | n20994 ;
  assign n20996 = n20995 ^ n303 ^ 1'b0 ;
  assign n20997 = ~n6447 & n19397 ;
  assign n20998 = n20997 ^ n17955 ^ 1'b0 ;
  assign n20999 = ~n3386 & n5586 ;
  assign n21000 = n20999 ^ n7121 ^ 1'b0 ;
  assign n21001 = n21000 ^ n20024 ^ n3459 ;
  assign n21002 = n9970 | n11548 ;
  assign n21003 = n21002 ^ n11165 ^ 1'b0 ;
  assign n21004 = n21003 ^ n14137 ^ x55 ;
  assign n21005 = n2785 & ~n9794 ;
  assign n21006 = n21005 ^ n20191 ^ 1'b0 ;
  assign n21007 = n2592 & ~n8572 ;
  assign n21008 = ~n21006 & n21007 ;
  assign n21011 = ~n2002 & n10775 ;
  assign n21012 = n1246 & n21011 ;
  assign n21013 = n21012 ^ n9561 ^ 1'b0 ;
  assign n21014 = n11151 | n21013 ;
  assign n21009 = n11524 ^ n11086 ^ 1'b0 ;
  assign n21010 = ~n247 & n21009 ;
  assign n21015 = n21014 ^ n21010 ^ 1'b0 ;
  assign n21016 = n14449 & ~n19334 ;
  assign n21017 = n4404 | n21016 ;
  assign n21018 = n8687 | n21017 ;
  assign n21026 = n4135 ^ n3418 ^ 1'b0 ;
  assign n21027 = n3699 | n21026 ;
  assign n21020 = n5457 ^ n274 ^ 1'b0 ;
  assign n21021 = n8707 & n21020 ;
  assign n21022 = n16418 ^ n1581 ^ 1'b0 ;
  assign n21023 = n8161 & ~n21022 ;
  assign n21024 = ( n12568 & n21021 ) | ( n12568 & n21023 ) | ( n21021 & n21023 ) ;
  assign n21025 = n14709 & n21024 ;
  assign n21028 = n21027 ^ n21025 ^ 1'b0 ;
  assign n21029 = n21028 ^ n7422 ^ n2237 ;
  assign n21019 = n10433 & n14762 ;
  assign n21030 = n21029 ^ n21019 ^ 1'b0 ;
  assign n21031 = n20300 | n21004 ;
  assign n21032 = n18321 ^ n1470 ^ 1'b0 ;
  assign n21033 = n21032 ^ n20951 ^ 1'b0 ;
  assign n21034 = n1090 & ~n7873 ;
  assign n21035 = n21034 ^ n10527 ^ 1'b0 ;
  assign n21036 = n21035 ^ n9831 ^ n7270 ;
  assign n21037 = n18649 ^ n4068 ^ 1'b0 ;
  assign n21038 = n6396 | n21037 ;
  assign n21039 = ( n1049 & n3999 ) | ( n1049 & ~n11444 ) | ( n3999 & ~n11444 ) ;
  assign n21040 = ( n6260 & n13432 ) | ( n6260 & ~n21039 ) | ( n13432 & ~n21039 ) ;
  assign n21041 = n11549 ^ n9262 ^ 1'b0 ;
  assign n21042 = ~n11779 & n21041 ;
  assign n21043 = n21004 | n21042 ;
  assign n21044 = n16091 ^ n8626 ^ 1'b0 ;
  assign n21045 = ~n3612 & n15614 ;
  assign n21046 = n21045 ^ n6713 ^ 1'b0 ;
  assign n21047 = ( ~n413 & n1058 ) | ( ~n413 & n2870 ) | ( n1058 & n2870 ) ;
  assign n21048 = n21047 ^ n11882 ^ n1485 ;
  assign n21049 = n21048 ^ n9925 ^ 1'b0 ;
  assign n21050 = n1004 & n9557 ;
  assign n21051 = n21050 ^ n17248 ^ 1'b0 ;
  assign n21052 = n6761 ^ n4216 ^ 1'b0 ;
  assign n21053 = n6442 & ~n21052 ;
  assign n21054 = n21053 ^ n4077 ^ 1'b0 ;
  assign n21055 = n3937 & ~n6632 ;
  assign n21056 = n19457 ^ n14127 ^ n6985 ;
  assign n21057 = ( n12263 & ~n21055 ) | ( n12263 & n21056 ) | ( ~n21055 & n21056 ) ;
  assign n21058 = n18364 | n21057 ;
  assign n21059 = n21054 & ~n21058 ;
  assign n21060 = n7400 & n12372 ;
  assign n21061 = n10465 | n21060 ;
  assign n21062 = n21061 ^ n17264 ^ 1'b0 ;
  assign n21065 = n16125 ^ n4404 ^ 1'b0 ;
  assign n21063 = n334 & n11625 ;
  assign n21064 = n15854 & n21063 ;
  assign n21066 = n21065 ^ n21064 ^ 1'b0 ;
  assign n21067 = n2021 & n5865 ;
  assign n21068 = n3230 ^ n2578 ^ 1'b0 ;
  assign n21069 = ~n21067 & n21068 ;
  assign n21070 = n5281 | n18932 ;
  assign n21071 = n21069 | n21070 ;
  assign n21072 = n7281 ^ n5888 ^ 1'b0 ;
  assign n21073 = n13195 ^ n12016 ^ 1'b0 ;
  assign n21074 = ~n17888 & n19014 ;
  assign n21075 = n8487 & n21074 ;
  assign n21076 = n15493 ^ n15440 ^ 1'b0 ;
  assign n21077 = ~n20561 & n21076 ;
  assign n21078 = ~n251 & n21077 ;
  assign n21079 = n18889 ^ n663 ^ 1'b0 ;
  assign n21080 = n1577 & n15795 ;
  assign n21081 = n467 & ~n21080 ;
  assign n21082 = ( ~n7437 & n21079 ) | ( ~n7437 & n21081 ) | ( n21079 & n21081 ) ;
  assign n21083 = ( n1897 & ~n7877 ) | ( n1897 & n11055 ) | ( ~n7877 & n11055 ) ;
  assign n21084 = ( ~n1246 & n9607 ) | ( ~n1246 & n21083 ) | ( n9607 & n21083 ) ;
  assign n21085 = n14843 ^ n8786 ^ n3765 ;
  assign n21086 = n21085 ^ n5661 ^ 1'b0 ;
  assign n21087 = n14073 & n21086 ;
  assign n21089 = n14338 ^ n3549 ^ 1'b0 ;
  assign n21088 = n9685 | n13514 ;
  assign n21090 = n21089 ^ n21088 ^ n13974 ;
  assign n21091 = n2260 ^ n2117 ^ 1'b0 ;
  assign n21092 = ~n19506 & n21091 ;
  assign n21093 = ~n17182 & n21092 ;
  assign n21094 = ~n1388 & n4667 ;
  assign n21095 = n9304 & n21094 ;
  assign n21096 = n21095 ^ n4941 ^ 1'b0 ;
  assign n21097 = n21009 & ~n21096 ;
  assign n21098 = n2695 & n21097 ;
  assign n21099 = n5387 | n8231 ;
  assign n21100 = n21099 ^ n5654 ^ 1'b0 ;
  assign n21101 = n5899 & ~n21100 ;
  assign n21102 = ~n3566 & n21101 ;
  assign n21103 = n10651 & n21102 ;
  assign n21104 = n9973 ^ n8258 ^ 1'b0 ;
  assign n21105 = ( ~n1700 & n4161 ) | ( ~n1700 & n10881 ) | ( n4161 & n10881 ) ;
  assign n21106 = n21105 ^ n3267 ^ 1'b0 ;
  assign n21107 = n21106 ^ n15068 ^ n7837 ;
  assign n21108 = ( n3449 & ~n8153 ) | ( n3449 & n13665 ) | ( ~n8153 & n13665 ) ;
  assign n21109 = n12622 ^ n2324 ^ 1'b0 ;
  assign n21110 = n16648 & ~n21109 ;
  assign n21113 = n16595 ^ n9170 ^ 1'b0 ;
  assign n21114 = ( ~n12636 & n18280 ) | ( ~n12636 & n21113 ) | ( n18280 & n21113 ) ;
  assign n21111 = ~x0 & n6521 ;
  assign n21112 = n21111 ^ n13696 ^ 1'b0 ;
  assign n21115 = n21114 ^ n21112 ^ n4382 ;
  assign n21116 = n21115 ^ n16813 ^ 1'b0 ;
  assign n21117 = n13469 & ~n21116 ;
  assign n21118 = n5107 & ~n5425 ;
  assign n21119 = n7938 ^ n1600 ^ 1'b0 ;
  assign n21120 = ( n15916 & n17734 ) | ( n15916 & n21119 ) | ( n17734 & n21119 ) ;
  assign n21121 = n7007 | n8780 ;
  assign n21122 = n2273 & ~n13363 ;
  assign n21124 = n740 & ~n10831 ;
  assign n21123 = n5753 | n16733 ;
  assign n21125 = n21124 ^ n21123 ^ 1'b0 ;
  assign n21126 = n6560 & ~n15402 ;
  assign n21127 = n21126 ^ n6810 ^ n4068 ;
  assign n21128 = ~n3446 & n21127 ;
  assign n21129 = ~n10186 & n21128 ;
  assign n21130 = n6654 ^ n4499 ^ 1'b0 ;
  assign n21131 = ~n7253 & n21130 ;
  assign n21132 = n21131 ^ n10177 ^ n9064 ;
  assign n21133 = ~n165 & n3912 ;
  assign n21134 = n8308 ^ n5747 ^ 1'b0 ;
  assign n21135 = n19640 & ~n21134 ;
  assign n21136 = n4687 ^ n408 ^ 1'b0 ;
  assign n21137 = n474 | n9855 ;
  assign n21138 = n5525 | n21137 ;
  assign n21139 = n17955 ^ n15213 ^ 1'b0 ;
  assign n21140 = n8065 & n21139 ;
  assign n21141 = n5050 & n8545 ;
  assign n21142 = ( n374 & n1323 ) | ( n374 & ~n21141 ) | ( n1323 & ~n21141 ) ;
  assign n21143 = ( ~n5854 & n12961 ) | ( ~n5854 & n21142 ) | ( n12961 & n21142 ) ;
  assign n21144 = ~n2599 & n11542 ;
  assign n21145 = n9105 ^ n2835 ^ 1'b0 ;
  assign n21146 = ~n331 & n8513 ;
  assign n21147 = n4777 & n6139 ;
  assign n21148 = n2669 & n17185 ;
  assign n21149 = n21148 ^ n5863 ^ 1'b0 ;
  assign n21150 = n17587 ^ n2578 ^ n937 ;
  assign n21151 = n14797 ^ n10620 ^ n3756 ;
  assign n21152 = n3828 ^ n3731 ^ 1'b0 ;
  assign n21153 = n2137 & n12312 ;
  assign n21154 = n21153 ^ n2984 ^ 1'b0 ;
  assign n21155 = n1436 & n5116 ;
  assign n21156 = n1895 & n21155 ;
  assign n21157 = n16393 & n21156 ;
  assign n21158 = ( ~n390 & n490 ) | ( ~n390 & n5170 ) | ( n490 & n5170 ) ;
  assign n21159 = ~n2597 & n2651 ;
  assign n21160 = ( ~n2708 & n3323 ) | ( ~n2708 & n8127 ) | ( n3323 & n8127 ) ;
  assign n21161 = n21160 ^ n19926 ^ 1'b0 ;
  assign n21162 = n12141 ^ n2308 ^ 1'b0 ;
  assign n21163 = n1669 & ~n9140 ;
  assign n21164 = n21163 ^ n915 ^ 1'b0 ;
  assign n21165 = ~n4795 & n20616 ;
  assign n21166 = n3850 & n21165 ;
  assign n21167 = n21166 ^ n2018 ^ n1515 ;
  assign n21168 = n7796 & n18084 ;
  assign n21169 = n17151 ^ n16249 ^ 1'b0 ;
  assign n21170 = ( n824 & n4321 ) | ( n824 & n8295 ) | ( n4321 & n8295 ) ;
  assign n21171 = n14584 | n21170 ;
  assign n21172 = n7489 & ~n9251 ;
  assign n21173 = n16411 ^ n12558 ^ 1'b0 ;
  assign n21174 = ( n4884 & ~n7432 ) | ( n4884 & n21173 ) | ( ~n7432 & n21173 ) ;
  assign n21175 = ( n5208 & ~n13564 ) | ( n5208 & n19427 ) | ( ~n13564 & n19427 ) ;
  assign n21176 = n6814 | n19131 ;
  assign n21177 = n21176 ^ n6462 ^ 1'b0 ;
  assign n21178 = n8985 | n19170 ;
  assign n21179 = n21178 ^ n164 ^ 1'b0 ;
  assign n21180 = n2661 & n5338 ;
  assign n21184 = ( n10118 & ~n11925 ) | ( n10118 & n14334 ) | ( ~n11925 & n14334 ) ;
  assign n21185 = n10030 & n21184 ;
  assign n21181 = ( ~n1864 & n2196 ) | ( ~n1864 & n4148 ) | ( n2196 & n4148 ) ;
  assign n21182 = ~n17321 & n21181 ;
  assign n21183 = ~n13014 & n21182 ;
  assign n21186 = n21185 ^ n21183 ^ n15699 ;
  assign n21189 = n16616 ^ n14341 ^ n13313 ;
  assign n21187 = n11407 & ~n18725 ;
  assign n21188 = n21187 ^ n13615 ^ 1'b0 ;
  assign n21190 = n21189 ^ n21188 ^ n365 ;
  assign n21191 = n11370 ^ n8667 ^ n4845 ;
  assign n21192 = n9856 & ~n20066 ;
  assign n21193 = n21191 & n21192 ;
  assign n21197 = n2521 & n17713 ;
  assign n21198 = n21197 ^ n17861 ^ 1'b0 ;
  assign n21199 = ( ~n1497 & n19375 ) | ( ~n1497 & n21198 ) | ( n19375 & n21198 ) ;
  assign n21194 = n20787 ^ n6247 ^ 1'b0 ;
  assign n21195 = ( ~n14126 & n19450 ) | ( ~n14126 & n21194 ) | ( n19450 & n21194 ) ;
  assign n21196 = n9125 | n21195 ;
  assign n21200 = n21199 ^ n21196 ^ 1'b0 ;
  assign n21201 = n13413 ^ n10881 ^ 1'b0 ;
  assign n21202 = ~n6180 & n21201 ;
  assign n21203 = ~n6019 & n7245 ;
  assign n21204 = n21203 ^ n1260 ^ 1'b0 ;
  assign n21205 = n6804 ^ n4479 ^ 1'b0 ;
  assign n21206 = n734 | n21205 ;
  assign n21207 = n21206 ^ n15469 ^ n10805 ;
  assign n21208 = n12001 ^ n5924 ^ 1'b0 ;
  assign n21209 = n4437 & n12402 ;
  assign n21211 = n8856 ^ n542 ^ 1'b0 ;
  assign n21210 = n7598 | n11940 ;
  assign n21212 = n21211 ^ n21210 ^ 1'b0 ;
  assign n21213 = ( n1230 & n3382 ) | ( n1230 & n6315 ) | ( n3382 & n6315 ) ;
  assign n21215 = n11348 ^ n7255 ^ 1'b0 ;
  assign n21214 = n831 | n11402 ;
  assign n21216 = n21215 ^ n21214 ^ 1'b0 ;
  assign n21217 = ~n14697 & n21216 ;
  assign n21218 = n3896 & ~n12316 ;
  assign n21219 = n6029 & n21218 ;
  assign n21220 = n21219 ^ n3102 ^ 1'b0 ;
  assign n21221 = ( n4774 & ~n6929 ) | ( n4774 & n18328 ) | ( ~n6929 & n18328 ) ;
  assign n21222 = n21221 ^ n13796 ^ 1'b0 ;
  assign n21223 = n10054 ^ n7614 ^ 1'b0 ;
  assign n21224 = n3077 | n3177 ;
  assign n21225 = n21224 ^ n1490 ^ 1'b0 ;
  assign n21226 = n7311 & ~n11287 ;
  assign n21227 = n20197 ^ n16141 ^ 1'b0 ;
  assign n21228 = ~n3928 & n21227 ;
  assign n21229 = n15087 ^ n10627 ^ n3655 ;
  assign n21230 = ~n10692 & n10831 ;
  assign n21231 = ( n5010 & n12714 ) | ( n5010 & ~n20167 ) | ( n12714 & ~n20167 ) ;
  assign n21232 = ~n2202 & n9357 ;
  assign n21233 = n12590 & n21232 ;
  assign n21234 = n10780 ^ n712 ^ 1'b0 ;
  assign n21235 = ~n21233 & n21234 ;
  assign n21236 = n13284 ^ n4407 ^ 1'b0 ;
  assign n21237 = ( n967 & n9279 ) | ( n967 & ~n21236 ) | ( n9279 & ~n21236 ) ;
  assign n21238 = ( ~n13215 & n14580 ) | ( ~n13215 & n14974 ) | ( n14580 & n14974 ) ;
  assign n21239 = n2740 & ~n21238 ;
  assign n21240 = ~n21237 & n21239 ;
  assign n21241 = ( ~n229 & n3532 ) | ( ~n229 & n18660 ) | ( n3532 & n18660 ) ;
  assign n21242 = n3455 & ~n21241 ;
  assign n21243 = n18878 & ~n19007 ;
  assign n21244 = n478 & n4302 ;
  assign n21245 = n21244 ^ n895 ^ 1'b0 ;
  assign n21246 = ( n5855 & n11733 ) | ( n5855 & n21245 ) | ( n11733 & n21245 ) ;
  assign n21247 = n21246 ^ n2670 ^ 1'b0 ;
  assign n21248 = n11386 | n21247 ;
  assign n21249 = n17398 ^ n916 ^ 1'b0 ;
  assign n21250 = ~n17420 & n21249 ;
  assign n21251 = ( n16040 & n20991 ) | ( n16040 & n21250 ) | ( n20991 & n21250 ) ;
  assign n21252 = n225 ^ x3 ^ 1'b0 ;
  assign n21253 = n9254 & ~n21252 ;
  assign n21254 = n21253 ^ n19548 ^ 1'b0 ;
  assign n21255 = n21254 ^ n5407 ^ 1'b0 ;
  assign n21256 = n18212 ^ n5773 ^ 1'b0 ;
  assign n21257 = n4121 | n19682 ;
  assign n21258 = n21257 ^ n2952 ^ 1'b0 ;
  assign n21259 = n905 & n21258 ;
  assign n21260 = ~n21256 & n21259 ;
  assign n21261 = n12940 & n14994 ;
  assign n21262 = ~n1126 & n21261 ;
  assign n21263 = n1230 | n3883 ;
  assign n21264 = n6409 & ~n7587 ;
  assign n21265 = n21263 & ~n21264 ;
  assign n21266 = n14639 & n21265 ;
  assign n21268 = n17387 ^ n16454 ^ n12554 ;
  assign n21267 = ~n1850 & n5159 ;
  assign n21269 = n21268 ^ n21267 ^ 1'b0 ;
  assign n21270 = n13970 ^ n11733 ^ 1'b0 ;
  assign n21271 = n3160 & n11916 ;
  assign n21272 = ~n4226 & n21271 ;
  assign n21273 = ~n21270 & n21272 ;
  assign n21274 = n21273 ^ n12897 ^ n12577 ;
  assign n21275 = n8985 ^ n1850 ^ 1'b0 ;
  assign n21276 = n12807 | n21275 ;
  assign n21277 = n4383 & ~n21276 ;
  assign n21278 = n3050 & n14154 ;
  assign n21279 = n20109 & n21278 ;
  assign n21280 = n19663 & ~n19686 ;
  assign n21281 = n1427 & ~n21280 ;
  assign n21282 = n21281 ^ n13336 ^ 1'b0 ;
  assign n21283 = n7137 ^ n4443 ^ 1'b0 ;
  assign n21284 = n16995 | n21283 ;
  assign n21285 = n1403 | n21284 ;
  assign n21286 = n3676 & ~n5681 ;
  assign n21287 = n21286 ^ n11392 ^ 1'b0 ;
  assign n21288 = n2497 & ~n20788 ;
  assign n21289 = n10699 & ~n21288 ;
  assign n21290 = n21287 & n21289 ;
  assign n21291 = n15380 ^ n7274 ^ 1'b0 ;
  assign n21292 = n1383 | n21291 ;
  assign n21293 = ( n1778 & n20364 ) | ( n1778 & ~n21292 ) | ( n20364 & ~n21292 ) ;
  assign n21294 = n21293 ^ n13458 ^ n990 ;
  assign n21297 = n11342 ^ n6675 ^ 1'b0 ;
  assign n21298 = ~n8972 & n21297 ;
  assign n21295 = n9298 | n12689 ;
  assign n21296 = n21295 ^ n10692 ^ 1'b0 ;
  assign n21299 = n21298 ^ n21296 ^ n240 ;
  assign n21300 = n21299 ^ n8511 ^ n3257 ;
  assign n21301 = n3914 | n4749 ;
  assign n21302 = n21301 ^ n7785 ^ 1'b0 ;
  assign n21303 = n4236 & n13096 ;
  assign n21304 = n16073 & n21303 ;
  assign n21305 = ( n17440 & ~n21302 ) | ( n17440 & n21304 ) | ( ~n21302 & n21304 ) ;
  assign n21306 = n21305 ^ n13466 ^ 1'b0 ;
  assign n21307 = ~n13872 & n16905 ;
  assign n21308 = n21307 ^ n1295 ^ 1'b0 ;
  assign n21311 = n5841 ^ n1598 ^ 1'b0 ;
  assign n21309 = ~n4852 & n8017 ;
  assign n21310 = n4419 & n21309 ;
  assign n21312 = n21311 ^ n21310 ^ 1'b0 ;
  assign n21313 = n9302 & n21312 ;
  assign n21314 = n21308 & n21313 ;
  assign n21315 = n247 & n4687 ;
  assign n21316 = n21315 ^ n13721 ^ 1'b0 ;
  assign n21317 = n1770 & ~n7973 ;
  assign n21318 = n11744 ^ n2460 ^ 1'b0 ;
  assign n21319 = ~n21317 & n21318 ;
  assign n21320 = n10813 ^ n3730 ^ 1'b0 ;
  assign n21321 = n6631 & ~n21320 ;
  assign n21322 = n21321 ^ n8225 ^ 1'b0 ;
  assign n21323 = n1343 | n21322 ;
  assign n21324 = n9764 | n21323 ;
  assign n21325 = n431 & n10698 ;
  assign n21326 = n21325 ^ n7900 ^ n1127 ;
  assign n21327 = n1049 & n15310 ;
  assign n21328 = n11391 | n21327 ;
  assign n21329 = ( ~n1890 & n3593 ) | ( ~n1890 & n21328 ) | ( n3593 & n21328 ) ;
  assign n21330 = n1903 | n18399 ;
  assign n21332 = n1709 & n5761 ;
  assign n21333 = ~n3326 & n21332 ;
  assign n21331 = n2855 & ~n16390 ;
  assign n21334 = n21333 ^ n21331 ^ 1'b0 ;
  assign n21335 = n11044 ^ n10795 ^ n222 ;
  assign n21336 = n1118 & n11617 ;
  assign n21337 = n6993 & n11822 ;
  assign n21338 = ( n2031 & n19916 ) | ( n2031 & ~n21337 ) | ( n19916 & ~n21337 ) ;
  assign n21339 = ( n761 & n2822 ) | ( n761 & ~n9268 ) | ( n2822 & ~n9268 ) ;
  assign n21340 = n21339 ^ n19059 ^ n4033 ;
  assign n21341 = ( ~n824 & n12686 ) | ( ~n824 & n13797 ) | ( n12686 & n13797 ) ;
  assign n21342 = n21341 ^ n2822 ^ 1'b0 ;
  assign n21343 = n3176 | n16485 ;
  assign n21344 = n12943 | n21343 ;
  assign n21345 = n13953 ^ n11509 ^ 1'b0 ;
  assign n21346 = n3807 & n21345 ;
  assign n21347 = n8361 ^ n4096 ^ 1'b0 ;
  assign n21348 = ~n12849 & n21347 ;
  assign n21349 = n21348 ^ n8482 ^ 1'b0 ;
  assign n21350 = n11802 & ~n15503 ;
  assign n21351 = n21350 ^ n10578 ^ 1'b0 ;
  assign n21352 = n15257 & ~n16195 ;
  assign n21353 = n21352 ^ n1794 ^ 1'b0 ;
  assign n21354 = n14141 ^ n10793 ^ 1'b0 ;
  assign n21355 = n21354 ^ n18208 ^ n5484 ;
  assign n21356 = n21355 ^ n20197 ^ n1588 ;
  assign n21357 = ( n6845 & ~n8376 ) | ( n6845 & n9075 ) | ( ~n8376 & n9075 ) ;
  assign n21358 = n5821 | n21357 ;
  assign n21359 = n11348 & ~n21358 ;
  assign n21360 = ~n11031 & n14700 ;
  assign n21361 = n1441 | n16649 ;
  assign n21362 = n11966 & ~n21361 ;
  assign n21363 = n1881 & ~n1911 ;
  assign n21364 = n5586 ^ n1196 ^ n210 ;
  assign n21365 = ( ~n9367 & n13612 ) | ( ~n9367 & n20441 ) | ( n13612 & n20441 ) ;
  assign n21366 = ( n3636 & n8029 ) | ( n3636 & n15301 ) | ( n8029 & n15301 ) ;
  assign n21367 = n13473 ^ n6419 ^ n2126 ;
  assign n21368 = ( ~n6537 & n10758 ) | ( ~n6537 & n21367 ) | ( n10758 & n21367 ) ;
  assign n21369 = ( x99 & ~n7939 ) | ( x99 & n21368 ) | ( ~n7939 & n21368 ) ;
  assign n21370 = n11595 ^ n9171 ^ 1'b0 ;
  assign n21371 = n21369 & ~n21370 ;
  assign n21372 = n10003 ^ n1959 ^ 1'b0 ;
  assign n21377 = ~n972 & n2342 ;
  assign n21378 = ~n2342 & n21377 ;
  assign n21373 = n1036 & n3015 ;
  assign n21374 = ~n3015 & n21373 ;
  assign n21375 = n586 & ~n21374 ;
  assign n21376 = ~n586 & n21375 ;
  assign n21379 = n21378 ^ n21376 ^ n5867 ;
  assign n21380 = n21379 ^ n14043 ^ 1'b0 ;
  assign n21381 = ( ~n3640 & n5849 ) | ( ~n3640 & n8145 ) | ( n5849 & n8145 ) ;
  assign n21382 = ( n2252 & n5559 ) | ( n2252 & n5868 ) | ( n5559 & n5868 ) ;
  assign n21383 = n21382 ^ n1544 ^ 1'b0 ;
  assign n21384 = ~n20310 & n21383 ;
  assign n21388 = n1249 & n5369 ;
  assign n21385 = ( ~x7 & n2991 ) | ( ~x7 & n4505 ) | ( n2991 & n4505 ) ;
  assign n21386 = n5881 & n21385 ;
  assign n21387 = n12751 & ~n21386 ;
  assign n21389 = n21388 ^ n21387 ^ 1'b0 ;
  assign n21390 = ( ~n3063 & n7996 ) | ( ~n3063 & n13984 ) | ( n7996 & n13984 ) ;
  assign n21391 = ( ~n10132 & n12225 ) | ( ~n10132 & n20533 ) | ( n12225 & n20533 ) ;
  assign n21392 = n4263 ^ n2300 ^ 1'b0 ;
  assign n21393 = n1751 & ~n21392 ;
  assign n21394 = n14389 ^ n8497 ^ n2310 ;
  assign n21395 = n21394 ^ n9682 ^ 1'b0 ;
  assign n21396 = n17341 | n21395 ;
  assign n21397 = n20865 ^ n10617 ^ 1'b0 ;
  assign n21398 = n3530 & n3610 ;
  assign n21399 = n7004 & ~n7565 ;
  assign n21400 = n18353 ^ n4095 ^ 1'b0 ;
  assign n21401 = n3006 & n21400 ;
  assign n21402 = ( ~n1697 & n9197 ) | ( ~n1697 & n19563 ) | ( n9197 & n19563 ) ;
  assign n21403 = n19104 ^ n684 ^ 1'b0 ;
  assign n21404 = n21402 & ~n21403 ;
  assign n21406 = ( ~n1554 & n4175 ) | ( ~n1554 & n5317 ) | ( n4175 & n5317 ) ;
  assign n21407 = n9277 ^ n6461 ^ 1'b0 ;
  assign n21408 = n21406 | n21407 ;
  assign n21405 = n4448 & n5878 ;
  assign n21409 = n21408 ^ n21405 ^ 1'b0 ;
  assign n21410 = n19348 ^ n12568 ^ n4538 ;
  assign n21411 = n17117 & n18023 ;
  assign n21412 = n8560 ^ n465 ^ 1'b0 ;
  assign n21413 = n21412 ^ n20700 ^ 1'b0 ;
  assign n21414 = n7343 | n21413 ;
  assign n21415 = n9659 ^ n3211 ^ 1'b0 ;
  assign n21416 = ~n6138 & n21415 ;
  assign n21417 = ~n2308 & n4476 ;
  assign n21418 = ( n356 & ~n17792 ) | ( n356 & n17955 ) | ( ~n17792 & n17955 ) ;
  assign n21420 = n14421 ^ n6460 ^ 1'b0 ;
  assign n21421 = n15304 ^ n13519 ^ 1'b0 ;
  assign n21422 = n7388 | n21421 ;
  assign n21423 = n21420 & ~n21422 ;
  assign n21419 = n8082 & n14994 ;
  assign n21424 = n21423 ^ n21419 ^ 1'b0 ;
  assign n21425 = ( n7878 & n18780 ) | ( n7878 & ~n21424 ) | ( n18780 & ~n21424 ) ;
  assign n21426 = n14759 ^ n14205 ^ 1'b0 ;
  assign n21427 = ~n2018 & n21426 ;
  assign n21428 = n19522 ^ n13466 ^ 1'b0 ;
  assign n21429 = ~n15811 & n21428 ;
  assign n21430 = n21177 ^ n9316 ^ 1'b0 ;
  assign n21431 = ~n257 & n21430 ;
  assign n21432 = n3296 ^ n2653 ^ 1'b0 ;
  assign n21433 = n2589 & ~n21432 ;
  assign n21434 = ~n15061 & n21433 ;
  assign n21435 = ( n3441 & n13751 ) | ( n3441 & ~n14338 ) | ( n13751 & ~n14338 ) ;
  assign n21436 = n8795 ^ n160 ^ 1'b0 ;
  assign n21437 = ~n1159 & n21436 ;
  assign n21438 = n21437 ^ n15752 ^ n10153 ;
  assign n21439 = n17550 ^ n14332 ^ n2534 ;
  assign n21440 = n21439 ^ n11031 ^ n575 ;
  assign n21441 = n289 & ~n6496 ;
  assign n21442 = ~n1160 & n21441 ;
  assign n21443 = n1035 & n9004 ;
  assign n21444 = ~n4043 & n21443 ;
  assign n21445 = x13 & n353 ;
  assign n21446 = n21445 ^ n11609 ^ n6456 ;
  assign n21447 = n13122 | n21446 ;
  assign n21448 = n10069 | n21447 ;
  assign n21449 = n21444 | n21448 ;
  assign n21450 = n21449 ^ n2417 ^ 1'b0 ;
  assign n21451 = n1871 ^ n1462 ^ 1'b0 ;
  assign n21452 = n5237 ^ n3972 ^ 1'b0 ;
  assign n21453 = n19014 & n21452 ;
  assign n21454 = n927 & n5792 ;
  assign n21455 = n21454 ^ n3720 ^ 1'b0 ;
  assign n21456 = ~n672 & n21455 ;
  assign n21457 = ( n2303 & ~n5731 ) | ( n2303 & n21456 ) | ( ~n5731 & n21456 ) ;
  assign n21458 = n4068 & n5736 ;
  assign n21459 = n15707 | n19031 ;
  assign n21460 = n2106 & ~n21459 ;
  assign n21461 = ( n5581 & ~n21458 ) | ( n5581 & n21460 ) | ( ~n21458 & n21460 ) ;
  assign n21462 = n1433 ^ n1215 ^ 1'b0 ;
  assign n21463 = n2542 & ~n10558 ;
  assign n21464 = n2997 & ~n8430 ;
  assign n21465 = n21464 ^ n20211 ^ n18015 ;
  assign n21466 = ( n21462 & n21463 ) | ( n21462 & ~n21465 ) | ( n21463 & ~n21465 ) ;
  assign n21470 = ( ~n12507 & n13122 ) | ( ~n12507 & n17939 ) | ( n13122 & n17939 ) ;
  assign n21471 = ( n1051 & ~n17541 ) | ( n1051 & n21470 ) | ( ~n17541 & n21470 ) ;
  assign n21467 = n279 | n2893 ;
  assign n21468 = n21467 ^ n3126 ^ 1'b0 ;
  assign n21469 = n10484 | n21468 ;
  assign n21472 = n21471 ^ n21469 ^ 1'b0 ;
  assign n21473 = n5661 & n21472 ;
  assign n21474 = n7032 & n21473 ;
  assign n21475 = n7022 ^ n5317 ^ 1'b0 ;
  assign n21476 = n20936 & ~n21475 ;
  assign n21477 = ~n14714 & n21476 ;
  assign n21478 = ~n3777 & n21477 ;
  assign n21479 = n9778 ^ n7030 ^ 1'b0 ;
  assign n21480 = ~n8140 & n21479 ;
  assign n21481 = n21480 ^ n13627 ^ 1'b0 ;
  assign n21482 = ~n9970 & n16165 ;
  assign n21483 = n8138 ^ n5333 ^ n824 ;
  assign n21484 = n3993 ^ n2714 ^ 1'b0 ;
  assign n21485 = n21483 & n21484 ;
  assign n21486 = ~n9209 & n21485 ;
  assign n21487 = n21486 ^ n1041 ^ 1'b0 ;
  assign n21488 = n21487 ^ n1438 ^ 1'b0 ;
  assign n21489 = ~n261 & n9514 ;
  assign n21491 = n5453 ^ n1341 ^ n579 ;
  assign n21492 = n21491 ^ n16305 ^ n1581 ;
  assign n21490 = n9742 ^ n7100 ^ 1'b0 ;
  assign n21493 = n21492 ^ n21490 ^ n3051 ;
  assign n21494 = ~n12027 & n14073 ;
  assign n21495 = n19767 ^ n12492 ^ 1'b0 ;
  assign n21496 = n8953 ^ x46 ^ 1'b0 ;
  assign n21497 = n1046 | n21496 ;
  assign n21500 = n6472 ^ n3104 ^ 1'b0 ;
  assign n21498 = n340 | n1403 ;
  assign n21499 = n4287 & ~n21498 ;
  assign n21501 = n21500 ^ n21499 ^ 1'b0 ;
  assign n21502 = n21501 ^ n5809 ^ 1'b0 ;
  assign n21503 = n11613 | n13545 ;
  assign n21504 = n21503 ^ n18576 ^ n5806 ;
  assign n21505 = n15851 ^ n9844 ^ 1'b0 ;
  assign n21506 = ( n3362 & n15656 ) | ( n3362 & n21505 ) | ( n15656 & n21505 ) ;
  assign n21507 = n21184 ^ n14347 ^ 1'b0 ;
  assign n21508 = n9850 | n21507 ;
  assign n21509 = n21506 & ~n21508 ;
  assign n21510 = n21509 ^ n20250 ^ n4856 ;
  assign n21511 = n3428 ^ n1648 ^ 1'b0 ;
  assign n21512 = n210 & n21511 ;
  assign n21513 = n4180 | n4995 ;
  assign n21514 = n21512 & n21513 ;
  assign n21515 = ~n11096 & n21514 ;
  assign n21516 = n8463 ^ n1671 ^ 1'b0 ;
  assign n21517 = ~n17158 & n21516 ;
  assign n21518 = n10843 & n21517 ;
  assign n21519 = n20310 ^ n18223 ^ 1'b0 ;
  assign n21520 = n2021 & n21519 ;
  assign n21521 = n7003 | n15515 ;
  assign n21522 = ( n1818 & n6652 ) | ( n1818 & n7415 ) | ( n6652 & n7415 ) ;
  assign n21523 = n7391 | n11106 ;
  assign n21524 = n16366 ^ n13823 ^ 1'b0 ;
  assign n21526 = ~n7560 & n9093 ;
  assign n21527 = n7323 & n10045 ;
  assign n21528 = ~n21526 & n21527 ;
  assign n21529 = n21528 ^ n1756 ^ 1'b0 ;
  assign n21525 = n8351 | n11032 ;
  assign n21530 = n21529 ^ n21525 ^ 1'b0 ;
  assign n21531 = n7707 & n19348 ;
  assign n21532 = n21531 ^ n9632 ^ 1'b0 ;
  assign n21533 = n21532 ^ n16887 ^ n5593 ;
  assign n21534 = n21533 ^ n7304 ^ 1'b0 ;
  assign n21535 = n12357 & ~n21534 ;
  assign n21536 = n6580 | n11320 ;
  assign n21537 = n21536 ^ n8474 ^ n5720 ;
  assign n21538 = n3252 & ~n6589 ;
  assign n21539 = n19916 & ~n21538 ;
  assign n21540 = ~n21537 & n21539 ;
  assign n21542 = ~n1643 & n4369 ;
  assign n21543 = n3103 & n21542 ;
  assign n21541 = n17695 ^ n15684 ^ n3120 ;
  assign n21544 = n21543 ^ n21541 ^ 1'b0 ;
  assign n21545 = ~n386 & n7694 ;
  assign n21546 = n21545 ^ n15625 ^ 1'b0 ;
  assign n21547 = ( n1374 & n11996 ) | ( n1374 & ~n18398 ) | ( n11996 & ~n18398 ) ;
  assign n21548 = n4544 ^ n3436 ^ 1'b0 ;
  assign n21549 = n19280 & ~n21548 ;
  assign n21550 = n2180 ^ n1431 ^ 1'b0 ;
  assign n21551 = n6555 & ~n21550 ;
  assign n21552 = x13 | n2217 ;
  assign n21553 = n21551 | n21552 ;
  assign n21554 = n8014 ^ n1855 ^ 1'b0 ;
  assign n21555 = n4778 & ~n21554 ;
  assign n21556 = n21555 ^ n9059 ^ n8268 ;
  assign n21559 = n3403 ^ n1441 ^ 1'b0 ;
  assign n21560 = n21559 ^ n6527 ^ 1'b0 ;
  assign n21561 = ~n4433 & n21560 ;
  assign n21558 = ( ~n740 & n756 ) | ( ~n740 & n2740 ) | ( n756 & n2740 ) ;
  assign n21557 = n11203 ^ n6138 ^ n4135 ;
  assign n21562 = n21561 ^ n21558 ^ n21557 ;
  assign n21563 = n9766 & ~n20356 ;
  assign n21564 = n21563 ^ n2712 ^ 1'b0 ;
  assign n21565 = ~n1271 & n8005 ;
  assign n21566 = ~n21564 & n21565 ;
  assign n21567 = ~n6971 & n21566 ;
  assign n21568 = n2957 | n14280 ;
  assign n21569 = ( ~n588 & n21567 ) | ( ~n588 & n21568 ) | ( n21567 & n21568 ) ;
  assign n21570 = n1351 | n20045 ;
  assign n21571 = n16417 ^ n15925 ^ n730 ;
  assign n21572 = n14952 ^ n12463 ^ 1'b0 ;
  assign n21573 = n21571 | n21572 ;
  assign n21574 = n20616 ^ n5348 ^ n922 ;
  assign n21575 = n8143 ^ n245 ^ 1'b0 ;
  assign n21576 = ( ~n9781 & n21574 ) | ( ~n9781 & n21575 ) | ( n21574 & n21575 ) ;
  assign n21577 = n21576 ^ n17508 ^ 1'b0 ;
  assign n21578 = x119 & ~n1113 ;
  assign n21579 = n21578 ^ n18437 ^ 1'b0 ;
  assign n21580 = n6025 ^ n5090 ^ 1'b0 ;
  assign n21581 = n13944 | n21580 ;
  assign n21582 = n21581 ^ n1285 ^ 1'b0 ;
  assign n21583 = n211 & n7859 ;
  assign n21584 = ( x106 & n776 ) | ( x106 & n7771 ) | ( n776 & n7771 ) ;
  assign n21585 = n12681 & n21584 ;
  assign n21586 = n13880 ^ n9762 ^ n2055 ;
  assign n21587 = n20986 ^ n19969 ^ n14313 ;
  assign n21588 = n4329 ^ n1162 ^ 1'b0 ;
  assign n21589 = n10044 | n21588 ;
  assign n21590 = n5170 | n7292 ;
  assign n21592 = n1782 & n16532 ;
  assign n21593 = n21592 ^ n2056 ^ 1'b0 ;
  assign n21591 = x119 & n17581 ;
  assign n21594 = n21593 ^ n21591 ^ 1'b0 ;
  assign n21595 = n21594 ^ n12071 ^ 1'b0 ;
  assign n21596 = n10840 ^ n4397 ^ n2331 ;
  assign n21597 = n21596 ^ n10341 ^ 1'b0 ;
  assign n21598 = n4020 & n18002 ;
  assign n21599 = ~n4616 & n21598 ;
  assign n21600 = n314 | n6428 ;
  assign n21601 = n11024 ^ n10776 ^ 1'b0 ;
  assign n21602 = n17053 & n21601 ;
  assign n21603 = n6899 & n21602 ;
  assign n21604 = n4414 | n12532 ;
  assign n21605 = n4710 | n21604 ;
  assign n21606 = n17686 ^ n16872 ^ n4871 ;
  assign n21607 = n21181 ^ n6225 ^ 1'b0 ;
  assign n21608 = ~n5032 & n21607 ;
  assign n21609 = n15758 ^ n2619 ^ n2421 ;
  assign n21610 = ( n5873 & n8043 ) | ( n5873 & ~n13822 ) | ( n8043 & ~n13822 ) ;
  assign n21611 = n21609 | n21610 ;
  assign n21612 = n187 & ~n1214 ;
  assign n21613 = n2245 & n21612 ;
  assign n21614 = n21613 ^ n3654 ^ 1'b0 ;
  assign n21615 = ~n719 & n9585 ;
  assign n21616 = n21615 ^ n4487 ^ 1'b0 ;
  assign n21617 = n5849 & n8742 ;
  assign n21618 = n21616 & n21617 ;
  assign n21619 = n4199 & ~n10603 ;
  assign n21620 = n16466 | n21619 ;
  assign n21621 = n21620 ^ n17155 ^ n599 ;
  assign n21622 = ( n9020 & n10734 ) | ( n9020 & ~n12754 ) | ( n10734 & ~n12754 ) ;
  assign n21623 = ~n2029 & n18729 ;
  assign n21624 = ( n362 & n2462 ) | ( n362 & ~n21623 ) | ( n2462 & ~n21623 ) ;
  assign n21626 = ~n5614 & n14316 ;
  assign n21625 = n2449 & ~n9356 ;
  assign n21627 = n21626 ^ n21625 ^ 1'b0 ;
  assign n21628 = n17557 ^ n1727 ^ 1'b0 ;
  assign n21629 = n21627 & ~n21628 ;
  assign n21630 = n4054 | n19789 ;
  assign n21631 = n6407 ^ n1061 ^ 1'b0 ;
  assign n21632 = n7221 & ~n21631 ;
  assign n21633 = n3953 & ~n10768 ;
  assign n21634 = ~n13032 & n21633 ;
  assign n21635 = n5536 | n21634 ;
  assign n21636 = n644 & ~n4463 ;
  assign n21637 = n21636 ^ n10974 ^ 1'b0 ;
  assign n21638 = n1414 & n7938 ;
  assign n21639 = n21638 ^ n13314 ^ 1'b0 ;
  assign n21640 = n21639 ^ n940 ^ n753 ;
  assign n21641 = n6055 ^ n4713 ^ 1'b0 ;
  assign n21642 = ( n1739 & ~n19405 ) | ( n1739 & n21641 ) | ( ~n19405 & n21641 ) ;
  assign n21643 = n9702 ^ n5607 ^ 1'b0 ;
  assign n21644 = n11211 | n17046 ;
  assign n21645 = n15813 ^ n575 ^ 1'b0 ;
  assign n21646 = n10805 | n21645 ;
  assign n21647 = n15050 & ~n19183 ;
  assign n21648 = n21646 & n21647 ;
  assign n21649 = n4384 | n18729 ;
  assign n21650 = n9613 & ~n21649 ;
  assign n21651 = ( ~n4653 & n6582 ) | ( ~n4653 & n6948 ) | ( n6582 & n6948 ) ;
  assign n21652 = n15403 & ~n21651 ;
  assign n21653 = n21652 ^ n3581 ^ 1'b0 ;
  assign n21654 = n16853 & ~n21653 ;
  assign n21655 = n21654 ^ n18167 ^ 1'b0 ;
  assign n21656 = n21650 | n21655 ;
  assign n21657 = ~n6541 & n13847 ;
  assign n21658 = ~n5037 & n21657 ;
  assign n21659 = n21658 ^ n13771 ^ n8918 ;
  assign n21660 = n13754 & n17945 ;
  assign n21661 = ( ~n1162 & n20453 ) | ( ~n1162 & n21660 ) | ( n20453 & n21660 ) ;
  assign n21662 = n6804 ^ n2259 ^ n802 ;
  assign n21663 = n12129 & ~n21662 ;
  assign n21664 = n21663 ^ n2437 ^ 1'b0 ;
  assign n21665 = n12636 ^ n11679 ^ 1'b0 ;
  assign n21666 = ~n2607 & n5399 ;
  assign n21667 = n21666 ^ n6207 ^ 1'b0 ;
  assign n21668 = ~n4300 & n21667 ;
  assign n21669 = ~n12966 & n21668 ;
  assign n21670 = ~n3884 & n21669 ;
  assign n21671 = ~n3604 & n5038 ;
  assign n21672 = ~n15919 & n21671 ;
  assign n21673 = n3198 & ~n21672 ;
  assign n21674 = n3212 & ~n9818 ;
  assign n21675 = n21674 ^ n5894 ^ 1'b0 ;
  assign n21676 = ( ~n1819 & n3022 ) | ( ~n1819 & n21675 ) | ( n3022 & n21675 ) ;
  assign n21677 = n4144 ^ n1175 ^ n1148 ;
  assign n21678 = n21677 ^ n10793 ^ n4458 ;
  assign n21679 = ( n1942 & ~n5329 ) | ( n1942 & n21678 ) | ( ~n5329 & n21678 ) ;
  assign n21680 = n18842 ^ n3931 ^ 1'b0 ;
  assign n21681 = n13183 ^ n3248 ^ 1'b0 ;
  assign n21682 = n1550 & ~n21681 ;
  assign n21685 = n932 & ~n6255 ;
  assign n21686 = n827 & n21685 ;
  assign n21687 = n4048 & ~n21686 ;
  assign n21683 = n10726 ^ n309 ^ 1'b0 ;
  assign n21684 = n7962 & n21683 ;
  assign n21688 = n21687 ^ n21684 ^ 1'b0 ;
  assign n21689 = n1974 ^ n209 ^ 1'b0 ;
  assign n21690 = ~n17567 & n21689 ;
  assign n21691 = n21057 ^ n1542 ^ 1'b0 ;
  assign n21692 = n620 | n9801 ;
  assign n21693 = n6140 & n21692 ;
  assign n21694 = n15492 ^ n12440 ^ 1'b0 ;
  assign n21695 = n21693 & n21694 ;
  assign n21702 = n10645 ^ n5317 ^ n1192 ;
  assign n21700 = n20375 ^ n12400 ^ n8027 ;
  assign n21701 = n21700 ^ n8471 ^ 1'b0 ;
  assign n21696 = x121 & n1770 ;
  assign n21697 = n5092 & n21696 ;
  assign n21698 = n3572 | n21697 ;
  assign n21699 = n5720 & ~n21698 ;
  assign n21703 = n21702 ^ n21701 ^ n21699 ;
  assign n21704 = ~n3678 & n7274 ;
  assign n21705 = n21704 ^ n13623 ^ 1'b0 ;
  assign n21706 = n21705 ^ n15975 ^ n15380 ;
  assign n21707 = n1308 ^ x0 ^ 1'b0 ;
  assign n21708 = ~n383 & n21707 ;
  assign n21709 = n5767 | n21708 ;
  assign n21710 = n21709 ^ n1374 ^ 1'b0 ;
  assign n21711 = ~n4094 & n21710 ;
  assign n21712 = n1622 & ~n6858 ;
  assign n21713 = n21712 ^ n10615 ^ n3659 ;
  assign n21714 = n1179 & ~n4385 ;
  assign n21715 = ~n447 & n21714 ;
  assign n21716 = n8853 | n21715 ;
  assign n21717 = n4542 & ~n21716 ;
  assign n21718 = n21713 & n21717 ;
  assign n21719 = n21718 ^ n19306 ^ 1'b0 ;
  assign n21720 = n9587 | n13357 ;
  assign n21721 = n21720 ^ n4306 ^ 1'b0 ;
  assign n21722 = n5836 & ~n21721 ;
  assign n21723 = n21722 ^ n2092 ^ 1'b0 ;
  assign n21724 = n10109 | n21619 ;
  assign n21725 = ( n2204 & n5873 ) | ( n2204 & ~n21724 ) | ( n5873 & ~n21724 ) ;
  assign n21726 = n18383 ^ n16339 ^ n2547 ;
  assign n21727 = n21726 ^ n18118 ^ n11071 ;
  assign n21728 = n4616 | n11137 ;
  assign n21729 = n20011 ^ n10824 ^ n1163 ;
  assign n21730 = n21729 ^ n10298 ^ 1'b0 ;
  assign n21731 = n5523 | n21730 ;
  assign n21732 = n21731 ^ n15725 ^ n11434 ;
  assign n21733 = n7291 | n12254 ;
  assign n21734 = ~n4861 & n21733 ;
  assign n21735 = n782 | n18703 ;
  assign n21736 = n21735 ^ n21065 ^ 1'b0 ;
  assign n21737 = n12339 ^ n4924 ^ 1'b0 ;
  assign n21738 = ~n16350 & n21737 ;
  assign n21739 = n21738 ^ n3402 ^ x114 ;
  assign n21740 = n4819 | n21739 ;
  assign n21741 = n8567 ^ n2731 ^ 1'b0 ;
  assign n21742 = n9140 | n21741 ;
  assign n21743 = n21742 ^ n17478 ^ n10643 ;
  assign n21744 = n2344 & ~n21743 ;
  assign n21745 = n8245 ^ n993 ^ n546 ;
  assign n21746 = n21745 ^ n16485 ^ n10584 ;
  assign n21747 = n4829 & n21746 ;
  assign n21748 = n2869 ^ n1311 ^ 1'b0 ;
  assign n21749 = n932 ^ x73 ^ 1'b0 ;
  assign n21750 = ~n8767 & n21749 ;
  assign n21751 = ( n580 & n4884 ) | ( n580 & ~n21750 ) | ( n4884 & ~n21750 ) ;
  assign n21752 = n2455 & ~n15943 ;
  assign n21753 = n21751 & n21752 ;
  assign n21754 = ~n12350 & n12485 ;
  assign n21755 = ~n11161 & n12472 ;
  assign n21756 = ( n15824 & n21754 ) | ( n15824 & n21755 ) | ( n21754 & n21755 ) ;
  assign n21757 = ~n7042 & n13453 ;
  assign n21758 = n21757 ^ n7177 ^ 1'b0 ;
  assign n21759 = n8715 & n21224 ;
  assign n21760 = ~n17002 & n21759 ;
  assign n21761 = n4617 ^ n4405 ^ 1'b0 ;
  assign n21762 = ~n5341 & n21761 ;
  assign n21767 = ~n8560 & n10591 ;
  assign n21764 = n8608 ^ n2419 ^ 1'b0 ;
  assign n21765 = n13198 & n21764 ;
  assign n21763 = n17188 ^ n6788 ^ 1'b0 ;
  assign n21766 = n21765 ^ n21763 ^ 1'b0 ;
  assign n21768 = n21767 ^ n21766 ^ 1'b0 ;
  assign n21769 = n8084 & ~n21768 ;
  assign n21770 = n4389 & n18128 ;
  assign n21771 = ~n21769 & n21770 ;
  assign n21772 = n589 & n11525 ;
  assign n21773 = n21772 ^ n3164 ^ 1'b0 ;
  assign n21774 = ( n5332 & n6426 ) | ( n5332 & n8254 ) | ( n6426 & n8254 ) ;
  assign n21775 = n7269 ^ n4341 ^ 1'b0 ;
  assign n21776 = n18197 ^ n8403 ^ 1'b0 ;
  assign n21777 = n21775 | n21776 ;
  assign n21778 = n1467 & ~n21777 ;
  assign n21779 = n21778 ^ n6953 ^ 1'b0 ;
  assign n21780 = n21779 ^ n631 ^ 1'b0 ;
  assign n21781 = n21774 & ~n21780 ;
  assign n21784 = n13148 ^ n11958 ^ 1'b0 ;
  assign n21785 = n2862 | n21784 ;
  assign n21786 = n4820 ^ n3756 ^ 1'b0 ;
  assign n21787 = n21785 | n21786 ;
  assign n21782 = n10523 & n15980 ;
  assign n21783 = ( n12632 & ~n15901 ) | ( n12632 & n21782 ) | ( ~n15901 & n21782 ) ;
  assign n21788 = n21787 ^ n21783 ^ n18948 ;
  assign n21789 = n21788 ^ n11949 ^ n10919 ;
  assign n21790 = ( n1358 & n1378 ) | ( n1358 & ~n11542 ) | ( n1378 & ~n11542 ) ;
  assign n21791 = n6205 ^ n1445 ^ 1'b0 ;
  assign n21792 = n6460 & n21791 ;
  assign n21793 = n21792 ^ n2863 ^ x48 ;
  assign n21794 = n12412 & n21793 ;
  assign n21795 = n21794 ^ n3373 ^ 1'b0 ;
  assign n21796 = ~n2845 & n16464 ;
  assign n21797 = n21796 ^ n2951 ^ 1'b0 ;
  assign n21798 = n7225 ^ n1833 ^ 1'b0 ;
  assign n21799 = n21797 & n21798 ;
  assign n21800 = ~n10394 & n11051 ;
  assign n21801 = n20691 ^ n5049 ^ 1'b0 ;
  assign n21802 = n14251 ^ n7481 ^ 1'b0 ;
  assign n21803 = ~n3951 & n21802 ;
  assign n21804 = n21803 ^ n14532 ^ 1'b0 ;
  assign n21806 = n17440 ^ n2272 ^ 1'b0 ;
  assign n21807 = n18115 & n21806 ;
  assign n21805 = n11684 ^ n8748 ^ n6376 ;
  assign n21808 = n21807 ^ n21805 ^ n21697 ;
  assign n21809 = n10875 ^ n6308 ^ 1'b0 ;
  assign n21810 = n6891 & ~n21809 ;
  assign n21811 = n9058 & n21810 ;
  assign n21814 = ( n11241 & n12682 ) | ( n11241 & ~n16339 ) | ( n12682 & ~n16339 ) ;
  assign n21815 = n20819 & n21814 ;
  assign n21816 = n21815 ^ n9358 ^ 1'b0 ;
  assign n21812 = n1477 | n13094 ;
  assign n21813 = n17149 & n21812 ;
  assign n21817 = n21816 ^ n21813 ^ 1'b0 ;
  assign n21818 = ~n6273 & n9982 ;
  assign n21819 = ( n11632 & ~n19129 ) | ( n11632 & n21818 ) | ( ~n19129 & n21818 ) ;
  assign n21820 = ( ~n3999 & n11645 ) | ( ~n3999 & n12516 ) | ( n11645 & n12516 ) ;
  assign n21821 = n15168 ^ n6152 ^ n1996 ;
  assign n21822 = n21821 ^ n18654 ^ 1'b0 ;
  assign n21823 = n21822 ^ n11707 ^ 1'b0 ;
  assign n21824 = n14334 ^ n10335 ^ 1'b0 ;
  assign n21825 = n21824 ^ n5747 ^ 1'b0 ;
  assign n21829 = n1577 & n15107 ;
  assign n21826 = n12317 & n13405 ;
  assign n21827 = n2640 & n21826 ;
  assign n21828 = n17914 | n21827 ;
  assign n21830 = n21829 ^ n21828 ^ 1'b0 ;
  assign n21831 = n1535 & n17636 ;
  assign n21832 = n10762 | n16350 ;
  assign n21833 = ( n7765 & n21831 ) | ( n7765 & n21832 ) | ( n21831 & n21832 ) ;
  assign n21834 = n2137 & ~n7226 ;
  assign n21835 = n21834 ^ n3472 ^ 1'b0 ;
  assign n21836 = ( ~n10539 & n17231 ) | ( ~n10539 & n21835 ) | ( n17231 & n21835 ) ;
  assign n21837 = ~n2008 & n8230 ;
  assign n21838 = n1112 & ~n2515 ;
  assign n21839 = ( n21836 & n21837 ) | ( n21836 & ~n21838 ) | ( n21837 & ~n21838 ) ;
  assign n21840 = n21839 ^ n19595 ^ n5907 ;
  assign n21841 = n6412 ^ n4865 ^ n522 ;
  assign n21842 = n10305 | n21841 ;
  assign n21843 = n3926 & ~n21842 ;
  assign n21844 = n21843 ^ n7643 ^ n820 ;
  assign n21845 = ~n4642 & n17432 ;
  assign n21846 = n21388 ^ n13244 ^ 1'b0 ;
  assign n21847 = n20237 & ~n21769 ;
  assign n21848 = n133 & n5108 ;
  assign n21849 = ~n17407 & n21848 ;
  assign n21850 = n6609 & ~n6717 ;
  assign n21851 = ~n1598 & n21850 ;
  assign n21852 = n4900 | n21851 ;
  assign n21853 = n21354 ^ n2961 ^ n2875 ;
  assign n21854 = ( n1199 & n4881 ) | ( n1199 & n10040 ) | ( n4881 & n10040 ) ;
  assign n21855 = n8731 & ~n10112 ;
  assign n21856 = n21855 ^ n5888 ^ 1'b0 ;
  assign n21857 = ( n8851 & n15093 ) | ( n8851 & ~n21856 ) | ( n15093 & ~n21856 ) ;
  assign n21858 = n16031 ^ n2879 ^ 1'b0 ;
  assign n21859 = n11266 & n21858 ;
  assign n21860 = n10097 & n21859 ;
  assign n21861 = n21860 ^ n10664 ^ n1674 ;
  assign n21862 = n11948 ^ n6671 ^ 1'b0 ;
  assign n21864 = n11410 ^ n11295 ^ x3 ;
  assign n21863 = ( ~n2206 & n9530 ) | ( ~n2206 & n13618 ) | ( n9530 & n13618 ) ;
  assign n21865 = n21864 ^ n21863 ^ n1723 ;
  assign n21866 = n17888 ^ n14151 ^ 1'b0 ;
  assign n21867 = n8543 & n21866 ;
  assign n21868 = n15475 | n15543 ;
  assign n21869 = n5155 & n16395 ;
  assign n21870 = n21869 ^ n609 ^ 1'b0 ;
  assign n21871 = ( n542 & n2653 ) | ( n542 & n3643 ) | ( n2653 & n3643 ) ;
  assign n21872 = n16182 ^ n9996 ^ 1'b0 ;
  assign n21873 = ( n4011 & ~n14612 ) | ( n4011 & n19506 ) | ( ~n14612 & n19506 ) ;
  assign n21874 = n6728 ^ n1644 ^ 1'b0 ;
  assign n21875 = ~n21873 & n21874 ;
  assign n21876 = ~n7189 & n21875 ;
  assign n21877 = n21876 ^ n1076 ^ 1'b0 ;
  assign n21878 = n9221 | n9670 ;
  assign n21879 = n21878 ^ n15491 ^ n6077 ;
  assign n21880 = ~n1673 & n4074 ;
  assign n21881 = n449 & n21880 ;
  assign n21882 = n12999 | n21881 ;
  assign n21883 = n2186 & ~n21882 ;
  assign n21886 = ( ~n705 & n12488 ) | ( ~n705 & n20421 ) | ( n12488 & n20421 ) ;
  assign n21884 = ( n9628 & n12849 ) | ( n9628 & n14247 ) | ( n12849 & n14247 ) ;
  assign n21885 = n10485 | n21884 ;
  assign n21887 = n21886 ^ n21885 ^ 1'b0 ;
  assign n21888 = n134 | n8100 ;
  assign n21889 = n9349 & ~n21888 ;
  assign n21890 = n18929 ^ n599 ^ 1'b0 ;
  assign n21891 = n21889 | n21890 ;
  assign n21892 = n20885 & ~n21708 ;
  assign n21893 = n2416 | n10180 ;
  assign n21894 = n3456 | n21893 ;
  assign n21895 = n1334 & ~n15786 ;
  assign n21896 = ( n8892 & n21894 ) | ( n8892 & n21895 ) | ( n21894 & n21895 ) ;
  assign n21897 = n18125 ^ n1233 ^ 1'b0 ;
  assign n21898 = n2282 | n8799 ;
  assign n21899 = n980 & ~n21898 ;
  assign n21900 = ( n710 & n4248 ) | ( n710 & n9982 ) | ( n4248 & n9982 ) ;
  assign n21901 = n10692 | n14620 ;
  assign n21902 = n21900 | n21901 ;
  assign n21903 = ~n21899 & n21902 ;
  assign n21904 = ~n16780 & n21903 ;
  assign n21905 = n1448 & n4867 ;
  assign n21906 = n10528 & ~n21905 ;
  assign n21907 = n21906 ^ n15851 ^ 1'b0 ;
  assign n21908 = ~n11509 & n21907 ;
  assign n21910 = n9976 | n21491 ;
  assign n21911 = n5080 | n21910 ;
  assign n21909 = n13359 | n13550 ;
  assign n21912 = n21911 ^ n21909 ^ 1'b0 ;
  assign n21913 = n20310 ^ n10605 ^ 1'b0 ;
  assign n21914 = n3766 & ~n21913 ;
  assign n21915 = ~n7201 & n15598 ;
  assign n21916 = n21915 ^ n10831 ^ n3143 ;
  assign n21917 = ~n20334 & n21916 ;
  assign n21921 = n5761 ^ n3469 ^ 1'b0 ;
  assign n21918 = ~n2243 & n3041 ;
  assign n21919 = ~n487 & n21918 ;
  assign n21920 = ~n17257 & n21919 ;
  assign n21922 = n21921 ^ n21920 ^ n5625 ;
  assign n21923 = n21922 ^ n9070 ^ n675 ;
  assign n21925 = ~n5032 & n9693 ;
  assign n21926 = n21925 ^ n9856 ^ 1'b0 ;
  assign n21924 = n3234 | n20313 ;
  assign n21927 = n21926 ^ n21924 ^ 1'b0 ;
  assign n21928 = n2724 & n6134 ;
  assign n21929 = ~n11534 & n21928 ;
  assign n21930 = n8204 & ~n8351 ;
  assign n21931 = n21930 ^ n2928 ^ 1'b0 ;
  assign n21932 = n6918 & n8598 ;
  assign n21933 = n21932 ^ n14144 ^ 1'b0 ;
  assign n21934 = n7574 | n8741 ;
  assign n21935 = n12640 | n21934 ;
  assign n21936 = ( n4498 & n13460 ) | ( n4498 & ~n21935 ) | ( n13460 & ~n21935 ) ;
  assign n21937 = n5396 ^ n3176 ^ 1'b0 ;
  assign n21938 = ( n7232 & n20683 ) | ( n7232 & n21937 ) | ( n20683 & n21937 ) ;
  assign n21939 = ~n2817 & n3440 ;
  assign n21940 = n21939 ^ n11293 ^ 1'b0 ;
  assign n21941 = n2527 & n10774 ;
  assign n21942 = n9820 & n21941 ;
  assign n21943 = n1452 ^ n641 ^ 1'b0 ;
  assign n21944 = ( n1534 & n4489 ) | ( n1534 & ~n10039 ) | ( n4489 & ~n10039 ) ;
  assign n21945 = n21944 ^ n3111 ^ 1'b0 ;
  assign n21946 = n10464 & n21945 ;
  assign n21947 = n21943 & n21946 ;
  assign n21948 = n17759 ^ n12490 ^ 1'b0 ;
  assign n21949 = ~n6421 & n21948 ;
  assign n21950 = n9590 & ~n19649 ;
  assign n21951 = n8038 & n21950 ;
  assign n21952 = n16568 ^ n9725 ^ n5049 ;
  assign n21953 = n21952 ^ n12325 ^ n6211 ;
  assign n21954 = ~n1953 & n15418 ;
  assign n21955 = n21954 ^ n19256 ^ 1'b0 ;
  assign n21956 = ( ~n2039 & n3553 ) | ( ~n2039 & n19143 ) | ( n3553 & n19143 ) ;
  assign n21957 = n6787 & n7964 ;
  assign n21958 = n21957 ^ n6410 ^ 1'b0 ;
  assign n21959 = n21767 | n21958 ;
  assign n21960 = n21956 | n21959 ;
  assign n21961 = n6709 & ~n8685 ;
  assign n21962 = n1532 & n21961 ;
  assign n21963 = n21926 ^ n1715 ^ 1'b0 ;
  assign n21964 = n1175 ^ n1073 ^ n391 ;
  assign n21965 = n21964 ^ n6166 ^ 1'b0 ;
  assign n21966 = n2371 | n18783 ;
  assign n21967 = n10435 | n21966 ;
  assign n21968 = ( n6630 & n18295 ) | ( n6630 & n21967 ) | ( n18295 & n21967 ) ;
  assign n21969 = n21965 & n21968 ;
  assign n21970 = n17171 ^ n11493 ^ n10153 ;
  assign n21971 = n825 & ~n11402 ;
  assign n21972 = ~n5213 & n21971 ;
  assign n21973 = n7718 & n20801 ;
  assign n21974 = n21973 ^ n626 ^ 1'b0 ;
  assign n21975 = n8869 & ~n9436 ;
  assign n21976 = n12445 ^ n7269 ^ 1'b0 ;
  assign n21977 = n2984 & n21976 ;
  assign n21978 = ~n5994 & n21977 ;
  assign n21981 = n15234 ^ n8013 ^ n4789 ;
  assign n21980 = n2094 | n15738 ;
  assign n21982 = n21981 ^ n21980 ^ n143 ;
  assign n21979 = n2434 & n12326 ;
  assign n21983 = n21982 ^ n21979 ^ 1'b0 ;
  assign n21984 = n5049 ^ n606 ^ 1'b0 ;
  assign n21985 = n14376 ^ n9231 ^ n2800 ;
  assign n21986 = n14119 ^ n7869 ^ 1'b0 ;
  assign n21987 = n3770 & ~n21986 ;
  assign n21988 = n782 | n10243 ;
  assign n21989 = n11095 & ~n21988 ;
  assign n21990 = ~n6394 & n21989 ;
  assign n21991 = ( n13052 & n21987 ) | ( n13052 & ~n21990 ) | ( n21987 & ~n21990 ) ;
  assign n21992 = ~n10633 & n10981 ;
  assign n21993 = n833 | n9571 ;
  assign n21994 = n21993 ^ n16890 ^ 1'b0 ;
  assign n21995 = n18524 ^ n6003 ^ n279 ;
  assign n21996 = n12981 & ~n21812 ;
  assign n21997 = n11049 ^ n8533 ^ 1'b0 ;
  assign n21998 = n8980 & ~n21997 ;
  assign n21999 = n1330 & n21998 ;
  assign n22000 = n19002 ^ n18741 ^ n6906 ;
  assign n22001 = n4420 | n7947 ;
  assign n22002 = n12682 ^ n8702 ^ 1'b0 ;
  assign n22003 = n19550 ^ n5801 ^ 1'b0 ;
  assign n22004 = n19330 ^ n6206 ^ 1'b0 ;
  assign n22005 = ( n2836 & n8809 ) | ( n2836 & ~n11935 ) | ( n8809 & ~n11935 ) ;
  assign n22006 = n22005 ^ n17548 ^ 1'b0 ;
  assign n22007 = n14370 ^ n9105 ^ 1'b0 ;
  assign n22008 = n7032 | n11292 ;
  assign n22009 = n22008 ^ n11979 ^ 1'b0 ;
  assign n22010 = n3673 & ~n4250 ;
  assign n22011 = ~n3951 & n22010 ;
  assign n22013 = n1123 | n11465 ;
  assign n22014 = n22013 ^ n12069 ^ n11160 ;
  assign n22015 = n22014 ^ x13 ^ 1'b0 ;
  assign n22012 = n11444 & n18129 ;
  assign n22016 = n22015 ^ n22012 ^ n12628 ;
  assign n22017 = n6512 & n19312 ;
  assign n22018 = ( n1470 & n8065 ) | ( n1470 & n12031 ) | ( n8065 & n12031 ) ;
  assign n22019 = ( n16937 & ~n18538 ) | ( n16937 & n22018 ) | ( ~n18538 & n22018 ) ;
  assign n22020 = ~n21616 & n22019 ;
  assign n22021 = n11779 & n22020 ;
  assign n22022 = n16127 ^ n11331 ^ n2927 ;
  assign n22027 = ( n654 & n2464 ) | ( n654 & n7766 ) | ( n2464 & n7766 ) ;
  assign n22028 = n8872 & ~n22027 ;
  assign n22024 = ~n1523 & n8867 ;
  assign n22025 = n22024 ^ n3187 ^ 1'b0 ;
  assign n22023 = n1998 & ~n5504 ;
  assign n22026 = n22025 ^ n22023 ^ n2191 ;
  assign n22029 = n22028 ^ n22026 ^ n5024 ;
  assign n22030 = x82 & n4713 ;
  assign n22031 = ~n397 & n7291 ;
  assign n22032 = n15044 ^ n7364 ^ 1'b0 ;
  assign n22033 = n22031 & n22032 ;
  assign n22034 = n22030 | n22033 ;
  assign n22035 = n17326 ^ n15920 ^ 1'b0 ;
  assign n22036 = ~n5958 & n22035 ;
  assign n22037 = n9218 ^ n5687 ^ 1'b0 ;
  assign n22038 = n22037 ^ n17653 ^ 1'b0 ;
  assign n22039 = ( n5625 & n6877 ) | ( n5625 & n22038 ) | ( n6877 & n22038 ) ;
  assign n22040 = n22039 ^ n19611 ^ 1'b0 ;
  assign n22041 = n16482 | n22040 ;
  assign n22042 = n21410 ^ n9426 ^ 1'b0 ;
  assign n22043 = n858 | n22042 ;
  assign n22044 = n8663 ^ n3873 ^ n1045 ;
  assign n22045 = n17666 ^ n14060 ^ 1'b0 ;
  assign n22046 = ~n1690 & n11471 ;
  assign n22047 = ~n5077 & n22046 ;
  assign n22048 = n19923 ^ n11693 ^ n1658 ;
  assign n22049 = n15221 & ~n22048 ;
  assign n22050 = n2886 | n4303 ;
  assign n22051 = n13116 & n22050 ;
  assign n22052 = n22049 & n22051 ;
  assign n22053 = n15456 ^ n3376 ^ 1'b0 ;
  assign n22054 = ( n2058 & ~n9707 ) | ( n2058 & n17044 ) | ( ~n9707 & n17044 ) ;
  assign n22055 = n7821 | n22054 ;
  assign n22056 = n1444 & ~n2933 ;
  assign n22057 = n22056 ^ n7293 ^ 1'b0 ;
  assign n22058 = n5677 ^ n2171 ^ 1'b0 ;
  assign n22059 = ~n22057 & n22058 ;
  assign n22060 = n20152 ^ n2933 ^ 1'b0 ;
  assign n22061 = n13682 & ~n22060 ;
  assign n22062 = n701 & ~n22061 ;
  assign n22063 = ( ~n4208 & n5107 ) | ( ~n4208 & n5789 ) | ( n5107 & n5789 ) ;
  assign n22064 = ( n1576 & ~n6370 ) | ( n1576 & n22063 ) | ( ~n6370 & n22063 ) ;
  assign n22065 = ( n7219 & ~n9461 ) | ( n7219 & n10806 ) | ( ~n9461 & n10806 ) ;
  assign n22066 = ( n3291 & ~n13177 ) | ( n3291 & n22065 ) | ( ~n13177 & n22065 ) ;
  assign n22067 = n2333 & n14550 ;
  assign n22068 = x22 & ~n824 ;
  assign n22069 = n11949 & ~n22068 ;
  assign n22070 = n11170 ^ n3943 ^ 1'b0 ;
  assign n22071 = ( n7375 & n9017 ) | ( n7375 & n11860 ) | ( n9017 & n11860 ) ;
  assign n22072 = n22071 ^ n1955 ^ 1'b0 ;
  assign n22073 = n22070 & ~n22072 ;
  assign n22074 = n4970 ^ n386 ^ 1'b0 ;
  assign n22075 = ~n2759 & n18856 ;
  assign n22076 = n22075 ^ n20140 ^ 1'b0 ;
  assign n22077 = n21512 ^ n14996 ^ n1621 ;
  assign n22078 = ( n4265 & ~n11856 ) | ( n4265 & n16419 ) | ( ~n11856 & n16419 ) ;
  assign n22079 = ~n10605 & n16684 ;
  assign n22080 = n11475 & ~n22079 ;
  assign n22081 = n7602 & ~n17994 ;
  assign n22082 = n22081 ^ n6226 ^ 1'b0 ;
  assign n22083 = n3538 | n10277 ;
  assign n22084 = n22083 ^ n2968 ^ 1'b0 ;
  assign n22085 = n20572 & ~n22084 ;
  assign n22086 = n18098 & n22085 ;
  assign n22087 = n9373 & n19758 ;
  assign n22088 = n22087 ^ n10464 ^ 1'b0 ;
  assign n22089 = n21003 ^ n12572 ^ 1'b0 ;
  assign n22090 = ~n20264 & n22089 ;
  assign n22091 = n16048 ^ n6288 ^ 1'b0 ;
  assign n22092 = n1715 & n4331 ;
  assign n22093 = ( n4571 & n6833 ) | ( n4571 & n12009 ) | ( n6833 & n12009 ) ;
  assign n22094 = n22093 ^ n8868 ^ n4586 ;
  assign n22095 = n9958 ^ n1687 ^ n1314 ;
  assign n22096 = n389 & n21559 ;
  assign n22097 = n2472 & n2635 ;
  assign n22098 = x96 & ~n5313 ;
  assign n22099 = ( ~n15515 & n15992 ) | ( ~n15515 & n17283 ) | ( n15992 & n17283 ) ;
  assign n22100 = n22099 ^ n12657 ^ n4521 ;
  assign n22101 = n299 | n5508 ;
  assign n22102 = n7308 & ~n22101 ;
  assign n22103 = ~n10309 & n22102 ;
  assign n22104 = n12519 ^ n3689 ^ 1'b0 ;
  assign n22105 = n21943 ^ n1218 ^ n201 ;
  assign n22106 = n22105 ^ n10992 ^ n4664 ;
  assign n22107 = n22106 ^ n10610 ^ 1'b0 ;
  assign n22108 = n15254 ^ n4644 ^ 1'b0 ;
  assign n22109 = ~n8557 & n22108 ;
  assign n22110 = n12805 & ~n19024 ;
  assign n22111 = n22110 ^ n8507 ^ 1'b0 ;
  assign n22112 = ~n7468 & n16109 ;
  assign n22114 = n20007 ^ n4749 ^ n1856 ;
  assign n22113 = ~n3113 & n8301 ;
  assign n22115 = n22114 ^ n22113 ^ n17096 ;
  assign n22116 = n17960 ^ n1343 ^ n528 ;
  assign n22117 = ~n661 & n21424 ;
  assign n22118 = n2109 & n3340 ;
  assign n22119 = n22118 ^ n5477 ^ n1680 ;
  assign n22120 = ~n9583 & n11751 ;
  assign n22121 = n5786 & n22120 ;
  assign n22122 = n3263 | n13612 ;
  assign n22123 = n12789 | n22122 ;
  assign n22124 = n12425 ^ n4239 ^ 1'b0 ;
  assign n22125 = ~n14744 & n22124 ;
  assign n22126 = n10352 ^ n7216 ^ 1'b0 ;
  assign n22127 = ( n7438 & n11061 ) | ( n7438 & ~n22126 ) | ( n11061 & ~n22126 ) ;
  assign n22128 = ( n576 & n8084 ) | ( n576 & ~n10376 ) | ( n8084 & ~n10376 ) ;
  assign n22129 = n19405 ^ n6198 ^ n1113 ;
  assign n22130 = n11125 | n15088 ;
  assign n22131 = n4010 ^ n1850 ^ n848 ;
  assign n22132 = ~n1952 & n22131 ;
  assign n22133 = n22130 & n22132 ;
  assign n22134 = n11631 ^ n5024 ^ 1'b0 ;
  assign n22135 = n3631 | n10652 ;
  assign n22136 = ~n15867 & n22135 ;
  assign n22137 = n867 & ~n22136 ;
  assign n22138 = n2195 & n13973 ;
  assign n22139 = n22138 ^ n13951 ^ 1'b0 ;
  assign n22140 = n1371 ^ n1143 ^ 1'b0 ;
  assign n22141 = ( n1438 & n11327 ) | ( n1438 & n21115 ) | ( n11327 & n21115 ) ;
  assign n22142 = n811 | n17072 ;
  assign n22143 = n7122 & ~n15695 ;
  assign n22144 = n22143 ^ n20139 ^ n14624 ;
  assign n22145 = n14469 | n22144 ;
  assign n22146 = n22145 ^ n3154 ^ 1'b0 ;
  assign n22147 = ~n8727 & n20305 ;
  assign n22148 = n22147 ^ n7001 ^ 1'b0 ;
  assign n22149 = n7782 ^ n1522 ^ 1'b0 ;
  assign n22150 = n22148 & n22149 ;
  assign n22151 = n22150 ^ n13088 ^ 1'b0 ;
  assign n22152 = n6751 & n16684 ;
  assign n22153 = n10173 ^ n2993 ^ 1'b0 ;
  assign n22154 = n10102 ^ n3572 ^ 1'b0 ;
  assign n22155 = n11499 & ~n22154 ;
  assign n22156 = n5289 & ~n7557 ;
  assign n22157 = n22156 ^ n12507 ^ n8936 ;
  assign n22158 = ~n4342 & n18731 ;
  assign n22159 = n22158 ^ n4870 ^ 1'b0 ;
  assign n22160 = n22159 ^ n7839 ^ 1'b0 ;
  assign n22161 = n22160 ^ n11947 ^ 1'b0 ;
  assign n22162 = n3414 & n22161 ;
  assign n22163 = n22162 ^ n3299 ^ 1'b0 ;
  assign n22164 = n1037 & ~n22163 ;
  assign n22165 = ( ~n21987 & n22157 ) | ( ~n21987 & n22164 ) | ( n22157 & n22164 ) ;
  assign n22166 = ~n7537 & n11181 ;
  assign n22167 = n22166 ^ n8138 ^ 1'b0 ;
  assign n22168 = ~n4211 & n22167 ;
  assign n22169 = n22168 ^ n18050 ^ 1'b0 ;
  assign n22170 = n10139 | n22169 ;
  assign n22171 = n12206 ^ n3856 ^ 1'b0 ;
  assign n22172 = ( n3448 & ~n8690 ) | ( n3448 & n22171 ) | ( ~n8690 & n22171 ) ;
  assign n22173 = ( n8826 & n10881 ) | ( n8826 & n15194 ) | ( n10881 & n15194 ) ;
  assign n22174 = ( n17407 & ~n22172 ) | ( n17407 & n22173 ) | ( ~n22172 & n22173 ) ;
  assign n22175 = n340 & n5174 ;
  assign n22176 = n8212 ^ n5834 ^ 1'b0 ;
  assign n22177 = n9252 & n22176 ;
  assign n22178 = n18882 ^ n12685 ^ 1'b0 ;
  assign n22179 = ~n3533 & n22178 ;
  assign n22180 = ( n16100 & n16957 ) | ( n16100 & ~n22179 ) | ( n16957 & ~n22179 ) ;
  assign n22181 = n423 & ~n1593 ;
  assign n22182 = ( n5812 & n8651 ) | ( n5812 & n22181 ) | ( n8651 & n22181 ) ;
  assign n22183 = n6925 | n8551 ;
  assign n22184 = n20782 | n22183 ;
  assign n22185 = n22184 ^ n17767 ^ n7473 ;
  assign n22186 = n18866 ^ n11515 ^ 1'b0 ;
  assign n22187 = n20842 | n22186 ;
  assign n22188 = n20097 ^ n19867 ^ 1'b0 ;
  assign n22189 = n4521 & n22188 ;
  assign n22190 = n18348 & n22189 ;
  assign n22191 = n22190 ^ n2954 ^ 1'b0 ;
  assign n22192 = n8299 ^ n4292 ^ 1'b0 ;
  assign n22193 = n8690 ^ n2617 ^ n1892 ;
  assign n22194 = n20782 ^ n5208 ^ 1'b0 ;
  assign n22195 = ( ~n6166 & n6830 ) | ( ~n6166 & n9814 ) | ( n6830 & n9814 ) ;
  assign n22196 = n22195 ^ n17523 ^ n1441 ;
  assign n22197 = ( n760 & n6483 ) | ( n760 & ~n11772 ) | ( n6483 & ~n11772 ) ;
  assign n22198 = n22197 ^ n15913 ^ 1'b0 ;
  assign n22199 = n21242 ^ n7184 ^ 1'b0 ;
  assign n22200 = ~n4618 & n22199 ;
  assign n22201 = n5986 | n17515 ;
  assign n22202 = n22201 ^ n6601 ^ 1'b0 ;
  assign n22203 = n8386 ^ n5161 ^ 1'b0 ;
  assign n22204 = n9284 ^ n1253 ^ 1'b0 ;
  assign n22205 = n22204 ^ n7182 ^ 1'b0 ;
  assign n22206 = n895 & ~n11259 ;
  assign n22207 = n4155 | n8482 ;
  assign n22208 = n22207 ^ n5992 ^ 1'b0 ;
  assign n22209 = n11682 | n22208 ;
  assign n22213 = n465 | n3332 ;
  assign n22210 = n11967 & ~n12764 ;
  assign n22211 = ~n2643 & n22210 ;
  assign n22212 = n22211 ^ n14641 ^ n3689 ;
  assign n22214 = n22213 ^ n22212 ^ n12689 ;
  assign n22215 = n22209 & ~n22214 ;
  assign n22216 = n3887 ^ n3703 ^ 1'b0 ;
  assign n22217 = n9528 | n15163 ;
  assign n22218 = n4596 & ~n22217 ;
  assign n22219 = n5926 ^ n4052 ^ 1'b0 ;
  assign n22220 = n5588 & ~n22219 ;
  assign n22221 = n22220 ^ n15035 ^ n2535 ;
  assign n22222 = n11876 | n22221 ;
  assign n22223 = n5315 & ~n22222 ;
  assign n22224 = n22213 & n22223 ;
  assign n22225 = n8691 ^ n7098 ^ 1'b0 ;
  assign n22226 = n22225 ^ n17096 ^ 1'b0 ;
  assign n22227 = ~n9676 & n22226 ;
  assign n22228 = n3824 ^ n1876 ^ 1'b0 ;
  assign n22229 = ~n18544 & n22228 ;
  assign n22230 = n14334 | n22229 ;
  assign n22231 = n3844 & ~n8176 ;
  assign n22232 = n22231 ^ n11999 ^ 1'b0 ;
  assign n22233 = ( n10012 & n15141 ) | ( n10012 & n22232 ) | ( n15141 & n22232 ) ;
  assign n22234 = n2375 ^ n2285 ^ 1'b0 ;
  assign n22235 = ~n4455 & n22234 ;
  assign n22236 = n22235 ^ n7975 ^ n4601 ;
  assign n22237 = ( n775 & n2381 ) | ( n775 & ~n7020 ) | ( n2381 & ~n7020 ) ;
  assign n22238 = ( n12244 & n22236 ) | ( n12244 & n22237 ) | ( n22236 & n22237 ) ;
  assign n22239 = n1002 | n14922 ;
  assign n22240 = n22239 ^ n12193 ^ 1'b0 ;
  assign n22245 = n5565 & n6675 ;
  assign n22246 = ~n4449 & n22245 ;
  assign n22243 = n9397 ^ n9234 ^ 1'b0 ;
  assign n22244 = ~n12366 & n22243 ;
  assign n22241 = ~n10305 & n10323 ;
  assign n22242 = n22241 ^ n2269 ^ 1'b0 ;
  assign n22247 = n22246 ^ n22244 ^ n22242 ;
  assign n22248 = ~n4839 & n22247 ;
  assign n22249 = n17741 ^ n1434 ^ 1'b0 ;
  assign n22250 = n7139 ^ n1515 ^ 1'b0 ;
  assign n22251 = n12043 | n22250 ;
  assign n22252 = n22251 ^ x101 ^ 1'b0 ;
  assign n22253 = n4372 | n22252 ;
  assign n22254 = n22253 ^ n15997 ^ n5573 ;
  assign n22255 = ~n12186 & n22254 ;
  assign n22256 = ( n846 & n14838 ) | ( n846 & ~n16131 ) | ( n14838 & ~n16131 ) ;
  assign n22257 = n13081 ^ n942 ^ 1'b0 ;
  assign n22258 = n182 & ~n22257 ;
  assign n22259 = n18420 ^ n17015 ^ n6605 ;
  assign n22260 = n16302 ^ n10010 ^ 1'b0 ;
  assign n22261 = ~n22259 & n22260 ;
  assign n22262 = ~n22258 & n22261 ;
  assign n22263 = ~n4881 & n19914 ;
  assign n22264 = ~n3850 & n15075 ;
  assign n22265 = n20334 ^ n11859 ^ 1'b0 ;
  assign n22266 = ( ~x123 & n4550 ) | ( ~x123 & n18618 ) | ( n4550 & n18618 ) ;
  assign n22267 = n12024 ^ n6191 ^ n3792 ;
  assign n22268 = ( n1839 & ~n3515 ) | ( n1839 & n3911 ) | ( ~n3515 & n3911 ) ;
  assign n22269 = ~n5439 & n22268 ;
  assign n22270 = n6785 & n7094 ;
  assign n22271 = ~n18674 & n22270 ;
  assign n22272 = n22271 ^ n9028 ^ 1'b0 ;
  assign n22273 = ~n3654 & n3939 ;
  assign n22274 = n1183 | n1990 ;
  assign n22275 = n22273 | n22274 ;
  assign n22276 = n22275 ^ n8673 ^ 1'b0 ;
  assign n22277 = n982 | n22276 ;
  assign n22278 = ~n13727 & n20215 ;
  assign n22279 = ~n9942 & n14598 ;
  assign n22280 = n22279 ^ n12847 ^ 1'b0 ;
  assign n22281 = n13813 | n16682 ;
  assign n22288 = n17811 ^ n13296 ^ n4742 ;
  assign n22283 = n1046 & n12463 ;
  assign n22284 = n3795 & ~n18051 ;
  assign n22285 = n9432 | n22284 ;
  assign n22286 = n22285 ^ n5293 ^ 1'b0 ;
  assign n22287 = ~n22283 & n22286 ;
  assign n22289 = n22288 ^ n22287 ^ 1'b0 ;
  assign n22282 = ~n11402 & n21292 ;
  assign n22290 = n22289 ^ n22282 ^ 1'b0 ;
  assign n22291 = n903 | n6394 ;
  assign n22292 = n8011 | n22291 ;
  assign n22293 = ( n1398 & ~n3019 ) | ( n1398 & n22292 ) | ( ~n3019 & n22292 ) ;
  assign n22294 = n2139 | n22293 ;
  assign n22295 = n22294 ^ n6471 ^ 1'b0 ;
  assign n22296 = n14457 & ~n20007 ;
  assign n22297 = n22296 ^ n3860 ^ 1'b0 ;
  assign n22299 = n15867 ^ n368 ^ 1'b0 ;
  assign n22298 = n5458 & ~n11604 ;
  assign n22300 = n22299 ^ n22298 ^ 1'b0 ;
  assign n22301 = n16728 ^ n5961 ^ 1'b0 ;
  assign n22302 = ~n20545 & n22301 ;
  assign n22303 = n14441 ^ n10515 ^ 1'b0 ;
  assign n22304 = n8253 & n22303 ;
  assign n22305 = n866 & n5987 ;
  assign n22306 = n22305 ^ n12697 ^ 1'b0 ;
  assign n22307 = n15594 ^ n14641 ^ 1'b0 ;
  assign n22308 = ( ~n10775 & n22306 ) | ( ~n10775 & n22307 ) | ( n22306 & n22307 ) ;
  assign n22309 = n7469 ^ n5036 ^ n3044 ;
  assign n22310 = n17901 | n22309 ;
  assign n22311 = n22310 ^ n21359 ^ 1'b0 ;
  assign n22312 = ~n5817 & n10154 ;
  assign n22313 = n22312 ^ n6587 ^ 1'b0 ;
  assign n22314 = n22313 ^ n7486 ^ 1'b0 ;
  assign n22315 = ~n1141 & n3418 ;
  assign n22316 = ~n22314 & n22315 ;
  assign n22319 = n1083 & ~n7255 ;
  assign n22320 = n22319 ^ n7953 ^ 1'b0 ;
  assign n22321 = n22320 ^ n5425 ^ n1610 ;
  assign n22322 = n9198 ^ n6955 ^ 1'b0 ;
  assign n22323 = n2361 & n22322 ;
  assign n22324 = ( n3173 & n22321 ) | ( n3173 & ~n22323 ) | ( n22321 & ~n22323 ) ;
  assign n22317 = n7549 & n9640 ;
  assign n22318 = n3945 & n22317 ;
  assign n22325 = n22324 ^ n22318 ^ 1'b0 ;
  assign n22326 = n8884 ^ n6544 ^ n5599 ;
  assign n22327 = n22326 ^ n6736 ^ 1'b0 ;
  assign n22328 = n663 & n22327 ;
  assign n22329 = n4731 ^ n1721 ^ 1'b0 ;
  assign n22330 = ~n3152 & n22329 ;
  assign n22331 = n18469 | n22330 ;
  assign n22333 = n9705 ^ n5421 ^ 1'b0 ;
  assign n22332 = n12786 & n19804 ;
  assign n22334 = n22333 ^ n22332 ^ 1'b0 ;
  assign n22335 = n7022 | n10149 ;
  assign n22338 = n1473 & n13609 ;
  assign n22339 = n22338 ^ n2290 ^ 1'b0 ;
  assign n22340 = n22339 ^ n9996 ^ 1'b0 ;
  assign n22341 = n10841 | n22340 ;
  assign n22336 = ~n7066 & n13389 ;
  assign n22337 = ~n20912 & n22336 ;
  assign n22342 = n22341 ^ n22337 ^ 1'b0 ;
  assign n22343 = n4634 & n22342 ;
  assign n22344 = n3836 & ~n15771 ;
  assign n22345 = n22344 ^ n8127 ^ 1'b0 ;
  assign n22351 = n11925 ^ n593 ^ 1'b0 ;
  assign n22352 = ~n9403 & n22351 ;
  assign n22353 = n22352 ^ n20351 ^ 1'b0 ;
  assign n22354 = n22353 ^ n9060 ^ 1'b0 ;
  assign n22346 = n2111 | n10083 ;
  assign n22347 = n22346 ^ n3320 ^ 1'b0 ;
  assign n22348 = n5783 & n14916 ;
  assign n22349 = n22348 ^ n11229 ^ 1'b0 ;
  assign n22350 = ~n22347 & n22349 ;
  assign n22355 = n22354 ^ n22350 ^ n16905 ;
  assign n22356 = ( ~n10841 & n17552 ) | ( ~n10841 & n22355 ) | ( n17552 & n22355 ) ;
  assign n22357 = n3483 ^ n809 ^ 1'b0 ;
  assign n22358 = ( n5214 & n12985 ) | ( n5214 & n22357 ) | ( n12985 & n22357 ) ;
  assign n22359 = n2512 & ~n3257 ;
  assign n22360 = ( ~n4783 & n12553 ) | ( ~n4783 & n22359 ) | ( n12553 & n22359 ) ;
  assign n22361 = n20098 ^ n3282 ^ 1'b0 ;
  assign n22362 = n6301 & n22361 ;
  assign n22363 = n4878 | n10543 ;
  assign n22364 = ~n10723 & n22363 ;
  assign n22365 = n22364 ^ n4689 ^ n1694 ;
  assign n22366 = n22365 ^ n6919 ^ n494 ;
  assign n22367 = ~n2670 & n7886 ;
  assign n22368 = n22367 ^ n15682 ^ 1'b0 ;
  assign n22369 = n22368 ^ n9923 ^ n9122 ;
  assign n22370 = n14122 ^ n8603 ^ n929 ;
  assign n22371 = ( n4448 & ~n6409 ) | ( n4448 & n22370 ) | ( ~n6409 & n22370 ) ;
  assign n22372 = n21385 ^ n19838 ^ 1'b0 ;
  assign n22373 = n4699 & ~n15303 ;
  assign n22374 = n1264 | n20525 ;
  assign n22375 = n22374 ^ x107 ^ 1'b0 ;
  assign n22376 = n22375 ^ n146 ^ 1'b0 ;
  assign n22377 = n3417 & ~n5186 ;
  assign n22378 = n21179 & n22377 ;
  assign n22379 = n11911 | n17341 ;
  assign n22380 = n16458 ^ n8716 ^ 1'b0 ;
  assign n22382 = n1126 ^ x110 ^ 1'b0 ;
  assign n22383 = x106 & n22382 ;
  assign n22384 = n22383 ^ n10562 ^ 1'b0 ;
  assign n22381 = n4837 | n5979 ;
  assign n22385 = n22384 ^ n22381 ^ n16149 ;
  assign n22386 = n15287 ^ n10867 ^ n3240 ;
  assign n22387 = n18340 & n22386 ;
  assign n22388 = n22387 ^ n15228 ^ 1'b0 ;
  assign n22389 = n22385 | n22388 ;
  assign n22390 = n4919 & ~n4962 ;
  assign n22391 = n2806 | n22390 ;
  assign n22392 = n11824 ^ n8914 ^ 1'b0 ;
  assign n22393 = n4720 & ~n22392 ;
  assign n22394 = n22393 ^ n2265 ^ 1'b0 ;
  assign n22395 = n2635 & ~n22394 ;
  assign n22396 = ~n665 & n10435 ;
  assign n22397 = n16228 ^ n4589 ^ 1'b0 ;
  assign n22398 = n21368 | n22397 ;
  assign n22399 = n22398 ^ n10878 ^ n3987 ;
  assign n22400 = n10769 ^ n7021 ^ 1'b0 ;
  assign n22401 = ~n551 & n22400 ;
  assign n22402 = ( ~n2176 & n14490 ) | ( ~n2176 & n22401 ) | ( n14490 & n22401 ) ;
  assign n22403 = n1960 & ~n4615 ;
  assign n22404 = n22402 | n22403 ;
  assign n22405 = n19185 ^ n936 ^ 1'b0 ;
  assign n22406 = ~n203 & n9362 ;
  assign n22407 = ~n18956 & n22406 ;
  assign n22408 = n21023 ^ n6775 ^ 1'b0 ;
  assign n22409 = n2440 & n22408 ;
  assign n22410 = n4552 | n6580 ;
  assign n22411 = n22410 ^ n10066 ^ n8487 ;
  assign n22412 = n22411 ^ n5789 ^ 1'b0 ;
  assign n22413 = n5384 & n22412 ;
  assign n22414 = n2965 & ~n10372 ;
  assign n22415 = n22414 ^ n11226 ^ n3376 ;
  assign n22418 = n14148 ^ n3136 ^ 1'b0 ;
  assign n22419 = n8858 & n22418 ;
  assign n22420 = ( n9892 & n12857 ) | ( n9892 & ~n22419 ) | ( n12857 & ~n22419 ) ;
  assign n22416 = n12779 ^ n641 ^ 1'b0 ;
  assign n22417 = n14803 & n22416 ;
  assign n22421 = n22420 ^ n22417 ^ 1'b0 ;
  assign n22422 = n7931 & ~n7981 ;
  assign n22423 = n12351 & n22422 ;
  assign n22424 = n18625 ^ n10698 ^ n1843 ;
  assign n22425 = n7692 ^ n477 ^ 1'b0 ;
  assign n22426 = n6376 ^ n5531 ^ 1'b0 ;
  assign n22427 = n10411 | n22426 ;
  assign n22428 = n22425 | n22427 ;
  assign n22429 = n16009 ^ n7437 ^ 1'b0 ;
  assign n22430 = n372 | n22429 ;
  assign n22431 = ( n10415 & n19282 ) | ( n10415 & n22430 ) | ( n19282 & n22430 ) ;
  assign n22432 = n13534 ^ n3122 ^ 1'b0 ;
  assign n22433 = n2151 & n5671 ;
  assign n22434 = n22433 ^ n7747 ^ 1'b0 ;
  assign n22435 = n494 | n6190 ;
  assign n22436 = n22434 | n22435 ;
  assign n22437 = n9418 & ~n16293 ;
  assign n22438 = n22437 ^ n15284 ^ 1'b0 ;
  assign n22439 = n20387 & ~n21767 ;
  assign n22440 = n15261 ^ n786 ^ 1'b0 ;
  assign n22441 = n20860 ^ n2121 ^ 1'b0 ;
  assign n22442 = n21635 | n22441 ;
  assign n22443 = n22440 & ~n22442 ;
  assign n22444 = n3279 & ~n18962 ;
  assign n22445 = ( n2000 & n3429 ) | ( n2000 & ~n22444 ) | ( n3429 & ~n22444 ) ;
  assign n22446 = n7551 & n9398 ;
  assign n22447 = n17882 & n22446 ;
  assign n22448 = ( ~n850 & n22445 ) | ( ~n850 & n22447 ) | ( n22445 & n22447 ) ;
  assign n22449 = n7087 ^ n850 ^ 1'b0 ;
  assign n22450 = n4158 ^ n928 ^ 1'b0 ;
  assign n22451 = n22283 ^ n3483 ^ 1'b0 ;
  assign n22452 = n22450 & ~n22451 ;
  assign n22453 = n1621 & ~n9385 ;
  assign n22454 = n1794 & n3193 ;
  assign n22455 = n21446 & n22454 ;
  assign n22456 = n1579 & ~n17803 ;
  assign n22457 = ( n6076 & ~n10305 ) | ( n6076 & n14239 ) | ( ~n10305 & n14239 ) ;
  assign n22458 = n18725 ^ n8166 ^ 1'b0 ;
  assign n22459 = ( ~n7296 & n19221 ) | ( ~n7296 & n22458 ) | ( n19221 & n22458 ) ;
  assign n22460 = n22459 ^ n15261 ^ n15259 ;
  assign n22461 = n2054 & n5993 ;
  assign n22462 = n22461 ^ n6030 ^ 1'b0 ;
  assign n22463 = n753 & n22462 ;
  assign n22464 = n1450 & ~n2575 ;
  assign n22465 = n15709 ^ n635 ^ 1'b0 ;
  assign n22466 = n1061 | n22465 ;
  assign n22467 = ( n3400 & n5029 ) | ( n3400 & ~n15189 ) | ( n5029 & ~n15189 ) ;
  assign n22468 = n13981 | n22467 ;
  assign n22469 = n181 & n4913 ;
  assign n22470 = ~n14462 & n22469 ;
  assign n22471 = n22470 ^ n20157 ^ 1'b0 ;
  assign n22472 = n10030 & ~n22471 ;
  assign n22473 = n9277 ^ n4452 ^ 1'b0 ;
  assign n22474 = ~n2169 & n22473 ;
  assign n22475 = ( n8574 & ~n13609 ) | ( n8574 & n22474 ) | ( ~n13609 & n22474 ) ;
  assign n22476 = n15194 ^ n7180 ^ n3805 ;
  assign n22477 = n22476 ^ n652 ^ 1'b0 ;
  assign n22478 = n4733 & ~n5078 ;
  assign n22479 = n11465 & n22478 ;
  assign n22480 = n770 & n3420 ;
  assign n22481 = n22480 ^ n20448 ^ 1'b0 ;
  assign n22482 = n22481 ^ n18924 ^ n7404 ;
  assign n22483 = n16294 ^ n5272 ^ 1'b0 ;
  assign n22484 = n22482 & n22483 ;
  assign n22485 = n22484 ^ n2991 ^ 1'b0 ;
  assign n22486 = n6547 ^ n1089 ^ 1'b0 ;
  assign n22487 = n15666 | n22486 ;
  assign n22488 = n22487 ^ n20381 ^ n8204 ;
  assign n22489 = n1917 & ~n22488 ;
  assign n22490 = n484 & n22489 ;
  assign n22491 = n14404 & ~n22490 ;
  assign n22492 = n22491 ^ n2397 ^ 1'b0 ;
  assign n22493 = n19880 ^ n8237 ^ n6818 ;
  assign n22494 = ( ~n2083 & n8550 ) | ( ~n2083 & n18772 ) | ( n8550 & n18772 ) ;
  assign n22495 = n13903 ^ n8517 ^ 1'b0 ;
  assign n22496 = n14329 ^ n2489 ^ 1'b0 ;
  assign n22497 = n3508 & n6070 ;
  assign n22498 = n22497 ^ n7945 ^ 1'b0 ;
  assign n22499 = n1556 | n22498 ;
  assign n22500 = n22499 ^ n5922 ^ 1'b0 ;
  assign n22501 = ( n617 & n8004 ) | ( n617 & n22500 ) | ( n8004 & n22500 ) ;
  assign n22502 = ~n13321 & n22501 ;
  assign n22503 = n6756 & ~n12367 ;
  assign n22504 = n9658 & n22503 ;
  assign n22505 = n22504 ^ n9201 ^ n8270 ;
  assign n22506 = n20036 & ~n22505 ;
  assign n22507 = n12665 ^ n3060 ^ 1'b0 ;
  assign n22508 = n20700 & ~n22507 ;
  assign n22509 = n18453 ^ n13878 ^ 1'b0 ;
  assign n22514 = n12195 ^ n256 ^ 1'b0 ;
  assign n22510 = n7605 ^ n422 ^ 1'b0 ;
  assign n22511 = n3718 & n22510 ;
  assign n22512 = n22511 ^ n9814 ^ n925 ;
  assign n22513 = n22512 ^ n15318 ^ n7958 ;
  assign n22515 = n22514 ^ n22513 ^ 1'b0 ;
  assign n22516 = n6667 | n11586 ;
  assign n22517 = n2990 & ~n22516 ;
  assign n22518 = n18942 ^ n9349 ^ n5793 ;
  assign n22519 = n22518 ^ n6591 ^ 1'b0 ;
  assign n22520 = n1137 | n1205 ;
  assign n22521 = n22520 ^ n7160 ^ n4370 ;
  assign n22522 = n5073 | n22521 ;
  assign n22523 = ~n6653 & n8837 ;
  assign n22524 = n16299 ^ n14149 ^ n3211 ;
  assign n22525 = ( n8929 & n22523 ) | ( n8929 & ~n22524 ) | ( n22523 & ~n22524 ) ;
  assign n22526 = n8777 & n14667 ;
  assign n22527 = n13480 | n13541 ;
  assign n22528 = n22527 ^ n10214 ^ 1'b0 ;
  assign n22529 = n22528 ^ n4742 ^ 1'b0 ;
  assign n22530 = n17130 ^ n8188 ^ 1'b0 ;
  assign n22531 = n19228 | n22530 ;
  assign n22532 = n19387 ^ n9034 ^ 1'b0 ;
  assign n22533 = n13291 & n22532 ;
  assign n22534 = n22533 ^ n10633 ^ 1'b0 ;
  assign n22535 = ~n22531 & n22534 ;
  assign n22536 = n372 | n4986 ;
  assign n22537 = n20592 ^ n2380 ^ 1'b0 ;
  assign n22538 = n22537 ^ n16340 ^ 1'b0 ;
  assign n22539 = n4657 ^ n892 ^ 1'b0 ;
  assign n22540 = ( n8138 & n13264 ) | ( n8138 & n22539 ) | ( n13264 & n22539 ) ;
  assign n22541 = n22540 ^ n19453 ^ 1'b0 ;
  assign n22542 = n10440 ^ n3978 ^ 1'b0 ;
  assign n22543 = n8845 ^ n4923 ^ n4768 ;
  assign n22544 = n12897 ^ n10438 ^ 1'b0 ;
  assign n22545 = ~n22543 & n22544 ;
  assign n22546 = ( n3847 & n11942 ) | ( n3847 & n20473 ) | ( n11942 & n20473 ) ;
  assign n22547 = n20655 & n22546 ;
  assign n22548 = n2687 | n10487 ;
  assign n22549 = n6846 | n22548 ;
  assign n22550 = x113 | n22549 ;
  assign n22551 = n18239 | n18503 ;
  assign n22552 = ~n3395 & n7928 ;
  assign n22553 = n14516 ^ n14175 ^ 1'b0 ;
  assign n22554 = n22552 & ~n22553 ;
  assign n22555 = n22554 ^ n12691 ^ n7040 ;
  assign n22556 = ( ~n1156 & n9458 ) | ( ~n1156 & n15777 ) | ( n9458 & n15777 ) ;
  assign n22557 = n2069 | n17051 ;
  assign n22558 = n1336 ^ n562 ^ 1'b0 ;
  assign n22559 = ~n1430 & n22558 ;
  assign n22560 = n13655 ^ n3074 ^ 1'b0 ;
  assign n22561 = n8304 | n22560 ;
  assign n22562 = n22559 | n22561 ;
  assign n22563 = n8838 & n12646 ;
  assign n22564 = n22563 ^ n1419 ^ 1'b0 ;
  assign n22565 = n15163 | n22564 ;
  assign n22566 = n22565 ^ n19393 ^ 1'b0 ;
  assign n22567 = ~n4486 & n22566 ;
  assign n22568 = ~n5329 & n21559 ;
  assign n22569 = n22568 ^ n3766 ^ 1'b0 ;
  assign n22570 = n12867 | n17339 ;
  assign n22571 = n15893 ^ n3146 ^ 1'b0 ;
  assign n22572 = ( n1436 & ~n21311 ) | ( n1436 & n22571 ) | ( ~n21311 & n22571 ) ;
  assign n22573 = n10212 ^ n7685 ^ n6156 ;
  assign n22574 = ( n4779 & n6821 ) | ( n4779 & ~n22573 ) | ( n6821 & ~n22573 ) ;
  assign n22575 = n10270 | n16272 ;
  assign n22576 = n6601 ^ n3337 ^ n1481 ;
  assign n22577 = n4505 & n22576 ;
  assign n22578 = n7055 & ~n22577 ;
  assign n22579 = n22578 ^ n20308 ^ 1'b0 ;
  assign n22580 = n3429 & ~n22579 ;
  assign n22581 = n20233 ^ n3931 ^ 1'b0 ;
  assign n22582 = n4854 & ~n22581 ;
  assign n22584 = n888 & n5801 ;
  assign n22585 = n19164 & n22584 ;
  assign n22586 = n16893 & ~n22585 ;
  assign n22587 = n22586 ^ n8010 ^ 1'b0 ;
  assign n22583 = n7217 & ~n15269 ;
  assign n22588 = n22587 ^ n22583 ^ 1'b0 ;
  assign n22589 = ( n4483 & n4574 ) | ( n4483 & ~n8366 ) | ( n4574 & ~n8366 ) ;
  assign n22590 = n22589 ^ n20247 ^ n6247 ;
  assign n22591 = ~n15187 & n22590 ;
  assign n22592 = n21476 ^ n18124 ^ n6108 ;
  assign n22593 = n17113 ^ n14810 ^ 1'b0 ;
  assign n22594 = n15886 ^ n8781 ^ 1'b0 ;
  assign n22595 = n22593 & ~n22594 ;
  assign n22596 = n3615 & n22595 ;
  assign n22597 = n10987 & ~n22596 ;
  assign n22598 = n22597 ^ n3578 ^ 1'b0 ;
  assign n22599 = n8668 ^ n5945 ^ 1'b0 ;
  assign n22600 = n13186 & n22599 ;
  assign n22601 = ~n6980 & n22600 ;
  assign n22602 = n14126 ^ n1936 ^ 1'b0 ;
  assign n22603 = ~n12329 & n16165 ;
  assign n22604 = ~n9983 & n13595 ;
  assign n22605 = n10959 | n22604 ;
  assign n22606 = n22605 ^ n17348 ^ n3550 ;
  assign n22607 = n6691 ^ n4884 ^ n2149 ;
  assign n22608 = n20796 ^ n270 ^ 1'b0 ;
  assign n22609 = n10317 ^ x89 ^ 1'b0 ;
  assign n22610 = n848 & ~n22609 ;
  assign n22611 = ~n148 & n22135 ;
  assign n22612 = n22611 ^ n6394 ^ 1'b0 ;
  assign n22613 = n22612 ^ n19832 ^ 1'b0 ;
  assign n22614 = n2787 ^ n878 ^ n433 ;
  assign n22615 = ( ~n12971 & n13646 ) | ( ~n12971 & n17079 ) | ( n13646 & n17079 ) ;
  assign n22616 = n3642 ^ n404 ^ 1'b0 ;
  assign n22617 = n3257 | n22616 ;
  assign n22618 = n22617 ^ n4107 ^ 1'b0 ;
  assign n22619 = n3352 & n9409 ;
  assign n22620 = n22619 ^ n5513 ^ 1'b0 ;
  assign n22621 = n770 & n22620 ;
  assign n22622 = ~n10974 & n22621 ;
  assign n22623 = n17573 & ~n18608 ;
  assign n22624 = n639 & ~n3011 ;
  assign n22625 = n22624 ^ n11836 ^ n11224 ;
  assign n22626 = n1850 & n19286 ;
  assign n22627 = n5750 & n22626 ;
  assign n22628 = n8780 | n22627 ;
  assign n22629 = n252 & n13658 ;
  assign n22630 = n3800 & n22629 ;
  assign n22631 = n13112 | n22630 ;
  assign n22632 = n22631 ^ n13457 ^ 1'b0 ;
  assign n22633 = n8686 & n22632 ;
  assign n22634 = n12612 ^ n1633 ^ 1'b0 ;
  assign n22635 = ~n16446 & n22634 ;
  assign n22636 = n19823 ^ n7663 ^ 1'b0 ;
  assign n22637 = ~n5931 & n22636 ;
  assign n22638 = n8501 & ~n21677 ;
  assign n22639 = ~n8466 & n22638 ;
  assign n22640 = n20671 ^ n16541 ^ n3874 ;
  assign n22641 = n9460 | n11693 ;
  assign n22642 = n22641 ^ n432 ^ 1'b0 ;
  assign n22643 = n3933 & n22642 ;
  assign n22644 = n22643 ^ x103 ^ 1'b0 ;
  assign n22645 = n22644 ^ n4919 ^ 1'b0 ;
  assign n22646 = n18840 ^ n12679 ^ n5301 ;
  assign n22647 = n5738 ^ n4542 ^ 1'b0 ;
  assign n22648 = n22647 ^ n3157 ^ 1'b0 ;
  assign n22649 = n5980 & ~n22648 ;
  assign n22650 = n10129 & ~n22649 ;
  assign n22651 = n8345 & ~n13565 ;
  assign n22652 = ~n12161 & n22651 ;
  assign n22653 = n3663 | n7842 ;
  assign n22654 = n22653 ^ n12664 ^ 1'b0 ;
  assign n22655 = ~n20223 & n22654 ;
  assign n22660 = n21874 ^ n2687 ^ 1'b0 ;
  assign n22661 = n2457 & ~n22660 ;
  assign n22656 = n20754 & n22229 ;
  assign n22657 = n7289 | n22656 ;
  assign n22658 = n10298 & ~n22657 ;
  assign n22659 = ( n8942 & ~n10854 ) | ( n8942 & n22658 ) | ( ~n10854 & n22658 ) ;
  assign n22662 = n22661 ^ n22659 ^ n9200 ;
  assign n22663 = n293 & ~n13575 ;
  assign n22664 = n17830 ^ n6996 ^ 1'b0 ;
  assign n22665 = n7765 & ~n13441 ;
  assign n22666 = ~n6225 & n22665 ;
  assign n22667 = ( n599 & n7725 ) | ( n599 & ~n22309 ) | ( n7725 & ~n22309 ) ;
  assign n22668 = ~n2741 & n22667 ;
  assign n22669 = n22668 ^ n7522 ^ 1'b0 ;
  assign n22670 = n19185 & n22669 ;
  assign n22671 = n14595 | n22630 ;
  assign n22672 = n13976 | n22671 ;
  assign n22673 = n22672 ^ n2586 ^ 1'b0 ;
  assign n22674 = ( n665 & n12223 ) | ( n665 & ~n21528 ) | ( n12223 & ~n21528 ) ;
  assign n22675 = n3179 & n12587 ;
  assign n22676 = n19801 & n22675 ;
  assign n22677 = n19372 ^ n911 ^ 1'b0 ;
  assign n22678 = n12297 & ~n22677 ;
  assign n22679 = n8630 ^ n3503 ^ 1'b0 ;
  assign n22680 = n8787 & n22679 ;
  assign n22681 = ( ~n868 & n2273 ) | ( ~n868 & n6260 ) | ( n2273 & n6260 ) ;
  assign n22682 = ( n4392 & n8302 ) | ( n4392 & ~n15174 ) | ( n8302 & ~n15174 ) ;
  assign n22683 = ( ~n6214 & n22681 ) | ( ~n6214 & n22682 ) | ( n22681 & n22682 ) ;
  assign n22684 = ~n4523 & n13173 ;
  assign n22685 = n22684 ^ n7059 ^ 1'b0 ;
  assign n22686 = ( n477 & ~n7022 ) | ( n477 & n22685 ) | ( ~n7022 & n22685 ) ;
  assign n22687 = n22686 ^ n17203 ^ n10951 ;
  assign n22690 = n12893 ^ n2580 ^ 1'b0 ;
  assign n22691 = n18011 | n22690 ;
  assign n22688 = ( n3044 & n9872 ) | ( n3044 & n13536 ) | ( n9872 & n13536 ) ;
  assign n22689 = ( n389 & ~n6912 ) | ( n389 & n22688 ) | ( ~n6912 & n22688 ) ;
  assign n22692 = n22691 ^ n22689 ^ n2898 ;
  assign n22693 = n22692 ^ n12830 ^ 1'b0 ;
  assign n22694 = ( ~n7638 & n11725 ) | ( ~n7638 & n22693 ) | ( n11725 & n22693 ) ;
  assign n22695 = n12768 ^ n7665 ^ n5955 ;
  assign n22696 = n5554 | n11350 ;
  assign n22697 = n18021 ^ n11150 ^ 1'b0 ;
  assign n22698 = n8528 & n22697 ;
  assign n22699 = n22698 ^ n8464 ^ 1'b0 ;
  assign n22700 = n20957 ^ n11327 ^ 1'b0 ;
  assign n22701 = n3845 | n8497 ;
  assign n22702 = n22701 ^ n2788 ^ 1'b0 ;
  assign n22703 = n1831 & n11269 ;
  assign n22705 = n21894 ^ n8603 ^ n2472 ;
  assign n22704 = n3132 & ~n3802 ;
  assign n22706 = n22705 ^ n22704 ^ 1'b0 ;
  assign n22707 = ( n7287 & n20778 ) | ( n7287 & ~n22357 ) | ( n20778 & ~n22357 ) ;
  assign n22708 = ( n2316 & n4118 ) | ( n2316 & n5370 ) | ( n4118 & n5370 ) ;
  assign n22709 = n2804 ^ n181 ^ 1'b0 ;
  assign n22710 = n15408 & ~n22709 ;
  assign n22711 = n2372 & ~n22710 ;
  assign n22712 = n22708 & n22711 ;
  assign n22713 = n8623 | n11815 ;
  assign n22714 = ~n12571 & n12750 ;
  assign n22715 = ( ~x52 & n16913 ) | ( ~x52 & n22714 ) | ( n16913 & n22714 ) ;
  assign n22716 = n9451 ^ n4478 ^ n1503 ;
  assign n22717 = n22715 | n22716 ;
  assign n22718 = ~n1819 & n3836 ;
  assign n22719 = ~n19397 & n22718 ;
  assign n22720 = ( ~n4035 & n6702 ) | ( ~n4035 & n16674 ) | ( n6702 & n16674 ) ;
  assign n22721 = n3987 | n15169 ;
  assign n22722 = n22721 ^ n8154 ^ 1'b0 ;
  assign n22723 = n14876 ^ n9495 ^ n2873 ;
  assign n22724 = n19909 ^ n7110 ^ n6272 ;
  assign n22725 = n6872 ^ n6551 ^ 1'b0 ;
  assign n22726 = n22725 ^ n12593 ^ n4878 ;
  assign n22727 = n20222 ^ n8347 ^ 1'b0 ;
  assign n22728 = n932 & ~n22727 ;
  assign n22734 = n4833 ^ n4787 ^ 1'b0 ;
  assign n22731 = n10794 ^ n9880 ^ 1'b0 ;
  assign n22732 = n2576 & n22731 ;
  assign n22729 = n5333 ^ n254 ^ 1'b0 ;
  assign n22730 = ~n3327 & n22729 ;
  assign n22733 = n22732 ^ n22730 ^ 1'b0 ;
  assign n22735 = n22734 ^ n22733 ^ 1'b0 ;
  assign n22736 = n16785 ^ n13912 ^ 1'b0 ;
  assign n22737 = ~n21788 & n22736 ;
  assign n22738 = n17567 ^ n11238 ^ 1'b0 ;
  assign n22739 = n9473 | n22738 ;
  assign n22741 = n3254 ^ n491 ^ 1'b0 ;
  assign n22742 = n1035 & ~n22741 ;
  assign n22743 = n22742 ^ n14697 ^ 1'b0 ;
  assign n22744 = ~n10519 & n22743 ;
  assign n22740 = ~n8523 & n16997 ;
  assign n22745 = n22744 ^ n22740 ^ 1'b0 ;
  assign n22746 = n5753 | n19649 ;
  assign n22747 = n16710 & ~n22746 ;
  assign n22748 = n21618 ^ n9193 ^ 1'b0 ;
  assign n22749 = n22747 | n22748 ;
  assign n22750 = ( n3006 & ~n4589 ) | ( n3006 & n12573 ) | ( ~n4589 & n12573 ) ;
  assign n22751 = n13025 ^ n9575 ^ 1'b0 ;
  assign n22752 = ~n22750 & n22751 ;
  assign n22753 = ~n21200 & n21766 ;
  assign n22754 = n6264 ^ n2146 ^ 1'b0 ;
  assign n22755 = n822 | n22754 ;
  assign n22756 = n13582 | n22755 ;
  assign n22757 = n22756 ^ n12805 ^ n10173 ;
  assign n22759 = n2949 & ~n6458 ;
  assign n22760 = n22759 ^ n2212 ^ 1'b0 ;
  assign n22758 = n5726 & n12845 ;
  assign n22761 = n22760 ^ n22758 ^ 1'b0 ;
  assign n22762 = n818 & n7508 ;
  assign n22763 = ~n10645 & n22762 ;
  assign n22764 = n22763 ^ n4768 ^ 1'b0 ;
  assign n22765 = n16056 | n22764 ;
  assign n22766 = n997 & n9116 ;
  assign n22767 = n12040 ^ x9 ^ 1'b0 ;
  assign n22768 = ~n22766 & n22767 ;
  assign n22769 = ~n11044 & n17868 ;
  assign n22770 = n22769 ^ n14455 ^ 1'b0 ;
  assign n22771 = n1917 & n5669 ;
  assign n22772 = n22771 ^ n18512 ^ n18125 ;
  assign n22777 = n1502 ^ n890 ^ n739 ;
  assign n22774 = n6744 | n11049 ;
  assign n22775 = n4567 | n22774 ;
  assign n22773 = n12706 ^ n2469 ^ n1696 ;
  assign n22776 = n22775 ^ n22773 ^ n5145 ;
  assign n22778 = n22777 ^ n22776 ^ n4326 ;
  assign n22779 = n22260 ^ n9743 ^ 1'b0 ;
  assign n22780 = ( n1107 & n3767 ) | ( n1107 & n4073 ) | ( n3767 & n4073 ) ;
  assign n22781 = n14591 & n22780 ;
  assign n22782 = n2047 & n8158 ;
  assign n22783 = n22782 ^ n11541 ^ 1'b0 ;
  assign n22784 = n22783 ^ n22474 ^ n10775 ;
  assign n22785 = n1943 ^ n1298 ^ 1'b0 ;
  assign n22786 = ~n22784 & n22785 ;
  assign n22787 = n8690 ^ n601 ^ 1'b0 ;
  assign n22788 = n1170 | n17395 ;
  assign n22789 = n7221 & ~n22788 ;
  assign n22790 = ~n15702 & n22789 ;
  assign n22791 = n22790 ^ n13262 ^ n7573 ;
  assign n22792 = n17203 & ~n20375 ;
  assign n22793 = ( n504 & n5246 ) | ( n504 & ~n5677 ) | ( n5246 & ~n5677 ) ;
  assign n22794 = n22793 ^ n21708 ^ n14338 ;
  assign n22795 = n11893 ^ n7582 ^ 1'b0 ;
  assign n22796 = n1116 & ~n1680 ;
  assign n22797 = n22713 ^ n579 ^ 1'b0 ;
  assign n22798 = n22796 & ~n22797 ;
  assign n22799 = ~n2106 & n5753 ;
  assign n22800 = n22799 ^ n12866 ^ 1'b0 ;
  assign n22801 = ( x40 & ~n14915 ) | ( x40 & n19853 ) | ( ~n14915 & n19853 ) ;
  assign n22802 = ( n6073 & n11182 ) | ( n6073 & ~n12687 ) | ( n11182 & ~n12687 ) ;
  assign n22803 = n8793 ^ n844 ^ 1'b0 ;
  assign n22804 = n5046 | n22803 ;
  assign n22805 = n22804 ^ n16157 ^ n3195 ;
  assign n22807 = n16678 ^ n16348 ^ n10859 ;
  assign n22806 = n11142 & n14187 ;
  assign n22808 = n22807 ^ n22806 ^ 1'b0 ;
  assign n22810 = n4065 & ~n9376 ;
  assign n22811 = n22810 ^ n4195 ^ 1'b0 ;
  assign n22812 = n6698 | n22811 ;
  assign n22813 = n21814 | n22812 ;
  assign n22814 = n7820 ^ n4158 ^ 1'b0 ;
  assign n22815 = n22813 & ~n22814 ;
  assign n22809 = n17253 | n20224 ;
  assign n22816 = n22815 ^ n22809 ^ 1'b0 ;
  assign n22817 = ~x58 & n9362 ;
  assign n22818 = n7130 & n21949 ;
  assign n22819 = n19976 & n22818 ;
  assign n22820 = n7395 & ~n15777 ;
  assign n22821 = n22820 ^ n2421 ^ 1'b0 ;
  assign n22822 = n18787 ^ n4223 ^ 1'b0 ;
  assign n22823 = ( n10765 & n13502 ) | ( n10765 & n20980 ) | ( n13502 & n20980 ) ;
  assign n22824 = ( n9655 & n22822 ) | ( n9655 & n22823 ) | ( n22822 & n22823 ) ;
  assign n22825 = n4007 & n17914 ;
  assign n22826 = n13897 ^ n9920 ^ 1'b0 ;
  assign n22827 = n6806 | n22826 ;
  assign n22828 = n22827 ^ n16007 ^ 1'b0 ;
  assign n22829 = ~n8671 & n22828 ;
  assign n22830 = n14136 ^ n1956 ^ 1'b0 ;
  assign n22831 = n5900 & n22830 ;
  assign n22832 = n22831 ^ n5043 ^ 1'b0 ;
  assign n22833 = ( n9850 & ~n10432 ) | ( n9850 & n22832 ) | ( ~n10432 & n22832 ) ;
  assign n22834 = n22420 & n22833 ;
  assign n22835 = ~n3395 & n15501 ;
  assign n22836 = n1436 | n14475 ;
  assign n22837 = n6150 & n10103 ;
  assign n22838 = ~n1132 & n22837 ;
  assign n22839 = n1545 & ~n10931 ;
  assign n22840 = n22838 & n22839 ;
  assign n22841 = n20086 ^ n2699 ^ 1'b0 ;
  assign n22842 = n9251 | n22841 ;
  assign n22843 = ( n9122 & n13014 ) | ( n9122 & n22842 ) | ( n13014 & n22842 ) ;
  assign n22845 = n865 ^ x103 ^ 1'b0 ;
  assign n22844 = ( n4094 & n8383 ) | ( n4094 & ~n17533 ) | ( n8383 & ~n17533 ) ;
  assign n22846 = n22845 ^ n22844 ^ n5467 ;
  assign n22847 = n152 & n5987 ;
  assign n22848 = n18326 ^ n17648 ^ 1'b0 ;
  assign n22849 = n383 | n22848 ;
  assign n22850 = n6380 | n20864 ;
  assign n22851 = n13517 & ~n22850 ;
  assign n22852 = n3123 & ~n5351 ;
  assign n22853 = n13635 & n22852 ;
  assign n22854 = ~n9928 & n17063 ;
  assign n22855 = n22854 ^ n10800 ^ 1'b0 ;
  assign n22856 = ( n6473 & n6934 ) | ( n6473 & n10562 ) | ( n6934 & n10562 ) ;
  assign n22859 = n5306 ^ n1854 ^ 1'b0 ;
  assign n22860 = n9044 ^ n1678 ^ 1'b0 ;
  assign n22861 = n22859 & ~n22860 ;
  assign n22857 = n5048 & n5074 ;
  assign n22858 = n17385 & n22857 ;
  assign n22862 = n22861 ^ n22858 ^ 1'b0 ;
  assign n22863 = n3935 & n11756 ;
  assign n22864 = ~n19075 & n22863 ;
  assign n22865 = ~n1528 & n13473 ;
  assign n22866 = ( n8395 & n13830 ) | ( n8395 & ~n15615 ) | ( n13830 & ~n15615 ) ;
  assign n22867 = ( ~n2867 & n5955 ) | ( ~n2867 & n15804 ) | ( n5955 & n15804 ) ;
  assign n22868 = n10391 | n22867 ;
  assign n22869 = n22868 ^ n17990 ^ n8897 ;
  assign n22870 = n22866 | n22869 ;
  assign n22871 = n22870 ^ n8656 ^ 1'b0 ;
  assign n22872 = n12534 ^ n867 ^ n865 ;
  assign n22873 = n22872 ^ n6663 ^ n431 ;
  assign n22874 = n10815 & ~n18481 ;
  assign n22875 = n22874 ^ n7995 ^ 1'b0 ;
  assign n22876 = n22875 ^ n2186 ^ 1'b0 ;
  assign n22877 = n14170 ^ n13433 ^ n3158 ;
  assign n22878 = n3931 & n4095 ;
  assign n22879 = n252 & n22878 ;
  assign n22880 = n6814 | n22879 ;
  assign n22881 = n20048 | n22880 ;
  assign n22882 = n4039 ^ n2976 ^ 1'b0 ;
  assign n22883 = n22882 ^ n17170 ^ n14459 ;
  assign n22884 = n2479 | n13242 ;
  assign n22885 = n22884 ^ n1629 ^ 1'b0 ;
  assign n22886 = n22885 ^ n3538 ^ 1'b0 ;
  assign n22887 = ~n22883 & n22886 ;
  assign n22888 = n11975 ^ n2406 ^ n1334 ;
  assign n22889 = n22888 ^ n17635 ^ 1'b0 ;
  assign n22890 = n10334 & n21023 ;
  assign n22891 = ~n7193 & n22890 ;
  assign n22892 = n22891 ^ n5740 ^ 1'b0 ;
  assign n22893 = ~n9858 & n18496 ;
  assign n22894 = n22893 ^ n7273 ^ 1'b0 ;
  assign n22895 = n2246 & ~n12872 ;
  assign n22896 = n10057 & ~n22895 ;
  assign n22897 = n21559 ^ n15930 ^ 1'b0 ;
  assign n22898 = ( n3616 & n6533 ) | ( n3616 & ~n16061 ) | ( n6533 & ~n16061 ) ;
  assign n22899 = n21092 ^ n9302 ^ n8007 ;
  assign n22900 = ( n6810 & ~n14759 ) | ( n6810 & n22899 ) | ( ~n14759 & n22899 ) ;
  assign n22901 = ~n1379 & n17215 ;
  assign n22902 = n6127 & n22901 ;
  assign n22903 = n3366 ^ n2940 ^ 1'b0 ;
  assign n22904 = ~n22902 & n22903 ;
  assign n22905 = ~n2815 & n5416 ;
  assign n22906 = n5171 ^ n296 ^ 1'b0 ;
  assign n22907 = n22905 | n22906 ;
  assign n22908 = n5439 ^ n5418 ^ 1'b0 ;
  assign n22909 = n7455 & n11553 ;
  assign n22910 = ( ~n1231 & n1732 ) | ( ~n1231 & n3035 ) | ( n1732 & n3035 ) ;
  assign n22911 = n12188 & n15067 ;
  assign n22912 = n7311 & ~n7657 ;
  assign n22913 = n22912 ^ n7466 ^ 1'b0 ;
  assign n22914 = n6053 | n10462 ;
  assign n22915 = n626 | n22914 ;
  assign n22916 = n22915 ^ n17168 ^ n13019 ;
  assign n22917 = n22913 & n22916 ;
  assign n22918 = n22913 ^ n21317 ^ n298 ;
  assign n22919 = n1882 & n4079 ;
  assign n22920 = ~n10841 & n22919 ;
  assign n22921 = n22920 ^ n9287 ^ 1'b0 ;
  assign n22922 = n22921 ^ n14759 ^ n872 ;
  assign n22923 = n2445 & n22922 ;
  assign n22924 = n22923 ^ n19760 ^ 1'b0 ;
  assign n22925 = n9380 & n22924 ;
  assign n22926 = n10277 & n22925 ;
  assign n22927 = ~n2039 & n12052 ;
  assign n22928 = ( n22918 & ~n22926 ) | ( n22918 & n22927 ) | ( ~n22926 & n22927 ) ;
  assign n22929 = n2783 & n5862 ;
  assign n22930 = n22929 ^ n5358 ^ 1'b0 ;
  assign n22931 = n22930 ^ n6611 ^ 1'b0 ;
  assign n22932 = n2645 | n11547 ;
  assign n22933 = n22932 ^ n2483 ^ 1'b0 ;
  assign n22934 = ( n18422 & ~n19698 ) | ( n18422 & n22933 ) | ( ~n19698 & n22933 ) ;
  assign n22935 = n5872 ^ n3143 ^ 1'b0 ;
  assign n22936 = n22935 ^ n10646 ^ 1'b0 ;
  assign n22937 = n20862 | n22936 ;
  assign n22938 = n3025 | n5367 ;
  assign n22939 = n19648 | n22938 ;
  assign n22940 = n16153 ^ n10795 ^ n721 ;
  assign n22941 = n11615 ^ n8931 ^ 1'b0 ;
  assign n22942 = ( ~n1754 & n19612 ) | ( ~n1754 & n22941 ) | ( n19612 & n22941 ) ;
  assign n22943 = n19430 ^ n16809 ^ n15650 ;
  assign n22944 = n20054 ^ n1188 ^ 1'b0 ;
  assign n22945 = n3594 & n5701 ;
  assign n22946 = n22945 ^ n3874 ^ 1'b0 ;
  assign n22947 = n2536 & ~n22946 ;
  assign n22948 = ~n14600 & n22947 ;
  assign n22949 = n18211 ^ n15654 ^ 1'b0 ;
  assign n22950 = n9476 & n14650 ;
  assign n22951 = n22950 ^ n5821 ^ 1'b0 ;
  assign n22952 = ( n7616 & ~n8032 ) | ( n7616 & n11562 ) | ( ~n8032 & n11562 ) ;
  assign n22953 = n7075 | n22952 ;
  assign n22955 = n17121 ^ n968 ^ 1'b0 ;
  assign n22956 = n17107 & n22955 ;
  assign n22954 = n11170 | n17548 ;
  assign n22957 = n22956 ^ n22954 ^ 1'b0 ;
  assign n22958 = n22957 ^ n11964 ^ 1'b0 ;
  assign n22959 = ~n22953 & n22958 ;
  assign n22960 = ~n299 & n3608 ;
  assign n22961 = ~n624 & n22780 ;
  assign n22962 = n22961 ^ n15867 ^ 1'b0 ;
  assign n22963 = n10618 ^ n7587 ^ 1'b0 ;
  assign n22964 = n4331 & ~n22963 ;
  assign n22965 = n22964 ^ n13488 ^ 1'b0 ;
  assign n22966 = ( ~n6166 & n22962 ) | ( ~n6166 & n22965 ) | ( n22962 & n22965 ) ;
  assign n22967 = n5743 & ~n11967 ;
  assign n22970 = x125 & n6242 ;
  assign n22971 = n22970 ^ n18963 ^ n3012 ;
  assign n22968 = n10678 ^ n4701 ^ 1'b0 ;
  assign n22969 = ~n5615 & n22968 ;
  assign n22972 = n22971 ^ n22969 ^ n14119 ;
  assign n22973 = n5500 ^ n2618 ^ 1'b0 ;
  assign n22974 = n6547 | n12053 ;
  assign n22975 = n6083 & ~n14694 ;
  assign n22976 = n22975 ^ n197 ^ 1'b0 ;
  assign n22977 = n22830 & ~n22976 ;
  assign n22978 = n20416 & n22977 ;
  assign n22979 = n1740 & ~n22978 ;
  assign n22982 = ~n10624 & n13929 ;
  assign n22983 = n22982 ^ n5646 ^ 1'b0 ;
  assign n22980 = ~n522 & n21114 ;
  assign n22981 = n6716 & ~n22980 ;
  assign n22984 = n22983 ^ n22981 ^ 1'b0 ;
  assign n22986 = n3604 & ~n3879 ;
  assign n22987 = n22986 ^ n10912 ^ 1'b0 ;
  assign n22985 = n3688 ^ n2136 ^ n1501 ;
  assign n22988 = n22987 ^ n22985 ^ 1'b0 ;
  assign n22989 = n9175 ^ n6705 ^ 1'b0 ;
  assign n22990 = n16261 ^ n2285 ^ 1'b0 ;
  assign n22991 = n18945 ^ n17784 ^ 1'b0 ;
  assign n22992 = ~n11836 & n22991 ;
  assign n22993 = ( ~n9439 & n13246 ) | ( ~n9439 & n16767 ) | ( n13246 & n16767 ) ;
  assign n22994 = ( n11048 & ~n12058 ) | ( n11048 & n17708 ) | ( ~n12058 & n17708 ) ;
  assign n22995 = n1132 & ~n2397 ;
  assign n22996 = n7932 & n8663 ;
  assign n22997 = n7456 & n8406 ;
  assign n22998 = n6255 & n22997 ;
  assign n22999 = n11752 ^ n10080 ^ 1'b0 ;
  assign n23000 = n3677 & ~n8210 ;
  assign n23001 = n23000 ^ n2928 ^ 1'b0 ;
  assign n23003 = n1480 & n15980 ;
  assign n23004 = n23003 ^ n3554 ^ 1'b0 ;
  assign n23005 = n3868 & n23004 ;
  assign n23006 = ~n4150 & n23005 ;
  assign n23002 = n14466 & ~n18437 ;
  assign n23007 = n23006 ^ n23002 ^ n10959 ;
  assign n23008 = n22235 ^ n14585 ^ 1'b0 ;
  assign n23009 = n3694 & n7581 ;
  assign n23010 = n15738 & ~n23009 ;
  assign n23011 = n23010 ^ n12307 ^ 1'b0 ;
  assign n23012 = x11 & n3658 ;
  assign n23013 = n2431 | n20646 ;
  assign n23014 = n7987 ^ n1268 ^ 1'b0 ;
  assign n23015 = n20237 & n23014 ;
  assign n23016 = n23015 ^ n4661 ^ 1'b0 ;
  assign n23017 = n3387 & ~n23016 ;
  assign n23018 = ( n6825 & n9841 ) | ( n6825 & n20100 ) | ( n9841 & n20100 ) ;
  assign n23021 = n1433 ^ x112 ^ 1'b0 ;
  assign n23022 = n1358 | n23021 ;
  assign n23023 = n23022 ^ n4935 ^ n4044 ;
  assign n23019 = n852 & ~n5741 ;
  assign n23020 = n17533 & n23019 ;
  assign n23024 = n23023 ^ n23020 ^ n1523 ;
  assign n23025 = ~n2467 & n8307 ;
  assign n23026 = n23025 ^ n12946 ^ n10132 ;
  assign n23027 = n2956 & ~n4792 ;
  assign n23028 = ~n10430 & n23027 ;
  assign n23029 = n7224 & ~n19762 ;
  assign n23030 = n3371 & ~n8426 ;
  assign n23031 = n9579 & n10498 ;
  assign n23032 = ~n1556 & n23031 ;
  assign n23033 = n23032 ^ n12930 ^ n2751 ;
  assign n23034 = n8018 | n13604 ;
  assign n23035 = ( n8523 & n23033 ) | ( n8523 & n23034 ) | ( n23033 & n23034 ) ;
  assign n23036 = n16183 ^ n4370 ^ 1'b0 ;
  assign n23037 = n1143 | n23036 ;
  assign n23038 = n23037 ^ n18703 ^ 1'b0 ;
  assign n23039 = ~n11599 & n14967 ;
  assign n23040 = n1349 & n23039 ;
  assign n23041 = n1818 & n11576 ;
  assign n23042 = ~n12174 & n23041 ;
  assign n23043 = n23042 ^ n4787 ^ 1'b0 ;
  assign n23044 = ~n4982 & n14418 ;
  assign n23045 = n2365 | n6454 ;
  assign n23046 = ~n10758 & n23045 ;
  assign n23047 = ~n23044 & n23046 ;
  assign n23048 = n6669 ^ n3636 ^ 1'b0 ;
  assign n23049 = n3349 & n23048 ;
  assign n23050 = ( n4144 & n4387 ) | ( n4144 & ~n9037 ) | ( n4387 & ~n9037 ) ;
  assign n23051 = ( n730 & n14691 ) | ( n730 & ~n23050 ) | ( n14691 & ~n23050 ) ;
  assign n23052 = ( ~n936 & n9119 ) | ( ~n936 & n10168 ) | ( n9119 & n10168 ) ;
  assign n23053 = n7512 ^ n340 ^ 1'b0 ;
  assign n23054 = n9961 ^ n7691 ^ 1'b0 ;
  assign n23055 = ~n771 & n23054 ;
  assign n23056 = ( n19001 & n20980 ) | ( n19001 & n23055 ) | ( n20980 & n23055 ) ;
  assign n23057 = x10 & n3398 ;
  assign n23058 = n21150 | n23057 ;
  assign n23059 = n23058 ^ n10831 ^ 1'b0 ;
  assign n23060 = n2098 & n9352 ;
  assign n23061 = n23060 ^ n22930 ^ 1'b0 ;
  assign n23062 = ~n11692 & n20611 ;
  assign n23063 = n23062 ^ n11165 ^ 1'b0 ;
  assign n23064 = ~n10952 & n23063 ;
  assign n23065 = ~n2128 & n23064 ;
  assign n23066 = n13283 ^ n7980 ^ 1'b0 ;
  assign n23067 = n1495 | n22792 ;
  assign n23068 = ( n3745 & ~n16221 ) | ( n3745 & n19937 ) | ( ~n16221 & n19937 ) ;
  assign n23071 = ~n5676 & n8908 ;
  assign n23072 = n23071 ^ n17603 ^ 1'b0 ;
  assign n23069 = n16458 & n22571 ;
  assign n23070 = n4719 & ~n23069 ;
  assign n23073 = n23072 ^ n23070 ^ n2128 ;
  assign n23074 = n4150 & ~n12720 ;
  assign n23075 = n10980 & n23074 ;
  assign n23076 = n21446 ^ n17890 ^ 1'b0 ;
  assign n23077 = n23076 ^ n8120 ^ 1'b0 ;
  assign n23078 = n7771 & n23077 ;
  assign n23079 = n14116 | n18015 ;
  assign n23080 = n18250 & ~n23079 ;
  assign n23081 = ( n146 & n4741 ) | ( n146 & n7859 ) | ( n4741 & n7859 ) ;
  assign n23082 = ( ~n3459 & n5013 ) | ( ~n3459 & n6172 ) | ( n5013 & n6172 ) ;
  assign n23083 = n4456 & ~n8045 ;
  assign n23084 = ( n23081 & ~n23082 ) | ( n23081 & n23083 ) | ( ~n23082 & n23083 ) ;
  assign n23085 = n15384 & n23084 ;
  assign n23086 = n2977 & n23085 ;
  assign n23087 = n15058 ^ n7164 ^ 1'b0 ;
  assign n23089 = ~n10360 & n13389 ;
  assign n23088 = n8154 | n13268 ;
  assign n23090 = n23089 ^ n23088 ^ n12472 ;
  assign n23091 = n5939 ^ n5811 ^ n2438 ;
  assign n23092 = n23091 ^ n8356 ^ n5400 ;
  assign n23093 = n16374 ^ n203 ^ 1'b0 ;
  assign n23094 = ~n13412 & n23093 ;
  assign n23095 = ( ~n12946 & n14620 ) | ( ~n12946 & n23094 ) | ( n14620 & n23094 ) ;
  assign n23096 = n9283 ^ n3968 ^ 1'b0 ;
  assign n23097 = n1712 & ~n23096 ;
  assign n23098 = n4607 & n23097 ;
  assign n23099 = n23098 ^ n18043 ^ 1'b0 ;
  assign n23100 = n10699 ^ n3046 ^ 1'b0 ;
  assign n23101 = n2153 & n8146 ;
  assign n23102 = n17154 | n18778 ;
  assign n23103 = n23101 | n23102 ;
  assign n23104 = n5236 ^ n4857 ^ 1'b0 ;
  assign n23105 = n11489 & ~n23104 ;
  assign n23106 = ( n1785 & n9481 ) | ( n1785 & ~n22326 ) | ( n9481 & ~n22326 ) ;
  assign n23107 = ( n18049 & n23105 ) | ( n18049 & ~n23106 ) | ( n23105 & ~n23106 ) ;
  assign n23109 = n15724 ^ n4253 ^ 1'b0 ;
  assign n23110 = ( n9262 & n12421 ) | ( n9262 & n23109 ) | ( n12421 & n23109 ) ;
  assign n23108 = ( n1680 & n7152 ) | ( n1680 & ~n12517 ) | ( n7152 & ~n12517 ) ;
  assign n23111 = n23110 ^ n23108 ^ n9376 ;
  assign n23112 = ~x127 & n14676 ;
  assign n23113 = n17736 & n23112 ;
  assign n23114 = n4950 & ~n23113 ;
  assign n23115 = n16649 ^ n3245 ^ 1'b0 ;
  assign n23116 = n23115 ^ n22393 ^ n10122 ;
  assign n23117 = n17157 ^ n7463 ^ 1'b0 ;
  assign n23118 = n12699 ^ n10940 ^ 1'b0 ;
  assign n23119 = n23117 & ~n23118 ;
  assign n23120 = ( ~n1011 & n4099 ) | ( ~n1011 & n16868 ) | ( n4099 & n16868 ) ;
  assign n23121 = n23120 ^ n4938 ^ 1'b0 ;
  assign n23122 = n19212 & ~n23121 ;
  assign n23123 = n2746 | n23122 ;
  assign n23124 = n4881 & ~n10732 ;
  assign n23125 = n19276 ^ n7432 ^ 1'b0 ;
  assign n23126 = n11564 & n23125 ;
  assign n23127 = n23126 ^ n19346 ^ n16722 ;
  assign n23128 = n1176 | n13473 ;
  assign n23129 = n23128 ^ n17555 ^ n10991 ;
  assign n23130 = n9562 ^ n247 ^ 1'b0 ;
  assign n23131 = n13221 & n20568 ;
  assign n23132 = n18778 | n22380 ;
  assign n23133 = n21043 | n23132 ;
  assign n23134 = n3027 | n7176 ;
  assign n23135 = n10040 ^ n8217 ^ 1'b0 ;
  assign n23136 = ~n5587 & n23135 ;
  assign n23137 = ~n21692 & n22320 ;
  assign n23138 = n10898 ^ n5911 ^ 1'b0 ;
  assign n23139 = n10588 & ~n23138 ;
  assign n23140 = n23139 ^ n12439 ^ 1'b0 ;
  assign n23141 = n12419 ^ n1585 ^ 1'b0 ;
  assign n23142 = n6404 & n23141 ;
  assign n23143 = ( ~n787 & n16982 ) | ( ~n787 & n23142 ) | ( n16982 & n23142 ) ;
  assign n23144 = ~n7672 & n11463 ;
  assign n23145 = ~n23143 & n23144 ;
  assign n23146 = n23145 ^ n21829 ^ n6312 ;
  assign n23147 = n2960 | n6445 ;
  assign n23148 = ( n5125 & ~n8947 ) | ( n5125 & n11430 ) | ( ~n8947 & n11430 ) ;
  assign n23149 = ~n9021 & n23148 ;
  assign n23150 = ( n3821 & n23147 ) | ( n3821 & ~n23149 ) | ( n23147 & ~n23149 ) ;
  assign n23151 = n16383 ^ n8748 ^ 1'b0 ;
  assign n23152 = n23151 ^ n1985 ^ 1'b0 ;
  assign n23153 = n5335 & ~n23152 ;
  assign n23154 = n13238 ^ n5818 ^ 1'b0 ;
  assign n23155 = n3303 & n4797 ;
  assign n23156 = n23155 ^ n5697 ^ 1'b0 ;
  assign n23157 = n6169 | n11049 ;
  assign n23158 = n23157 ^ n3592 ^ 1'b0 ;
  assign n23159 = n23158 ^ n14449 ^ n2497 ;
  assign n23160 = ( ~n1982 & n8793 ) | ( ~n1982 & n23159 ) | ( n8793 & n23159 ) ;
  assign n23161 = n21944 ^ n13953 ^ n506 ;
  assign n23162 = n1770 & n15058 ;
  assign n23163 = n23162 ^ n19699 ^ 1'b0 ;
  assign n23164 = n3730 | n6969 ;
  assign n23165 = n23164 ^ n16918 ^ 1'b0 ;
  assign n23166 = n5960 & ~n17172 ;
  assign n23167 = n17047 & n23166 ;
  assign n23168 = n8894 ^ n6918 ^ 1'b0 ;
  assign n23169 = n10068 & ~n23168 ;
  assign n23170 = n10146 & n23169 ;
  assign n23171 = n7355 ^ n2055 ^ n1029 ;
  assign n23172 = n12918 & ~n23171 ;
  assign n23173 = ~n2560 & n23172 ;
  assign n23174 = n2177 ^ n1196 ^ 1'b0 ;
  assign n23175 = n20826 & ~n23174 ;
  assign n23176 = n1918 | n3134 ;
  assign n23177 = n1591 & ~n23176 ;
  assign n23178 = n12631 & n17143 ;
  assign n23179 = n23177 & n23178 ;
  assign n23180 = ( n5269 & n20014 ) | ( n5269 & ~n23179 ) | ( n20014 & ~n23179 ) ;
  assign n23181 = ( n2247 & ~n3688 ) | ( n2247 & n20495 ) | ( ~n3688 & n20495 ) ;
  assign n23182 = n16371 ^ n3125 ^ 1'b0 ;
  assign n23183 = ~n3751 & n23182 ;
  assign n23184 = n8114 & n17072 ;
  assign n23185 = ~n4409 & n8785 ;
  assign n23186 = ~n157 & n23185 ;
  assign n23187 = n17576 & n23186 ;
  assign n23188 = n9199 & ~n16219 ;
  assign n23189 = n12493 & n23188 ;
  assign n23190 = n2470 | n23189 ;
  assign n23191 = n1728 | n23190 ;
  assign n23192 = n9605 ^ n4925 ^ 1'b0 ;
  assign n23193 = n1795 | n17057 ;
  assign n23194 = ~n22387 & n23193 ;
  assign n23195 = n12747 ^ n4450 ^ 1'b0 ;
  assign n23196 = ~n4749 & n23195 ;
  assign n23197 = ~n1091 & n13682 ;
  assign n23198 = n23197 ^ n14763 ^ 1'b0 ;
  assign n23199 = n5438 ^ n4355 ^ 1'b0 ;
  assign n23200 = n14479 & n23199 ;
  assign n23201 = n23200 ^ n4088 ^ 1'b0 ;
  assign n23202 = ( ~n528 & n10114 ) | ( ~n528 & n23201 ) | ( n10114 & n23201 ) ;
  assign n23203 = n6114 | n15676 ;
  assign n23204 = n12350 ^ n9329 ^ 1'b0 ;
  assign n23205 = ~n5687 & n23204 ;
  assign n23206 = n2773 & n23205 ;
  assign n23207 = n23206 ^ n2493 ^ 1'b0 ;
  assign n23208 = n3622 & ~n23207 ;
  assign n23209 = n23208 ^ n21839 ^ n4978 ;
  assign n23210 = n5550 | n13830 ;
  assign n23211 = n23210 ^ n13153 ^ 1'b0 ;
  assign n23212 = n6003 | n23211 ;
  assign n23213 = n10575 ^ n1929 ^ 1'b0 ;
  assign n23214 = n7618 & ~n23213 ;
  assign n23215 = n23214 ^ n5642 ^ 1'b0 ;
  assign n23216 = n10888 & n23215 ;
  assign n23217 = n8477 & n23216 ;
  assign n23218 = n5462 & ~n7739 ;
  assign n23219 = ~n9580 & n23218 ;
  assign n23220 = n9487 & n16932 ;
  assign n23224 = n13515 ^ n5404 ^ 1'b0 ;
  assign n23221 = n12901 ^ n5406 ^ 1'b0 ;
  assign n23222 = n10011 & ~n23221 ;
  assign n23223 = ( n2932 & n4915 ) | ( n2932 & n23222 ) | ( n4915 & n23222 ) ;
  assign n23225 = n23224 ^ n23223 ^ n12942 ;
  assign n23226 = n9926 ^ n9751 ^ 1'b0 ;
  assign n23227 = ( n7130 & n18230 ) | ( n7130 & ~n23226 ) | ( n18230 & ~n23226 ) ;
  assign n23228 = n20341 ^ n6012 ^ 1'b0 ;
  assign n23229 = n9173 | n23228 ;
  assign n23230 = ~n2699 & n11067 ;
  assign n23231 = n23230 ^ n18659 ^ n13132 ;
  assign n23232 = n3791 | n16320 ;
  assign n23233 = n6872 | n23232 ;
  assign n23234 = n18057 ^ n9751 ^ n9068 ;
  assign n23235 = n7636 & n23234 ;
  assign n23236 = n23235 ^ n9354 ^ 1'b0 ;
  assign n23237 = n23236 ^ n7179 ^ 1'b0 ;
  assign n23238 = n4717 ^ n2637 ^ 1'b0 ;
  assign n23239 = n958 ^ n328 ^ 1'b0 ;
  assign n23240 = n23239 ^ n9163 ^ n7837 ;
  assign n23241 = n8854 ^ n3090 ^ n2986 ;
  assign n23242 = n5655 & ~n20558 ;
  assign n23243 = n7497 & n23242 ;
  assign n23244 = ( n18058 & n23241 ) | ( n18058 & n23243 ) | ( n23241 & n23243 ) ;
  assign n23245 = ~n17486 & n23244 ;
  assign n23246 = n7177 ^ n578 ^ 1'b0 ;
  assign n23247 = ~n4574 & n7953 ;
  assign n23248 = ( n5217 & n21797 ) | ( n5217 & n23247 ) | ( n21797 & n23247 ) ;
  assign n23249 = ~n7294 & n23248 ;
  assign n23250 = n23249 ^ n6203 ^ 1'b0 ;
  assign n23251 = ( n2706 & n13232 ) | ( n2706 & n19053 ) | ( n13232 & n19053 ) ;
  assign n23252 = n16485 ^ n15056 ^ 1'b0 ;
  assign n23253 = n725 | n23252 ;
  assign n23254 = n23253 ^ n8857 ^ 1'b0 ;
  assign n23255 = n9639 & n22922 ;
  assign n23256 = n23255 ^ n10006 ^ 1'b0 ;
  assign n23257 = ~n10085 & n16457 ;
  assign n23258 = ~n9712 & n23257 ;
  assign n23259 = ( n13262 & n17451 ) | ( n13262 & ~n23258 ) | ( n17451 & ~n23258 ) ;
  assign n23260 = n16368 | n18538 ;
  assign n23261 = ( n5431 & ~n13328 ) | ( n5431 & n22717 ) | ( ~n13328 & n22717 ) ;
  assign n23262 = n4505 ^ n3574 ^ n609 ;
  assign n23263 = ( x78 & n2386 ) | ( x78 & n23262 ) | ( n2386 & n23262 ) ;
  assign n23264 = n3933 & n23263 ;
  assign n23265 = ~n13290 & n23264 ;
  assign n23266 = n23265 ^ n225 ^ 1'b0 ;
  assign n23267 = n16632 & n23266 ;
  assign n23268 = ~n6295 & n8005 ;
  assign n23269 = n5272 | n7209 ;
  assign n23270 = n6530 ^ n641 ^ 1'b0 ;
  assign n23271 = ( n15358 & n22149 ) | ( n15358 & n23270 ) | ( n22149 & n23270 ) ;
  assign n23272 = n4341 & n17115 ;
  assign n23273 = n23272 ^ n10720 ^ 1'b0 ;
  assign n23274 = ( ~n6852 & n8166 ) | ( ~n6852 & n23273 ) | ( n8166 & n23273 ) ;
  assign n23276 = ( n815 & n4336 ) | ( n815 & n18218 ) | ( n4336 & n18218 ) ;
  assign n23275 = n19247 ^ n17290 ^ 1'b0 ;
  assign n23277 = n23276 ^ n23275 ^ n7431 ;
  assign n23278 = n1723 & n13604 ;
  assign n23279 = n18033 ^ n5988 ^ 1'b0 ;
  assign n23280 = ~n23278 & n23279 ;
  assign n23281 = n12419 ^ n841 ^ 1'b0 ;
  assign n23282 = ( ~x91 & n3157 ) | ( ~x91 & n7291 ) | ( n3157 & n7291 ) ;
  assign n23283 = n16157 & ~n23282 ;
  assign n23284 = n6722 & n22761 ;
  assign n23285 = n5696 & n23284 ;
  assign n23286 = n10800 ^ n4828 ^ 1'b0 ;
  assign n23287 = n1440 | n23286 ;
  assign n23288 = n15291 ^ n4380 ^ 1'b0 ;
  assign n23289 = n17945 & n23288 ;
  assign n23290 = ( n5857 & n17692 ) | ( n5857 & ~n19000 ) | ( n17692 & ~n19000 ) ;
  assign n23291 = n23290 ^ n12637 ^ 1'b0 ;
  assign n23292 = n4361 | n6408 ;
  assign n23293 = n23292 ^ n9186 ^ 1'b0 ;
  assign n23294 = n23293 ^ n5822 ^ 1'b0 ;
  assign n23295 = n5504 | n17550 ;
  assign n23296 = n3710 & ~n9942 ;
  assign n23297 = ~n1971 & n23296 ;
  assign n23298 = n4649 & n10562 ;
  assign n23299 = n17398 ^ n3418 ^ 1'b0 ;
  assign n23300 = n4286 ^ n3803 ^ 1'b0 ;
  assign n23303 = n6646 | n21512 ;
  assign n23304 = n791 & n23303 ;
  assign n23305 = n9304 & n23304 ;
  assign n23306 = n12831 | n23305 ;
  assign n23307 = n11850 & ~n23306 ;
  assign n23301 = n21443 ^ n17057 ^ n7958 ;
  assign n23302 = n13864 & ~n23301 ;
  assign n23308 = n23307 ^ n23302 ^ 1'b0 ;
  assign n23309 = ( ~n6398 & n15222 ) | ( ~n6398 & n23308 ) | ( n15222 & n23308 ) ;
  assign n23310 = n11199 ^ n8290 ^ 1'b0 ;
  assign n23311 = n23310 ^ n234 ^ 1'b0 ;
  assign n23312 = n7715 & n23311 ;
  assign n23313 = n2595 & ~n8654 ;
  assign n23314 = ~n6638 & n12096 ;
  assign n23315 = n14957 & n23314 ;
  assign n23316 = n9170 ^ n1314 ^ n1207 ;
  assign n23317 = n23070 ^ n3694 ^ 1'b0 ;
  assign n23319 = x117 & ~n12558 ;
  assign n23320 = n23319 ^ n5973 ^ 1'b0 ;
  assign n23318 = ~n4601 & n11215 ;
  assign n23321 = n23320 ^ n23318 ^ 1'b0 ;
  assign n23322 = n345 & n8424 ;
  assign n23323 = n2767 & n23322 ;
  assign n23324 = n13702 & ~n23323 ;
  assign n23325 = n8608 ^ n7813 ^ 1'b0 ;
  assign n23326 = n256 & n23325 ;
  assign n23327 = n7918 & ~n23326 ;
  assign n23328 = ( n10553 & ~n11082 ) | ( n10553 & n23327 ) | ( ~n11082 & n23327 ) ;
  assign n23329 = n5417 ^ n3027 ^ n145 ;
  assign n23330 = n1710 | n2106 ;
  assign n23331 = n1914 & ~n20883 ;
  assign n23332 = n23331 ^ n803 ^ 1'b0 ;
  assign n23333 = n16649 ^ n8150 ^ 1'b0 ;
  assign n23334 = n15738 & n23333 ;
  assign n23335 = n22182 ^ x77 ^ 1'b0 ;
  assign n23336 = n9371 & n20936 ;
  assign n23337 = n23336 ^ n4150 ^ 1'b0 ;
  assign n23338 = ~n2668 & n5239 ;
  assign n23339 = n23338 ^ n3807 ^ 1'b0 ;
  assign n23340 = n23339 ^ n16165 ^ 1'b0 ;
  assign n23341 = n6594 & ~n23340 ;
  assign n23342 = ( n2974 & n12858 ) | ( n2974 & n13933 ) | ( n12858 & n13933 ) ;
  assign n23343 = ~n3092 & n23342 ;
  assign n23344 = n23343 ^ n5289 ^ 1'b0 ;
  assign n23345 = n12381 & ~n23344 ;
  assign n23346 = n23345 ^ n16877 ^ 1'b0 ;
  assign n23347 = n23346 ^ n21767 ^ n1563 ;
  assign n23348 = n3672 & ~n8695 ;
  assign n23349 = n2808 & n6993 ;
  assign n23350 = n23349 ^ n16393 ^ 1'b0 ;
  assign n23351 = n23350 ^ n6724 ^ n203 ;
  assign n23352 = ~n4901 & n7421 ;
  assign n23358 = n10503 ^ n1579 ^ 1'b0 ;
  assign n23353 = n10457 ^ n6239 ^ 1'b0 ;
  assign n23354 = n5312 | n23353 ;
  assign n23355 = n6591 & ~n23354 ;
  assign n23356 = ~n2927 & n23355 ;
  assign n23357 = n10644 | n23356 ;
  assign n23359 = n23358 ^ n23357 ^ 1'b0 ;
  assign n23360 = ~n882 & n14172 ;
  assign n23361 = n16470 ^ n7905 ^ 1'b0 ;
  assign n23362 = ~n14378 & n23361 ;
  assign n23363 = n23362 ^ n630 ^ 1'b0 ;
  assign n23364 = n9005 | n23363 ;
  assign n23365 = ( ~n2335 & n2872 ) | ( ~n2335 & n6179 ) | ( n2872 & n6179 ) ;
  assign n23366 = ( n5245 & n5660 ) | ( n5245 & n23365 ) | ( n5660 & n23365 ) ;
  assign n23367 = ( n5178 & n15121 ) | ( n5178 & n23366 ) | ( n15121 & n23366 ) ;
  assign n23368 = n3389 & n12552 ;
  assign n23371 = n9481 ^ n8708 ^ n4091 ;
  assign n23372 = ( ~n2193 & n6601 ) | ( ~n2193 & n23371 ) | ( n6601 & n23371 ) ;
  assign n23369 = n7455 & ~n15480 ;
  assign n23370 = n23369 ^ n22099 ^ 1'b0 ;
  assign n23373 = n23372 ^ n23370 ^ n20182 ;
  assign n23374 = n272 & ~n7986 ;
  assign n23375 = ~n14431 & n17410 ;
  assign n23376 = n23375 ^ n9878 ^ 1'b0 ;
  assign n23377 = n1996 & ~n18231 ;
  assign n23378 = n23377 ^ n12499 ^ 1'b0 ;
  assign n23379 = n4473 & n10775 ;
  assign n23383 = n1297 | n4893 ;
  assign n23384 = n11560 ^ n4175 ^ 1'b0 ;
  assign n23385 = n11665 & n23384 ;
  assign n23386 = ( ~n16384 & n23383 ) | ( ~n16384 & n23385 ) | ( n23383 & n23385 ) ;
  assign n23380 = n6022 & n6751 ;
  assign n23381 = n6304 & n23380 ;
  assign n23382 = ( ~n12118 & n18948 ) | ( ~n12118 & n23381 ) | ( n18948 & n23381 ) ;
  assign n23387 = n23386 ^ n23382 ^ n17610 ;
  assign n23388 = n10172 & ~n18835 ;
  assign n23389 = n1397 | n10190 ;
  assign n23390 = n10040 ^ n9738 ^ 1'b0 ;
  assign n23391 = n6110 & ~n20182 ;
  assign n23392 = n23391 ^ n9131 ^ 1'b0 ;
  assign n23393 = ~n8705 & n13246 ;
  assign n23394 = n1935 & n23393 ;
  assign n23395 = n23394 ^ n11327 ^ n5260 ;
  assign n23396 = n23395 ^ n9823 ^ 1'b0 ;
  assign n23397 = n4033 | n10499 ;
  assign n23398 = n20585 ^ n4050 ^ 1'b0 ;
  assign n23399 = n571 & ~n23398 ;
  assign n23400 = ~n7437 & n23399 ;
  assign n23401 = n12788 ^ n3767 ^ 1'b0 ;
  assign n23402 = n529 & ~n3329 ;
  assign n23403 = n23402 ^ n14429 ^ 1'b0 ;
  assign n23404 = n23403 ^ n21988 ^ 1'b0 ;
  assign n23405 = n15580 & n20280 ;
  assign n23406 = ( n6593 & ~n19653 ) | ( n6593 & n20136 ) | ( ~n19653 & n20136 ) ;
  assign n23407 = n23406 ^ n16921 ^ 1'b0 ;
  assign n23408 = n23044 ^ n12264 ^ 1'b0 ;
  assign n23409 = n925 | n23408 ;
  assign n23410 = n9461 | n17719 ;
  assign n23411 = n4637 | n23410 ;
  assign n23412 = n14812 & n15316 ;
  assign n23413 = n3671 ^ n387 ^ 1'b0 ;
  assign n23414 = n13232 & n23413 ;
  assign n23415 = n23414 ^ n15546 ^ 1'b0 ;
  assign n23416 = n7551 ^ n1984 ^ 1'b0 ;
  assign n23417 = n11539 ^ n9318 ^ 1'b0 ;
  assign n23418 = n13734 ^ n576 ^ 1'b0 ;
  assign n23419 = ~n23417 & n23418 ;
  assign n23420 = n23419 ^ n11625 ^ n10502 ;
  assign n23421 = n470 | n14197 ;
  assign n23422 = n23421 ^ n16673 ^ 1'b0 ;
  assign n23423 = n8478 ^ n5337 ^ x83 ;
  assign n23424 = ( n1514 & n23422 ) | ( n1514 & n23423 ) | ( n23422 & n23423 ) ;
  assign n23425 = ( n14469 & n14978 ) | ( n14469 & n18608 ) | ( n14978 & n18608 ) ;
  assign n23426 = n9240 ^ n6070 ^ 1'b0 ;
  assign n23427 = ~n3449 & n23426 ;
  assign n23428 = n10264 ^ n7184 ^ 1'b0 ;
  assign n23429 = n1384 & ~n6851 ;
  assign n23430 = ~n23428 & n23429 ;
  assign n23431 = n193 | n11560 ;
  assign n23432 = n5048 | n23431 ;
  assign n23433 = n23432 ^ n3357 ^ 1'b0 ;
  assign n23434 = n23430 | n23433 ;
  assign n23435 = n2406 & ~n5163 ;
  assign n23436 = n10323 & n23435 ;
  assign n23437 = ( n5915 & n13276 ) | ( n5915 & ~n23436 ) | ( n13276 & ~n23436 ) ;
  assign n23438 = n12357 | n14067 ;
  assign n23439 = ~n3626 & n12631 ;
  assign n23440 = n3984 & ~n23439 ;
  assign n23441 = n23440 ^ n21874 ^ 1'b0 ;
  assign n23442 = ( ~n13233 & n18128 ) | ( ~n13233 & n18363 ) | ( n18128 & n18363 ) ;
  assign n23443 = ~n11940 & n23442 ;
  assign n23444 = n4230 & n23443 ;
  assign n23445 = n4687 & n5665 ;
  assign n23446 = n19433 ^ n5293 ^ 1'b0 ;
  assign n23447 = n10732 | n23446 ;
  assign n23448 = ~x102 & n9416 ;
  assign n23449 = ( n11808 & ~n18481 ) | ( n11808 & n23448 ) | ( ~n18481 & n23448 ) ;
  assign n23450 = n7505 | n23449 ;
  assign n23451 = n23450 ^ n19227 ^ 1'b0 ;
  assign n23452 = n5643 | n9313 ;
  assign n23453 = n23451 & ~n23452 ;
  assign n23454 = n9225 ^ n7506 ^ 1'b0 ;
  assign n23455 = n152 | n23454 ;
  assign n23456 = n15204 ^ n1135 ^ 1'b0 ;
  assign n23457 = n23455 | n23456 ;
  assign n23458 = n23457 ^ n17170 ^ 1'b0 ;
  assign n23459 = n8366 ^ n7605 ^ 1'b0 ;
  assign n23460 = n8991 ^ n2055 ^ n298 ;
  assign n23461 = ( n11391 & n21352 ) | ( n11391 & n23460 ) | ( n21352 & n23460 ) ;
  assign n23462 = n15193 ^ n8165 ^ n4521 ;
  assign n23463 = n11522 & ~n12706 ;
  assign n23464 = n23463 ^ n14908 ^ n7656 ;
  assign n23465 = n193 & ~n4934 ;
  assign n23466 = n4882 ^ n2589 ^ 1'b0 ;
  assign n23467 = n2026 & ~n23466 ;
  assign n23468 = ~n6875 & n23467 ;
  assign n23469 = n6645 ^ n5591 ^ 1'b0 ;
  assign n23470 = n23468 & ~n23469 ;
  assign n23471 = n23470 ^ n438 ^ 1'b0 ;
  assign n23472 = n2026 & n18236 ;
  assign n23473 = n14578 & n23472 ;
  assign n23474 = n21280 ^ n157 ^ 1'b0 ;
  assign n23475 = n23474 ^ n15783 ^ n788 ;
  assign n23476 = ( n2860 & n15501 ) | ( n2860 & n16131 ) | ( n15501 & n16131 ) ;
  assign n23477 = ~n22286 & n23476 ;
  assign n23478 = n5784 | n14606 ;
  assign n23479 = n18147 & ~n23478 ;
  assign n23480 = n13160 ^ n1491 ^ 1'b0 ;
  assign n23481 = ~n4498 & n7318 ;
  assign n23482 = ( n6761 & n8028 ) | ( n6761 & n23481 ) | ( n8028 & n23481 ) ;
  assign n23483 = n23482 ^ n14921 ^ 1'b0 ;
  assign n23484 = n11555 & ~n23483 ;
  assign n23485 = ~n23480 & n23484 ;
  assign n23486 = n7587 ^ n2940 ^ 1'b0 ;
  assign n23487 = ~n9769 & n23486 ;
  assign n23488 = ~n1238 & n23487 ;
  assign n23489 = ~n1690 & n3931 ;
  assign n23490 = n23489 ^ n7255 ^ 1'b0 ;
  assign n23491 = ( n9169 & ~n23488 ) | ( n9169 & n23490 ) | ( ~n23488 & n23490 ) ;
  assign n23492 = n12382 ^ n3086 ^ 1'b0 ;
  assign n23493 = n23491 & n23492 ;
  assign n23494 = n23493 ^ n4300 ^ 1'b0 ;
  assign n23495 = n6552 & ~n10975 ;
  assign n23496 = n3276 ^ n2374 ^ 1'b0 ;
  assign n23497 = ( ~n6442 & n15439 ) | ( ~n6442 & n23496 ) | ( n15439 & n23496 ) ;
  assign n23498 = n3948 & ~n3967 ;
  assign n23499 = n11946 & n23498 ;
  assign n23500 = n2836 & ~n23499 ;
  assign n23501 = n23500 ^ n18827 ^ n13552 ;
  assign n23502 = n10640 & ~n18390 ;
  assign n23503 = n17900 ^ n4717 ^ 1'b0 ;
  assign n23504 = n3744 & ~n23503 ;
  assign n23505 = ( n5999 & n12576 ) | ( n5999 & n23504 ) | ( n12576 & n23504 ) ;
  assign n23506 = n23502 & n23505 ;
  assign n23507 = n731 | n13833 ;
  assign n23508 = n23507 ^ n10435 ^ 1'b0 ;
  assign n23509 = n2110 | n3876 ;
  assign n23510 = ~n6695 & n9366 ;
  assign n23511 = n23509 & n23510 ;
  assign n23512 = n12547 & ~n23511 ;
  assign n23513 = n16768 | n23512 ;
  assign n23514 = n23513 ^ n3586 ^ 1'b0 ;
  assign n23516 = n14612 ^ n10757 ^ n3485 ;
  assign n23515 = n2858 | n3072 ;
  assign n23517 = n23516 ^ n23515 ^ 1'b0 ;
  assign n23518 = n4646 & ~n20739 ;
  assign n23519 = n1591 & n23518 ;
  assign n23520 = ~n8413 & n17780 ;
  assign n23521 = n23519 & n23520 ;
  assign n23522 = ~n3552 & n6380 ;
  assign n23523 = n21287 ^ n2163 ^ 1'b0 ;
  assign n23524 = n2264 | n23523 ;
  assign n23525 = n21638 & ~n23524 ;
  assign n23526 = ( n2110 & ~n7706 ) | ( n2110 & n16330 ) | ( ~n7706 & n16330 ) ;
  assign n23527 = n7402 ^ n5196 ^ 1'b0 ;
  assign n23528 = n14300 ^ n6875 ^ 1'b0 ;
  assign n23529 = n19511 | n23528 ;
  assign n23530 = ( n8801 & n19133 ) | ( n8801 & n23529 ) | ( n19133 & n23529 ) ;
  assign n23531 = n9747 ^ n7076 ^ n5934 ;
  assign n23532 = n1002 & ~n15248 ;
  assign n23533 = n23532 ^ n9072 ^ 1'b0 ;
  assign n23534 = n12321 & ~n16817 ;
  assign n23535 = n23534 ^ n16310 ^ 1'b0 ;
  assign n23536 = n8118 ^ n4802 ^ 1'b0 ;
  assign n23537 = n23535 & ~n23536 ;
  assign n23538 = ~n4483 & n17852 ;
  assign n23539 = n23538 ^ n3372 ^ 1'b0 ;
  assign n23540 = n16632 | n22840 ;
  assign n23541 = n23540 ^ n21197 ^ 1'b0 ;
  assign n23542 = n17939 ^ n5278 ^ 1'b0 ;
  assign n23543 = ( n2304 & ~n3568 ) | ( n2304 & n23542 ) | ( ~n3568 & n23542 ) ;
  assign n23544 = n1770 & ~n3850 ;
  assign n23545 = n13970 ^ n11489 ^ 1'b0 ;
  assign n23546 = ( n15275 & n23544 ) | ( n15275 & ~n23545 ) | ( n23544 & ~n23545 ) ;
  assign n23547 = n2912 & n10172 ;
  assign n23548 = n7274 & n23547 ;
  assign n23549 = n23548 ^ n8539 ^ 1'b0 ;
  assign n23550 = n5252 & ~n22393 ;
  assign n23551 = n22401 ^ n16868 ^ n8337 ;
  assign n23552 = n23551 ^ n7723 ^ 1'b0 ;
  assign n23553 = n169 & ~n588 ;
  assign n23554 = n23553 ^ n15580 ^ n2422 ;
  assign n23555 = n18786 ^ n2590 ^ 1'b0 ;
  assign n23556 = ( n12442 & n14826 ) | ( n12442 & ~n23555 ) | ( n14826 & ~n23555 ) ;
  assign n23557 = ~n13250 & n23556 ;
  assign n23558 = n20169 ^ n6607 ^ 1'b0 ;
  assign n23559 = ~n1622 & n7936 ;
  assign n23560 = n23559 ^ n7778 ^ 1'b0 ;
  assign n23561 = n5317 ^ n584 ^ 1'b0 ;
  assign n23562 = n4135 | n23561 ;
  assign n23563 = ~n9716 & n23562 ;
  assign n23564 = ~x16 & n2445 ;
  assign n23565 = n18054 ^ n7621 ^ 1'b0 ;
  assign n23566 = n5586 & ~n23565 ;
  assign n23567 = n9184 ^ n9144 ^ 1'b0 ;
  assign n23568 = n11400 | n23567 ;
  assign n23569 = n11071 ^ n4207 ^ 1'b0 ;
  assign n23570 = n2822 & ~n23569 ;
  assign n23571 = n4941 ^ n4751 ^ 1'b0 ;
  assign n23572 = n8304 | n23571 ;
  assign n23573 = ( ~n17308 & n23570 ) | ( ~n17308 & n23572 ) | ( n23570 & n23572 ) ;
  assign n23574 = n12307 & n13625 ;
  assign n23575 = n6394 | n6808 ;
  assign n23576 = n23575 ^ n6379 ^ 1'b0 ;
  assign n23577 = n23576 ^ n14978 ^ n11967 ;
  assign n23578 = n9381 & ~n20705 ;
  assign n23579 = n630 | n9164 ;
  assign n23580 = n13929 & ~n16504 ;
  assign n23581 = n23580 ^ n4800 ^ 1'b0 ;
  assign n23582 = ~n895 & n12706 ;
  assign n23583 = n2891 & n8444 ;
  assign n23584 = n13702 & n23583 ;
  assign n23585 = ~n4085 & n15053 ;
  assign n23586 = ~n10036 & n23585 ;
  assign n23587 = n3707 | n23586 ;
  assign n23588 = ~n2426 & n23587 ;
  assign n23589 = n18091 | n20817 ;
  assign n23590 = n13337 & ~n22742 ;
  assign n23592 = n7346 | n15239 ;
  assign n23593 = n23592 ^ n16650 ^ 1'b0 ;
  assign n23591 = n614 & n1036 ;
  assign n23594 = n23593 ^ n23591 ^ 1'b0 ;
  assign n23595 = n2296 ^ n1456 ^ 1'b0 ;
  assign n23596 = n3718 & n9619 ;
  assign n23597 = n23596 ^ n14412 ^ 1'b0 ;
  assign n23598 = n22528 ^ n7937 ^ 1'b0 ;
  assign n23599 = n23597 & n23598 ;
  assign n23600 = n11153 ^ n3587 ^ 1'b0 ;
  assign n23601 = n5155 & n23600 ;
  assign n23602 = ( n891 & ~n1259 ) | ( n891 & n5177 ) | ( ~n1259 & n5177 ) ;
  assign n23603 = n4664 & ~n23602 ;
  assign n23608 = n9557 ^ n9345 ^ 1'b0 ;
  assign n23609 = n775 & ~n17061 ;
  assign n23610 = ~n23608 & n23609 ;
  assign n23604 = ~n14551 & n20427 ;
  assign n23605 = n23604 ^ n8487 ^ 1'b0 ;
  assign n23606 = ~n3011 & n23605 ;
  assign n23607 = n23606 ^ n7537 ^ 1'b0 ;
  assign n23611 = n23610 ^ n23607 ^ n16151 ;
  assign n23612 = n4170 | n23611 ;
  assign n23613 = ( ~n2363 & n5899 ) | ( ~n2363 & n15937 ) | ( n5899 & n15937 ) ;
  assign n23615 = ~n8901 & n11893 ;
  assign n23614 = n6315 & ~n11813 ;
  assign n23616 = n23615 ^ n23614 ^ 1'b0 ;
  assign n23617 = n5378 & ~n20368 ;
  assign n23618 = ~n3025 & n23617 ;
  assign n23619 = n6905 ^ n6775 ^ n2962 ;
  assign n23625 = n8342 ^ n1573 ^ 1'b0 ;
  assign n23620 = n23033 ^ n3806 ^ 1'b0 ;
  assign n23621 = ~n9135 & n23620 ;
  assign n23622 = n6199 & n23621 ;
  assign n23623 = n23622 ^ n19615 ^ 1'b0 ;
  assign n23624 = ( n8575 & ~n10988 ) | ( n8575 & n23623 ) | ( ~n10988 & n23623 ) ;
  assign n23626 = n23625 ^ n23624 ^ n20976 ;
  assign n23627 = n17155 ^ n16864 ^ 1'b0 ;
  assign n23628 = n8417 | n9114 ;
  assign n23629 = ~n5029 & n23628 ;
  assign n23630 = n23629 ^ n7123 ^ 1'b0 ;
  assign n23631 = n17318 ^ n9647 ^ 1'b0 ;
  assign n23632 = n19943 ^ n18684 ^ n5453 ;
  assign n23633 = n4132 ^ n3745 ^ 1'b0 ;
  assign n23634 = ( n1796 & ~n2744 ) | ( n1796 & n23633 ) | ( ~n2744 & n23633 ) ;
  assign n23635 = n15835 ^ n7594 ^ n4234 ;
  assign n23636 = n23635 ^ n7324 ^ n7010 ;
  assign n23637 = n23636 ^ n5370 ^ n1470 ;
  assign n23638 = n23637 ^ n3242 ^ 1'b0 ;
  assign n23639 = ~n1718 & n8618 ;
  assign n23640 = n23639 ^ n12729 ^ 1'b0 ;
  assign n23641 = n6366 | n17134 ;
  assign n23642 = n23641 ^ n21894 ^ 1'b0 ;
  assign n23643 = n4724 & n23642 ;
  assign n23644 = n6191 ^ n3568 ^ n3389 ;
  assign n23645 = n8669 | n13593 ;
  assign n23646 = n23645 ^ n9483 ^ n295 ;
  assign n23647 = n9215 ^ n8173 ^ 1'b0 ;
  assign n23648 = n10756 & n23647 ;
  assign n23649 = n23648 ^ n10980 ^ n4402 ;
  assign n23650 = n12278 ^ n3698 ^ 1'b0 ;
  assign n23651 = ~n3452 & n5177 ;
  assign n23652 = n23651 ^ n7837 ^ 1'b0 ;
  assign n23653 = n3515 & ~n15392 ;
  assign n23654 = ~n1554 & n23653 ;
  assign n23655 = n6858 & n23654 ;
  assign n23659 = ( n2965 & ~n4513 ) | ( n2965 & n13853 ) | ( ~n4513 & n13853 ) ;
  assign n23660 = n23659 ^ n21921 ^ 1'b0 ;
  assign n23661 = ( n2425 & n2949 ) | ( n2425 & ~n15665 ) | ( n2949 & ~n15665 ) ;
  assign n23662 = n7508 & ~n23661 ;
  assign n23663 = n23660 & n23662 ;
  assign n23656 = n4424 ^ x34 ^ 1'b0 ;
  assign n23657 = n12016 & n23656 ;
  assign n23658 = n2239 & n23657 ;
  assign n23664 = n23663 ^ n23658 ^ 1'b0 ;
  assign n23665 = n6017 & n16604 ;
  assign n23666 = n19469 ^ n16799 ^ 1'b0 ;
  assign n23667 = n23665 & n23666 ;
  assign n23671 = n3450 & ~n4915 ;
  assign n23672 = n23671 ^ n4026 ^ 1'b0 ;
  assign n23670 = ( n4088 & n4394 ) | ( n4088 & ~n13298 ) | ( n4394 & ~n13298 ) ;
  assign n23668 = n14313 ^ n7910 ^ n3011 ;
  assign n23669 = ( n7546 & n21763 ) | ( n7546 & ~n23668 ) | ( n21763 & ~n23668 ) ;
  assign n23673 = n23672 ^ n23670 ^ n23669 ;
  assign n23674 = n5092 & ~n17524 ;
  assign n23677 = n12127 ^ n6986 ^ 1'b0 ;
  assign n23676 = ( n2690 & ~n10790 ) | ( n2690 & n16244 ) | ( ~n10790 & n16244 ) ;
  assign n23678 = n23677 ^ n23676 ^ n14413 ;
  assign n23675 = ~n423 & n6367 ;
  assign n23679 = n23678 ^ n23675 ^ 1'b0 ;
  assign n23680 = n13114 & n23679 ;
  assign n23681 = n23680 ^ n6220 ^ 1'b0 ;
  assign n23682 = n313 & ~n808 ;
  assign n23683 = n23682 ^ n14109 ^ 1'b0 ;
  assign n23684 = n15994 ^ n10342 ^ 1'b0 ;
  assign n23685 = ~n8904 & n23684 ;
  assign n23686 = ( n12558 & n13237 ) | ( n12558 & n23685 ) | ( n13237 & n23685 ) ;
  assign n23687 = ( n5392 & ~n6148 ) | ( n5392 & n8611 ) | ( ~n6148 & n8611 ) ;
  assign n23688 = ( ~n941 & n4149 ) | ( ~n941 & n23687 ) | ( n4149 & n23687 ) ;
  assign n23689 = n23688 ^ n5421 ^ x2 ;
  assign n23690 = n11331 ^ n10424 ^ 1'b0 ;
  assign n23691 = ~n6479 & n11873 ;
  assign n23692 = ~n4261 & n23691 ;
  assign n23693 = n21923 & ~n23692 ;
  assign n23694 = ~n10158 & n23693 ;
  assign n23695 = n11433 ^ n7614 ^ n2641 ;
  assign n23696 = n17919 & n23695 ;
  assign n23697 = ~n206 & n23696 ;
  assign n23698 = n11693 | n18583 ;
  assign n23699 = n23698 ^ n7060 ^ 1'b0 ;
  assign n23700 = x113 & ~n2304 ;
  assign n23701 = n895 | n6638 ;
  assign n23702 = n2272 & ~n23701 ;
  assign n23703 = ( n324 & n11693 ) | ( n324 & n13532 ) | ( n11693 & n13532 ) ;
  assign n23704 = n23703 ^ n4634 ^ n4472 ;
  assign n23705 = ~n4050 & n23704 ;
  assign n23706 = n17518 & n23705 ;
  assign n23707 = n13876 & n23706 ;
  assign n23708 = ( ~n992 & n19956 ) | ( ~n992 & n23707 ) | ( n19956 & n23707 ) ;
  assign n23709 = ( n3486 & ~n4487 ) | ( n3486 & n7083 ) | ( ~n4487 & n7083 ) ;
  assign n23710 = n5634 | n18286 ;
  assign n23711 = n9087 | n23710 ;
  assign n23712 = n23709 | n23711 ;
  assign n23713 = n2377 & n6701 ;
  assign n23714 = n23713 ^ n6741 ^ 1'b0 ;
  assign n23715 = n9477 | n23714 ;
  assign n23716 = n20066 ^ n12942 ^ 1'b0 ;
  assign n23717 = n19877 & ~n23716 ;
  assign n23718 = n6865 & n8569 ;
  assign n23719 = ( ~n7486 & n12215 ) | ( ~n7486 & n22754 ) | ( n12215 & n22754 ) ;
  assign n23720 = n17260 ^ n4126 ^ 1'b0 ;
  assign n23721 = n23720 ^ n7379 ^ 1'b0 ;
  assign n23722 = n23719 | n23721 ;
  assign n23727 = n3932 ^ n2011 ^ 1'b0 ;
  assign n23728 = n3016 & ~n23727 ;
  assign n23724 = n5191 ^ n4618 ^ n2464 ;
  assign n23723 = n594 & n16425 ;
  assign n23725 = n23724 ^ n23723 ^ 1'b0 ;
  assign n23726 = n23725 ^ n21233 ^ n3789 ;
  assign n23729 = n23728 ^ n23726 ^ 1'b0 ;
  assign n23730 = n8578 ^ n5823 ^ 1'b0 ;
  assign n23731 = n13539 ^ n9042 ^ 1'b0 ;
  assign n23732 = n23731 ^ n10515 ^ n10036 ;
  assign n23734 = ( n478 & n1080 ) | ( n478 & n1173 ) | ( n1080 & n1173 ) ;
  assign n23735 = n23734 ^ n2776 ^ n1649 ;
  assign n23733 = ( ~n1898 & n14048 ) | ( ~n1898 & n18958 ) | ( n14048 & n18958 ) ;
  assign n23736 = n23735 ^ n23733 ^ n2743 ;
  assign n23737 = ( n4434 & n6560 ) | ( n4434 & n23736 ) | ( n6560 & n23736 ) ;
  assign n23738 = n23737 ^ n18572 ^ 1'b0 ;
  assign n23739 = ~n6671 & n23738 ;
  assign n23740 = ( n8601 & n14671 ) | ( n8601 & n17242 ) | ( n14671 & n17242 ) ;
  assign n23741 = ( n1143 & n22623 ) | ( n1143 & n22823 ) | ( n22623 & n22823 ) ;
  assign n23742 = n18919 ^ n377 ^ 1'b0 ;
  assign n23744 = ~n5798 & n14519 ;
  assign n23745 = n23744 ^ n6527 ^ 1'b0 ;
  assign n23743 = n10127 & ~n17893 ;
  assign n23746 = n23745 ^ n23743 ^ 1'b0 ;
  assign n23747 = n23746 ^ n19144 ^ n4122 ;
  assign n23748 = n3436 | n23747 ;
  assign n23749 = ( n5113 & n8776 ) | ( n5113 & ~n12874 ) | ( n8776 & ~n12874 ) ;
  assign n23750 = n23749 ^ n10101 ^ 1'b0 ;
  assign n23751 = n23750 ^ n8717 ^ 1'b0 ;
  assign n23752 = n11186 & ~n21543 ;
  assign n23753 = n23752 ^ n252 ^ 1'b0 ;
  assign n23754 = ~n1343 & n11572 ;
  assign n23755 = n23754 ^ n4601 ^ 1'b0 ;
  assign n23756 = n19919 ^ n3094 ^ 1'b0 ;
  assign n23757 = ~n14307 & n19618 ;
  assign n23758 = n11301 & n23757 ;
  assign n23759 = n13699 ^ n4049 ^ n1441 ;
  assign n23760 = n2159 & n5938 ;
  assign n23761 = ~n2159 & n23760 ;
  assign n23762 = n5310 | n23761 ;
  assign n23763 = n15121 | n23762 ;
  assign n23764 = n9667 | n9933 ;
  assign n23765 = n23763 | n23764 ;
  assign n23766 = ~n8430 & n23765 ;
  assign n23767 = n23766 ^ n23310 ^ 1'b0 ;
  assign n23768 = n2176 | n23767 ;
  assign n23769 = n9393 | n23768 ;
  assign n23770 = ( n12472 & n21743 ) | ( n12472 & n23769 ) | ( n21743 & n23769 ) ;
  assign n23771 = n20352 & ~n23273 ;
  assign n23772 = n12656 & n17553 ;
  assign n23773 = n1610 & n23772 ;
  assign n23774 = n5545 ^ n4065 ^ 1'b0 ;
  assign n23775 = ~n9633 & n23774 ;
  assign n23776 = n10387 ^ n2454 ^ 1'b0 ;
  assign n23777 = n23776 ^ n4778 ^ 1'b0 ;
  assign n23778 = n7552 | n23777 ;
  assign n23779 = n3983 ^ n2106 ^ 1'b0 ;
  assign n23780 = n23779 ^ n10949 ^ n9443 ;
  assign n23781 = n22630 ^ n1776 ^ 1'b0 ;
  assign n23782 = n23780 & n23781 ;
  assign n23783 = n19624 ^ n2233 ^ 1'b0 ;
  assign n23784 = n18021 ^ n7091 ^ 1'b0 ;
  assign n23785 = ~n3615 & n5263 ;
  assign n23786 = n23785 ^ n4695 ^ 1'b0 ;
  assign n23787 = n4216 & ~n23786 ;
  assign n23788 = ~n16344 & n23787 ;
  assign n23789 = n4588 & ~n14424 ;
  assign n23790 = ~n16835 & n23789 ;
  assign n23791 = n11676 ^ n2893 ^ 1'b0 ;
  assign n23792 = n18569 | n23791 ;
  assign n23793 = n12561 ^ n238 ^ 1'b0 ;
  assign n23794 = n5548 & n23793 ;
  assign n23795 = n2717 & n23794 ;
  assign n23796 = n20128 ^ n11514 ^ 1'b0 ;
  assign n23797 = ( ~n7254 & n10956 ) | ( ~n7254 & n14221 ) | ( n10956 & n14221 ) ;
  assign n23798 = n23797 ^ n21394 ^ 1'b0 ;
  assign n23799 = ~n10757 & n13291 ;
  assign n23800 = n23799 ^ n6978 ^ 1'b0 ;
  assign n23801 = n23800 ^ n2318 ^ 1'b0 ;
  assign n23802 = n5851 & ~n6544 ;
  assign n23803 = n23801 & n23802 ;
  assign n23804 = n6837 ^ n4620 ^ 1'b0 ;
  assign n23805 = ~n4430 & n23804 ;
  assign n23806 = n5784 & ~n11384 ;
  assign n23807 = ~n23805 & n23806 ;
  assign n23808 = n453 & n10737 ;
  assign n23809 = n23808 ^ n8047 ^ 1'b0 ;
  assign n23811 = n3350 ^ n1211 ^ 1'b0 ;
  assign n23812 = ( n11539 & n15421 ) | ( n11539 & ~n23811 ) | ( n15421 & ~n23811 ) ;
  assign n23810 = n9850 | n22479 ;
  assign n23813 = n23812 ^ n23810 ^ 1'b0 ;
  assign n23814 = n3989 | n12896 ;
  assign n23815 = n23814 ^ n1434 ^ 1'b0 ;
  assign n23816 = n23815 ^ n14257 ^ n7076 ;
  assign n23817 = n13905 ^ x67 ^ 1'b0 ;
  assign n23818 = n23817 ^ n17057 ^ n4248 ;
  assign n23819 = n20047 ^ n5092 ^ 1'b0 ;
  assign n23820 = n23819 ^ n19855 ^ n2200 ;
  assign n23821 = n18513 ^ n10074 ^ n8532 ;
  assign n23822 = x66 & ~n16703 ;
  assign n23823 = n5104 | n9111 ;
  assign n23824 = n23823 ^ n6278 ^ 1'b0 ;
  assign n23825 = n23824 ^ n3657 ^ 1'b0 ;
  assign n23826 = n2621 & n23825 ;
  assign n23827 = n5102 & n6982 ;
  assign n23828 = n4479 | n7027 ;
  assign n23829 = n10334 & ~n14415 ;
  assign n23830 = ~n23828 & n23829 ;
  assign n23831 = ~n7162 & n23830 ;
  assign n23832 = ~n1629 & n23831 ;
  assign n23833 = n1515 & n23832 ;
  assign n23834 = ~n5673 & n23833 ;
  assign n23836 = n17901 ^ n12512 ^ n7580 ;
  assign n23835 = n12511 | n15046 ;
  assign n23837 = n23836 ^ n23835 ^ 1'b0 ;
  assign n23838 = ( n19111 & n21422 ) | ( n19111 & ~n23837 ) | ( n21422 & ~n23837 ) ;
  assign n23839 = ~n9821 & n13494 ;
  assign n23840 = n23839 ^ n10824 ^ 1'b0 ;
  assign n23841 = ~n1937 & n7457 ;
  assign n23842 = n23840 & n23841 ;
  assign n23843 = n20231 & ~n23842 ;
  assign n23844 = n10661 ^ n6007 ^ 1'b0 ;
  assign n23845 = n17171 | n23844 ;
  assign n23846 = ~n10462 & n17257 ;
  assign n23847 = n12013 & ~n23846 ;
  assign n23848 = n7809 ^ n1610 ^ 1'b0 ;
  assign n23849 = n10466 & ~n23848 ;
  assign n23850 = ( n5389 & ~n8450 ) | ( n5389 & n23849 ) | ( ~n8450 & n23849 ) ;
  assign n23851 = n23850 ^ n8864 ^ n2979 ;
  assign n23852 = ( n3025 & ~n14111 ) | ( n3025 & n23851 ) | ( ~n14111 & n23851 ) ;
  assign n23853 = ( n1514 & n3027 ) | ( n1514 & n14877 ) | ( n3027 & n14877 ) ;
  assign n23854 = n5003 ^ n3816 ^ 1'b0 ;
  assign n23855 = n3745 & n23854 ;
  assign n23856 = n21240 ^ n20699 ^ 1'b0 ;
  assign n23857 = n20212 ^ n11789 ^ n5686 ;
  assign n23858 = n23857 ^ n5143 ^ n3522 ;
  assign n23859 = n1414 | n8272 ;
  assign n23860 = ( n1532 & ~n7709 ) | ( n1532 & n23859 ) | ( ~n7709 & n23859 ) ;
  assign n23861 = n12014 & ~n23860 ;
  assign n23862 = ~n18400 & n23861 ;
  assign n23863 = n19211 | n21236 ;
  assign n23864 = n3771 & n20513 ;
  assign n23865 = ~n23863 & n23864 ;
  assign n23866 = n1199 | n13358 ;
  assign n23867 = n18065 & ~n23866 ;
  assign n23868 = n3040 ^ n2663 ^ 1'b0 ;
  assign n23869 = n6949 ^ n4746 ^ 1'b0 ;
  assign n23870 = n3082 & ~n23869 ;
  assign n23871 = n20515 | n23870 ;
  assign n23872 = ( n4558 & n6385 ) | ( n4558 & n8700 ) | ( n6385 & n8700 ) ;
  assign n23873 = n8810 & n23872 ;
  assign n23874 = n23873 ^ n6058 ^ 1'b0 ;
  assign n23875 = n471 | n21454 ;
  assign n23876 = n23875 ^ n16271 ^ 1'b0 ;
  assign n23877 = n938 | n1402 ;
  assign n23878 = n23877 ^ n3887 ^ 1'b0 ;
  assign n23879 = n18878 ^ n521 ^ 1'b0 ;
  assign n23880 = ~n23878 & n23879 ;
  assign n23881 = n2865 & n4687 ;
  assign n23882 = n23881 ^ n9403 ^ 1'b0 ;
  assign n23883 = ( n3378 & n14204 ) | ( n3378 & n14362 ) | ( n14204 & n14362 ) ;
  assign n23884 = n8356 & ~n23883 ;
  assign n23885 = n3051 ^ n2415 ^ 1'b0 ;
  assign n23886 = n14560 | n23885 ;
  assign n23887 = n10496 & n20242 ;
  assign n23888 = n9205 & n23887 ;
  assign n23889 = n11165 ^ n10526 ^ n6983 ;
  assign n23890 = n16230 & n18623 ;
  assign n23891 = n23890 ^ n11776 ^ n5387 ;
  assign n23892 = n12636 ^ n5854 ^ 1'b0 ;
  assign n23894 = n143 & ~n3029 ;
  assign n23895 = ~n8004 & n23894 ;
  assign n23893 = n4329 & ~n20252 ;
  assign n23896 = n23895 ^ n23893 ^ 1'b0 ;
  assign n23897 = n9327 | n10147 ;
  assign n23898 = n23177 ^ n14907 ^ n5602 ;
  assign n23899 = ~n6317 & n23898 ;
  assign n23900 = n23899 ^ n17161 ^ 1'b0 ;
  assign n23901 = n5966 & n14265 ;
  assign n23903 = n223 & n9502 ;
  assign n23902 = x63 & ~n12497 ;
  assign n23904 = n23903 ^ n23902 ^ 1'b0 ;
  assign n23905 = ~n2873 & n23904 ;
  assign n23906 = n23901 & n23905 ;
  assign n23907 = n23906 ^ n18252 ^ 1'b0 ;
  assign n23908 = n23189 ^ n8644 ^ n3802 ;
  assign n23909 = n23270 ^ n5219 ^ n1060 ;
  assign n23910 = ~n2406 & n21337 ;
  assign n23911 = n251 & ~n1970 ;
  assign n23912 = n23911 ^ n5847 ^ 1'b0 ;
  assign n23913 = ( ~n8021 & n23910 ) | ( ~n8021 & n23912 ) | ( n23910 & n23912 ) ;
  assign n23914 = ~n2137 & n8637 ;
  assign n23915 = n2504 ^ n1221 ^ 1'b0 ;
  assign n23916 = n22131 & n23915 ;
  assign n23920 = n16995 & ~n20136 ;
  assign n23917 = n12785 & ~n16031 ;
  assign n23918 = n23917 ^ n4013 ^ 1'b0 ;
  assign n23919 = n1967 | n23918 ;
  assign n23921 = n23920 ^ n23919 ^ 1'b0 ;
  assign n23922 = n14620 | n22897 ;
  assign n23923 = n23922 ^ n11709 ^ 1'b0 ;
  assign n23924 = ( ~n2669 & n2731 ) | ( ~n2669 & n16025 ) | ( n2731 & n16025 ) ;
  assign n23925 = ( n5717 & n7318 ) | ( n5717 & n16312 ) | ( n7318 & n16312 ) ;
  assign n23926 = n9085 ^ n1331 ^ n279 ;
  assign n23927 = n4392 | n8731 ;
  assign n23928 = n20018 | n23927 ;
  assign n23929 = n2344 | n23928 ;
  assign n23930 = n16587 ^ n6806 ^ 1'b0 ;
  assign n23931 = n3752 | n23930 ;
  assign n23932 = n17377 ^ n12778 ^ 1'b0 ;
  assign n23933 = n17841 ^ n15781 ^ 1'b0 ;
  assign n23934 = n21769 ^ n20572 ^ n17154 ;
  assign n23935 = n15208 ^ n8140 ^ 1'b0 ;
  assign n23936 = ( ~n2597 & n13693 ) | ( ~n2597 & n17107 ) | ( n13693 & n17107 ) ;
  assign n23937 = n12612 & n23936 ;
  assign n23938 = n23937 ^ n2927 ^ 1'b0 ;
  assign n23939 = n7986 & ~n23938 ;
  assign n23940 = n11374 ^ n5022 ^ 1'b0 ;
  assign n23941 = n23265 & n23940 ;
  assign n23942 = n6460 & ~n9158 ;
  assign n23943 = n23942 ^ n13827 ^ 1'b0 ;
  assign n23944 = n5569 & ~n7616 ;
  assign n23946 = n12882 ^ n8176 ^ n3403 ;
  assign n23945 = n1022 & n1984 ;
  assign n23947 = n23946 ^ n23945 ^ 1'b0 ;
  assign n23948 = n13916 & n14311 ;
  assign n23949 = n4414 & n18753 ;
  assign n23950 = n10850 ^ n10594 ^ n4155 ;
  assign n23951 = n22015 ^ n3582 ^ n620 ;
  assign n23952 = n6481 & n16462 ;
  assign n23953 = n23952 ^ n11633 ^ 1'b0 ;
  assign n23954 = n14375 & n23953 ;
  assign n23955 = n6555 & n6872 ;
  assign n23956 = n23955 ^ n5559 ^ 1'b0 ;
  assign n23957 = n5299 ^ x87 ^ 1'b0 ;
  assign n23958 = ~n3088 & n11072 ;
  assign n23959 = n5169 & ~n19663 ;
  assign n23960 = n23959 ^ n21998 ^ 1'b0 ;
  assign n23961 = ( ~n1654 & n23958 ) | ( ~n1654 & n23960 ) | ( n23958 & n23960 ) ;
  assign n23962 = ~n3826 & n23961 ;
  assign n23963 = n21783 & n23962 ;
  assign n23964 = n2499 & n12099 ;
  assign n23965 = n13700 ^ n170 ^ 1'b0 ;
  assign n23966 = n5597 & ~n23965 ;
  assign n23967 = ~n23964 & n23966 ;
  assign n23968 = n3800 & ~n11467 ;
  assign n23969 = n23968 ^ n19805 ^ n4190 ;
  assign n23970 = ~n23967 & n23969 ;
  assign n23971 = ~n15093 & n23970 ;
  assign n23972 = n771 | n20643 ;
  assign n23973 = n7656 & ~n23972 ;
  assign n23974 = n8334 ^ n225 ^ 1'b0 ;
  assign n23975 = ~n12807 & n17666 ;
  assign n23976 = n7798 & n23975 ;
  assign n23977 = n22620 & n23976 ;
  assign n23978 = n23977 ^ n18958 ^ n9628 ;
  assign n23979 = n9928 | n10769 ;
  assign n23980 = ( ~n9487 & n23504 ) | ( ~n9487 & n23979 ) | ( n23504 & n23979 ) ;
  assign n23981 = ( n1528 & n18821 ) | ( n1528 & n23980 ) | ( n18821 & n23980 ) ;
  assign n23982 = n23981 ^ n3729 ^ 1'b0 ;
  assign n23984 = ~n5598 & n6511 ;
  assign n23985 = n14435 & n23984 ;
  assign n23986 = n8477 ^ x40 ^ 1'b0 ;
  assign n23987 = ( n9321 & ~n23985 ) | ( n9321 & n23986 ) | ( ~n23985 & n23986 ) ;
  assign n23983 = n11198 | n11811 ;
  assign n23988 = n23987 ^ n23983 ^ 1'b0 ;
  assign n23992 = ~n1196 & n8810 ;
  assign n23993 = n22427 & n23992 ;
  assign n23989 = n7581 & n13753 ;
  assign n23990 = n23989 ^ n6214 ^ 1'b0 ;
  assign n23991 = n11559 | n23990 ;
  assign n23994 = n23993 ^ n23991 ^ 1'b0 ;
  assign n23995 = n10609 ^ n6609 ^ n1763 ;
  assign n23996 = n23995 ^ n1249 ^ 1'b0 ;
  assign n23997 = ( n8229 & ~n9163 ) | ( n8229 & n14208 ) | ( ~n9163 & n14208 ) ;
  assign n23998 = n11589 ^ n10645 ^ n603 ;
  assign n23999 = n23997 | n23998 ;
  assign n24000 = n23996 & ~n23999 ;
  assign n24001 = n260 | n2687 ;
  assign n24002 = n15697 | n16621 ;
  assign n24003 = n673 & n9683 ;
  assign n24004 = ( ~n16480 & n21195 ) | ( ~n16480 & n24003 ) | ( n21195 & n24003 ) ;
  assign n24005 = n16028 ^ n9685 ^ 1'b0 ;
  assign n24006 = ( n2760 & ~n7444 ) | ( n2760 & n24005 ) | ( ~n7444 & n24005 ) ;
  assign n24007 = n1470 & ~n1868 ;
  assign n24008 = n24007 ^ n20264 ^ n9149 ;
  assign n24009 = n15250 ^ n2751 ^ 1'b0 ;
  assign n24010 = ( n6819 & n10016 ) | ( n6819 & ~n13898 ) | ( n10016 & ~n13898 ) ;
  assign n24011 = n24010 ^ n15974 ^ 1'b0 ;
  assign n24012 = n21702 | n24011 ;
  assign n24013 = n17039 ^ n12277 ^ 1'b0 ;
  assign n24014 = n7053 & n24013 ;
  assign n24016 = n12872 ^ n2241 ^ 1'b0 ;
  assign n24017 = n2544 | n2937 ;
  assign n24018 = n24016 & ~n24017 ;
  assign n24015 = n7631 & n8157 ;
  assign n24019 = n24018 ^ n24015 ^ 1'b0 ;
  assign n24020 = n24019 ^ n22578 ^ n5557 ;
  assign n24021 = ( ~n6203 & n10050 ) | ( ~n6203 & n15965 ) | ( n10050 & n15965 ) ;
  assign n24022 = n7232 & n19376 ;
  assign n24023 = n24022 ^ n20034 ^ 1'b0 ;
  assign n24024 = ~n18777 & n24023 ;
  assign n24025 = n3821 & n10421 ;
  assign n24026 = n24025 ^ n8501 ^ 1'b0 ;
  assign n24027 = n14464 ^ n7565 ^ n4703 ;
  assign n24028 = ( n3910 & n24026 ) | ( n3910 & ~n24027 ) | ( n24026 & ~n24027 ) ;
  assign n24029 = n18177 ^ n1710 ^ 1'b0 ;
  assign n24030 = n3094 & n24029 ;
  assign n24031 = n9514 & n16238 ;
  assign n24032 = n13503 & n24031 ;
  assign n24033 = n12691 ^ n4301 ^ 1'b0 ;
  assign n24037 = n6974 ^ n5874 ^ 1'b0 ;
  assign n24034 = n2926 ^ n1224 ^ 1'b0 ;
  assign n24035 = n9610 & n24034 ;
  assign n24036 = n19533 & n24035 ;
  assign n24038 = n24037 ^ n24036 ^ 1'b0 ;
  assign n24039 = n19345 ^ n14183 ^ 1'b0 ;
  assign n24040 = ~n11934 & n24039 ;
  assign n24041 = n19142 & n24040 ;
  assign n24042 = ~n8769 & n24041 ;
  assign n24043 = ~n3176 & n10095 ;
  assign n24044 = n19231 ^ n11827 ^ 1'b0 ;
  assign n24045 = n24043 & ~n24044 ;
  assign n24046 = ~n15588 & n17326 ;
  assign n24047 = ~n9946 & n24046 ;
  assign n24048 = n12916 ^ n1445 ^ n298 ;
  assign n24049 = n6914 ^ n2202 ^ 1'b0 ;
  assign n24050 = ~n9251 & n24049 ;
  assign n24051 = n24050 ^ n6376 ^ n1528 ;
  assign n24052 = n3965 | n11418 ;
  assign n24053 = n17391 ^ n10180 ^ x0 ;
  assign n24054 = ~n1904 & n7203 ;
  assign n24055 = n24054 ^ n5884 ^ 1'b0 ;
  assign n24056 = ~n10837 & n24055 ;
  assign n24057 = n16526 & ~n24056 ;
  assign n24058 = n23628 & ~n24057 ;
  assign n24059 = ~n11150 & n24058 ;
  assign n24060 = n13425 ^ n3383 ^ n2055 ;
  assign n24061 = n14949 & ~n24060 ;
  assign n24062 = n17199 & n24061 ;
  assign n24063 = n9786 ^ n1034 ^ 1'b0 ;
  assign n24064 = n13380 & ~n18126 ;
  assign n24065 = n6077 & n24064 ;
  assign n24066 = n5601 ^ n2324 ^ 1'b0 ;
  assign n24067 = ~n3811 & n24066 ;
  assign n24068 = n3704 & n24067 ;
  assign n24069 = n3914 & ~n24068 ;
  assign n24070 = n11501 & n20319 ;
  assign n24071 = n14698 ^ n8433 ^ n1567 ;
  assign n24072 = n24071 ^ n14772 ^ n14314 ;
  assign n24073 = n20137 ^ n16474 ^ n4415 ;
  assign n24074 = n3564 ^ n1723 ^ 1'b0 ;
  assign n24075 = n10836 | n24074 ;
  assign n24076 = ( n6781 & ~n20693 ) | ( n6781 & n24075 ) | ( ~n20693 & n24075 ) ;
  assign n24077 = n24076 ^ n16693 ^ 1'b0 ;
  assign n24078 = n8060 & ~n24077 ;
  assign n24079 = n6720 ^ n597 ^ 1'b0 ;
  assign n24080 = n9020 & n21559 ;
  assign n24081 = n24079 & n24080 ;
  assign n24082 = n24081 ^ n5986 ^ 1'b0 ;
  assign n24083 = ~n10959 & n24082 ;
  assign n24084 = n1558 & n2846 ;
  assign n24085 = n24084 ^ n7121 ^ 1'b0 ;
  assign n24086 = n10633 ^ n384 ^ 1'b0 ;
  assign n24087 = n12553 & ~n24086 ;
  assign n24088 = n4501 & n9328 ;
  assign n24089 = n24088 ^ n17128 ^ 1'b0 ;
  assign n24090 = n24089 ^ n2364 ^ n1881 ;
  assign n24091 = n6684 ^ n923 ^ 1'b0 ;
  assign n24092 = n7339 & n24091 ;
  assign n24093 = n15048 & ~n24092 ;
  assign n24097 = n2551 | n2559 ;
  assign n24098 = n1135 & ~n24097 ;
  assign n24099 = n7508 ^ n4166 ^ 1'b0 ;
  assign n24100 = n2815 & ~n24099 ;
  assign n24101 = n24098 | n24100 ;
  assign n24102 = n24101 ^ n12104 ^ n5226 ;
  assign n24094 = n2357 | n7248 ;
  assign n24095 = n8967 & ~n24094 ;
  assign n24096 = n5728 | n24095 ;
  assign n24103 = n24102 ^ n24096 ^ 1'b0 ;
  assign n24104 = n11096 & n23385 ;
  assign n24105 = ~n16154 & n24104 ;
  assign n24110 = n19539 ^ n18250 ^ n2276 ;
  assign n24106 = n6249 | n7289 ;
  assign n24107 = n24106 ^ n11137 ^ 1'b0 ;
  assign n24108 = n15836 ^ n1694 ^ n1046 ;
  assign n24109 = n24107 & ~n24108 ;
  assign n24111 = n24110 ^ n24109 ^ 1'b0 ;
  assign n24112 = ~n1102 & n6206 ;
  assign n24113 = n24112 ^ n8491 ^ 1'b0 ;
  assign n24114 = n5130 & ~n13566 ;
  assign n24115 = n24114 ^ n20716 ^ 1'b0 ;
  assign n24116 = n24115 ^ n7469 ^ 1'b0 ;
  assign n24117 = n2355 | n9092 ;
  assign n24118 = n24117 ^ n10342 ^ 1'b0 ;
  assign n24119 = n13367 & ~n16302 ;
  assign n24120 = n24119 ^ n8793 ^ n3159 ;
  assign n24121 = ( ~n1398 & n1552 ) | ( ~n1398 & n1733 ) | ( n1552 & n1733 ) ;
  assign n24122 = n5885 & ~n24121 ;
  assign n24123 = n9106 | n12120 ;
  assign n24124 = n24123 ^ n1349 ^ 1'b0 ;
  assign n24125 = ~n927 & n10342 ;
  assign n24126 = n24125 ^ n23817 ^ 1'b0 ;
  assign n24127 = n1121 & ~n1383 ;
  assign n24128 = ~n432 & n24127 ;
  assign n24129 = n20454 ^ n6383 ^ 1'b0 ;
  assign n24130 = n24128 | n24129 ;
  assign n24131 = n3824 & ~n16840 ;
  assign n24132 = ( ~n1588 & n10142 ) | ( ~n1588 & n14853 ) | ( n10142 & n14853 ) ;
  assign n24133 = n14469 ^ n8947 ^ 1'b0 ;
  assign n24134 = n10211 & n24133 ;
  assign n24135 = n1542 & n3308 ;
  assign n24137 = n20112 ^ n5772 ^ 1'b0 ;
  assign n24138 = ~n15611 & n24137 ;
  assign n24136 = n3883 | n7116 ;
  assign n24139 = n24138 ^ n24136 ^ 1'b0 ;
  assign n24140 = n3688 & ~n15221 ;
  assign n24141 = n24140 ^ n14307 ^ 1'b0 ;
  assign n24142 = n24141 ^ n8013 ^ 1'b0 ;
  assign n24143 = n7392 ^ n4178 ^ n259 ;
  assign n24144 = n24143 ^ n20712 ^ n10859 ;
  assign n24145 = n6140 & n22131 ;
  assign n24146 = n10502 & n24145 ;
  assign n24147 = n9310 & n21558 ;
  assign n24148 = ( n22293 & n24146 ) | ( n22293 & n24147 ) | ( n24146 & n24147 ) ;
  assign n24149 = ( n3552 & n10177 ) | ( n3552 & n17792 ) | ( n10177 & n17792 ) ;
  assign n24150 = n14915 & n19468 ;
  assign n24151 = ~n10432 & n24150 ;
  assign n24152 = n24149 & n24151 ;
  assign n24153 = n11834 ^ n3505 ^ 1'b0 ;
  assign n24154 = ~n24152 & n24153 ;
  assign n24155 = n2130 & ~n8959 ;
  assign n24156 = ~n21906 & n24155 ;
  assign n24157 = n10676 ^ n4100 ^ 1'b0 ;
  assign n24158 = n2815 ^ n1692 ^ 1'b0 ;
  assign n24159 = n16214 | n20913 ;
  assign n24160 = n24159 ^ n16328 ^ 1'b0 ;
  assign n24161 = n7852 ^ n1902 ^ x4 ;
  assign n24162 = n2025 | n4362 ;
  assign n24163 = n24161 | n24162 ;
  assign n24164 = n8609 & n10808 ;
  assign n24165 = ~n24163 & n24164 ;
  assign n24166 = n3845 & n14043 ;
  assign n24167 = n9225 ^ n5652 ^ n1756 ;
  assign n24168 = x25 & ~n24167 ;
  assign n24169 = n20336 & ~n24168 ;
  assign n24170 = ( n11482 & n11920 ) | ( n11482 & n15168 ) | ( n11920 & n15168 ) ;
  assign n24171 = n24170 ^ n9133 ^ n8564 ;
  assign n24172 = ( ~n1510 & n1623 ) | ( ~n1510 & n22915 ) | ( n1623 & n22915 ) ;
  assign n24173 = n14858 ^ n14380 ^ n7125 ;
  assign n24174 = ~n181 & n21080 ;
  assign n24175 = n13889 ^ n11292 ^ n4052 ;
  assign n24176 = n11158 | n24175 ;
  assign n24177 = ~n1825 & n24176 ;
  assign n24178 = n19368 & n19387 ;
  assign n24179 = ~n2340 & n16686 ;
  assign n24180 = ( n3461 & n9539 ) | ( n3461 & ~n10962 ) | ( n9539 & ~n10962 ) ;
  assign n24181 = n15856 ^ n10244 ^ 1'b0 ;
  assign n24182 = n12867 & n24181 ;
  assign n24183 = ~n15919 & n24182 ;
  assign n24184 = ~n24180 & n24183 ;
  assign n24185 = n9004 ^ n2547 ^ 1'b0 ;
  assign n24186 = n16851 | n24185 ;
  assign n24187 = ( n18127 & n23293 ) | ( n18127 & n24186 ) | ( n23293 & n24186 ) ;
  assign n24188 = n15179 ^ n10117 ^ 1'b0 ;
  assign n24190 = n11934 ^ n9481 ^ 1'b0 ;
  assign n24189 = n16150 ^ n4320 ^ 1'b0 ;
  assign n24191 = n24190 ^ n24189 ^ n19306 ;
  assign n24192 = n6295 ^ n800 ^ 1'b0 ;
  assign n24193 = n20654 ^ n15905 ^ 1'b0 ;
  assign n24194 = n13339 | n24193 ;
  assign n24195 = x13 & ~n10693 ;
  assign n24196 = ~n2815 & n24195 ;
  assign n24197 = n5872 ^ n1466 ^ 1'b0 ;
  assign n24198 = n8978 & ~n24197 ;
  assign n24199 = n19348 ^ n10553 ^ 1'b0 ;
  assign n24200 = n4028 & ~n5423 ;
  assign n24201 = ~n550 & n24200 ;
  assign n24202 = n24199 & ~n24201 ;
  assign n24203 = ~n24198 & n24202 ;
  assign n24204 = n17404 ^ n13006 ^ n3349 ;
  assign n24205 = ( n7522 & n12704 ) | ( n7522 & ~n24204 ) | ( n12704 & ~n24204 ) ;
  assign n24206 = ( n2497 & ~n3214 ) | ( n2497 & n4206 ) | ( ~n3214 & n4206 ) ;
  assign n24207 = ( ~n4302 & n6741 ) | ( ~n4302 & n24206 ) | ( n6741 & n24206 ) ;
  assign n24208 = ( ~n19944 & n22512 ) | ( ~n19944 & n24207 ) | ( n22512 & n24207 ) ;
  assign n24209 = n5446 & ~n24128 ;
  assign n24210 = n24209 ^ n6239 ^ 1'b0 ;
  assign n24211 = n24210 ^ n16139 ^ 1'b0 ;
  assign n24212 = n3368 | n18033 ;
  assign n24213 = n24212 ^ n12618 ^ 1'b0 ;
  assign n24214 = n484 | n7332 ;
  assign n24215 = n13108 & ~n18593 ;
  assign n24216 = n24215 ^ n732 ^ 1'b0 ;
  assign n24217 = n5483 & ~n10905 ;
  assign n24218 = ( n5436 & n12168 ) | ( n5436 & ~n22039 ) | ( n12168 & ~n22039 ) ;
  assign n24219 = n1488 & ~n1855 ;
  assign n24220 = n24219 ^ n10107 ^ n4317 ;
  assign n24221 = n3483 ^ n2029 ^ 1'b0 ;
  assign n24222 = n24220 | n24221 ;
  assign n24223 = n4576 | n16247 ;
  assign n24224 = n24223 ^ n13711 ^ 1'b0 ;
  assign n24225 = n6824 & ~n24224 ;
  assign n24226 = n5314 & n24225 ;
  assign n24227 = ~n23244 & n24226 ;
  assign n24228 = n8408 & n9767 ;
  assign n24232 = ( n6444 & n7554 ) | ( n6444 & n14976 ) | ( n7554 & n14976 ) ;
  assign n24229 = n10122 & ~n18170 ;
  assign n24230 = n24229 ^ n418 ^ 1'b0 ;
  assign n24231 = n2898 & ~n24230 ;
  assign n24233 = n24232 ^ n24231 ^ 1'b0 ;
  assign n24234 = n4929 ^ n3850 ^ n1133 ;
  assign n24235 = n24234 ^ n15955 ^ x57 ;
  assign n24237 = ~n7695 & n7923 ;
  assign n24236 = n3111 & n15143 ;
  assign n24238 = n24237 ^ n24236 ^ n11343 ;
  assign n24239 = n2464 & ~n10076 ;
  assign n24240 = ( n14234 & ~n16189 ) | ( n14234 & n24239 ) | ( ~n16189 & n24239 ) ;
  assign n24241 = n2617 & ~n11331 ;
  assign n24242 = ~n11836 & n19577 ;
  assign n24243 = ~n2077 & n24242 ;
  assign n24244 = n337 & n9080 ;
  assign n24245 = n8193 ^ n6544 ^ n1167 ;
  assign n24246 = ( n4120 & ~n24244 ) | ( n4120 & n24245 ) | ( ~n24244 & n24245 ) ;
  assign n24247 = n3613 ^ n2931 ^ n1156 ;
  assign n24248 = n4491 | n9303 ;
  assign n24249 = n9349 & ~n24248 ;
  assign n24250 = n1324 | n24249 ;
  assign n24251 = n3123 & n21660 ;
  assign n24252 = ( n3866 & n3880 ) | ( n3866 & ~n6168 ) | ( n3880 & ~n6168 ) ;
  assign n24253 = n3442 ^ n1600 ^ 1'b0 ;
  assign n24254 = n24252 | n24253 ;
  assign n24255 = n1675 | n24254 ;
  assign n24256 = ~n7343 & n24255 ;
  assign n24257 = ~n10360 & n24256 ;
  assign n24258 = n8130 ^ n3682 ^ 1'b0 ;
  assign n24259 = n2483 & n24258 ;
  assign n24260 = ~n4938 & n10644 ;
  assign n24261 = n24260 ^ n4344 ^ n968 ;
  assign n24262 = n20919 ^ n19688 ^ 1'b0 ;
  assign n24263 = n6512 & ~n6901 ;
  assign n24264 = n2737 & n24263 ;
  assign n24265 = ~n10008 & n24264 ;
  assign n24266 = ( n433 & n1108 ) | ( n433 & n3163 ) | ( n1108 & n3163 ) ;
  assign n24267 = n24266 ^ n8623 ^ 1'b0 ;
  assign n24268 = n5726 & n7794 ;
  assign n24269 = n24268 ^ n22852 ^ 1'b0 ;
  assign n24270 = ( ~n5846 & n19366 ) | ( ~n5846 & n24269 ) | ( n19366 & n24269 ) ;
  assign n24271 = n1046 & ~n3275 ;
  assign n24272 = ( ~n817 & n8955 ) | ( ~n817 & n24271 ) | ( n8955 & n24271 ) ;
  assign n24273 = n6555 & ~n8033 ;
  assign n24274 = n24273 ^ n9812 ^ n3724 ;
  assign n24275 = x45 & n21179 ;
  assign n24276 = n21773 | n23819 ;
  assign n24277 = ~n6313 & n7217 ;
  assign n24278 = n24277 ^ n4940 ^ 1'b0 ;
  assign n24279 = ( n4236 & n16317 ) | ( n4236 & n24278 ) | ( n16317 & n24278 ) ;
  assign n24280 = n12263 ^ n11275 ^ 1'b0 ;
  assign n24281 = ~n15323 & n24280 ;
  assign n24282 = ~n6429 & n12918 ;
  assign n24283 = n24282 ^ n15570 ^ 1'b0 ;
  assign n24284 = ( ~n5475 & n15705 ) | ( ~n5475 & n24283 ) | ( n15705 & n24283 ) ;
  assign n24285 = ( ~n4369 & n12001 ) | ( ~n4369 & n20540 ) | ( n12001 & n20540 ) ;
  assign n24286 = n4312 | n12470 ;
  assign n24287 = n24286 ^ n5250 ^ 1'b0 ;
  assign n24288 = n24287 ^ n6429 ^ n5361 ;
  assign n24289 = n13286 & ~n24288 ;
  assign n24290 = n24289 ^ n4900 ^ n1682 ;
  assign n24291 = n6764 ^ n3703 ^ 1'b0 ;
  assign n24292 = n23973 | n24291 ;
  assign n24293 = n24292 ^ n742 ^ 1'b0 ;
  assign n24294 = n5221 ^ x96 ^ 1'b0 ;
  assign n24295 = n4345 & n9157 ;
  assign n24296 = n24294 & ~n24295 ;
  assign n24297 = n24296 ^ n580 ^ 1'b0 ;
  assign n24298 = n8383 & n24297 ;
  assign n24299 = n5910 & ~n11721 ;
  assign n24300 = ~n7079 & n24299 ;
  assign n24301 = ~n5178 & n24300 ;
  assign n24302 = n18702 & n24301 ;
  assign n24303 = n22867 ^ n10223 ^ 1'b0 ;
  assign n24304 = n15036 ^ n12844 ^ n3025 ;
  assign n24305 = n10617 | n14269 ;
  assign n24306 = n24305 ^ n13786 ^ n13660 ;
  assign n24307 = n24306 ^ n14963 ^ 1'b0 ;
  assign n24308 = ~n5523 & n24307 ;
  assign n24309 = ( n5181 & ~n11873 ) | ( n5181 & n22246 ) | ( ~n11873 & n22246 ) ;
  assign n24310 = n24309 ^ n10030 ^ 1'b0 ;
  assign n24311 = ~n10732 & n12234 ;
  assign n24312 = n24311 ^ n13339 ^ 1'b0 ;
  assign n24313 = n24310 & ~n24312 ;
  assign n24314 = n7140 & ~n22548 ;
  assign n24315 = n5548 & n24314 ;
  assign n24316 = n24315 ^ n14322 ^ 1'b0 ;
  assign n24317 = n13843 ^ n5512 ^ 1'b0 ;
  assign n24318 = ~n13932 & n24317 ;
  assign n24319 = n20073 ^ n4342 ^ 1'b0 ;
  assign n24320 = ~n11695 & n24319 ;
  assign n24321 = n2912 & n4915 ;
  assign n24322 = n13016 & n23742 ;
  assign n24323 = n24321 & n24322 ;
  assign n24324 = n15676 & n24323 ;
  assign n24325 = n2131 | n23819 ;
  assign n24326 = n2081 | n12492 ;
  assign n24327 = n21807 | n24326 ;
  assign n24328 = ( n3946 & n8184 ) | ( n3946 & n13769 ) | ( n8184 & n13769 ) ;
  assign n24329 = ~n6019 & n9441 ;
  assign n24330 = ~n7918 & n24329 ;
  assign n24331 = n24328 & ~n24330 ;
  assign n24332 = ( n5956 & ~n11095 ) | ( n5956 & n16284 ) | ( ~n11095 & n16284 ) ;
  assign n24333 = n21634 ^ n18427 ^ n1865 ;
  assign n24334 = n4706 ^ n4314 ^ 1'b0 ;
  assign n24335 = n11858 | n24334 ;
  assign n24336 = n4914 | n24335 ;
  assign n24337 = n24336 ^ n13137 ^ 1'b0 ;
  assign n24338 = n2462 & n9540 ;
  assign n24339 = n24338 ^ n9101 ^ 1'b0 ;
  assign n24340 = n8536 | n10396 ;
  assign n24341 = n24340 ^ n4592 ^ 1'b0 ;
  assign n24342 = n5207 & ~n14317 ;
  assign n24343 = n20352 ^ n4548 ^ 1'b0 ;
  assign n24344 = ( n1057 & n11376 ) | ( n1057 & ~n24343 ) | ( n11376 & ~n24343 ) ;
  assign n24345 = n12343 ^ n7925 ^ n6332 ;
  assign n24346 = ( n11183 & n12796 ) | ( n11183 & ~n23403 ) | ( n12796 & ~n23403 ) ;
  assign n24347 = n16243 ^ n6435 ^ 1'b0 ;
  assign n24348 = n14859 & n24347 ;
  assign n24349 = n14738 ^ n13382 ^ 1'b0 ;
  assign n24350 = n24348 & n24349 ;
  assign n24351 = n7052 & n13985 ;
  assign n24352 = n24351 ^ n10943 ^ 1'b0 ;
  assign n24353 = n9924 | n24352 ;
  assign n24354 = n24353 ^ n4318 ^ 1'b0 ;
  assign n24355 = n24350 | n24354 ;
  assign n24356 = n2007 & ~n6256 ;
  assign n24357 = ~n19909 & n24356 ;
  assign n24358 = n7955 & ~n10975 ;
  assign n24359 = n24358 ^ n3760 ^ 1'b0 ;
  assign n24360 = n22987 ^ n9678 ^ 1'b0 ;
  assign n24361 = ~n16272 & n24360 ;
  assign n24362 = n9955 ^ n8426 ^ n7621 ;
  assign n24363 = n24362 ^ n6968 ^ 1'b0 ;
  assign n24364 = n4170 & ~n17552 ;
  assign n24365 = n24364 ^ n17053 ^ 1'b0 ;
  assign n24366 = ( n212 & n24363 ) | ( n212 & n24365 ) | ( n24363 & n24365 ) ;
  assign n24367 = n9275 ^ n6309 ^ 1'b0 ;
  assign n24368 = n22420 ^ n131 ^ 1'b0 ;
  assign n24369 = n24367 | n24368 ;
  assign n24370 = n24369 ^ n6045 ^ n514 ;
  assign n24371 = n10910 | n13731 ;
  assign n24372 = n8592 ^ n2900 ^ 1'b0 ;
  assign n24373 = n15975 | n24372 ;
  assign n24375 = n4370 & n9185 ;
  assign n24376 = ~n5984 & n24375 ;
  assign n24374 = n2630 & ~n12884 ;
  assign n24377 = n24376 ^ n24374 ^ 1'b0 ;
  assign n24378 = n10602 ^ n10515 ^ 1'b0 ;
  assign n24379 = ( n408 & n8089 ) | ( n408 & n19946 ) | ( n8089 & n19946 ) ;
  assign n24380 = ~n5011 & n23749 ;
  assign n24381 = ~n11101 & n24380 ;
  assign n24382 = n10540 ^ n10485 ^ n4741 ;
  assign n24383 = n24381 & ~n24382 ;
  assign n24385 = n23326 ^ n10602 ^ 1'b0 ;
  assign n24386 = n4567 & ~n24385 ;
  assign n24384 = x23 & ~n18422 ;
  assign n24387 = n24386 ^ n24384 ^ 1'b0 ;
  assign n24388 = n11589 ^ n6435 ^ 1'b0 ;
  assign n24389 = n10241 & n20379 ;
  assign n24390 = n24388 & n24389 ;
  assign n24391 = n3218 ^ n2896 ^ 1'b0 ;
  assign n24392 = ~n1253 & n24391 ;
  assign n24393 = n746 & n24392 ;
  assign n24394 = n8151 ^ n535 ^ 1'b0 ;
  assign n24395 = n6686 | n24217 ;
  assign n24396 = n24394 & ~n24395 ;
  assign n24397 = n9321 ^ n8035 ^ n4778 ;
  assign n24398 = n9622 ^ n4645 ^ 1'b0 ;
  assign n24399 = ~n24397 & n24398 ;
  assign n24400 = ( ~n3088 & n4172 ) | ( ~n3088 & n7697 ) | ( n4172 & n7697 ) ;
  assign n24401 = ( n8601 & ~n8814 ) | ( n8601 & n24400 ) | ( ~n8814 & n24400 ) ;
  assign n24402 = ( n16251 & ~n20038 ) | ( n16251 & n23006 ) | ( ~n20038 & n23006 ) ;
  assign n24403 = n24402 ^ n289 ^ 1'b0 ;
  assign n24404 = ( n18090 & n21472 ) | ( n18090 & n24403 ) | ( n21472 & n24403 ) ;
  assign n24405 = n12046 ^ n11176 ^ n4665 ;
  assign n24406 = n3939 ^ n2110 ^ 1'b0 ;
  assign n24407 = n4172 | n24406 ;
  assign n24408 = n24407 ^ n7674 ^ 1'b0 ;
  assign n24409 = n11187 | n24408 ;
  assign n24410 = n1257 | n24409 ;
  assign n24411 = n13380 ^ n6816 ^ n5262 ;
  assign n24412 = n17342 | n24411 ;
  assign n24413 = n8541 & n9607 ;
  assign n24414 = n24412 & n24413 ;
  assign n24415 = n10984 ^ n2723 ^ 1'b0 ;
  assign n24416 = n4338 & ~n24415 ;
  assign n24417 = n10576 & n24416 ;
  assign n24418 = n1709 & n12785 ;
  assign n24419 = n24417 & n24418 ;
  assign n24420 = ( ~n360 & n1710 ) | ( ~n360 & n3062 ) | ( n1710 & n3062 ) ;
  assign n24421 = n7708 | n24420 ;
  assign n24422 = n13025 & ~n24421 ;
  assign n24423 = n5544 & n17656 ;
  assign n24424 = n9850 ^ n9628 ^ n6429 ;
  assign n24425 = ~n8532 & n21253 ;
  assign n24426 = n6182 | n24425 ;
  assign n24427 = n11418 ^ n10132 ^ 1'b0 ;
  assign n24428 = n17607 ^ n16177 ^ 1'b0 ;
  assign n24429 = ~n24427 & n24428 ;
  assign n24430 = n5839 & ~n14506 ;
  assign n24431 = n7929 ^ n6834 ^ 1'b0 ;
  assign n24432 = n4724 & n24431 ;
  assign n24433 = x61 | n24432 ;
  assign n24434 = n1487 & n16603 ;
  assign n24435 = n12813 ^ n12279 ^ 1'b0 ;
  assign n24436 = n7574 & n24435 ;
  assign n24437 = n2847 | n13536 ;
  assign n24438 = n3564 & ~n24437 ;
  assign n24439 = n3584 & ~n3792 ;
  assign n24440 = n24439 ^ n22023 ^ 1'b0 ;
  assign n24441 = n4714 & n24440 ;
  assign n24442 = n7916 | n10157 ;
  assign n24443 = n18961 ^ n12703 ^ n10418 ;
  assign n24444 = n24442 & ~n24443 ;
  assign n24445 = n13856 ^ n9921 ^ 1'b0 ;
  assign n24446 = n17147 ^ n14314 ^ 1'b0 ;
  assign n24447 = n14582 ^ n12239 ^ 1'b0 ;
  assign n24448 = n2417 & ~n24447 ;
  assign n24450 = n225 | n16142 ;
  assign n24449 = n15989 | n17811 ;
  assign n24451 = n24450 ^ n24449 ^ 1'b0 ;
  assign n24452 = ~n16233 & n24451 ;
  assign n24453 = n6421 & n24452 ;
  assign n24454 = n10223 ^ n9324 ^ 1'b0 ;
  assign n24455 = n8063 | n24454 ;
  assign n24456 = ( ~n730 & n2308 ) | ( ~n730 & n7312 ) | ( n2308 & n7312 ) ;
  assign n24457 = n24455 | n24456 ;
  assign n24458 = n247 & ~n1199 ;
  assign n24459 = n10204 & n15667 ;
  assign n24460 = ~n24458 & n24459 ;
  assign n24463 = n6173 ^ n5965 ^ 1'b0 ;
  assign n24464 = n566 & ~n24463 ;
  assign n24465 = n13231 & n24464 ;
  assign n24466 = n24465 ^ n1734 ^ 1'b0 ;
  assign n24461 = n242 & n9528 ;
  assign n24462 = ( n14239 & n16603 ) | ( n14239 & n24461 ) | ( n16603 & n24461 ) ;
  assign n24467 = n24466 ^ n24462 ^ n21769 ;
  assign n24468 = n5417 ^ n5040 ^ 1'b0 ;
  assign n24469 = n13718 & n24468 ;
  assign n24470 = ( n2416 & n6946 ) | ( n2416 & n16971 ) | ( n6946 & n16971 ) ;
  assign n24471 = ~n2574 & n20639 ;
  assign n24472 = n17670 & n24471 ;
  assign n24473 = ~n18053 & n20853 ;
  assign n24474 = n24473 ^ n7717 ^ 1'b0 ;
  assign n24475 = n420 & ~n15937 ;
  assign n24476 = n24475 ^ n9223 ^ 1'b0 ;
  assign n24482 = n7649 ^ n7554 ^ 1'b0 ;
  assign n24477 = n4979 ^ n1089 ^ 1'b0 ;
  assign n24478 = n163 & ~n24477 ;
  assign n24479 = n10777 ^ n8117 ^ x123 ;
  assign n24480 = n6433 & ~n24479 ;
  assign n24481 = n24478 & n24480 ;
  assign n24483 = n24482 ^ n24481 ^ 1'b0 ;
  assign n24484 = n721 & ~n24483 ;
  assign n24485 = ~n3390 & n12922 ;
  assign n24486 = n7468 & n24485 ;
  assign n24487 = n24484 & n24486 ;
  assign n24488 = n10118 & n15748 ;
  assign n24489 = n24488 ^ n13914 ^ 1'b0 ;
  assign n24490 = n4256 | n5112 ;
  assign n24491 = n24489 & ~n24490 ;
  assign n24492 = n8036 | n24491 ;
  assign n24494 = n11485 ^ n4498 ^ n3935 ;
  assign n24493 = n6223 & ~n18338 ;
  assign n24495 = n24494 ^ n24493 ^ n478 ;
  assign n24496 = n17407 ^ n14703 ^ 1'b0 ;
  assign n24497 = n3751 | n24496 ;
  assign n24498 = ( n4993 & n15061 ) | ( n4993 & n24497 ) | ( n15061 & n24497 ) ;
  assign n24499 = ~n11365 & n16980 ;
  assign n24500 = n24498 & n24499 ;
  assign n24501 = n475 | n15002 ;
  assign n24502 = n17120 | n24501 ;
  assign n24503 = ( n2128 & ~n2645 ) | ( n2128 & n5651 ) | ( ~n2645 & n5651 ) ;
  assign n24504 = n4719 & ~n24503 ;
  assign n24505 = n10005 & ~n24504 ;
  assign n24506 = n8294 & n24505 ;
  assign n24507 = n6196 | n11707 ;
  assign n24508 = n20772 ^ n18846 ^ n915 ;
  assign n24509 = n732 & n24508 ;
  assign n24510 = ~n24507 & n24509 ;
  assign n24511 = n2478 | n13143 ;
  assign n24512 = n10661 & ~n24511 ;
  assign n24513 = n265 & ~n890 ;
  assign n24514 = n15237 & n24513 ;
  assign n24515 = n5331 & ~n24455 ;
  assign n24516 = n12018 ^ n5425 ^ n2554 ;
  assign n24517 = ( n214 & n4210 ) | ( n214 & ~n10341 ) | ( n4210 & ~n10341 ) ;
  assign n24518 = n21256 ^ n16790 ^ n6876 ;
  assign n24519 = n13966 ^ n2306 ^ n992 ;
  assign n24520 = n24519 ^ n6125 ^ 1'b0 ;
  assign n24521 = n24520 ^ n23006 ^ n22181 ;
  assign n24522 = n19115 ^ n3030 ^ 1'b0 ;
  assign n24523 = ~n631 & n3466 ;
  assign n24524 = n24523 ^ n5826 ^ 1'b0 ;
  assign n24525 = n24524 ^ n11320 ^ 1'b0 ;
  assign n24526 = n4119 & ~n24525 ;
  assign n24527 = ~n10136 & n24526 ;
  assign n24528 = n4853 ^ n2678 ^ 1'b0 ;
  assign n24529 = n5425 & ~n24528 ;
  assign n24530 = n24529 ^ n11584 ^ n8346 ;
  assign n24531 = n24530 ^ n16849 ^ n2815 ;
  assign n24532 = n9744 ^ n6747 ^ n925 ;
  assign n24533 = n24532 ^ n13763 ^ n6858 ;
  assign n24534 = n23243 ^ n18961 ^ n15469 ;
  assign n24535 = n12513 & n24534 ;
  assign n24537 = n15495 ^ n2016 ^ 1'b0 ;
  assign n24538 = ~n14878 & n24537 ;
  assign n24539 = n3845 & n24538 ;
  assign n24536 = n5965 | n21012 ;
  assign n24540 = n24539 ^ n24536 ^ 1'b0 ;
  assign n24541 = n19882 ^ n15231 ^ 1'b0 ;
  assign n24542 = n11581 ^ n161 ^ 1'b0 ;
  assign n24543 = n14855 & ~n24542 ;
  assign n24544 = ( ~n1436 & n4455 ) | ( ~n1436 & n11261 ) | ( n4455 & n11261 ) ;
  assign n24545 = n24544 ^ n804 ^ n227 ;
  assign n24546 = n960 | n24545 ;
  assign n24548 = n5687 ^ n3883 ^ 1'b0 ;
  assign n24549 = n1869 & n24548 ;
  assign n24550 = n24549 ^ n18048 ^ 1'b0 ;
  assign n24551 = n858 | n24550 ;
  assign n24547 = n1925 | n14319 ;
  assign n24552 = n24551 ^ n24547 ^ 1'b0 ;
  assign n24553 = ( ~n15088 & n15387 ) | ( ~n15088 & n24552 ) | ( n15387 & n24552 ) ;
  assign n24555 = n13869 ^ n193 ^ x103 ;
  assign n24554 = n16913 ^ n5928 ^ n4340 ;
  assign n24556 = n24555 ^ n24554 ^ n7113 ;
  assign n24557 = n22283 ^ n10541 ^ 1'b0 ;
  assign n24558 = n1871 & n10153 ;
  assign n24559 = n1113 & n5347 ;
  assign n24561 = n19287 ^ n2285 ^ 1'b0 ;
  assign n24562 = n12418 & n24561 ;
  assign n24563 = n24562 ^ n21843 ^ 1'b0 ;
  assign n24560 = n7211 & ~n21343 ;
  assign n24564 = n24563 ^ n24560 ^ 1'b0 ;
  assign n24566 = n8253 ^ n1260 ^ 1'b0 ;
  assign n24567 = n3950 & ~n24566 ;
  assign n24565 = n16346 | n21984 ;
  assign n24568 = n24567 ^ n24565 ^ 1'b0 ;
  assign n24569 = n5557 ^ n2416 ^ 1'b0 ;
  assign n24570 = ( n6669 & n13628 ) | ( n6669 & ~n18893 ) | ( n13628 & ~n18893 ) ;
  assign n24571 = n21206 ^ n15564 ^ 1'b0 ;
  assign n24572 = n9318 ^ n4020 ^ 1'b0 ;
  assign n24573 = n10298 ^ n929 ^ 1'b0 ;
  assign n24574 = n3038 & n24573 ;
  assign n24575 = n24572 & n24574 ;
  assign n24576 = n12240 ^ n5675 ^ 1'b0 ;
  assign n24577 = ( ~n4956 & n16261 ) | ( ~n4956 & n24576 ) | ( n16261 & n24576 ) ;
  assign n24578 = n14343 ^ n5813 ^ 1'b0 ;
  assign n24579 = n4601 & ~n24578 ;
  assign n24580 = ~n22819 & n24341 ;
  assign n24581 = n24580 ^ n3777 ^ 1'b0 ;
  assign n24582 = ~n12198 & n20441 ;
  assign n24583 = n24582 ^ n10028 ^ 1'b0 ;
  assign n24584 = n16935 ^ n8027 ^ n726 ;
  assign n24585 = n1297 | n24584 ;
  assign n24586 = n24585 ^ n1673 ^ 1'b0 ;
  assign n24588 = ~n11329 & n11460 ;
  assign n24589 = ~n7298 & n24588 ;
  assign n24587 = n11475 & ~n12120 ;
  assign n24590 = n24589 ^ n24587 ^ 1'b0 ;
  assign n24591 = n24590 ^ n18350 ^ n15420 ;
  assign n24592 = n6294 & n18040 ;
  assign n24593 = n24592 ^ n5502 ^ 1'b0 ;
  assign n24594 = n8817 ^ n1850 ^ n965 ;
  assign n24595 = n10036 | n24594 ;
  assign n24596 = ~n14014 & n24595 ;
  assign n24597 = ~n24593 & n24596 ;
  assign n24598 = ( n3636 & ~n5828 ) | ( n3636 & n10869 ) | ( ~n5828 & n10869 ) ;
  assign n24599 = n2611 & ~n20080 ;
  assign n24600 = ( n1205 & n24598 ) | ( n1205 & n24599 ) | ( n24598 & n24599 ) ;
  assign n24601 = n3788 & ~n22048 ;
  assign n24602 = n21675 & n24601 ;
  assign n24603 = n9810 & n24182 ;
  assign n24604 = ~n7189 & n24603 ;
  assign n24605 = n4697 & ~n18454 ;
  assign n24606 = n2844 | n15452 ;
  assign n24607 = n24606 ^ n1158 ^ 1'b0 ;
  assign n24608 = n14143 | n23819 ;
  assign n24609 = n24608 ^ n21716 ^ 1'b0 ;
  assign n24613 = ~n474 & n5214 ;
  assign n24614 = ~n2868 & n24613 ;
  assign n24610 = n3912 ^ n2702 ^ 1'b0 ;
  assign n24611 = n293 | n24610 ;
  assign n24612 = n24611 ^ n15421 ^ 1'b0 ;
  assign n24615 = n24614 ^ n24612 ^ n1648 ;
  assign n24618 = n20336 ^ n8914 ^ n206 ;
  assign n24616 = ( n4256 & n5085 ) | ( n4256 & n10212 ) | ( n5085 & n10212 ) ;
  assign n24617 = ~n23269 & n24616 ;
  assign n24619 = n24618 ^ n24617 ^ 1'b0 ;
  assign n24620 = n14612 ^ n8101 ^ 1'b0 ;
  assign n24621 = n16907 | n24620 ;
  assign n24626 = n18094 ^ n6611 ^ n608 ;
  assign n24627 = n19834 | n24626 ;
  assign n24628 = n14245 & ~n24627 ;
  assign n24629 = n442 | n24628 ;
  assign n24622 = n14859 & ~n16011 ;
  assign n24623 = ~n19814 & n24622 ;
  assign n24624 = n1029 & n24623 ;
  assign n24625 = n2201 & ~n24624 ;
  assign n24630 = n24629 ^ n24625 ^ 1'b0 ;
  assign n24631 = ( n7217 & n9434 ) | ( n7217 & n16314 ) | ( n9434 & n16314 ) ;
  assign n24632 = n3044 & n24631 ;
  assign n24633 = n323 & ~n7844 ;
  assign n24634 = n7914 | n24633 ;
  assign n24635 = n23063 | n24634 ;
  assign n24638 = n4847 | n12768 ;
  assign n24639 = n9925 & ~n24638 ;
  assign n24636 = n13812 ^ n2207 ^ 1'b0 ;
  assign n24637 = n4376 & n24636 ;
  assign n24640 = n24639 ^ n24637 ^ n23906 ;
  assign n24641 = n11040 ^ n5527 ^ 1'b0 ;
  assign n24642 = ( n2028 & ~n13715 ) | ( n2028 & n22708 ) | ( ~n13715 & n22708 ) ;
  assign n24643 = n16202 & n24642 ;
  assign n24645 = n21337 ^ n4387 ^ 1'b0 ;
  assign n24646 = n1141 | n24645 ;
  assign n24644 = x92 & ~n1997 ;
  assign n24647 = n24646 ^ n24644 ^ 1'b0 ;
  assign n24648 = n5999 ^ n5037 ^ 1'b0 ;
  assign n24649 = n24647 & n24648 ;
  assign n24650 = ~n3019 & n6013 ;
  assign n24651 = ~n5815 & n24650 ;
  assign n24652 = n23586 & n24651 ;
  assign n24653 = ~n15456 & n18954 ;
  assign n24654 = n24653 ^ n11045 ^ 1'b0 ;
  assign n24655 = n5143 | n9572 ;
  assign n24656 = n24655 ^ n12031 ^ 1'b0 ;
  assign n24657 = n9359 ^ n1230 ^ 1'b0 ;
  assign n24658 = n175 & ~n13659 ;
  assign n24659 = ( n1010 & n4429 ) | ( n1010 & n24658 ) | ( n4429 & n24658 ) ;
  assign n24660 = n2687 & n13099 ;
  assign n24661 = n993 | n13953 ;
  assign n24662 = n5561 & n6641 ;
  assign n24663 = n24662 ^ n5281 ^ 1'b0 ;
  assign n24664 = n24663 ^ n5715 ^ 1'b0 ;
  assign n24665 = n24664 ^ n937 ^ 1'b0 ;
  assign n24666 = n22905 | n24665 ;
  assign n24667 = n20744 ^ n12507 ^ 1'b0 ;
  assign n24668 = n1046 | n3850 ;
  assign n24669 = n24668 ^ n9426 ^ n1610 ;
  assign n24670 = n24669 ^ n10794 ^ 1'b0 ;
  assign n24671 = n5537 | n24670 ;
  assign n24672 = n8241 | n24671 ;
  assign n24673 = n8532 & ~n15945 ;
  assign n24674 = n1251 ^ n800 ^ 1'b0 ;
  assign n24675 = n2307 & ~n2680 ;
  assign n24676 = n24675 ^ n17209 ^ n7270 ;
  assign n24677 = n6965 & ~n12801 ;
  assign n24678 = n3438 & n10287 ;
  assign n24679 = n965 & n12138 ;
  assign n24680 = n4416 ^ n1461 ^ 1'b0 ;
  assign n24681 = n3305 | n24680 ;
  assign n24682 = n24681 ^ n18051 ^ 1'b0 ;
  assign n24683 = n24682 ^ n1314 ^ 1'b0 ;
  assign n24684 = n20885 & n24683 ;
  assign n24685 = n24537 ^ n4414 ^ 1'b0 ;
  assign n24686 = n7449 & ~n24685 ;
  assign n24687 = n16595 ^ n6055 ^ n4778 ;
  assign n24688 = ~n10664 & n24687 ;
  assign n24689 = n24688 ^ n1974 ^ 1'b0 ;
  assign n24690 = ( ~n2074 & n3582 ) | ( ~n2074 & n4385 ) | ( n3582 & n4385 ) ;
  assign n24691 = n4383 & ~n18660 ;
  assign n24692 = n24691 ^ n10235 ^ 1'b0 ;
  assign n24693 = ( n4150 & n24690 ) | ( n4150 & n24692 ) | ( n24690 & n24692 ) ;
  assign n24694 = n15471 ^ n9792 ^ 1'b0 ;
  assign n24695 = n579 | n14095 ;
  assign n24696 = n24695 ^ n8668 ^ 1'b0 ;
  assign n24698 = n940 & n17196 ;
  assign n24697 = n2122 & ~n11440 ;
  assign n24699 = n24698 ^ n24697 ^ 1'b0 ;
  assign n24700 = n12885 ^ n9571 ^ 1'b0 ;
  assign n24701 = ( n5403 & ~n6145 ) | ( n5403 & n7199 ) | ( ~n6145 & n7199 ) ;
  assign n24702 = n23967 & n24701 ;
  assign n24703 = n313 & ~n16621 ;
  assign n24704 = ~n15781 & n24703 ;
  assign n24705 = ~n16303 & n24704 ;
  assign n24706 = n22348 ^ n18115 ^ 1'b0 ;
  assign n24707 = ~n11081 & n24706 ;
  assign n24708 = ~n794 & n14891 ;
  assign n24709 = n24708 ^ n11312 ^ 1'b0 ;
  assign n24710 = n24709 ^ n2413 ^ 1'b0 ;
  assign n24711 = n16721 & n24710 ;
  assign n24712 = n2698 & n24711 ;
  assign n24713 = n15179 ^ n4753 ^ 1'b0 ;
  assign n24714 = ( ~n8335 & n19831 ) | ( ~n8335 & n24713 ) | ( n19831 & n24713 ) ;
  assign n24715 = n23208 ^ x106 ^ 1'b0 ;
  assign n24716 = n3961 & n6997 ;
  assign n24717 = ~n3726 & n24716 ;
  assign n24718 = n11461 ^ n4296 ^ n165 ;
  assign n24719 = ( n11507 & ~n24717 ) | ( n11507 & n24718 ) | ( ~n24717 & n24718 ) ;
  assign n24720 = ~n3671 & n24719 ;
  assign n24721 = n19907 ^ n18771 ^ n15474 ;
  assign n24722 = n436 & ~n12509 ;
  assign n24723 = n10620 | n12284 ;
  assign n24724 = n24723 ^ n4132 ^ 1'b0 ;
  assign n24725 = n23636 & ~n24724 ;
  assign n24726 = n5196 | n24725 ;
  assign n24727 = ( n2598 & n17294 ) | ( n2598 & ~n24726 ) | ( n17294 & ~n24726 ) ;
  assign n24728 = ~n1594 & n21434 ;
  assign n24729 = n24728 ^ n16753 ^ 1'b0 ;
  assign n24730 = n11802 ^ n10456 ^ 1'b0 ;
  assign n24731 = n24343 | n24730 ;
  assign n24732 = n11271 & ~n24455 ;
  assign n24733 = n12386 & n24732 ;
  assign n24734 = n20842 & ~n24733 ;
  assign n24735 = n2772 & ~n24734 ;
  assign n24736 = n3770 & n9548 ;
  assign n24737 = n1485 & n24736 ;
  assign n24738 = n24737 ^ n4099 ^ n3440 ;
  assign n24739 = x51 & ~n24738 ;
  assign n24740 = n24739 ^ n423 ^ n145 ;
  assign n24741 = ( ~n1020 & n7071 ) | ( ~n1020 & n9473 ) | ( n7071 & n9473 ) ;
  assign n24742 = x103 & ~n6340 ;
  assign n24743 = n10497 & n24742 ;
  assign n24744 = n24743 ^ n4521 ^ n254 ;
  assign n24745 = ( ~n2961 & n7108 ) | ( ~n2961 & n17450 ) | ( n7108 & n17450 ) ;
  assign n24746 = n10891 & ~n24745 ;
  assign n24747 = n24746 ^ n9873 ^ 1'b0 ;
  assign n24748 = n14587 & n15622 ;
  assign n24749 = n1696 & ~n18490 ;
  assign n24750 = n13437 ^ n3865 ^ 1'b0 ;
  assign n24751 = n7593 & n24750 ;
  assign n24752 = n17771 ^ n9766 ^ 1'b0 ;
  assign n24753 = n4204 & ~n24752 ;
  assign n24754 = n20681 | n24753 ;
  assign n24755 = n21258 ^ n19451 ^ 1'b0 ;
  assign n24756 = ( n12981 & ~n16398 ) | ( n12981 & n21787 ) | ( ~n16398 & n21787 ) ;
  assign n24757 = n1442 & ~n15736 ;
  assign n24758 = n12473 & n24757 ;
  assign n24759 = n1651 ^ n1569 ^ 1'b0 ;
  assign n24760 = ( n1871 & ~n4332 ) | ( n1871 & n24759 ) | ( ~n4332 & n24759 ) ;
  assign n24761 = n24760 ^ n20642 ^ 1'b0 ;
  assign n24762 = n13285 ^ n2009 ^ 1'b0 ;
  assign n24763 = n20489 & n24762 ;
  assign n24764 = n19539 ^ n6256 ^ 1'b0 ;
  assign n24765 = n6410 & ~n24764 ;
  assign n24766 = ( ~n3279 & n7598 ) | ( ~n3279 & n11616 ) | ( n7598 & n11616 ) ;
  assign n24767 = ~n10941 & n22241 ;
  assign n24768 = n24767 ^ n18139 ^ 1'b0 ;
  assign n24769 = n5473 ^ n5278 ^ 1'b0 ;
  assign n24770 = n24503 & ~n24769 ;
  assign n24771 = n298 & n24770 ;
  assign n24772 = ( n6034 & ~n12572 ) | ( n6034 & n24146 ) | ( ~n12572 & n24146 ) ;
  assign n24773 = n24772 ^ n4797 ^ 1'b0 ;
  assign n24774 = ~n1974 & n24773 ;
  assign n24775 = ~n3968 & n24774 ;
  assign n24776 = ~n9971 & n14821 ;
  assign n24777 = n24776 ^ n8232 ^ 1'b0 ;
  assign n24778 = n14821 ^ n3403 ^ 1'b0 ;
  assign n24779 = n22604 & n24778 ;
  assign n24780 = n11524 ^ n10591 ^ 1'b0 ;
  assign n24781 = n2481 & n24780 ;
  assign n24782 = n13573 ^ n3896 ^ 1'b0 ;
  assign n24783 = n24781 & ~n24782 ;
  assign n24784 = n5205 & n9441 ;
  assign n24785 = n24784 ^ n6053 ^ 1'b0 ;
  assign n24786 = n24785 ^ n23245 ^ 1'b0 ;
  assign n24787 = n24783 & n24786 ;
  assign n24788 = n10539 ^ n1774 ^ 1'b0 ;
  assign n24789 = n12240 ^ n10716 ^ n8677 ;
  assign n24790 = ( ~n10704 & n24788 ) | ( ~n10704 & n24789 ) | ( n24788 & n24789 ) ;
  assign n24791 = x91 & n2444 ;
  assign n24792 = ~n7594 & n24791 ;
  assign n24793 = ( n10980 & n11422 ) | ( n10980 & n24792 ) | ( n11422 & n24792 ) ;
  assign n24794 = ( ~n9343 & n14245 ) | ( ~n9343 & n24793 ) | ( n14245 & n24793 ) ;
  assign n24795 = ( n11723 & n19172 ) | ( n11723 & ~n24180 ) | ( n19172 & ~n24180 ) ;
  assign n24796 = n24795 ^ n17672 ^ n4231 ;
  assign n24797 = n734 & ~n2072 ;
  assign n24798 = n887 & ~n2893 ;
  assign n24799 = ~n17947 & n24798 ;
  assign n24800 = ~n432 & n14985 ;
  assign n24801 = n5361 & n24800 ;
  assign n24802 = n24801 ^ n22521 ^ 1'b0 ;
  assign n24803 = n4649 ^ n1965 ^ n211 ;
  assign n24804 = n19371 ^ n11019 ^ 1'b0 ;
  assign n24805 = n24803 & n24804 ;
  assign n24806 = n24544 ^ n6427 ^ 1'b0 ;
  assign n24807 = ( ~n18149 & n24805 ) | ( ~n18149 & n24806 ) | ( n24805 & n24806 ) ;
  assign n24808 = n12685 | n24807 ;
  assign n24809 = n8250 & ~n14448 ;
  assign n24810 = ~n3930 & n24809 ;
  assign n24811 = n21589 ^ n17614 ^ 1'b0 ;
  assign n24812 = n10024 | n24811 ;
  assign n24813 = n14667 ^ n1455 ^ n490 ;
  assign n24814 = n9557 & ~n9655 ;
  assign n24815 = n24814 ^ n23148 ^ n10309 ;
  assign n24816 = ~n4603 & n4730 ;
  assign n24817 = n7130 & n8852 ;
  assign n24818 = ( n8926 & ~n24816 ) | ( n8926 & n24817 ) | ( ~n24816 & n24817 ) ;
  assign n24819 = ( ~n1096 & n24815 ) | ( ~n1096 & n24818 ) | ( n24815 & n24818 ) ;
  assign n24820 = n4681 ^ n1803 ^ 1'b0 ;
  assign n24821 = n10987 ^ n7963 ^ 1'b0 ;
  assign n24822 = ~n1927 & n24821 ;
  assign n24823 = n491 | n24822 ;
  assign n24824 = n8392 & ~n19937 ;
  assign n24825 = ~n11155 & n24824 ;
  assign n24826 = n2171 & ~n24048 ;
  assign n24827 = n7784 & n24826 ;
  assign n24828 = n8780 | n12277 ;
  assign n24829 = n11464 | n20385 ;
  assign n24830 = n24829 ^ n11000 ^ 1'b0 ;
  assign n24831 = n24830 ^ n18758 ^ 1'b0 ;
  assign n24832 = n4290 & ~n15076 ;
  assign n24833 = n13937 ^ n6344 ^ 1'b0 ;
  assign n24834 = n1192 & n24833 ;
  assign n24835 = n10088 | n14526 ;
  assign n24836 = ~n1644 & n7665 ;
  assign n24837 = n16708 & n24836 ;
  assign n24838 = n5836 & ~n11042 ;
  assign n24839 = n24838 ^ n23665 ^ 1'b0 ;
  assign n24840 = n19880 ^ n12999 ^ 1'b0 ;
  assign n24841 = ~n1345 & n24840 ;
  assign n24842 = n2058 & n13430 ;
  assign n24843 = n24842 ^ n1043 ^ n798 ;
  assign n24844 = ( n10920 & n16621 ) | ( n10920 & ~n20280 ) | ( n16621 & ~n20280 ) ;
  assign n24845 = ( n330 & n22624 ) | ( n330 & ~n24844 ) | ( n22624 & ~n24844 ) ;
  assign n24846 = n5685 & ~n24845 ;
  assign n24847 = n24843 & ~n24846 ;
  assign n24848 = ( n14368 & n18581 ) | ( n14368 & ~n20216 ) | ( n18581 & ~n20216 ) ;
  assign n24849 = n13032 ^ n6447 ^ n1999 ;
  assign n24850 = n1022 & ~n10880 ;
  assign n24851 = n24850 ^ n23990 ^ 1'b0 ;
  assign n24852 = n24851 ^ n20683 ^ n16151 ;
  assign n24853 = n11409 & n11882 ;
  assign n24854 = n24853 ^ n1244 ^ 1'b0 ;
  assign n24855 = n8972 ^ n2637 ^ 1'b0 ;
  assign n24856 = ~n24854 & n24855 ;
  assign n24857 = n6209 ^ n4073 ^ 1'b0 ;
  assign n24858 = n10231 & ~n14440 ;
  assign n24859 = n24858 ^ n3566 ^ 1'b0 ;
  assign n24860 = n24859 ^ n3863 ^ 1'b0 ;
  assign n24861 = ~n9482 & n24860 ;
  assign n24862 = n13129 & ~n24861 ;
  assign n24863 = n22430 ^ n741 ^ 1'b0 ;
  assign n24864 = n21352 ^ n881 ^ 1'b0 ;
  assign n24865 = ~n24863 & n24864 ;
  assign n24866 = n5445 & ~n7216 ;
  assign n24867 = n24122 ^ n8209 ^ 1'b0 ;
  assign n24868 = n11845 | n24867 ;
  assign n24869 = n9776 | n19620 ;
  assign n24870 = ( ~n4873 & n12425 ) | ( ~n4873 & n17092 ) | ( n12425 & n17092 ) ;
  assign n24871 = n23093 ^ n20585 ^ 1'b0 ;
  assign n24872 = ~n3240 & n24305 ;
  assign n24873 = n22890 & ~n24872 ;
  assign n24874 = n13441 & n22286 ;
  assign n24875 = n4294 | n24874 ;
  assign n24876 = n7098 & ~n14305 ;
  assign n24877 = ~n1495 & n15653 ;
  assign n24878 = n24877 ^ n11070 ^ 1'b0 ;
  assign n24879 = n24876 & ~n24878 ;
  assign n24880 = ~n17238 & n24879 ;
  assign n24881 = ( n6110 & n8741 ) | ( n6110 & n10061 ) | ( n8741 & n10061 ) ;
  assign n24882 = ( ~n8991 & n15561 ) | ( ~n8991 & n24881 ) | ( n15561 & n24881 ) ;
  assign n24883 = n11766 ^ n6079 ^ n4605 ;
  assign n24884 = n24883 ^ n17906 ^ 1'b0 ;
  assign n24885 = n24882 & n24884 ;
  assign n24886 = n24885 ^ n6906 ^ 1'b0 ;
  assign n24887 = ~n11898 & n24886 ;
  assign n24888 = n12101 & n15396 ;
  assign n24889 = ~n17992 & n24888 ;
  assign n24890 = n24889 ^ n8090 ^ 1'b0 ;
  assign n24891 = ( n1652 & n1992 ) | ( n1652 & ~n24890 ) | ( n1992 & ~n24890 ) ;
  assign n24892 = n24891 ^ n11951 ^ n725 ;
  assign n24893 = ~n9522 & n11110 ;
  assign n24894 = n138 & n24893 ;
  assign n24895 = ( n12143 & ~n18026 ) | ( n12143 & n24894 ) | ( ~n18026 & n24894 ) ;
  assign n24896 = n24895 ^ n12068 ^ n8328 ;
  assign n24897 = n24896 ^ n19947 ^ n14665 ;
  assign n24898 = n23819 ^ n6935 ^ n2290 ;
  assign n24899 = n7308 | n15131 ;
  assign n24900 = n2233 | n6409 ;
  assign n24901 = n21416 ^ n13240 ^ 1'b0 ;
  assign n24902 = n6717 | n24901 ;
  assign n24903 = n22309 ^ n20455 ^ 1'b0 ;
  assign n24904 = ~n24299 & n24903 ;
  assign n24905 = ( n6303 & n6908 ) | ( n6303 & ~n24904 ) | ( n6908 & ~n24904 ) ;
  assign n24906 = n3395 & ~n17550 ;
  assign n24907 = n24906 ^ n18221 ^ n9722 ;
  assign n24908 = n13054 ^ n5609 ^ 1'b0 ;
  assign n24909 = ~n19340 & n24908 ;
  assign n24910 = n24909 ^ n22905 ^ 1'b0 ;
  assign n24911 = n11673 ^ n1673 ^ 1'b0 ;
  assign n24912 = n11022 & n24911 ;
  assign n24913 = n1972 | n9729 ;
  assign n24915 = n3659 | n12101 ;
  assign n24914 = ( ~n1162 & n7905 ) | ( ~n1162 & n20271 ) | ( n7905 & n20271 ) ;
  assign n24916 = n24915 ^ n24914 ^ n14762 ;
  assign n24918 = n3974 ^ n356 ^ 1'b0 ;
  assign n24917 = n8607 & n9618 ;
  assign n24919 = n24918 ^ n24917 ^ n21288 ;
  assign n24920 = ( n9033 & n9547 ) | ( n9033 & ~n19694 ) | ( n9547 & ~n19694 ) ;
  assign n24921 = n13458 ^ n2149 ^ 1'b0 ;
  assign n24922 = ~n3763 & n24921 ;
  assign n24923 = n11189 & n18574 ;
  assign n24924 = n24923 ^ n19852 ^ 1'b0 ;
  assign n24925 = ( n1297 & n3463 ) | ( n1297 & n5166 ) | ( n3463 & n5166 ) ;
  assign n24926 = n16443 | n24925 ;
  assign n24927 = n5589 & n12082 ;
  assign n24928 = n24927 ^ n14221 ^ 1'b0 ;
  assign n24929 = ( n3854 & n4303 ) | ( n3854 & ~n17130 ) | ( n4303 & ~n17130 ) ;
  assign n24930 = ( n7894 & ~n10627 ) | ( n7894 & n24929 ) | ( ~n10627 & n24929 ) ;
  assign n24931 = n24930 ^ n6387 ^ 1'b0 ;
  assign n24932 = n17197 & n24931 ;
  assign n24933 = n3345 | n9521 ;
  assign n24934 = n24932 | n24933 ;
  assign n24935 = n24934 ^ n9047 ^ 1'b0 ;
  assign n24936 = n24928 & n24935 ;
  assign n24937 = n18583 ^ n4430 ^ 1'b0 ;
  assign n24938 = ~n22744 & n24937 ;
  assign n24939 = n1335 ^ n1230 ^ 1'b0 ;
  assign n24940 = n24939 ^ n7333 ^ n3632 ;
  assign n24941 = n22554 ^ n19705 ^ n8392 ;
  assign n24942 = n23385 ^ n15900 ^ n6429 ;
  assign n24943 = n24942 ^ n2597 ^ 1'b0 ;
  assign n24944 = n9646 & n24943 ;
  assign n24945 = n24944 ^ n7021 ^ 1'b0 ;
  assign n24946 = ( n18289 & ~n19719 ) | ( n18289 & n24945 ) | ( ~n19719 & n24945 ) ;
  assign n24947 = n4709 | n4742 ;
  assign n24948 = n24947 ^ n14346 ^ 1'b0 ;
  assign n24949 = n5956 | n24948 ;
  assign n24950 = n11238 | n24949 ;
  assign n24952 = n8415 ^ n5017 ^ n4022 ;
  assign n24951 = n16356 & ~n20796 ;
  assign n24953 = n24952 ^ n24951 ^ 1'b0 ;
  assign n24954 = ~n6475 & n6635 ;
  assign n24955 = n1984 & ~n3390 ;
  assign n24956 = n24955 ^ n11789 ^ n5384 ;
  assign n24957 = n13473 ^ n7803 ^ n1652 ;
  assign n24958 = n288 | n23417 ;
  assign n24959 = n24958 ^ n17123 ^ 1'b0 ;
  assign n24960 = n8050 ^ n7549 ^ 1'b0 ;
  assign n24961 = n24959 & ~n24960 ;
  assign n24962 = n24961 ^ n24068 ^ n5093 ;
  assign n24963 = n15384 | n15724 ;
  assign n24964 = n24583 ^ n8567 ^ 1'b0 ;
  assign n24965 = ~n2126 & n24964 ;
  assign n24966 = n5855 & n7573 ;
  assign n24967 = n17456 ^ n8676 ^ 1'b0 ;
  assign n24968 = n16379 & ~n24967 ;
  assign n24969 = ~n10851 & n24968 ;
  assign n24970 = ~n8952 & n22612 ;
  assign n24971 = n2827 & ~n14484 ;
  assign n24972 = n24971 ^ n8947 ^ n4380 ;
  assign n24973 = ( x45 & ~n9441 ) | ( x45 & n24972 ) | ( ~n9441 & n24972 ) ;
  assign n24974 = n18704 ^ n11207 ^ 1'b0 ;
  assign n24975 = n1491 & ~n9432 ;
  assign n24976 = n24975 ^ n16176 ^ 1'b0 ;
  assign n24977 = n2740 & ~n4088 ;
  assign n24978 = n24977 ^ n6168 ^ 1'b0 ;
  assign n24979 = n10474 & ~n17854 ;
  assign n24980 = n9719 & ~n19052 ;
  assign n24981 = n24980 ^ n12952 ^ 1'b0 ;
  assign n24982 = n16320 | n24981 ;
  assign n24983 = n1582 | n11123 ;
  assign n24984 = n24982 & ~n24983 ;
  assign n24985 = n4021 & ~n6142 ;
  assign n24986 = ~n3106 & n24985 ;
  assign n24987 = n24986 ^ n10290 ^ 1'b0 ;
  assign n24988 = ~n3917 & n15238 ;
  assign n24989 = ~n7625 & n24988 ;
  assign n24994 = n13433 ^ n3471 ^ 1'b0 ;
  assign n24993 = ~n9255 & n12662 ;
  assign n24995 = n24994 ^ n24993 ^ 1'b0 ;
  assign n24990 = n8071 | n18407 ;
  assign n24991 = n22501 | n24990 ;
  assign n24992 = n11415 & n24991 ;
  assign n24996 = n24995 ^ n24992 ^ 1'b0 ;
  assign n24998 = n4942 ^ n1502 ^ n755 ;
  assign n24999 = n7289 | n24998 ;
  assign n25000 = n5490 | n24999 ;
  assign n25001 = n2640 | n25000 ;
  assign n24997 = n5641 | n8736 ;
  assign n25002 = n25001 ^ n24997 ^ 1'b0 ;
  assign n25003 = n20991 ^ n6332 ^ 1'b0 ;
  assign n25004 = ( ~n9655 & n11142 ) | ( ~n9655 & n11730 ) | ( n11142 & n11730 ) ;
  assign n25005 = n9722 ^ n9302 ^ 1'b0 ;
  assign n25006 = n1745 & n25005 ;
  assign n25007 = n20646 ^ n2651 ^ 1'b0 ;
  assign n25008 = n25006 & ~n25007 ;
  assign n25009 = n7775 ^ n2663 ^ 1'b0 ;
  assign n25010 = ( n10484 & n25008 ) | ( n10484 & n25009 ) | ( n25008 & n25009 ) ;
  assign n25013 = n1776 ^ n800 ^ 1'b0 ;
  assign n25014 = n3836 | n25013 ;
  assign n25011 = n5851 ^ n3195 ^ x34 ;
  assign n25012 = n25011 ^ n12779 ^ n1784 ;
  assign n25015 = n25014 ^ n25012 ^ n9782 ;
  assign n25016 = ( ~n12918 & n25010 ) | ( ~n12918 & n25015 ) | ( n25010 & n25015 ) ;
  assign n25017 = n8833 ^ n4993 ^ 1'b0 ;
  assign n25018 = n5530 ^ n1726 ^ 1'b0 ;
  assign n25019 = n8510 & n25018 ;
  assign n25020 = ~n5361 & n20212 ;
  assign n25021 = ~n5436 & n25020 ;
  assign n25022 = n25021 ^ n12250 ^ 1'b0 ;
  assign n25023 = n15781 ^ n10154 ^ 1'b0 ;
  assign n25024 = n8229 | n25023 ;
  assign n25025 = ( ~n8172 & n8668 ) | ( ~n8172 & n25024 ) | ( n8668 & n25024 ) ;
  assign n25026 = n9625 & n24612 ;
  assign n25027 = ~n25025 & n25026 ;
  assign n25028 = ( n6061 & n6890 ) | ( n6061 & ~n14212 ) | ( n6890 & ~n14212 ) ;
  assign n25029 = n1234 | n25028 ;
  assign n25030 = n24843 | n25029 ;
  assign n25031 = n951 & n9625 ;
  assign n25032 = n25031 ^ n7694 ^ 1'b0 ;
  assign n25033 = n11450 | n25032 ;
  assign n25034 = n16246 ^ n12844 ^ 1'b0 ;
  assign n25035 = ~n10929 & n25034 ;
  assign n25036 = n12622 & n25035 ;
  assign n25042 = n1096 ^ n525 ^ 1'b0 ;
  assign n25040 = n2517 & n18249 ;
  assign n25041 = n25040 ^ n4173 ^ 1'b0 ;
  assign n25038 = n13909 ^ n5259 ^ n2144 ;
  assign n25037 = n14556 ^ n13856 ^ 1'b0 ;
  assign n25039 = n25038 ^ n25037 ^ n14957 ;
  assign n25043 = n25042 ^ n25041 ^ n25039 ;
  assign n25045 = ~n6084 & n14186 ;
  assign n25046 = n4310 & n25045 ;
  assign n25047 = n25046 ^ n11095 ^ 1'b0 ;
  assign n25044 = ~n12986 & n16384 ;
  assign n25048 = n25047 ^ n25044 ^ 1'b0 ;
  assign n25049 = n7568 & ~n11913 ;
  assign n25050 = n798 & n25049 ;
  assign n25051 = ~n11291 & n20048 ;
  assign n25052 = n9296 | n12314 ;
  assign n25053 = n4787 ^ n3434 ^ 1'b0 ;
  assign n25054 = n7425 & ~n25053 ;
  assign n25055 = n12571 & n25054 ;
  assign n25056 = n25055 ^ n1745 ^ 1'b0 ;
  assign n25057 = n25056 ^ n20559 ^ n20182 ;
  assign n25058 = ( n15380 & ~n25052 ) | ( n15380 & n25057 ) | ( ~n25052 & n25057 ) ;
  assign n25059 = n4113 ^ n2049 ^ 1'b0 ;
  assign n25060 = n8955 ^ n5536 ^ n1226 ;
  assign n25061 = ( n14240 & n25059 ) | ( n14240 & ~n25060 ) | ( n25059 & ~n25060 ) ;
  assign n25062 = n1264 & ~n4765 ;
  assign n25063 = ( n8009 & n16157 ) | ( n8009 & ~n25062 ) | ( n16157 & ~n25062 ) ;
  assign n25065 = ~n3771 & n8717 ;
  assign n25064 = n3063 & ~n6761 ;
  assign n25066 = n25065 ^ n25064 ^ n18427 ;
  assign n25067 = n19550 ^ n5530 ^ 1'b0 ;
  assign n25068 = n21759 | n25067 ;
  assign n25069 = n8787 & ~n21869 ;
  assign n25070 = n6235 & n8609 ;
  assign n25071 = n839 & n25070 ;
  assign n25072 = n24219 ^ n7148 ^ 1'b0 ;
  assign n25073 = n946 | n8433 ;
  assign n25074 = n12714 | n15379 ;
  assign n25075 = n25074 ^ n3592 ^ 1'b0 ;
  assign n25076 = ( n162 & n8716 ) | ( n162 & ~n17209 ) | ( n8716 & ~n17209 ) ;
  assign n25077 = ~n18903 & n25076 ;
  assign n25078 = n10900 | n25077 ;
  assign n25079 = n4203 | n22015 ;
  assign n25080 = n23151 | n25079 ;
  assign n25081 = ( n3154 & ~n13041 ) | ( n3154 & n25080 ) | ( ~n13041 & n25080 ) ;
  assign n25082 = ~n822 & n14866 ;
  assign n25083 = ~n17661 & n20154 ;
  assign n25084 = n25082 & n25083 ;
  assign n25085 = n25084 ^ n15396 ^ n6614 ;
  assign n25086 = ~n1825 & n4746 ;
  assign n25087 = n25086 ^ n6570 ^ 1'b0 ;
  assign n25088 = n25087 ^ n20338 ^ n3144 ;
  assign n25089 = n25088 ^ n12386 ^ n3637 ;
  assign n25090 = n15925 ^ n10244 ^ 1'b0 ;
  assign n25091 = n25090 ^ n18496 ^ 1'b0 ;
  assign n25092 = n395 | n17267 ;
  assign n25093 = n18235 | n25092 ;
  assign n25095 = n8302 ^ n3961 ^ 1'b0 ;
  assign n25094 = ~n1819 & n15683 ;
  assign n25096 = n25095 ^ n25094 ^ 1'b0 ;
  assign n25097 = n14326 ^ n13865 ^ n222 ;
  assign n25098 = n17971 ^ n14551 ^ n10154 ;
  assign n25099 = n25098 ^ n3469 ^ 1'b0 ;
  assign n25100 = n25097 | n25099 ;
  assign n25101 = n14697 ^ n1242 ^ 1'b0 ;
  assign n25102 = ( n6808 & n8573 ) | ( n6808 & n15642 ) | ( n8573 & n15642 ) ;
  assign n25103 = n25102 ^ n473 ^ 1'b0 ;
  assign n25104 = x75 & ~n3294 ;
  assign n25105 = ~n7592 & n25104 ;
  assign n25106 = ( ~n4724 & n24816 ) | ( ~n4724 & n25105 ) | ( n24816 & n25105 ) ;
  assign n25107 = n3626 | n25106 ;
  assign n25108 = n25107 ^ n820 ^ 1'b0 ;
  assign n25109 = n25108 ^ n11734 ^ n7095 ;
  assign n25110 = n1285 ^ n862 ^ 1'b0 ;
  assign n25111 = ( ~n14517 & n23115 ) | ( ~n14517 & n25110 ) | ( n23115 & n25110 ) ;
  assign n25112 = n2782 & n7029 ;
  assign n25113 = n25112 ^ n17698 ^ n484 ;
  assign n25114 = n9405 & n13618 ;
  assign n25115 = n4180 & n25114 ;
  assign n25116 = n2516 & ~n3610 ;
  assign n25117 = ~n12112 & n25116 ;
  assign n25118 = n24830 ^ n22334 ^ 1'b0 ;
  assign n25119 = ~n1834 & n12706 ;
  assign n25120 = n6228 & n8007 ;
  assign n25121 = n25120 ^ n1104 ^ 1'b0 ;
  assign n25122 = n4927 & n5131 ;
  assign n25123 = n6424 ^ x98 ^ 1'b0 ;
  assign n25124 = n25123 ^ n4956 ^ 1'b0 ;
  assign n25125 = n180 | n20280 ;
  assign n25126 = n6126 & ~n25125 ;
  assign n25127 = n2912 & ~n7216 ;
  assign n25128 = n16621 & n25127 ;
  assign n25129 = n9409 ^ n5703 ^ 1'b0 ;
  assign n25132 = n2960 | n7616 ;
  assign n25130 = ~n474 & n6117 ;
  assign n25131 = n25130 ^ n5422 ^ n3636 ;
  assign n25133 = n25132 ^ n25131 ^ n11246 ;
  assign n25134 = n11046 ^ n4739 ^ 1'b0 ;
  assign n25135 = n3988 & n6570 ;
  assign n25136 = n11478 & n16526 ;
  assign n25137 = n25135 & n25136 ;
  assign n25138 = n8830 & n10071 ;
  assign n25139 = n5950 & n25138 ;
  assign n25147 = n614 & ~n1074 ;
  assign n25148 = ~n5458 & n25147 ;
  assign n25149 = ( n3293 & ~n10873 ) | ( n3293 & n25148 ) | ( ~n10873 & n25148 ) ;
  assign n25143 = n9572 | n16350 ;
  assign n25144 = n10808 | n25143 ;
  assign n25140 = n4840 | n6830 ;
  assign n25141 = n25140 ^ n903 ^ 1'b0 ;
  assign n25142 = n10304 & n25141 ;
  assign n25145 = n25144 ^ n25142 ^ n1323 ;
  assign n25146 = n11697 | n25145 ;
  assign n25150 = n25149 ^ n25146 ^ 1'b0 ;
  assign n25151 = ( n1022 & n16131 ) | ( n1022 & n17185 ) | ( n16131 & n17185 ) ;
  assign n25152 = n25151 ^ n19775 ^ n17694 ;
  assign n25153 = n16733 ^ n11960 ^ n9086 ;
  assign n25154 = n9628 & ~n16096 ;
  assign n25155 = n25154 ^ n6052 ^ 1'b0 ;
  assign n25156 = n25155 ^ n2617 ^ 1'b0 ;
  assign n25157 = n6652 & n10885 ;
  assign n25158 = ( ~n2965 & n8731 ) | ( ~n2965 & n25157 ) | ( n8731 & n25157 ) ;
  assign n25159 = ( ~n1463 & n16079 ) | ( ~n1463 & n17231 ) | ( n16079 & n17231 ) ;
  assign n25160 = n12325 | n25159 ;
  assign n25161 = n12381 ^ n5119 ^ 1'b0 ;
  assign n25162 = n4817 | n25161 ;
  assign n25163 = ( n2296 & n19640 ) | ( n2296 & ~n24709 ) | ( n19640 & ~n24709 ) ;
  assign n25165 = n20047 & ~n20738 ;
  assign n25164 = n7332 | n18595 ;
  assign n25166 = n25165 ^ n25164 ^ 1'b0 ;
  assign n25167 = n15750 | n25166 ;
  assign n25168 = n3261 & ~n10484 ;
  assign n25169 = ( n3027 & ~n3634 ) | ( n3027 & n25168 ) | ( ~n3634 & n25168 ) ;
  assign n25170 = ~n8050 & n19061 ;
  assign n25171 = n24945 ^ n11937 ^ 1'b0 ;
  assign n25172 = n10903 ^ n8306 ^ 1'b0 ;
  assign n25173 = n15342 & ~n25172 ;
  assign n25174 = n14655 ^ n2870 ^ 1'b0 ;
  assign n25175 = n1061 & n10658 ;
  assign n25176 = n20093 ^ n1368 ^ 1'b0 ;
  assign n25177 = n11531 ^ n10994 ^ 1'b0 ;
  assign n25178 = n3264 | n3358 ;
  assign n25179 = n25178 ^ n21619 ^ 1'b0 ;
  assign n25180 = n2265 | n25179 ;
  assign n25181 = n11309 ^ n10300 ^ 1'b0 ;
  assign n25182 = n7410 | n12550 ;
  assign n25183 = n25182 ^ n7614 ^ 1'b0 ;
  assign n25184 = n4633 ^ x22 ^ 1'b0 ;
  assign n25185 = n18627 | n24481 ;
  assign n25186 = n25185 ^ n10131 ^ 1'b0 ;
  assign n25187 = n312 & ~n17014 ;
  assign n25188 = n1441 & n15570 ;
  assign n25189 = ( n12187 & n24872 ) | ( n12187 & n25188 ) | ( n24872 & n25188 ) ;
  assign n25190 = ( ~n362 & n8056 ) | ( ~n362 & n25189 ) | ( n8056 & n25189 ) ;
  assign n25191 = n11179 | n14166 ;
  assign n25192 = ~n1795 & n9448 ;
  assign n25193 = n25192 ^ n16903 ^ 1'b0 ;
  assign n25194 = n1608 & ~n8639 ;
  assign n25195 = ~n2501 & n25194 ;
  assign n25196 = n14455 ^ n9313 ^ 1'b0 ;
  assign n25197 = ~n25195 & n25196 ;
  assign n25198 = n1035 & ~n5615 ;
  assign n25199 = n10431 & n25198 ;
  assign n25200 = ~n14531 & n18340 ;
  assign n25201 = n845 | n5796 ;
  assign n25202 = n25201 ^ n8516 ^ 1'b0 ;
  assign n25203 = n313 & n4501 ;
  assign n25204 = ~n7393 & n25203 ;
  assign n25205 = n2012 & n17036 ;
  assign n25206 = n1611 & n25205 ;
  assign n25207 = n6451 & ~n11114 ;
  assign n25208 = n25207 ^ n9367 ^ 1'b0 ;
  assign n25209 = n1285 & ~n25208 ;
  assign n25210 = n11971 & n20772 ;
  assign n25211 = n25210 ^ n5880 ^ 1'b0 ;
  assign n25212 = n25211 ^ n5691 ^ 1'b0 ;
  assign n25213 = ~n1062 & n18198 ;
  assign n25214 = n11444 ^ n4489 ^ 1'b0 ;
  assign n25215 = n10502 & n20654 ;
  assign n25216 = n16264 & n25215 ;
  assign n25217 = n11786 ^ n6687 ^ n4283 ;
  assign n25218 = ~n4239 & n8255 ;
  assign n25219 = n25218 ^ n11345 ^ 1'b0 ;
  assign n25220 = n5448 & ~n25219 ;
  assign n25221 = n18707 & n25220 ;
  assign n25222 = n16611 & ~n21280 ;
  assign n25223 = n10177 & n25222 ;
  assign n25224 = n13822 ^ n5723 ^ 1'b0 ;
  assign n25225 = ( n6808 & ~n8114 ) | ( n6808 & n14012 ) | ( ~n8114 & n14012 ) ;
  assign n25226 = n19211 | n25225 ;
  assign n25227 = n3717 & ~n4600 ;
  assign n25228 = n25227 ^ n21254 ^ n16703 ;
  assign n25229 = n25228 ^ n17333 ^ 1'b0 ;
  assign n25230 = ( ~n12727 & n15676 ) | ( ~n12727 & n21447 ) | ( n15676 & n21447 ) ;
  assign n25231 = n17071 ^ n2054 ^ 1'b0 ;
  assign n25232 = n16042 & n25231 ;
  assign n25233 = ~n3027 & n16291 ;
  assign n25234 = ~n2041 & n25233 ;
  assign n25235 = n12219 | n24589 ;
  assign n25236 = n6332 ^ n4356 ^ 1'b0 ;
  assign n25237 = n12765 & ~n13222 ;
  assign n25238 = n25237 ^ n14438 ^ 1'b0 ;
  assign n25239 = ~n1631 & n8910 ;
  assign n25240 = n4591 & n9116 ;
  assign n25241 = n9818 & n25240 ;
  assign n25242 = n22028 & n25241 ;
  assign n25243 = ( n9548 & n10065 ) | ( n9548 & n24100 ) | ( n10065 & n24100 ) ;
  assign n25244 = ~n5461 & n25243 ;
  assign n25245 = n14149 ^ n6146 ^ n1461 ;
  assign n25246 = n25245 ^ n11870 ^ n6199 ;
  assign n25247 = n19522 ^ n5861 ^ n3090 ;
  assign n25248 = n6820 & ~n25247 ;
  assign n25249 = ~n7964 & n25248 ;
  assign n25250 = n360 & ~n2158 ;
  assign n25251 = ( ~n22326 & n25249 ) | ( ~n22326 & n25250 ) | ( n25249 & n25250 ) ;
  assign n25252 = n24986 ^ n11292 ^ 1'b0 ;
  assign n25253 = n3781 & n25252 ;
  assign n25254 = n17766 | n19641 ;
  assign n25255 = n25254 ^ n18187 ^ n3450 ;
  assign n25256 = n7054 | n10651 ;
  assign n25257 = n25256 ^ n20646 ^ 1'b0 ;
  assign n25258 = n18731 ^ n1752 ^ 1'b0 ;
  assign n25259 = ( n4452 & n5306 ) | ( n4452 & n25258 ) | ( n5306 & n25258 ) ;
  assign n25260 = ~n4550 & n5338 ;
  assign n25261 = ~n25259 & n25260 ;
  assign n25262 = n9619 ^ n3847 ^ 1'b0 ;
  assign n25263 = n704 | n25262 ;
  assign n25264 = n8201 ^ n4591 ^ 1'b0 ;
  assign n25265 = n24477 ^ n2854 ^ 1'b0 ;
  assign n25266 = n1842 & ~n11737 ;
  assign n25267 = ~n25265 & n25266 ;
  assign n25268 = n4839 | n10553 ;
  assign n25269 = n11432 ^ n4713 ^ n3230 ;
  assign n25270 = n22714 & n23530 ;
  assign n25271 = n3391 ^ n1712 ^ 1'b0 ;
  assign n25272 = ~n3388 & n25271 ;
  assign n25273 = n7303 & n20421 ;
  assign n25274 = n25273 ^ n8064 ^ 1'b0 ;
  assign n25276 = n11365 ^ n7189 ^ 1'b0 ;
  assign n25277 = n4365 | n25276 ;
  assign n25275 = n5772 & ~n19762 ;
  assign n25278 = n25277 ^ n25275 ^ 1'b0 ;
  assign n25279 = n15205 ^ n12646 ^ n4318 ;
  assign n25280 = n7989 ^ n4417 ^ 1'b0 ;
  assign n25281 = n3836 ^ n858 ^ 1'b0 ;
  assign n25282 = n25280 & n25281 ;
  assign n25283 = ~n13989 & n25282 ;
  assign n25284 = n5890 | n11035 ;
  assign n25285 = x2 | n25284 ;
  assign n25287 = ( ~n1558 & n8805 ) | ( ~n1558 & n16398 ) | ( n8805 & n16398 ) ;
  assign n25286 = n6787 & n10815 ;
  assign n25288 = n25287 ^ n25286 ^ 1'b0 ;
  assign n25289 = n25288 ^ n10074 ^ 1'b0 ;
  assign n25290 = n3533 | n25289 ;
  assign n25291 = n14546 | n21447 ;
  assign n25292 = n24803 ^ n5053 ^ 1'b0 ;
  assign n25293 = n20801 ^ n10992 ^ 1'b0 ;
  assign n25294 = ~n20730 & n25293 ;
  assign n25295 = n8477 & ~n13983 ;
  assign n25296 = n11572 ^ n6659 ^ 1'b0 ;
  assign n25297 = n9275 ^ n2534 ^ 1'b0 ;
  assign n25298 = n4911 & ~n25297 ;
  assign n25299 = n14631 ^ n3564 ^ 1'b0 ;
  assign n25300 = n11616 ^ n4032 ^ 1'b0 ;
  assign n25301 = ( n25298 & ~n25299 ) | ( n25298 & n25300 ) | ( ~n25299 & n25300 ) ;
  assign n25302 = n9492 ^ n3722 ^ 1'b0 ;
  assign n25303 = n25302 ^ n11035 ^ 1'b0 ;
  assign n25304 = n17127 ^ n7284 ^ n1864 ;
  assign n25305 = n5642 ^ n841 ^ 1'b0 ;
  assign n25306 = n25304 & ~n25305 ;
  assign n25307 = ~n6858 & n25306 ;
  assign n25308 = n18509 ^ n3012 ^ n815 ;
  assign n25309 = n25307 & n25308 ;
  assign n25310 = n6300 | n25309 ;
  assign n25311 = n8787 & n16393 ;
  assign n25312 = n2106 & n25311 ;
  assign n25313 = n4658 & n5403 ;
  assign n25314 = ~n25312 & n25313 ;
  assign n25315 = n9759 ^ n6935 ^ 1'b0 ;
  assign n25316 = n2568 | n25315 ;
  assign n25317 = n8192 ^ n8027 ^ n1971 ;
  assign n25318 = ~n2224 & n23041 ;
  assign n25324 = n1515 & ~n5274 ;
  assign n25319 = n21708 ^ n10260 ^ n7348 ;
  assign n25320 = n1198 | n2077 ;
  assign n25321 = n25319 | n25320 ;
  assign n25322 = n25321 ^ n9850 ^ 1'b0 ;
  assign n25323 = n7147 | n25322 ;
  assign n25325 = n25324 ^ n25323 ^ 1'b0 ;
  assign n25326 = ( n6808 & ~n20546 ) | ( n6808 & n23953 ) | ( ~n20546 & n23953 ) ;
  assign n25329 = n4679 & n5225 ;
  assign n25330 = n2095 & n25329 ;
  assign n25331 = n4122 | n6897 ;
  assign n25332 = n25330 & ~n25331 ;
  assign n25327 = x52 | n1137 ;
  assign n25328 = ( n1231 & n6480 ) | ( n1231 & ~n25327 ) | ( n6480 & ~n25327 ) ;
  assign n25333 = n25332 ^ n25328 ^ 1'b0 ;
  assign n25334 = n14275 & n25333 ;
  assign n25335 = n21059 ^ n11665 ^ 1'b0 ;
  assign n25336 = n571 & ~n19368 ;
  assign n25337 = n12542 ^ n6243 ^ 1'b0 ;
  assign n25338 = n2432 & n3933 ;
  assign n25339 = n7702 & n15234 ;
  assign n25340 = n18253 ^ n4394 ^ n2515 ;
  assign n25341 = n7592 & n9983 ;
  assign n25342 = n4679 & n25341 ;
  assign n25343 = n25342 ^ n14150 ^ 1'b0 ;
  assign n25344 = n13386 | n20760 ;
  assign n25345 = n4234 | n25344 ;
  assign n25346 = n6003 & n10753 ;
  assign n25354 = ( n1034 & n16180 ) | ( n1034 & ~n20850 ) | ( n16180 & ~n20850 ) ;
  assign n25347 = n6908 & n12027 ;
  assign n25348 = ~n20676 & n25347 ;
  assign n25349 = n5761 & n6890 ;
  assign n25350 = n25349 ^ n6668 ^ 1'b0 ;
  assign n25351 = n25350 ^ n18227 ^ 1'b0 ;
  assign n25352 = n25348 | n25351 ;
  assign n25353 = n25352 ^ n14782 ^ 1'b0 ;
  assign n25355 = n25354 ^ n25353 ^ 1'b0 ;
  assign n25357 = ( n1528 & ~n10593 ) | ( n1528 & n10783 ) | ( ~n10593 & n10783 ) ;
  assign n25356 = n15804 ^ n10971 ^ 1'b0 ;
  assign n25358 = n25357 ^ n25356 ^ n14066 ;
  assign n25359 = n6851 ^ n5658 ^ n1874 ;
  assign n25360 = n7747 & n11805 ;
  assign n25361 = n6299 & n25360 ;
  assign n25362 = n9379 ^ n1371 ^ 1'b0 ;
  assign n25363 = ~n20698 & n23026 ;
  assign n25364 = ( ~n25361 & n25362 ) | ( ~n25361 & n25363 ) | ( n25362 & n25363 ) ;
  assign n25365 = n6774 ^ n4529 ^ 1'b0 ;
  assign n25366 = n3459 & n25365 ;
  assign n25367 = n25366 ^ n19445 ^ 1'b0 ;
  assign n25368 = n4562 | n15068 ;
  assign n25369 = n25368 ^ n17761 ^ n14462 ;
  assign n25370 = n4404 | n25369 ;
  assign n25371 = n25370 ^ n18348 ^ 1'b0 ;
  assign n25372 = n13623 | n17717 ;
  assign n25373 = ~n9855 & n13832 ;
  assign n25374 = ( n19506 & n23706 ) | ( n19506 & n25373 ) | ( n23706 & n25373 ) ;
  assign n25375 = ~n25372 & n25374 ;
  assign n25376 = ~n9560 & n21416 ;
  assign n25377 = n25376 ^ n10021 ^ 1'b0 ;
  assign n25378 = n15259 & n24066 ;
  assign n25379 = n2226 & n4349 ;
  assign n25380 = n25379 ^ n5060 ^ 1'b0 ;
  assign n25381 = ~n13340 & n18436 ;
  assign n25382 = n25380 & n25381 ;
  assign n25383 = ( n3098 & n20721 ) | ( n3098 & ~n25382 ) | ( n20721 & ~n25382 ) ;
  assign n25384 = x113 & ~n12280 ;
  assign n25385 = n8814 ^ n459 ^ 1'b0 ;
  assign n25386 = n1104 & ~n25385 ;
  assign n25387 = n6966 | n18687 ;
  assign n25388 = n2200 & ~n25387 ;
  assign n25389 = n11576 ^ n8036 ^ 1'b0 ;
  assign n25390 = ( n10713 & n18846 ) | ( n10713 & ~n20515 ) | ( n18846 & ~n20515 ) ;
  assign n25391 = n8126 ^ n4139 ^ x58 ;
  assign n25392 = n9436 ^ n9359 ^ n5358 ;
  assign n25393 = n9573 | n22140 ;
  assign n25394 = n25392 | n25393 ;
  assign n25395 = n10913 ^ n6357 ^ 1'b0 ;
  assign n25396 = n19659 & ~n25395 ;
  assign n25397 = ~n19219 & n19674 ;
  assign n25398 = ~n12430 & n25397 ;
  assign n25399 = n25149 ^ n22390 ^ 1'b0 ;
  assign n25400 = ~n6084 & n21294 ;
  assign n25401 = n25400 ^ n14630 ^ 1'b0 ;
  assign n25402 = n19876 ^ n8709 ^ n701 ;
  assign n25403 = ( n815 & n10074 ) | ( n815 & n18109 ) | ( n10074 & n18109 ) ;
  assign n25404 = n25403 ^ n23413 ^ n15827 ;
  assign n25405 = ~n2902 & n25404 ;
  assign n25406 = n24717 ^ n6560 ^ 1'b0 ;
  assign n25407 = n16835 ^ n5484 ^ 1'b0 ;
  assign n25408 = n20293 ^ n18324 ^ n15743 ;
  assign n25409 = n11044 | n25408 ;
  assign n25410 = n13830 & ~n25409 ;
  assign n25411 = n6720 ^ n3984 ^ n2698 ;
  assign n25412 = n25411 ^ n22668 ^ 1'b0 ;
  assign n25413 = n18196 | n25412 ;
  assign n25415 = n6042 | n14228 ;
  assign n25416 = n5154 & ~n25415 ;
  assign n25414 = ~n1918 & n19640 ;
  assign n25417 = n25416 ^ n25414 ^ 1'b0 ;
  assign n25419 = n8819 | n17061 ;
  assign n25420 = n25419 ^ n10878 ^ 1'b0 ;
  assign n25418 = n4966 & ~n9751 ;
  assign n25421 = n25420 ^ n25418 ^ 1'b0 ;
  assign n25422 = n25421 ^ n13824 ^ 1'b0 ;
  assign n25423 = n12822 & n25422 ;
  assign n25424 = n22136 & ~n23422 ;
  assign n25425 = n25424 ^ n13587 ^ 1'b0 ;
  assign n25426 = n7311 & ~n16565 ;
  assign n25427 = n25426 ^ n353 ^ 1'b0 ;
  assign n25428 = n13806 ^ n5212 ^ 1'b0 ;
  assign n25429 = ( x26 & ~n25427 ) | ( x26 & n25428 ) | ( ~n25427 & n25428 ) ;
  assign n25430 = n25429 ^ n19089 ^ n1640 ;
  assign n25431 = n10607 & ~n14490 ;
  assign n25432 = ~n2064 & n7962 ;
  assign n25433 = n7274 & n10908 ;
  assign n25434 = n24746 ^ n1099 ^ 1'b0 ;
  assign n25435 = n25433 & n25434 ;
  assign n25436 = n15880 ^ n195 ^ 1'b0 ;
  assign n25437 = n6393 | n13892 ;
  assign n25438 = n630 & n25437 ;
  assign n25439 = n17124 & n25438 ;
  assign n25440 = n2746 | n5399 ;
  assign n25441 = n13423 & ~n25440 ;
  assign n25442 = n9772 & ~n25441 ;
  assign n25443 = n25442 ^ n22595 ^ n17342 ;
  assign n25444 = n1669 & ~n8243 ;
  assign n25445 = ~n6426 & n25444 ;
  assign n25446 = n7131 | n16995 ;
  assign n25447 = n25446 ^ n1047 ^ 1'b0 ;
  assign n25448 = n25447 ^ n5395 ^ 1'b0 ;
  assign n25449 = n25448 ^ n23717 ^ 1'b0 ;
  assign n25450 = n16056 ^ n4224 ^ n803 ;
  assign n25451 = n6651 ^ x47 ^ 1'b0 ;
  assign n25452 = ( n1903 & ~n2855 ) | ( n1903 & n5807 ) | ( ~n2855 & n5807 ) ;
  assign n25453 = ~n7586 & n25452 ;
  assign n25454 = n7504 & ~n11856 ;
  assign n25455 = n340 & n25454 ;
  assign n25456 = n5984 | n23057 ;
  assign n25457 = n25456 ^ n14599 ^ 1'b0 ;
  assign n25458 = ( n13719 & ~n25455 ) | ( n13719 & n25457 ) | ( ~n25455 & n25457 ) ;
  assign n25459 = n25458 ^ n25149 ^ 1'b0 ;
  assign n25460 = n10360 ^ n4777 ^ 1'b0 ;
  assign n25461 = n13110 ^ n12618 ^ 1'b0 ;
  assign n25462 = ~n13772 & n20852 ;
  assign n25463 = n25462 ^ n13904 ^ 1'b0 ;
  assign n25464 = n4678 & ~n12535 ;
  assign n25465 = n25464 ^ n22589 ^ n10014 ;
  assign n25466 = n14560 ^ n4760 ^ n4133 ;
  assign n25467 = n25466 ^ n16053 ^ n3630 ;
  assign n25468 = ( n2028 & ~n14763 ) | ( n2028 & n17430 ) | ( ~n14763 & n17430 ) ;
  assign n25469 = n13972 ^ n4749 ^ 1'b0 ;
  assign n25470 = ~n8423 & n25469 ;
  assign n25471 = ~n6679 & n12280 ;
  assign n25472 = n18958 ^ n3887 ^ 1'b0 ;
  assign n25473 = ~n25471 & n25472 ;
  assign n25474 = n13984 & ~n15187 ;
  assign n25475 = n7273 & n25474 ;
  assign n25476 = n5287 | n25475 ;
  assign n25477 = n25476 ^ n12804 ^ 1'b0 ;
  assign n25478 = n3254 & ~n9807 ;
  assign n25479 = ~n16548 & n25478 ;
  assign n25480 = n25479 ^ n22313 ^ 1'b0 ;
  assign n25481 = ( n13425 & n21726 ) | ( n13425 & ~n25480 ) | ( n21726 & ~n25480 ) ;
  assign n25482 = n2868 ^ n1212 ^ 1'b0 ;
  assign n25483 = n7141 ^ n1589 ^ 1'b0 ;
  assign n25484 = ( ~n4583 & n24878 ) | ( ~n4583 & n25483 ) | ( n24878 & n25483 ) ;
  assign n25485 = ~n7798 & n10467 ;
  assign n25486 = n25485 ^ n24863 ^ 1'b0 ;
  assign n25487 = n20381 ^ n746 ^ 1'b0 ;
  assign n25488 = n14039 | n25487 ;
  assign n25489 = n17139 ^ n5438 ^ 1'b0 ;
  assign n25490 = ~n5855 & n25489 ;
  assign n25491 = n3341 & ~n22165 ;
  assign n25492 = n25491 ^ n4211 ^ 1'b0 ;
  assign n25493 = n16770 ^ n3436 ^ 1'b0 ;
  assign n25494 = ~n2095 & n25493 ;
  assign n25495 = n7060 ^ n5533 ^ 1'b0 ;
  assign n25496 = n162 & n25495 ;
  assign n25497 = ~n23481 & n25496 ;
  assign n25498 = ( n2728 & ~n6950 ) | ( n2728 & n25497 ) | ( ~n6950 & n25497 ) ;
  assign n25501 = ~n1136 & n15418 ;
  assign n25502 = n25501 ^ n20954 ^ 1'b0 ;
  assign n25499 = n387 & n6826 ;
  assign n25500 = n25499 ^ n4188 ^ 1'b0 ;
  assign n25503 = n25502 ^ n25500 ^ n15381 ;
  assign n25504 = n2657 | n9168 ;
  assign n25505 = n25504 ^ n12264 ^ 1'b0 ;
  assign n25506 = n25505 ^ n14981 ^ n2628 ;
  assign n25508 = n10598 | n13782 ;
  assign n25507 = ~n303 & n18781 ;
  assign n25509 = n25508 ^ n25507 ^ 1'b0 ;
  assign n25510 = n2554 | n6052 ;
  assign n25511 = n4214 & ~n9587 ;
  assign n25512 = ~n21561 & n25511 ;
  assign n25514 = n219 & ~n1325 ;
  assign n25513 = n6412 & n15972 ;
  assign n25515 = n25514 ^ n25513 ^ 1'b0 ;
  assign n25516 = ( ~n584 & n6915 ) | ( ~n584 & n9554 ) | ( n6915 & n9554 ) ;
  assign n25517 = n10959 ^ n9778 ^ n6196 ;
  assign n25518 = n6124 | n22612 ;
  assign n25519 = n15414 | n15822 ;
  assign n25520 = ( ~n1086 & n1259 ) | ( ~n1086 & n1893 ) | ( n1259 & n1893 ) ;
  assign n25521 = n25520 ^ n19634 ^ 1'b0 ;
  assign n25522 = n15075 | n25521 ;
  assign n25523 = n8227 | n25522 ;
  assign n25524 = n25523 ^ n20366 ^ 1'b0 ;
  assign n25525 = n5681 | n6549 ;
  assign n25526 = n1227 ^ n365 ^ 1'b0 ;
  assign n25527 = ( n5032 & n17313 ) | ( n5032 & ~n25526 ) | ( n17313 & ~n25526 ) ;
  assign n25528 = n21491 ^ n13219 ^ n5528 ;
  assign n25529 = n25528 ^ n15707 ^ n13328 ;
  assign n25530 = n25529 ^ n20527 ^ 1'b0 ;
  assign n25531 = n14755 ^ n8137 ^ 1'b0 ;
  assign n25532 = n4687 & n19173 ;
  assign n25533 = n25532 ^ n6159 ^ 1'b0 ;
  assign n25534 = n12442 & n19044 ;
  assign n25535 = n19483 ^ n4610 ^ 1'b0 ;
  assign n25536 = ~n1410 & n25535 ;
  assign n25537 = n1129 & ~n21280 ;
  assign n25538 = ( n153 & n478 ) | ( n153 & n2219 ) | ( n478 & n2219 ) ;
  assign n25539 = n10567 | n13827 ;
  assign n25540 = n25538 | n25539 ;
  assign n25541 = ~n6717 & n25540 ;
  assign n25542 = n6717 & n25541 ;
  assign n25543 = n25542 ^ n10398 ^ 1'b0 ;
  assign n25544 = n3050 ^ n1057 ^ 1'b0 ;
  assign n25545 = n25543 & n25544 ;
  assign n25546 = n25545 ^ n6425 ^ n5565 ;
  assign n25547 = ( n13742 & ~n19021 ) | ( n13742 & n25546 ) | ( ~n19021 & n25546 ) ;
  assign n25549 = ( ~n1347 & n4596 ) | ( ~n1347 & n6447 ) | ( n4596 & n6447 ) ;
  assign n25548 = n6274 ^ n4826 ^ 1'b0 ;
  assign n25550 = n25549 ^ n25548 ^ n1871 ;
  assign n25551 = n14585 & n25550 ;
  assign n25552 = ~n8870 & n25551 ;
  assign n25554 = ~n6859 & n13246 ;
  assign n25555 = n4884 ^ n3578 ^ 1'b0 ;
  assign n25556 = n23840 | n25555 ;
  assign n25557 = n25554 & ~n25556 ;
  assign n25553 = n16702 & n18488 ;
  assign n25558 = n25557 ^ n25553 ^ 1'b0 ;
  assign n25559 = n25558 ^ n22933 ^ 1'b0 ;
  assign n25560 = ( n265 & n13168 ) | ( n265 & n21460 ) | ( n13168 & n21460 ) ;
  assign n25561 = n25560 ^ n17966 ^ 1'b0 ;
  assign n25562 = n25561 ^ n10758 ^ 1'b0 ;
  assign n25563 = n20970 & ~n25562 ;
  assign n25564 = n21023 ^ n3620 ^ 1'b0 ;
  assign n25565 = ~n13541 & n25564 ;
  assign n25566 = n4065 ^ n154 ^ 1'b0 ;
  assign n25567 = n15634 | n25566 ;
  assign n25568 = n7219 & ~n25567 ;
  assign n25569 = ~n9734 & n21596 ;
  assign n25570 = n17474 & n25569 ;
  assign n25571 = ~n11966 & n20442 ;
  assign n25572 = n25570 & n25571 ;
  assign n25573 = n653 & ~n23767 ;
  assign n25574 = n6966 & n25573 ;
  assign n25575 = n5702 & ~n25038 ;
  assign n25576 = n12666 & n25575 ;
  assign n25577 = ( n846 & n6834 ) | ( n846 & n25576 ) | ( n6834 & n25576 ) ;
  assign n25578 = n7406 ^ n7189 ^ 1'b0 ;
  assign n25579 = n21843 ^ n9912 ^ 1'b0 ;
  assign n25580 = ( n9651 & ~n25578 ) | ( n9651 & n25579 ) | ( ~n25578 & n25579 ) ;
  assign n25581 = n14064 ^ n4926 ^ n933 ;
  assign n25582 = ~n17758 & n23428 ;
  assign n25583 = n25582 ^ n15300 ^ 1'b0 ;
  assign n25584 = n25581 & n25583 ;
  assign n25585 = n22063 ^ n393 ^ 1'b0 ;
  assign n25586 = n18689 ^ n9226 ^ 1'b0 ;
  assign n25587 = n10387 ^ n3745 ^ n2811 ;
  assign n25588 = n20516 & n25587 ;
  assign n25589 = ~n635 & n25588 ;
  assign n25591 = n18683 ^ n8177 ^ 1'b0 ;
  assign n25590 = n13853 ^ n1000 ^ 1'b0 ;
  assign n25592 = n25591 ^ n25590 ^ n18340 ;
  assign n25593 = n2029 & n4871 ;
  assign n25594 = n23687 ^ n3384 ^ n1023 ;
  assign n25595 = n25594 ^ n4063 ^ n2306 ;
  assign n25596 = ( ~n12264 & n15283 ) | ( ~n12264 & n25595 ) | ( n15283 & n25595 ) ;
  assign n25597 = n10369 | n11296 ;
  assign n25598 = n25597 ^ n24767 ^ 1'b0 ;
  assign n25599 = n8511 ^ n1341 ^ 1'b0 ;
  assign n25600 = n9606 | n12788 ;
  assign n25601 = n25600 ^ n3666 ^ 1'b0 ;
  assign n25602 = ~n5421 & n8785 ;
  assign n25603 = n22825 & ~n25602 ;
  assign n25604 = ~n18058 & n25603 ;
  assign n25605 = n7170 | n16667 ;
  assign n25606 = ~n1634 & n12154 ;
  assign n25607 = n25606 ^ n11136 ^ 1'b0 ;
  assign n25608 = n1298 & n19877 ;
  assign n25609 = n19891 ^ n7104 ^ 1'b0 ;
  assign n25610 = ( n5863 & ~n13515 ) | ( n5863 & n16667 ) | ( ~n13515 & n16667 ) ;
  assign n25611 = n7956 ^ n5940 ^ 1'b0 ;
  assign n25612 = n1778 & ~n25611 ;
  assign n25613 = ( n589 & ~n12372 ) | ( n589 & n25612 ) | ( ~n12372 & n25612 ) ;
  assign n25614 = n15339 ^ n3980 ^ n207 ;
  assign n25615 = n2621 | n25614 ;
  assign n25616 = n17771 | n25615 ;
  assign n25617 = n25616 ^ n2155 ^ 1'b0 ;
  assign n25618 = n25617 ^ n4415 ^ 1'b0 ;
  assign n25619 = n21915 ^ n20352 ^ n10931 ;
  assign n25620 = n25619 ^ n14191 ^ 1'b0 ;
  assign n25621 = n22273 & n25620 ;
  assign n25622 = n12358 | n15388 ;
  assign n25623 = n25622 ^ n13019 ^ 1'b0 ;
  assign n25624 = n12584 ^ n5669 ^ n3753 ;
  assign n25625 = ~n14612 & n25624 ;
  assign n25626 = n23177 ^ n11241 ^ 1'b0 ;
  assign n25627 = n12071 & n12657 ;
  assign n25628 = n25627 ^ n20533 ^ n12734 ;
  assign n25629 = n12206 | n12780 ;
  assign n25630 = n11302 & ~n25629 ;
  assign n25631 = ( ~n24753 & n25628 ) | ( ~n24753 & n25630 ) | ( n25628 & n25630 ) ;
  assign n25632 = n4828 | n17482 ;
  assign n25633 = n25632 ^ n15660 ^ 1'b0 ;
  assign n25634 = n5306 & n8209 ;
  assign n25635 = ~n3147 & n25634 ;
  assign n25636 = n20429 & ~n25635 ;
  assign n25637 = n25636 ^ n3111 ^ 1'b0 ;
  assign n25638 = ~n9358 & n9888 ;
  assign n25639 = n13475 ^ n8126 ^ n7016 ;
  assign n25640 = n16274 & ~n18202 ;
  assign n25641 = n25639 & ~n25640 ;
  assign n25642 = ( n2552 & n16489 ) | ( n2552 & n18353 ) | ( n16489 & n18353 ) ;
  assign n25644 = ( ~n4742 & n5747 ) | ( ~n4742 & n21824 ) | ( n5747 & n21824 ) ;
  assign n25643 = n4476 & ~n10008 ;
  assign n25645 = n25644 ^ n25643 ^ 1'b0 ;
  assign n25646 = n25645 ^ n15786 ^ n14572 ;
  assign n25647 = n6070 | n10177 ;
  assign n25648 = n21427 & n25647 ;
  assign n25649 = n25648 ^ n17346 ^ 1'b0 ;
  assign n25652 = n5093 ^ n3575 ^ 1'b0 ;
  assign n25650 = n6948 & ~n25624 ;
  assign n25651 = ~n11127 & n25650 ;
  assign n25653 = n25652 ^ n25651 ^ 1'b0 ;
  assign n25654 = n22308 ^ n20819 ^ x99 ;
  assign n25655 = n3699 | n25654 ;
  assign n25656 = n11946 & ~n15841 ;
  assign n25657 = n25656 ^ n11103 ^ 1'b0 ;
  assign n25658 = n5857 | n25657 ;
  assign n25659 = n22337 ^ n5394 ^ 1'b0 ;
  assign n25660 = n22498 | n25659 ;
  assign n25661 = n25660 ^ n15824 ^ 1'b0 ;
  assign n25662 = n16489 & n21258 ;
  assign n25663 = n6933 | n11213 ;
  assign n25664 = n25663 ^ n19405 ^ 1'b0 ;
  assign n25665 = n9862 ^ n2491 ^ 1'b0 ;
  assign n25666 = n18279 ^ n17890 ^ 1'b0 ;
  assign n25667 = n22363 ^ n19322 ^ 1'b0 ;
  assign n25668 = n16328 | n24690 ;
  assign n25669 = ( n361 & n12553 ) | ( n361 & ~n23032 ) | ( n12553 & ~n23032 ) ;
  assign n25671 = n6826 ^ n3827 ^ 1'b0 ;
  assign n25670 = ~n5488 & n10972 ;
  assign n25672 = n25671 ^ n25670 ^ 1'b0 ;
  assign n25673 = ~n8719 & n17832 ;
  assign n25674 = n10435 ^ n6950 ^ 1'b0 ;
  assign n25675 = n1224 | n21744 ;
  assign n25676 = n25675 ^ n6743 ^ 1'b0 ;
  assign n25677 = n477 | n7125 ;
  assign n25678 = n25677 ^ n17152 ^ 1'b0 ;
  assign n25679 = n5761 ^ n2924 ^ 1'b0 ;
  assign n25680 = ( ~n3103 & n11957 ) | ( ~n3103 & n21503 ) | ( n11957 & n21503 ) ;
  assign n25681 = ~n2430 & n13519 ;
  assign n25685 = ~n11566 & n13850 ;
  assign n25686 = n25685 ^ n12342 ^ 1'b0 ;
  assign n25683 = n14551 ^ n9258 ^ 1'b0 ;
  assign n25682 = ( n10808 & n16842 ) | ( n10808 & n24443 ) | ( n16842 & n24443 ) ;
  assign n25684 = n25683 ^ n25682 ^ n6419 ;
  assign n25687 = n25686 ^ n25684 ^ n6741 ;
  assign n25688 = ( ~n2788 & n25681 ) | ( ~n2788 & n25687 ) | ( n25681 & n25687 ) ;
  assign n25689 = n9591 ^ n9475 ^ 1'b0 ;
  assign n25690 = n3166 & ~n22941 ;
  assign n25692 = n21310 ^ n8585 ^ 1'b0 ;
  assign n25693 = n3707 & n25692 ;
  assign n25691 = n14738 | n22717 ;
  assign n25694 = n25693 ^ n25691 ^ 1'b0 ;
  assign n25698 = ( n2785 & n14866 ) | ( n2785 & n16743 ) | ( n14866 & n16743 ) ;
  assign n25695 = n13630 ^ n850 ^ 1'b0 ;
  assign n25696 = n6410 & n25695 ;
  assign n25697 = n21835 & n25696 ;
  assign n25699 = n25698 ^ n25697 ^ 1'b0 ;
  assign n25700 = n10453 & ~n25699 ;
  assign n25701 = n21712 ^ n20951 ^ 1'b0 ;
  assign n25702 = n8941 | n25701 ;
  assign n25704 = ~n14802 & n22888 ;
  assign n25703 = ~n4041 & n5283 ;
  assign n25705 = n25704 ^ n25703 ^ 1'b0 ;
  assign n25706 = n8075 & ~n20667 ;
  assign n25707 = n25706 ^ n13019 ^ 1'b0 ;
  assign n25708 = n23413 ^ n285 ^ 1'b0 ;
  assign n25709 = n16890 & n25708 ;
  assign n25710 = ( n3953 & n8240 ) | ( n3953 & n25709 ) | ( n8240 & n25709 ) ;
  assign n25711 = n25424 ^ n8239 ^ 1'b0 ;
  assign n25712 = n25711 ^ n21250 ^ n3238 ;
  assign n25713 = n286 ^ n272 ^ 1'b0 ;
  assign n25714 = ( n10986 & n18626 ) | ( n10986 & ~n25713 ) | ( n18626 & ~n25713 ) ;
  assign n25715 = n11356 ^ n5571 ^ 1'b0 ;
  assign n25716 = ( x58 & ~n2198 ) | ( x58 & n7962 ) | ( ~n2198 & n7962 ) ;
  assign n25717 = n25716 ^ n16310 ^ 1'b0 ;
  assign n25718 = n1000 & ~n25717 ;
  assign n25719 = n9791 | n20017 ;
  assign n25720 = n25718 | n25719 ;
  assign n25721 = n17745 ^ n13192 ^ 1'b0 ;
  assign n25722 = n25721 ^ n9837 ^ 1'b0 ;
  assign n25723 = ~n13553 & n25722 ;
  assign n25724 = n3357 | n25466 ;
  assign n25725 = ( n1071 & n4026 ) | ( n1071 & ~n9184 ) | ( n4026 & ~n9184 ) ;
  assign n25726 = n723 & ~n23432 ;
  assign n25727 = n15177 ^ n5341 ^ 1'b0 ;
  assign n25728 = n7177 & ~n13359 ;
  assign n25729 = n25728 ^ n13203 ^ 1'b0 ;
  assign n25730 = n10413 & ~n24666 ;
  assign n25731 = n25730 ^ n4414 ^ 1'b0 ;
  assign n25732 = n5186 ^ n992 ^ 1'b0 ;
  assign n25733 = n16893 & n25732 ;
  assign n25734 = n9234 ^ n4607 ^ n2078 ;
  assign n25735 = ( n18053 & ~n19077 ) | ( n18053 & n19547 ) | ( ~n19077 & n19547 ) ;
  assign n25736 = ~n458 & n11124 ;
  assign n25737 = n13281 ^ n4094 ^ 1'b0 ;
  assign n25738 = n10164 ^ n5186 ^ 1'b0 ;
  assign n25739 = n25737 & ~n25738 ;
  assign n25740 = n25739 ^ n18413 ^ 1'b0 ;
  assign n25741 = n25736 & ~n25740 ;
  assign n25742 = n25735 | n25741 ;
  assign n25743 = n276 & ~n1209 ;
  assign n25744 = n1613 & n24456 ;
  assign n25745 = ~n15300 & n25744 ;
  assign n25746 = n8350 | n20317 ;
  assign n25747 = n25746 ^ n18233 ^ 1'b0 ;
  assign n25748 = n10839 ^ n225 ^ 1'b0 ;
  assign n25749 = n25747 & n25748 ;
  assign n25750 = n13077 & n23541 ;
  assign n25755 = n1382 | n1984 ;
  assign n25754 = n1389 & ~n9327 ;
  assign n25756 = n25755 ^ n25754 ^ 1'b0 ;
  assign n25751 = n10483 ^ n2265 ^ 1'b0 ;
  assign n25752 = n12143 | n25751 ;
  assign n25753 = ( n8254 & n13258 ) | ( n8254 & ~n25752 ) | ( n13258 & ~n25752 ) ;
  assign n25757 = n25756 ^ n25753 ^ 1'b0 ;
  assign n25758 = n5044 & ~n11911 ;
  assign n25759 = ~n10003 & n25758 ;
  assign n25760 = n7280 | n25759 ;
  assign n25761 = n24489 | n25760 ;
  assign n25762 = ( ~n5499 & n7377 ) | ( ~n5499 & n25761 ) | ( n7377 & n25761 ) ;
  assign n25763 = ( n7794 & n11767 ) | ( n7794 & ~n12242 ) | ( n11767 & ~n12242 ) ;
  assign n25764 = n2044 & ~n25763 ;
  assign n25765 = n1171 & n6686 ;
  assign n25766 = n25765 ^ n25087 ^ 1'b0 ;
  assign n25767 = n25766 ^ n18269 ^ n16890 ;
  assign n25768 = n7470 & ~n22910 ;
  assign n25769 = n15064 ^ n1720 ^ 1'b0 ;
  assign n25770 = n7908 & n17643 ;
  assign n25771 = ~n763 & n24043 ;
  assign n25772 = n25771 ^ n316 ^ 1'b0 ;
  assign n25773 = n21433 ^ n6486 ^ 1'b0 ;
  assign n25774 = n25773 ^ n6214 ^ n3886 ;
  assign n25775 = ( n2141 & n5798 ) | ( n2141 & ~n23623 ) | ( n5798 & ~n23623 ) ;
  assign n25776 = n9591 & ~n10065 ;
  assign n25777 = ( ~n3572 & n4027 ) | ( ~n3572 & n25776 ) | ( n4027 & n25776 ) ;
  assign n25778 = n21417 ^ n8011 ^ 1'b0 ;
  assign n25779 = n8332 | n25778 ;
  assign n25780 = n22312 ^ n7071 ^ 1'b0 ;
  assign n25781 = ~n10607 & n25780 ;
  assign n25782 = ~n5392 & n25781 ;
  assign n25783 = n13246 & n22625 ;
  assign n25784 = ~n8523 & n25272 ;
  assign n25785 = n8985 & n25784 ;
  assign n25786 = n17473 ^ n3016 ^ n2835 ;
  assign n25787 = n25786 ^ n13480 ^ n2167 ;
  assign n25788 = n9422 ^ n7709 ^ 1'b0 ;
  assign n25789 = n7660 & ~n25788 ;
  assign n25790 = ~n872 & n9788 ;
  assign n25791 = n25790 ^ n25361 ^ n8432 ;
  assign n25792 = n2323 | n6794 ;
  assign n25793 = ( n3482 & ~n3822 ) | ( n3482 & n25792 ) | ( ~n3822 & n25792 ) ;
  assign n25794 = n14731 ^ n12799 ^ 1'b0 ;
  assign n25795 = n9752 & ~n14119 ;
  assign n25796 = ( n701 & ~n14326 ) | ( n701 & n20515 ) | ( ~n14326 & n20515 ) ;
  assign n25797 = n8004 | n25796 ;
  assign n25799 = n1708 | n5106 ;
  assign n25800 = n25799 ^ n3467 ^ 1'b0 ;
  assign n25798 = n3831 | n7839 ;
  assign n25801 = n25800 ^ n25798 ^ 1'b0 ;
  assign n25802 = n16412 ^ n10890 ^ 1'b0 ;
  assign n25803 = n12209 ^ n7817 ^ n599 ;
  assign n25804 = n11863 & ~n14511 ;
  assign n25805 = n25804 ^ n4530 ^ 1'b0 ;
  assign n25806 = x107 & n1652 ;
  assign n25807 = n7045 & n25806 ;
  assign n25808 = n21298 ^ n6560 ^ 1'b0 ;
  assign n25809 = ~n19395 & n25808 ;
  assign n25810 = n7438 ^ n3299 ^ n1502 ;
  assign n25811 = ( n4433 & n7537 ) | ( n4433 & n8528 ) | ( n7537 & n8528 ) ;
  assign n25812 = n17181 ^ n2156 ^ 1'b0 ;
  assign n25813 = n7381 | n25812 ;
  assign n25814 = ( n3701 & n7068 ) | ( n3701 & ~n25813 ) | ( n7068 & ~n25813 ) ;
  assign n25815 = n25814 ^ n8669 ^ 1'b0 ;
  assign n25816 = n2445 & ~n17842 ;
  assign n25817 = n19162 ^ n8049 ^ 1'b0 ;
  assign n25818 = n23947 ^ n3050 ^ 1'b0 ;
  assign n25819 = n1893 | n25818 ;
  assign n25820 = n12461 ^ n5135 ^ n686 ;
  assign n25821 = ~n12717 & n25820 ;
  assign n25822 = ( n2579 & ~n2889 ) | ( n2579 & n10264 ) | ( ~n2889 & n10264 ) ;
  assign n25823 = n885 | n25822 ;
  assign n25824 = n25821 & ~n25823 ;
  assign n25825 = n23105 ^ n3530 ^ 1'b0 ;
  assign n25826 = n25824 | n25825 ;
  assign n25827 = n19888 ^ n2460 ^ 1'b0 ;
  assign n25828 = n2192 | n25827 ;
  assign n25829 = ( n5513 & n6660 ) | ( n5513 & n11164 ) | ( n6660 & n11164 ) ;
  assign n25830 = ~n25828 & n25829 ;
  assign n25831 = n18856 ^ n11632 ^ n2520 ;
  assign n25832 = ( ~n1466 & n2457 ) | ( ~n1466 & n5925 ) | ( n2457 & n5925 ) ;
  assign n25833 = n25832 ^ n16121 ^ 1'b0 ;
  assign n25834 = n23933 ^ n23223 ^ n5696 ;
  assign n25835 = n786 | n20839 ;
  assign n25836 = n16948 & n25835 ;
  assign n25837 = n13597 ^ n6345 ^ 1'b0 ;
  assign n25838 = n25836 | n25837 ;
  assign n25839 = n25838 ^ n24783 ^ n14002 ;
  assign n25840 = n10204 | n16294 ;
  assign n25841 = n21611 ^ n16985 ^ 1'b0 ;
  assign n25842 = ~n411 & n17288 ;
  assign n25843 = n25115 & n25842 ;
  assign n25844 = n5530 | n8375 ;
  assign n25845 = n23964 | n25844 ;
  assign n25846 = ~n4753 & n25845 ;
  assign n25847 = n3478 & n12401 ;
  assign n25849 = n4739 | n15492 ;
  assign n25848 = n14111 ^ n10066 ^ 1'b0 ;
  assign n25850 = n25849 ^ n25848 ^ 1'b0 ;
  assign n25851 = n3828 & n6214 ;
  assign n25852 = ~n1947 & n25851 ;
  assign n25853 = x100 & n740 ;
  assign n25854 = ( ~n1532 & n15299 ) | ( ~n1532 & n19952 ) | ( n15299 & n19952 ) ;
  assign n25855 = ( ~n866 & n25853 ) | ( ~n866 & n25854 ) | ( n25853 & n25854 ) ;
  assign n25856 = n25855 ^ n6966 ^ n5935 ;
  assign n25857 = n15989 ^ n11123 ^ n2869 ;
  assign n25858 = ~n858 & n24050 ;
  assign n25859 = ~n6796 & n25858 ;
  assign n25860 = n24942 & ~n25859 ;
  assign n25861 = n3503 ^ n535 ^ 1'b0 ;
  assign n25862 = n1373 & n13966 ;
  assign n25863 = n25862 ^ n2653 ^ 1'b0 ;
  assign n25864 = ~n25861 & n25863 ;
  assign n25865 = ~n231 & n25864 ;
  assign n25866 = n9015 ^ n7152 ^ 1'b0 ;
  assign n25867 = n13302 & n25866 ;
  assign n25868 = ( n8350 & n10520 ) | ( n8350 & ~n25867 ) | ( n10520 & ~n25867 ) ;
  assign n25869 = n3597 & ~n4906 ;
  assign n25870 = n4213 & n25869 ;
  assign n25871 = n16769 & n17282 ;
  assign n25872 = n25870 & ~n25871 ;
  assign n25873 = ( n1800 & n12647 ) | ( n1800 & n18269 ) | ( n12647 & n18269 ) ;
  assign n25874 = n25873 ^ n21357 ^ n441 ;
  assign n25875 = n2312 & ~n3463 ;
  assign n25876 = n25875 ^ n5370 ^ 1'b0 ;
  assign n25877 = n24121 ^ n3261 ^ 1'b0 ;
  assign n25878 = n6148 | n25877 ;
  assign n25879 = n20883 | n25878 ;
  assign n25880 = n25879 ^ n3739 ^ 1'b0 ;
  assign n25881 = n2167 | n25880 ;
  assign n25882 = n9927 | n15217 ;
  assign n25883 = n14801 & ~n25882 ;
  assign n25884 = n8838 & ~n25883 ;
  assign n25885 = ~n8626 & n25884 ;
  assign n25886 = n11836 ^ n5185 ^ 1'b0 ;
  assign n25887 = ~n19052 & n25886 ;
  assign n25888 = n5257 & ~n13956 ;
  assign n25889 = n18623 ^ n4610 ^ 1'b0 ;
  assign n25890 = n4137 & n25889 ;
  assign n25891 = ~n25888 & n25890 ;
  assign n25892 = n12208 ^ n7144 ^ 1'b0 ;
  assign n25893 = n4044 & ~n25892 ;
  assign n25894 = n11531 | n25893 ;
  assign n25895 = n131 & n11601 ;
  assign n25896 = n25895 ^ n20982 ^ n5223 ;
  assign n25897 = n19394 ^ n11872 ^ 1'b0 ;
  assign n25898 = ( ~n5113 & n17046 ) | ( ~n5113 & n20838 ) | ( n17046 & n20838 ) ;
  assign n25899 = ~n11813 & n25898 ;
  assign n25900 = ( n13138 & ~n16195 ) | ( n13138 & n25899 ) | ( ~n16195 & n25899 ) ;
  assign n25901 = ~n4190 & n9439 ;
  assign n25902 = n25901 ^ n20237 ^ 1'b0 ;
  assign n25903 = n25902 ^ n18488 ^ 1'b0 ;
  assign n25904 = n17143 ^ n8086 ^ 1'b0 ;
  assign n25905 = ~n2279 & n9807 ;
  assign n25906 = n25905 ^ n8231 ^ 1'b0 ;
  assign n25907 = n18960 ^ n3382 ^ 1'b0 ;
  assign n25908 = n6254 & n25907 ;
  assign n25909 = n1633 | n18753 ;
  assign n25910 = n16158 | n25909 ;
  assign n25911 = ( n3949 & ~n12765 ) | ( n3949 & n25910 ) | ( ~n12765 & n25910 ) ;
  assign n25912 = ( ~n8519 & n17408 ) | ( ~n8519 & n25911 ) | ( n17408 & n25911 ) ;
  assign n25913 = ~n4887 & n12666 ;
  assign n25918 = n3044 & n8338 ;
  assign n25919 = n25918 ^ n6801 ^ 1'b0 ;
  assign n25914 = ( n443 & n1476 ) | ( n443 & ~n2471 ) | ( n1476 & ~n2471 ) ;
  assign n25915 = n1051 & ~n25914 ;
  assign n25916 = ( n3667 & n11232 ) | ( n3667 & ~n25915 ) | ( n11232 & ~n25915 ) ;
  assign n25917 = n25916 ^ n12149 ^ n2990 ;
  assign n25920 = n25919 ^ n25917 ^ n1123 ;
  assign n25921 = n4273 ^ n1555 ^ 1'b0 ;
  assign n25922 = n25921 ^ n3553 ^ n3279 ;
  assign n25923 = n178 & n9648 ;
  assign n25924 = n10840 & ~n16828 ;
  assign n25925 = n25924 ^ n1617 ^ 1'b0 ;
  assign n25926 = n25923 & n25925 ;
  assign n25927 = n25926 ^ n2253 ^ 1'b0 ;
  assign n25928 = n4896 & n25829 ;
  assign n25929 = ~n7350 & n14548 ;
  assign n25930 = ~n10158 & n25929 ;
  assign n25931 = ~n10608 & n17398 ;
  assign n25932 = ~n1201 & n7154 ;
  assign n25933 = ~n1221 & n1535 ;
  assign n25934 = n24108 ^ n3312 ^ 1'b0 ;
  assign n25935 = n17727 ^ n10464 ^ 1'b0 ;
  assign n25936 = n2598 & ~n25935 ;
  assign n25937 = n16492 ^ n11595 ^ n2709 ;
  assign n25938 = n471 & n10523 ;
  assign n25939 = n2264 & n25938 ;
  assign n25940 = ( n25936 & ~n25937 ) | ( n25936 & n25939 ) | ( ~n25937 & n25939 ) ;
  assign n25941 = n5735 & n13118 ;
  assign n25942 = n25941 ^ n25466 ^ 1'b0 ;
  assign n25943 = n4739 | n6768 ;
  assign n25944 = n16480 | n25943 ;
  assign n25945 = n1718 ^ n236 ^ 1'b0 ;
  assign n25946 = ~n19834 & n25945 ;
  assign n25959 = n10809 ^ n8945 ^ n3771 ;
  assign n25952 = x37 & n225 ;
  assign n25953 = ~x37 & n25952 ;
  assign n25954 = n1022 & n25953 ;
  assign n25955 = n1133 | n25954 ;
  assign n25956 = n25954 & ~n25955 ;
  assign n25949 = n820 | n946 ;
  assign n25950 = n946 & ~n25949 ;
  assign n25951 = n5407 | n25950 ;
  assign n25947 = ~n6457 & n6752 ;
  assign n25948 = n6457 & n25947 ;
  assign n25957 = n25956 ^ n25951 ^ n25948 ;
  assign n25958 = ( n4682 & n10734 ) | ( n4682 & n25957 ) | ( n10734 & n25957 ) ;
  assign n25960 = n25959 ^ n25958 ^ 1'b0 ;
  assign n25961 = n16070 | n22930 ;
  assign n25962 = n25961 ^ n13129 ^ n974 ;
  assign n25963 = n25962 ^ n24161 ^ n1940 ;
  assign n25964 = n8067 ^ n5987 ^ 1'b0 ;
  assign n25965 = n4210 & n5867 ;
  assign n25966 = n7310 & n25965 ;
  assign n25967 = n10452 ^ n1523 ^ 1'b0 ;
  assign n25968 = n13278 & n25967 ;
  assign n25969 = n6197 | n25968 ;
  assign n25970 = ~n2746 & n12773 ;
  assign n25971 = n7686 | n16955 ;
  assign n25972 = n25970 | n25971 ;
  assign n25973 = n22299 ^ n19702 ^ n5573 ;
  assign n25975 = n5435 ^ n1645 ^ 1'b0 ;
  assign n25974 = ~n12483 & n14119 ;
  assign n25976 = n25975 ^ n25974 ^ 1'b0 ;
  assign n25977 = n4819 | n20454 ;
  assign n25978 = n25976 & ~n25977 ;
  assign n25979 = n4699 | n18072 ;
  assign n25980 = n25979 ^ n19969 ^ n6631 ;
  assign n25981 = n25980 ^ n15495 ^ 1'b0 ;
  assign n25982 = ( n578 & ~n4318 ) | ( n578 & n25696 ) | ( ~n4318 & n25696 ) ;
  assign n25983 = n16531 ^ n5066 ^ n2934 ;
  assign n25984 = ( n998 & n4286 ) | ( n998 & n25983 ) | ( n4286 & n25983 ) ;
  assign n25985 = n7366 | n25984 ;
  assign n25986 = n25985 ^ n19547 ^ n17523 ;
  assign n25988 = n9168 | n12419 ;
  assign n25989 = n4293 | n25988 ;
  assign n25987 = n3538 | n3749 ;
  assign n25990 = n25989 ^ n25987 ^ 1'b0 ;
  assign n25991 = ~n5078 & n11365 ;
  assign n25992 = n9131 & n10255 ;
  assign n25993 = n13242 & n25992 ;
  assign n25994 = n2599 & ~n8111 ;
  assign n25995 = n25994 ^ n1902 ^ 1'b0 ;
  assign n25996 = n25995 ^ n12640 ^ 1'b0 ;
  assign n25997 = ~n6736 & n22424 ;
  assign n25998 = n17412 ^ n6874 ^ 1'b0 ;
  assign n25999 = ~n146 & n16698 ;
  assign n26000 = ~n25998 & n25999 ;
  assign n26001 = ( n5543 & n7105 ) | ( n5543 & n20320 ) | ( n7105 & n20320 ) ;
  assign n26002 = n26001 ^ n2767 ^ 1'b0 ;
  assign n26003 = ( n9746 & n22276 ) | ( n9746 & ~n26002 ) | ( n22276 & ~n26002 ) ;
  assign n26004 = n12644 ^ n8865 ^ 1'b0 ;
  assign n26005 = n19511 | n26004 ;
  assign n26006 = n26005 ^ n25483 ^ n14647 ;
  assign n26010 = ( n5059 & n8987 ) | ( n5059 & n9516 ) | ( n8987 & n9516 ) ;
  assign n26008 = ( n5011 & n8810 ) | ( n5011 & ~n19238 ) | ( n8810 & ~n19238 ) ;
  assign n26007 = n1415 & ~n20579 ;
  assign n26009 = n26008 ^ n26007 ^ 1'b0 ;
  assign n26011 = n26010 ^ n26009 ^ n7312 ;
  assign n26012 = n1784 ^ n1527 ^ 1'b0 ;
  assign n26013 = n22016 ^ n13146 ^ 1'b0 ;
  assign n26014 = ~n26012 & n26013 ;
  assign n26015 = n3883 & n17573 ;
  assign n26016 = ~n210 & n26015 ;
  assign n26017 = n1143 | n2986 ;
  assign n26018 = n26017 ^ n25910 ^ 1'b0 ;
  assign n26019 = ~n6925 & n16693 ;
  assign n26020 = ~n25820 & n26019 ;
  assign n26021 = n5582 | n6876 ;
  assign n26022 = n20233 & ~n26021 ;
  assign n26023 = n11532 ^ n6668 ^ 1'b0 ;
  assign n26024 = n26023 ^ n12687 ^ 1'b0 ;
  assign n26027 = n712 & ~n3345 ;
  assign n26028 = ~n7368 & n26027 ;
  assign n26025 = n4308 & ~n4661 ;
  assign n26026 = ~n22401 & n26025 ;
  assign n26029 = n26028 ^ n26026 ^ n279 ;
  assign n26031 = n3077 ^ n2767 ^ n2500 ;
  assign n26030 = n23608 ^ n3900 ^ 1'b0 ;
  assign n26032 = n26031 ^ n26030 ^ n3177 ;
  assign n26033 = ( n2304 & ~n4495 ) | ( n2304 & n26032 ) | ( ~n4495 & n26032 ) ;
  assign n26034 = n7101 | n8367 ;
  assign n26035 = n26034 ^ n11757 ^ 1'b0 ;
  assign n26036 = n17698 & n26035 ;
  assign n26037 = n19300 ^ n10636 ^ n5430 ;
  assign n26038 = n3949 | n26037 ;
  assign n26039 = n10106 ^ n4940 ^ n3688 ;
  assign n26040 = ~n7813 & n17546 ;
  assign n26041 = n1797 ^ n775 ^ 1'b0 ;
  assign n26042 = n9013 & n26041 ;
  assign n26043 = ~n10544 & n26042 ;
  assign n26044 = n3484 ^ n1459 ^ 1'b0 ;
  assign n26045 = ( n1460 & n3347 ) | ( n1460 & n6239 ) | ( n3347 & n6239 ) ;
  assign n26046 = n10002 & ~n12835 ;
  assign n26047 = n18687 | n26046 ;
  assign n26049 = n10398 ^ n3910 ^ 1'b0 ;
  assign n26048 = n24803 ^ n16179 ^ n12357 ;
  assign n26050 = n26049 ^ n26048 ^ 1'b0 ;
  assign n26051 = n15111 & n18343 ;
  assign n26052 = n26051 ^ n1516 ^ 1'b0 ;
  assign n26053 = n8730 | n26052 ;
  assign n26054 = n26050 & ~n26053 ;
  assign n26055 = n11496 & n24481 ;
  assign n26056 = n3847 & n4969 ;
  assign n26057 = n26056 ^ n9367 ^ 1'b0 ;
  assign n26058 = n1166 | n16918 ;
  assign n26059 = ( n8294 & ~n10444 ) | ( n8294 & n17017 ) | ( ~n10444 & n17017 ) ;
  assign n26060 = n26059 ^ n3669 ^ 1'b0 ;
  assign n26061 = n26058 & ~n26060 ;
  assign n26062 = n18338 ^ n11612 ^ 1'b0 ;
  assign n26063 = n15384 & n26062 ;
  assign n26064 = ~n771 & n9790 ;
  assign n26065 = n11974 & n26064 ;
  assign n26066 = n787 | n8487 ;
  assign n26067 = n15665 | n26066 ;
  assign n26068 = n8507 & n23763 ;
  assign n26069 = n26067 & n26068 ;
  assign n26070 = ( n11841 & n12280 ) | ( n11841 & ~n18246 ) | ( n12280 & ~n18246 ) ;
  assign n26076 = n8082 ^ n4161 ^ 1'b0 ;
  assign n26077 = n3933 & ~n26076 ;
  assign n26074 = n7169 & ~n10569 ;
  assign n26075 = n17311 & n26074 ;
  assign n26078 = n26077 ^ n26075 ^ n13008 ;
  assign n26071 = n5781 & n12718 ;
  assign n26072 = n4529 & n26071 ;
  assign n26073 = ( n3065 & ~n16520 ) | ( n3065 & n26072 ) | ( ~n16520 & n26072 ) ;
  assign n26079 = n26078 ^ n26073 ^ n2079 ;
  assign n26080 = n11750 ^ n913 ^ 1'b0 ;
  assign n26081 = n26080 ^ n8539 ^ 1'b0 ;
  assign n26082 = n162 & ~n9372 ;
  assign n26083 = n26082 ^ n11204 ^ 1'b0 ;
  assign n26084 = n6427 & ~n26083 ;
  assign n26085 = n19366 & n26084 ;
  assign n26086 = n5180 ^ n4984 ^ 1'b0 ;
  assign n26087 = n408 & n26086 ;
  assign n26088 = n9697 & ~n14276 ;
  assign n26089 = ~n26087 & n26088 ;
  assign n26090 = n7216 | n9618 ;
  assign n26091 = n12186 ^ n6989 ^ 1'b0 ;
  assign n26092 = ~n6903 & n26091 ;
  assign n26093 = n15788 ^ n15551 ^ 1'b0 ;
  assign n26094 = n26093 ^ n22775 ^ n7027 ;
  assign n26095 = n1515 | n8213 ;
  assign n26096 = n3139 & ~n26095 ;
  assign n26097 = n19811 & n25989 ;
  assign n26098 = n26097 ^ n5792 ^ 1'b0 ;
  assign n26099 = ~n26096 & n26098 ;
  assign n26100 = ( n10139 & n12488 ) | ( n10139 & n23120 ) | ( n12488 & n23120 ) ;
  assign n26101 = n9772 | n26100 ;
  assign n26102 = n26101 ^ n14647 ^ n11433 ;
  assign n26103 = n1928 | n7669 ;
  assign n26104 = n26103 ^ n6372 ^ 1'b0 ;
  assign n26105 = n7396 | n26104 ;
  assign n26106 = n26105 ^ n11944 ^ 1'b0 ;
  assign n26107 = ~n25166 & n25944 ;
  assign n26108 = ~n7373 & n26107 ;
  assign n26109 = ~n510 & n11132 ;
  assign n26110 = ~n3888 & n26109 ;
  assign n26111 = n22191 & n26110 ;
  assign n26112 = n8432 & ~n17339 ;
  assign n26113 = n26112 ^ n4748 ^ 1'b0 ;
  assign n26114 = n26113 ^ n24208 ^ n23719 ;
  assign n26115 = ~n14501 & n19467 ;
  assign n26116 = n26115 ^ n9137 ^ 1'b0 ;
  assign n26117 = n2699 | n10065 ;
  assign n26118 = n26117 ^ n15395 ^ 1'b0 ;
  assign n26119 = ( ~n932 & n26116 ) | ( ~n932 & n26118 ) | ( n26116 & n26118 ) ;
  assign n26120 = n1188 | n19466 ;
  assign n26121 = ( ~n2868 & n12542 ) | ( ~n2868 & n26120 ) | ( n12542 & n26120 ) ;
  assign n26122 = n20362 ^ n14180 ^ n5492 ;
  assign n26123 = ~n1015 & n20907 ;
  assign n26124 = n14392 ^ n3886 ^ 1'b0 ;
  assign n26125 = n2682 & n11347 ;
  assign n26126 = ~n16207 & n26125 ;
  assign n26127 = ~n10789 & n26126 ;
  assign n26128 = n15499 ^ n6250 ^ 1'b0 ;
  assign n26129 = n26128 ^ n13586 ^ n383 ;
  assign n26130 = n15058 ^ n12756 ^ n7377 ;
  assign n26131 = n26129 & n26130 ;
  assign n26132 = n663 & ~n26131 ;
  assign n26133 = n20052 ^ n19558 ^ 1'b0 ;
  assign n26134 = n3751 & ~n11673 ;
  assign n26135 = n1168 | n26134 ;
  assign n26136 = ~n5208 & n6214 ;
  assign n26137 = n10646 ^ n2246 ^ 1'b0 ;
  assign n26138 = ~n13866 & n22919 ;
  assign n26139 = ~n25362 & n26138 ;
  assign n26140 = n6668 & ~n26139 ;
  assign n26141 = n19873 ^ n13409 ^ 1'b0 ;
  assign n26142 = n26140 & n26141 ;
  assign n26143 = ~n2824 & n12068 ;
  assign n26144 = n20618 & n26143 ;
  assign n26145 = ~n13478 & n26144 ;
  assign n26146 = n925 | n10789 ;
  assign n26147 = ( n6140 & n15226 ) | ( n6140 & ~n26146 ) | ( n15226 & ~n26146 ) ;
  assign n26148 = n10266 & ~n10857 ;
  assign n26149 = n26148 ^ n13264 ^ 1'b0 ;
  assign n26150 = n6191 ^ n2377 ^ 1'b0 ;
  assign n26151 = n22048 | n26150 ;
  assign n26152 = n22756 ^ n1633 ^ 1'b0 ;
  assign n26153 = n7256 | n26152 ;
  assign n26154 = n15355 ^ n11881 ^ 1'b0 ;
  assign n26155 = n17349 & n26154 ;
  assign n26156 = ( n1326 & n3730 ) | ( n1326 & ~n23352 ) | ( n3730 & ~n23352 ) ;
  assign n26157 = n4864 & ~n26156 ;
  assign n26158 = n15839 ^ n5247 ^ 1'b0 ;
  assign n26159 = n9118 & ~n26158 ;
  assign n26160 = n13823 ^ n10747 ^ 1'b0 ;
  assign n26161 = ( ~n12414 & n26159 ) | ( ~n12414 & n26160 ) | ( n26159 & n26160 ) ;
  assign n26164 = n1935 & ~n17171 ;
  assign n26163 = n5088 | n5421 ;
  assign n26162 = n4764 & ~n18296 ;
  assign n26165 = n26164 ^ n26163 ^ n26162 ;
  assign n26166 = ~n5621 & n7833 ;
  assign n26167 = n1327 & n26166 ;
  assign n26168 = n26167 ^ n17638 ^ 1'b0 ;
  assign n26169 = n4207 & ~n10649 ;
  assign n26170 = n26169 ^ n20545 ^ 1'b0 ;
  assign n26171 = n26170 ^ n736 ^ 1'b0 ;
  assign n26172 = n17672 & n26171 ;
  assign n26173 = n26168 & n26172 ;
  assign n26174 = n12154 & n16378 ;
  assign n26175 = n26174 ^ n16767 ^ 1'b0 ;
  assign n26176 = ~n24175 & n26175 ;
  assign n26177 = n19668 ^ n3724 ^ 1'b0 ;
  assign n26178 = n26177 ^ n21043 ^ 1'b0 ;
  assign n26179 = ~n980 & n26178 ;
  assign n26180 = n3403 & n9618 ;
  assign n26181 = ~n6872 & n26180 ;
  assign n26182 = n12629 ^ n4075 ^ n3195 ;
  assign n26183 = n26182 ^ n458 ^ x4 ;
  assign n26184 = n5335 & ~n23910 ;
  assign n26185 = n26184 ^ n8482 ^ 1'b0 ;
  assign n26186 = n26185 ^ n23976 ^ n10268 ;
  assign n26187 = ( n5814 & ~n7338 ) | ( n5814 & n13966 ) | ( ~n7338 & n13966 ) ;
  assign n26188 = n4975 & ~n14916 ;
  assign n26189 = n26188 ^ n16565 ^ 1'b0 ;
  assign n26190 = n26187 & n26189 ;
  assign n26191 = n26190 ^ n3284 ^ 1'b0 ;
  assign n26192 = n10515 | n26191 ;
  assign n26193 = n2650 & ~n9436 ;
  assign n26194 = n26192 & n26193 ;
  assign n26195 = ( n18207 & ~n23842 ) | ( n18207 & n26194 ) | ( ~n23842 & n26194 ) ;
  assign n26196 = ( x86 & n18945 ) | ( x86 & n24945 ) | ( n18945 & n24945 ) ;
  assign n26197 = n24316 ^ n3905 ^ 1'b0 ;
  assign n26198 = n15574 & ~n26197 ;
  assign n26199 = n4147 ^ n3041 ^ n1784 ;
  assign n26200 = n4061 & ~n8716 ;
  assign n26201 = n26199 & n26200 ;
  assign n26202 = n8557 & ~n18830 ;
  assign n26203 = ( n12759 & ~n20820 ) | ( n12759 & n26202 ) | ( ~n20820 & n26202 ) ;
  assign n26204 = n15283 ^ n5247 ^ 1'b0 ;
  assign n26205 = n3136 & ~n26204 ;
  assign n26206 = n26205 ^ n17270 ^ n4917 ;
  assign n26207 = n7152 & ~n9821 ;
  assign n26208 = n26207 ^ n13545 ^ 1'b0 ;
  assign n26209 = n26208 ^ n16090 ^ n2300 ;
  assign n26210 = n5104 | n13160 ;
  assign n26211 = n25682 & ~n26210 ;
  assign n26212 = n18964 ^ n14028 ^ 1'b0 ;
  assign n26213 = n17688 | n26212 ;
  assign n26214 = n26213 ^ n10440 ^ 1'b0 ;
  assign n26215 = ~n14678 & n17242 ;
  assign n26216 = ~n17563 & n26215 ;
  assign n26217 = n3766 & n6946 ;
  assign n26218 = n26217 ^ n2085 ^ 1'b0 ;
  assign n26219 = n26218 ^ n1955 ^ 1'b0 ;
  assign n26220 = n14902 ^ n11106 ^ 1'b0 ;
  assign n26221 = ( n3549 & n9354 ) | ( n3549 & n18249 ) | ( n9354 & n18249 ) ;
  assign n26222 = ( n24223 & n26220 ) | ( n24223 & n26221 ) | ( n26220 & n26221 ) ;
  assign n26224 = n1327 & ~n23633 ;
  assign n26223 = n7045 | n12884 ;
  assign n26225 = n26224 ^ n26223 ^ 1'b0 ;
  assign n26226 = n13131 ^ n11906 ^ 1'b0 ;
  assign n26227 = ~n15878 & n26226 ;
  assign n26228 = n16728 ^ n15805 ^ 1'b0 ;
  assign n26229 = n18572 ^ n14012 ^ 1'b0 ;
  assign n26230 = n26229 ^ n15193 ^ n6055 ;
  assign n26231 = n22554 ^ n20373 ^ 1'b0 ;
  assign n26239 = n5737 & n6022 ;
  assign n26232 = n2831 ^ n210 ^ 1'b0 ;
  assign n26233 = n7936 & n26232 ;
  assign n26234 = n2826 | n18829 ;
  assign n26235 = n15316 & n26234 ;
  assign n26236 = n26235 ^ n13772 ^ 1'b0 ;
  assign n26237 = ( ~n8063 & n26233 ) | ( ~n8063 & n26236 ) | ( n26233 & n26236 ) ;
  assign n26238 = n2880 & n26237 ;
  assign n26240 = n26239 ^ n26238 ^ 1'b0 ;
  assign n26241 = ( n5171 & n5551 ) | ( n5171 & n6247 ) | ( n5551 & n6247 ) ;
  assign n26242 = n11313 & n26241 ;
  assign n26243 = n26240 & n26242 ;
  assign n26244 = n26056 ^ n24844 ^ 1'b0 ;
  assign n26245 = n13262 | n26244 ;
  assign n26246 = n21873 & ~n26245 ;
  assign n26247 = n18107 ^ n13075 ^ 1'b0 ;
  assign n26248 = n2724 | n26247 ;
  assign n26249 = n11261 | n14221 ;
  assign n26250 = n15594 | n26249 ;
  assign n26251 = n26250 ^ n6832 ^ 1'b0 ;
  assign n26252 = n24872 ^ n4867 ^ n982 ;
  assign n26253 = n584 & n25619 ;
  assign n26254 = n15299 ^ n12399 ^ n9480 ;
  assign n26255 = n4345 ^ n1307 ^ 1'b0 ;
  assign n26256 = n13831 ^ n3471 ^ 1'b0 ;
  assign n26257 = n26233 & n26256 ;
  assign n26258 = ( n10330 & n10755 ) | ( n10330 & ~n21067 ) | ( n10755 & ~n21067 ) ;
  assign n26259 = n9482 & ~n26258 ;
  assign n26260 = n3731 | n16842 ;
  assign n26261 = n1473 ^ n363 ^ 1'b0 ;
  assign n26263 = ~n3943 & n23342 ;
  assign n26262 = n9970 ^ n7130 ^ 1'b0 ;
  assign n26264 = n26263 ^ n26262 ^ n9683 ;
  assign n26265 = n6412 ^ n1244 ^ n561 ;
  assign n26266 = n9435 & n26265 ;
  assign n26267 = n26266 ^ n6028 ^ 1'b0 ;
  assign n26268 = n14101 | n26267 ;
  assign n26269 = ~n1532 & n5402 ;
  assign n26270 = n4364 & n26269 ;
  assign n26271 = n20866 ^ n1651 ^ n620 ;
  assign n26272 = ( ~n6220 & n26270 ) | ( ~n6220 & n26271 ) | ( n26270 & n26271 ) ;
  assign n26273 = ( n12579 & n19465 ) | ( n12579 & n22068 ) | ( n19465 & n22068 ) ;
  assign n26274 = ~n648 & n2441 ;
  assign n26275 = n26273 & n26274 ;
  assign n26276 = ( ~n8776 & n10687 ) | ( ~n8776 & n11971 ) | ( n10687 & n11971 ) ;
  assign n26277 = n17161 | n26276 ;
  assign n26278 = ( n7369 & n8957 ) | ( n7369 & ~n13723 ) | ( n8957 & ~n13723 ) ;
  assign n26279 = n26278 ^ n5131 ^ 1'b0 ;
  assign n26280 = n17128 ^ n5734 ^ n1545 ;
  assign n26281 = n4137 & n8639 ;
  assign n26282 = n26280 | n26281 ;
  assign n26283 = n26282 ^ n2816 ^ 1'b0 ;
  assign n26284 = n26283 ^ n20201 ^ 1'b0 ;
  assign n26285 = n10458 & ~n26284 ;
  assign n26286 = ( n617 & ~n11282 ) | ( n617 & n14505 ) | ( ~n11282 & n14505 ) ;
  assign n26287 = n26286 ^ n22552 ^ 1'b0 ;
  assign n26288 = n19067 | n19509 ;
  assign n26289 = n8677 & n14741 ;
  assign n26290 = n26289 ^ n19031 ^ 1'b0 ;
  assign n26291 = ~n9357 & n10038 ;
  assign n26292 = n26291 ^ n21839 ^ n21238 ;
  assign n26293 = ( n782 & n10011 ) | ( n782 & ~n10623 ) | ( n10011 & ~n10623 ) ;
  assign n26294 = ~n22206 & n23545 ;
  assign n26295 = n26293 & n26294 ;
  assign n26296 = ~n20836 & n23628 ;
  assign n26297 = ~n12514 & n26296 ;
  assign n26298 = ~n661 & n8321 ;
  assign n26299 = ~n17656 & n26298 ;
  assign n26300 = n9130 | n26299 ;
  assign n26301 = n26300 ^ n3613 ^ 1'b0 ;
  assign n26302 = n3128 | n7888 ;
  assign n26303 = n26302 ^ n12962 ^ 1'b0 ;
  assign n26304 = n22875 ^ n16296 ^ n2746 ;
  assign n26305 = n24567 ^ n2909 ^ 1'b0 ;
  assign n26306 = n26305 ^ n25265 ^ n5348 ;
  assign n26307 = n15519 ^ n6475 ^ 1'b0 ;
  assign n26308 = n7032 & ~n26307 ;
  assign n26309 = n12553 & ~n20373 ;
  assign n26310 = n22337 ^ n1365 ^ 1'b0 ;
  assign n26311 = x81 & ~n5367 ;
  assign n26312 = n26311 ^ n7254 ^ 1'b0 ;
  assign n26313 = n9702 & n26312 ;
  assign n26314 = ~n6412 & n26313 ;
  assign n26315 = n8870 ^ n7428 ^ 1'b0 ;
  assign n26316 = n22292 & ~n26315 ;
  assign n26317 = n18286 ^ n4975 ^ 1'b0 ;
  assign n26318 = n26316 & ~n26317 ;
  assign n26319 = n24134 ^ n641 ^ 1'b0 ;
  assign n26320 = n584 | n11584 ;
  assign n26321 = n26320 ^ n1654 ^ 1'b0 ;
  assign n26322 = n8564 ^ n2215 ^ 1'b0 ;
  assign n26323 = ~n26321 & n26322 ;
  assign n26324 = ~n5750 & n26323 ;
  assign n26325 = n20824 & n26324 ;
  assign n26326 = ~n1918 & n12787 ;
  assign n26327 = ~n8199 & n26326 ;
  assign n26328 = n8926 | n26327 ;
  assign n26329 = n12535 & ~n26328 ;
  assign n26330 = ~n12103 & n14625 ;
  assign n26331 = n18593 | n26330 ;
  assign n26332 = n5928 & n12171 ;
  assign n26333 = n26332 ^ n5291 ^ 1'b0 ;
  assign n26334 = n3910 & n11103 ;
  assign n26335 = n16111 & n26334 ;
  assign n26336 = n9354 & n9825 ;
  assign n26337 = n26336 ^ n17495 ^ 1'b0 ;
  assign n26338 = n11483 & ~n26337 ;
  assign n26339 = n665 & n26338 ;
  assign n26340 = n4358 & n19716 ;
  assign n26341 = n12133 ^ n7310 ^ 1'b0 ;
  assign n26342 = n21305 | n26341 ;
  assign n26343 = n4898 ^ n2590 ^ 1'b0 ;
  assign n26344 = n21513 & n26343 ;
  assign n26345 = n25129 ^ n23812 ^ 1'b0 ;
  assign n26346 = n26344 & ~n26345 ;
  assign n26347 = n870 ^ n607 ^ 1'b0 ;
  assign n26348 = n10486 & ~n26347 ;
  assign n26349 = ( ~n491 & n5824 ) | ( ~n491 & n10658 ) | ( n5824 & n10658 ) ;
  assign n26350 = n608 | n3413 ;
  assign n26351 = n26350 ^ n17523 ^ n16194 ;
  assign n26352 = n13209 ^ n7158 ^ 1'b0 ;
  assign n26353 = ( n26349 & n26351 ) | ( n26349 & n26352 ) | ( n26351 & n26352 ) ;
  assign n26354 = n19572 ^ n6117 ^ 1'b0 ;
  assign n26355 = n9657 | n14721 ;
  assign n26356 = ( n22033 & n26028 ) | ( n22033 & n26355 ) | ( n26028 & n26355 ) ;
  assign n26357 = n20409 & ~n21412 ;
  assign n26358 = n26357 ^ n3604 ^ 1'b0 ;
  assign n26359 = n6942 | n22265 ;
  assign n26360 = n2435 | n26359 ;
  assign n26361 = n690 | n10312 ;
  assign n26362 = n26361 ^ n18453 ^ 1'b0 ;
  assign n26363 = n19465 ^ n11507 ^ 1'b0 ;
  assign n26364 = n11176 & ~n26363 ;
  assign n26365 = n20222 | n26364 ;
  assign n26366 = ~n3447 & n8184 ;
  assign n26367 = ~n18389 & n26366 ;
  assign n26368 = n26367 ^ n16857 ^ n2448 ;
  assign n26369 = n22385 & n26368 ;
  assign n26370 = n9840 & n11756 ;
  assign n26371 = ( n3378 & ~n5719 ) | ( n3378 & n10125 ) | ( ~n5719 & n10125 ) ;
  assign n26372 = ~n21814 & n22612 ;
  assign n26373 = n26372 ^ n25587 ^ n22819 ;
  assign n26374 = n21766 ^ n15247 ^ n8730 ;
  assign n26375 = n26374 ^ n13198 ^ n4267 ;
  assign n26376 = ~n24737 & n26375 ;
  assign n26377 = n3894 & n26376 ;
  assign n26378 = n26377 ^ n13002 ^ 1'b0 ;
  assign n26379 = n18403 ^ n1376 ^ 1'b0 ;
  assign n26380 = n16698 & n26379 ;
  assign n26381 = n4768 & n13853 ;
  assign n26382 = ~n7987 & n26381 ;
  assign n26383 = n2454 | n26382 ;
  assign n26384 = ~n3649 & n26383 ;
  assign n26385 = n10709 & n26384 ;
  assign n26386 = n7657 | n10298 ;
  assign n26387 = n26386 ^ n5213 ^ 1'b0 ;
  assign n26388 = n2279 | n26387 ;
  assign n26389 = n15140 ^ n8872 ^ n4472 ;
  assign n26390 = n26388 & n26389 ;
  assign n26391 = n11035 & n15053 ;
  assign n26392 = n26391 ^ n19585 ^ n14389 ;
  assign n26393 = n26392 ^ n8231 ^ x6 ;
  assign n26394 = n25357 ^ n4767 ^ n4175 ;
  assign n26395 = n13311 & ~n26394 ;
  assign n26396 = n20397 ^ n9502 ^ n5061 ;
  assign n26397 = ( ~n1588 & n3887 ) | ( ~n1588 & n12888 ) | ( n3887 & n12888 ) ;
  assign n26398 = n19387 ^ n4483 ^ 1'b0 ;
  assign n26399 = n8884 | n26398 ;
  assign n26400 = n744 & ~n6411 ;
  assign n26401 = n26399 & n26400 ;
  assign n26402 = n1066 & n12068 ;
  assign n26403 = ~n6180 & n26402 ;
  assign n26404 = n599 & n3423 ;
  assign n26405 = n26404 ^ n24040 ^ 1'b0 ;
  assign n26406 = ~n16812 & n22697 ;
  assign n26407 = n26406 ^ n21743 ^ 1'b0 ;
  assign n26408 = n17635 & ~n26407 ;
  assign n26409 = n458 & n26408 ;
  assign n26410 = ( n11539 & n13700 ) | ( n11539 & ~n19243 ) | ( n13700 & ~n19243 ) ;
  assign n26411 = n24781 ^ n18444 ^ n11047 ;
  assign n26412 = n23903 | n26411 ;
  assign n26413 = ( n756 & n13323 ) | ( n756 & n26412 ) | ( n13323 & n26412 ) ;
  assign n26414 = n2363 ^ n1745 ^ n517 ;
  assign n26415 = n26414 ^ n25590 ^ n561 ;
  assign n26416 = n4447 | n4891 ;
  assign n26417 = n16842 ^ n3989 ^ 1'b0 ;
  assign n26418 = ( ~n15725 & n26416 ) | ( ~n15725 & n26417 ) | ( n26416 & n26417 ) ;
  assign n26419 = n26418 ^ n15522 ^ 1'b0 ;
  assign n26420 = n23432 ^ n10054 ^ n4646 ;
  assign n26421 = n23936 ^ n18647 ^ 1'b0 ;
  assign n26422 = n8041 ^ n1177 ^ 1'b0 ;
  assign n26423 = n26421 | n26422 ;
  assign n26424 = ~n1127 & n11189 ;
  assign n26425 = ~n4761 & n26424 ;
  assign n26428 = n5832 ^ n4709 ^ 1'b0 ;
  assign n26429 = n13430 & n26428 ;
  assign n26430 = ~n14102 & n26429 ;
  assign n26431 = n26430 ^ n10335 ^ n4373 ;
  assign n26432 = n26431 ^ n22160 ^ n15980 ;
  assign n26433 = n26432 ^ n5458 ^ 1'b0 ;
  assign n26434 = n5984 & n26433 ;
  assign n26426 = n8176 & n9588 ;
  assign n26427 = n26426 ^ n15519 ^ 1'b0 ;
  assign n26435 = n26434 ^ n26427 ^ 1'b0 ;
  assign n26436 = ~n2416 & n11634 ;
  assign n26437 = ~n8047 & n8719 ;
  assign n26438 = n26437 ^ n2822 ^ 1'b0 ;
  assign n26439 = ( n3615 & n15660 ) | ( n3615 & n23205 ) | ( n15660 & n23205 ) ;
  assign n26440 = n26439 ^ n3062 ^ n917 ;
  assign n26441 = n25483 ^ n16227 ^ 1'b0 ;
  assign n26442 = ( n5435 & ~n10432 ) | ( n5435 & n22333 ) | ( ~n10432 & n22333 ) ;
  assign n26444 = n10406 ^ n6408 ^ n6271 ;
  assign n26443 = n8005 | n16824 ;
  assign n26445 = n26444 ^ n26443 ^ 1'b0 ;
  assign n26446 = n23801 & n26445 ;
  assign n26447 = n20884 ^ n652 ^ 1'b0 ;
  assign n26448 = n10154 | n15283 ;
  assign n26449 = ~n1923 & n7984 ;
  assign n26450 = ~n26448 & n26449 ;
  assign n26451 = n13684 ^ n11226 ^ n1560 ;
  assign n26452 = n21087 | n26451 ;
  assign n26455 = n15671 ^ n14955 ^ 1'b0 ;
  assign n26456 = n3771 & n26455 ;
  assign n26453 = ~n1305 & n26355 ;
  assign n26454 = n26453 ^ n16450 ^ 1'b0 ;
  assign n26457 = n26456 ^ n26454 ^ n17981 ;
  assign n26458 = n19180 ^ n13102 ^ 1'b0 ;
  assign n26459 = ( ~n12349 & n18206 ) | ( ~n12349 & n21964 ) | ( n18206 & n21964 ) ;
  assign n26460 = n26459 ^ n16073 ^ n1593 ;
  assign n26461 = ( n3246 & ~n6117 ) | ( n3246 & n8826 ) | ( ~n6117 & n8826 ) ;
  assign n26462 = n5495 | n14283 ;
  assign n26463 = n26461 | n26462 ;
  assign n26464 = n8560 & ~n10471 ;
  assign n26465 = n17063 | n26464 ;
  assign n26466 = n26465 ^ n2977 ^ 1'b0 ;
  assign n26467 = n22057 ^ n6693 ^ 1'b0 ;
  assign n26468 = ~n1582 & n26467 ;
  assign n26469 = x123 & ~n6712 ;
  assign n26470 = n13160 ^ n3975 ^ n956 ;
  assign n26471 = n14177 | n24350 ;
  assign n26472 = n26470 | n26471 ;
  assign n26473 = ( n4533 & n20603 ) | ( n4533 & n26472 ) | ( n20603 & n26472 ) ;
  assign n26475 = n827 | n2124 ;
  assign n26474 = ( n4437 & ~n18560 ) | ( n4437 & n23724 ) | ( ~n18560 & n23724 ) ;
  assign n26476 = n26475 ^ n26474 ^ n1880 ;
  assign n26479 = n6370 ^ n5852 ^ n3628 ;
  assign n26480 = n1233 | n1894 ;
  assign n26481 = n26480 ^ n10120 ^ 1'b0 ;
  assign n26482 = n10322 & ~n26481 ;
  assign n26483 = n26482 ^ n1491 ^ 1'b0 ;
  assign n26484 = ~n26479 & n26483 ;
  assign n26477 = n9526 | n21166 ;
  assign n26478 = n2628 & ~n26477 ;
  assign n26485 = n26484 ^ n26478 ^ n21357 ;
  assign n26486 = n2268 & n7091 ;
  assign n26487 = n26486 ^ n3945 ^ 1'b0 ;
  assign n26488 = n14698 ^ n4123 ^ 1'b0 ;
  assign n26489 = n6139 & n26488 ;
  assign n26490 = n7950 & n26489 ;
  assign n26491 = n26490 ^ n23943 ^ 1'b0 ;
  assign n26492 = n19161 ^ n3958 ^ 1'b0 ;
  assign n26493 = ~n17544 & n26492 ;
  assign n26494 = n4110 & n26493 ;
  assign n26495 = n26494 ^ n12638 ^ 1'b0 ;
  assign n26496 = n25826 ^ n10666 ^ 1'b0 ;
  assign n26497 = ( n557 & n6187 ) | ( n557 & n9607 ) | ( n6187 & n9607 ) ;
  assign n26498 = n26497 ^ n1036 ^ 1'b0 ;
  assign n26499 = n22022 & ~n26498 ;
  assign n26500 = n26499 ^ n24186 ^ 1'b0 ;
  assign n26501 = n917 & ~n5944 ;
  assign n26502 = ~n2724 & n26501 ;
  assign n26503 = n24400 ^ n8712 ^ n6530 ;
  assign n26504 = n12647 & n26503 ;
  assign n26505 = ( ~n1370 & n7257 ) | ( ~n1370 & n20197 ) | ( n7257 & n20197 ) ;
  assign n26506 = n10914 & n18469 ;
  assign n26507 = n26506 ^ n25060 ^ 1'b0 ;
  assign n26508 = ( n3837 & n16485 ) | ( n3837 & n26507 ) | ( n16485 & n26507 ) ;
  assign n26509 = n1240 & n14083 ;
  assign n26510 = n16503 & n16603 ;
  assign n26511 = n16913 ^ n16153 ^ 1'b0 ;
  assign n26512 = n13659 ^ n5930 ^ 1'b0 ;
  assign n26513 = n26512 ^ n25975 ^ 1'b0 ;
  assign n26514 = n4895 ^ n803 ^ 1'b0 ;
  assign n26515 = n7839 & ~n9970 ;
  assign n26516 = n26515 ^ n16579 ^ 1'b0 ;
  assign n26517 = n26516 ^ n16117 ^ n10645 ;
  assign n26518 = n26517 ^ n18817 ^ 1'b0 ;
  assign n26519 = x84 & ~n26518 ;
  assign n26520 = n26519 ^ n24718 ^ n24252 ;
  assign n26521 = n20128 ^ n16531 ^ n5613 ;
  assign n26522 = n26521 ^ n16493 ^ 1'b0 ;
  assign n26523 = n12850 ^ n11562 ^ n6017 ;
  assign n26524 = n19052 ^ n7273 ^ n236 ;
  assign n26525 = ( n2180 & n15612 ) | ( n2180 & ~n26524 ) | ( n15612 & ~n26524 ) ;
  assign n26526 = n12718 ^ n5977 ^ 1'b0 ;
  assign n26527 = n2303 & ~n26526 ;
  assign n26528 = n19430 & n26527 ;
  assign n26529 = n26528 ^ n11532 ^ 1'b0 ;
  assign n26530 = n19675 & n26529 ;
  assign n26531 = ~n2400 & n9610 ;
  assign n26532 = n26531 ^ n18861 ^ 1'b0 ;
  assign n26533 = n4144 ^ n2258 ^ 1'b0 ;
  assign n26534 = n11723 ^ n3919 ^ 1'b0 ;
  assign n26535 = x118 & ~n26534 ;
  assign n26536 = ~n892 & n26535 ;
  assign n26537 = ~n26533 & n26536 ;
  assign n26538 = n15469 ^ n3159 ^ 1'b0 ;
  assign n26539 = n12866 | n25905 ;
  assign n26540 = ~n6356 & n26539 ;
  assign n26541 = n3945 & n7733 ;
  assign n26542 = ( ~n697 & n16336 ) | ( ~n697 & n26357 ) | ( n16336 & n26357 ) ;
  assign n26543 = ( n10687 & n19017 ) | ( n10687 & n26542 ) | ( n19017 & n26542 ) ;
  assign n26544 = n10071 | n24664 ;
  assign n26546 = n616 & ~n1450 ;
  assign n26545 = n1696 & n19239 ;
  assign n26547 = n26546 ^ n26545 ^ 1'b0 ;
  assign n26548 = n14196 & ~n21793 ;
  assign n26549 = n23798 & ~n26548 ;
  assign n26550 = n6178 & n26549 ;
  assign n26551 = n13105 ^ n6552 ^ 1'b0 ;
  assign n26552 = n11666 & ~n26551 ;
  assign n26553 = ~n15740 & n17173 ;
  assign n26554 = ~n11856 & n22360 ;
  assign n26555 = n6573 | n13819 ;
  assign n26556 = n26555 ^ n3834 ^ 1'b0 ;
  assign n26557 = n21705 & n26556 ;
  assign n26558 = n9996 | n26557 ;
  assign n26559 = n19270 & ~n26558 ;
  assign n26560 = n24116 ^ n17383 ^ 1'b0 ;
  assign n26561 = n4170 & n26560 ;
  assign n26562 = ( n5537 & ~n11967 ) | ( n5537 & n26561 ) | ( ~n11967 & n26561 ) ;
  assign n26564 = n7053 ^ n2555 ^ n2139 ;
  assign n26563 = n6228 & n19234 ;
  assign n26565 = n26564 ^ n26563 ^ 1'b0 ;
  assign n26566 = n26565 ^ n2731 ^ 1'b0 ;
  assign n26567 = n2654 & ~n6543 ;
  assign n26568 = n11572 & n26567 ;
  assign n26569 = n10608 | n24641 ;
  assign n26570 = n553 & n19368 ;
  assign n26571 = n26570 ^ n15044 ^ 1'b0 ;
  assign n26573 = ~n1871 & n22057 ;
  assign n26574 = ( ~n14163 & n24206 ) | ( ~n14163 & n25287 ) | ( n24206 & n25287 ) ;
  assign n26575 = ( n11998 & n26573 ) | ( n11998 & n26574 ) | ( n26573 & n26574 ) ;
  assign n26572 = n2107 | n12198 ;
  assign n26576 = n26575 ^ n26572 ^ 1'b0 ;
  assign n26577 = ~n250 & n6614 ;
  assign n26578 = n19872 ^ n18507 ^ n9730 ;
  assign n26579 = n12782 ^ n9483 ^ 1'b0 ;
  assign n26580 = n26579 ^ n9688 ^ 1'b0 ;
  assign n26581 = ~n11158 & n12553 ;
  assign n26582 = ~n16780 & n26581 ;
  assign n26583 = n12751 ^ n10458 ^ n2451 ;
  assign n26584 = n2334 & ~n7133 ;
  assign n26585 = n26584 ^ n384 ^ 1'b0 ;
  assign n26586 = ~n11954 & n26585 ;
  assign n26587 = n12706 ^ n10338 ^ 1'b0 ;
  assign n26588 = n8605 ^ n3048 ^ 1'b0 ;
  assign n26589 = n26587 | n26588 ;
  assign n26590 = ~n8106 & n21596 ;
  assign n26591 = n18932 & n26590 ;
  assign n26592 = ( n4605 & ~n8204 ) | ( n4605 & n15410 ) | ( ~n8204 & n15410 ) ;
  assign n26593 = n7548 ^ n5938 ^ n1502 ;
  assign n26594 = n26593 ^ n12787 ^ 1'b0 ;
  assign n26595 = ~n15717 & n26594 ;
  assign n26596 = n760 & n6524 ;
  assign n26597 = n17597 | n26596 ;
  assign n26598 = n2060 & n8944 ;
  assign n26599 = ( ~n5734 & n8421 ) | ( ~n5734 & n26598 ) | ( n8421 & n26598 ) ;
  assign n26600 = n26599 ^ n16383 ^ 1'b0 ;
  assign n26601 = n23933 ^ n1199 ^ 1'b0 ;
  assign n26602 = n19394 & ~n26601 ;
  assign n26604 = n2692 & n11455 ;
  assign n26605 = n26604 ^ n2576 ^ 1'b0 ;
  assign n26606 = n26605 ^ n7206 ^ 1'b0 ;
  assign n26607 = ~n8453 & n26606 ;
  assign n26603 = n3240 & n24698 ;
  assign n26608 = n26607 ^ n26603 ^ n25101 ;
  assign n26609 = n10352 ^ n7526 ^ n7097 ;
  assign n26610 = ( n5239 & n20508 ) | ( n5239 & n21357 ) | ( n20508 & n21357 ) ;
  assign n26611 = n8240 & ~n25902 ;
  assign n26612 = n3854 & ~n14067 ;
  assign n26613 = n22879 ^ n431 ^ 1'b0 ;
  assign n26614 = n22213 | n26613 ;
  assign n26615 = ~n2763 & n7697 ;
  assign n26616 = n26615 ^ n11235 ^ 1'b0 ;
  assign n26617 = n3449 | n7176 ;
  assign n26618 = n3240 & n8212 ;
  assign n26619 = n13715 ^ n2349 ^ n618 ;
  assign n26620 = ~n2818 & n3986 ;
  assign n26621 = n21063 ^ n6537 ^ 1'b0 ;
  assign n26622 = ~n3180 & n25039 ;
  assign n26623 = n26622 ^ n22344 ^ 1'b0 ;
  assign n26624 = n9673 & ~n14772 ;
  assign n26625 = ~n16182 & n26624 ;
  assign n26626 = n4156 & n6285 ;
  assign n26627 = n3240 & n26626 ;
  assign n26628 = n146 | n4561 ;
  assign n26629 = n26628 ^ n9177 ^ 1'b0 ;
  assign n26630 = ( n6878 & n11048 ) | ( n6878 & n26629 ) | ( n11048 & n26629 ) ;
  assign n26631 = n23112 ^ n4314 ^ n2792 ;
  assign n26632 = n15819 & n26631 ;
  assign n26633 = ~n6265 & n26632 ;
  assign n26634 = n26633 ^ n23958 ^ n22320 ;
  assign n26635 = n26634 ^ n15524 ^ n1112 ;
  assign n26636 = n8198 ^ n4697 ^ n1695 ;
  assign n26637 = n19220 ^ n4593 ^ 1'b0 ;
  assign n26638 = n1483 ^ n1209 ^ n1076 ;
  assign n26639 = ~n13296 & n21352 ;
  assign n26640 = ~n5773 & n26639 ;
  assign n26641 = n26638 | n26640 ;
  assign n26642 = n21651 ^ n8093 ^ n5517 ;
  assign n26643 = n9329 ^ n972 ^ 1'b0 ;
  assign n26644 = n4707 & n26643 ;
  assign n26645 = n19932 ^ n13186 ^ n7839 ;
  assign n26646 = ( n22488 & n26644 ) | ( n22488 & ~n26645 ) | ( n26644 & ~n26645 ) ;
  assign n26647 = n26642 & ~n26646 ;
  assign n26648 = n2265 & n26647 ;
  assign n26650 = n3961 ^ n1200 ^ n594 ;
  assign n26651 = n26650 ^ n11470 ^ 1'b0 ;
  assign n26649 = n19967 ^ n4154 ^ 1'b0 ;
  assign n26652 = n26651 ^ n26649 ^ 1'b0 ;
  assign n26653 = ( n9473 & ~n12035 ) | ( n9473 & n17632 ) | ( ~n12035 & n17632 ) ;
  assign n26654 = n19491 ^ n17200 ^ n2406 ;
  assign n26655 = n24718 ^ n22760 ^ n8321 ;
  assign n26656 = n12600 & n20669 ;
  assign n26657 = n16092 & n26656 ;
  assign n26658 = n13004 ^ n584 ^ 1'b0 ;
  assign n26659 = n9013 & n26658 ;
  assign n26660 = n20559 ^ n3525 ^ 1'b0 ;
  assign n26661 = n1776 | n26660 ;
  assign n26662 = n16162 & n17381 ;
  assign n26663 = ( n5484 & n5554 ) | ( n5484 & ~n15863 ) | ( n5554 & ~n15863 ) ;
  assign n26664 = ( n13441 & ~n16801 ) | ( n13441 & n22189 ) | ( ~n16801 & n22189 ) ;
  assign n26665 = n16105 ^ n15647 ^ n427 ;
  assign n26666 = n1754 | n9358 ;
  assign n26667 = n26666 ^ n15159 ^ n2984 ;
  assign n26668 = ( n2884 & n22259 ) | ( n2884 & n26667 ) | ( n22259 & n26667 ) ;
  assign n26670 = n2851 | n16610 ;
  assign n26669 = n19380 ^ n3366 ^ 1'b0 ;
  assign n26671 = n26670 ^ n26669 ^ n6256 ;
  assign n26672 = n6252 & n26671 ;
  assign n26673 = ( n1331 & n20423 ) | ( n1331 & ~n20443 ) | ( n20423 & ~n20443 ) ;
  assign n26674 = n18885 & n26673 ;
  assign n26675 = n21843 & n26674 ;
  assign n26676 = n1854 | n11715 ;
  assign n26679 = n2834 & n20380 ;
  assign n26677 = n3049 ^ n746 ^ 1'b0 ;
  assign n26678 = n8288 & n26677 ;
  assign n26680 = n26679 ^ n26678 ^ 1'b0 ;
  assign n26681 = ( n3074 & n11793 ) | ( n3074 & n15061 ) | ( n11793 & n15061 ) ;
  assign n26682 = n17460 ^ n8038 ^ n5664 ;
  assign n26683 = ( ~n5115 & n8154 ) | ( ~n5115 & n26682 ) | ( n8154 & n26682 ) ;
  assign n26684 = ( n3830 & ~n5583 ) | ( n3830 & n13332 ) | ( ~n5583 & n13332 ) ;
  assign n26685 = n3916 & n26684 ;
  assign n26686 = n26685 ^ n620 ^ 1'b0 ;
  assign n26687 = n11686 & ~n19959 ;
  assign n26688 = n19486 & ~n26687 ;
  assign n26689 = ~n26644 & n26688 ;
  assign n26690 = n14095 ^ n9085 ^ 1'b0 ;
  assign n26691 = n20873 ^ n9919 ^ n6522 ;
  assign n26692 = n26690 & n26691 ;
  assign n26693 = n14630 ^ n2933 ^ 1'b0 ;
  assign n26694 = n25090 ^ n21738 ^ n12112 ;
  assign n26695 = n21936 ^ n9164 ^ 1'b0 ;
  assign n26696 = n2021 & n8565 ;
  assign n26697 = ~n2183 & n5126 ;
  assign n26698 = ~n8609 & n26697 ;
  assign n26699 = n26698 ^ n1678 ^ 1'b0 ;
  assign n26700 = n26696 | n26699 ;
  assign n26701 = n1365 | n14086 ;
  assign n26706 = n7805 & n15291 ;
  assign n26705 = n6614 & ~n11402 ;
  assign n26707 = n26706 ^ n26705 ^ 1'b0 ;
  assign n26702 = n13052 & ~n18593 ;
  assign n26703 = ~n2378 & n26702 ;
  assign n26704 = n7003 | n26703 ;
  assign n26708 = n26707 ^ n26704 ^ 1'b0 ;
  assign n26709 = n16813 ^ n15854 ^ n1200 ;
  assign n26710 = n2547 | n10527 ;
  assign n26711 = n22879 & ~n26710 ;
  assign n26712 = n26711 ^ n21483 ^ n146 ;
  assign n26713 = n13460 ^ n13108 ^ 1'b0 ;
  assign n26714 = n15000 | n22431 ;
  assign n26715 = n26713 | n26714 ;
  assign n26716 = n3758 & ~n14727 ;
  assign n26717 = n24760 & n26716 ;
  assign n26718 = n6220 ^ n3383 ^ n270 ;
  assign n26719 = n5655 & ~n26718 ;
  assign n26720 = n1626 & n26719 ;
  assign n26721 = n20643 ^ n14778 ^ 1'b0 ;
  assign n26722 = n9349 & ~n26721 ;
  assign n26723 = ~n393 & n16603 ;
  assign n26724 = ~n7450 & n26723 ;
  assign n26725 = ~n6183 & n24255 ;
  assign n26726 = n26725 ^ n5247 ^ 1'b0 ;
  assign n26727 = n2705 & ~n16518 ;
  assign n26728 = n26727 ^ n5317 ^ 1'b0 ;
  assign n26729 = n8970 | n26728 ;
  assign n26730 = n21119 ^ n17515 ^ n6908 ;
  assign n26735 = n14998 ^ n11412 ^ n7581 ;
  assign n26734 = n10981 & ~n13475 ;
  assign n26732 = ~n2956 & n12937 ;
  assign n26731 = n6811 & ~n13449 ;
  assign n26733 = n26732 ^ n26731 ^ 1'b0 ;
  assign n26736 = n26735 ^ n26734 ^ n26733 ;
  assign n26737 = n8221 & n19539 ;
  assign n26738 = n24998 & n26737 ;
  assign n26739 = n26738 ^ n3513 ^ 1'b0 ;
  assign n26740 = n1845 ^ x104 ^ 1'b0 ;
  assign n26741 = ~n11566 & n26740 ;
  assign n26742 = n19293 ^ n10932 ^ 1'b0 ;
  assign n26743 = n22114 ^ n1060 ^ 1'b0 ;
  assign n26744 = n9054 & ~n26743 ;
  assign n26747 = n4871 & ~n14201 ;
  assign n26748 = n18958 & n26747 ;
  assign n26749 = n26748 ^ n339 ^ 1'b0 ;
  assign n26745 = n4891 | n15396 ;
  assign n26746 = n11227 & ~n26745 ;
  assign n26750 = n26749 ^ n26746 ^ 1'b0 ;
  assign n26751 = n20189 ^ n511 ^ 1'b0 ;
  assign n26752 = n26751 ^ n15107 ^ n8342 ;
  assign n26753 = ( ~n7232 & n7284 ) | ( ~n7232 & n8942 ) | ( n7284 & n8942 ) ;
  assign n26754 = ( n6818 & ~n10875 ) | ( n6818 & n12428 ) | ( ~n10875 & n12428 ) ;
  assign n26755 = n2216 & ~n15419 ;
  assign n26756 = n26755 ^ n6191 ^ 1'b0 ;
  assign n26757 = n26756 ^ n2849 ^ 1'b0 ;
  assign n26758 = ~n19200 & n26757 ;
  assign n26759 = ~n7103 & n11160 ;
  assign n26760 = n26759 ^ n1003 ^ 1'b0 ;
  assign n26761 = n20830 | n26760 ;
  assign n26762 = n2085 | n26761 ;
  assign n26763 = n12014 & ~n22213 ;
  assign n26764 = n16539 & n26763 ;
  assign n26765 = n10885 & n16023 ;
  assign n26766 = n469 | n25357 ;
  assign n26767 = ~n14137 & n26766 ;
  assign n26768 = n26767 ^ n13973 ^ 1'b0 ;
  assign n26769 = n26497 ^ n8795 ^ 1'b0 ;
  assign n26770 = ~n2039 & n21156 ;
  assign n26771 = n2567 & ~n8783 ;
  assign n26772 = ( n1736 & n5174 ) | ( n1736 & n7760 ) | ( n5174 & n7760 ) ;
  assign n26773 = n10597 ^ n358 ^ x122 ;
  assign n26774 = n16775 ^ n10967 ^ 1'b0 ;
  assign n26775 = ~n16568 & n26774 ;
  assign n26776 = n26775 ^ n25350 ^ n7377 ;
  assign n26777 = n18969 ^ n14521 ^ 1'b0 ;
  assign n26778 = n17348 | n26056 ;
  assign n26779 = n22428 ^ n948 ^ 1'b0 ;
  assign n26780 = ~n15888 & n26779 ;
  assign n26781 = ~n14622 & n19512 ;
  assign n26782 = n26781 ^ n4185 ^ 1'b0 ;
  assign n26783 = ( ~n9766 & n10483 ) | ( ~n9766 & n15496 ) | ( n10483 & n15496 ) ;
  assign n26784 = ~n5915 & n9898 ;
  assign n26785 = ~n26783 & n26784 ;
  assign n26786 = n26785 ^ n16111 ^ 1'b0 ;
  assign n26787 = n4271 ^ n2171 ^ 1'b0 ;
  assign n26788 = ~n5387 & n23535 ;
  assign n26789 = n11464 & n26788 ;
  assign n26790 = n12773 ^ n12464 ^ n12115 ;
  assign n26791 = ~n10165 & n19509 ;
  assign n26792 = ( n17021 & ~n17177 ) | ( n17021 & n26791 ) | ( ~n17177 & n26791 ) ;
  assign n26794 = ( ~n6327 & n13626 ) | ( ~n6327 & n22023 ) | ( n13626 & n22023 ) ;
  assign n26793 = n20351 ^ n17399 ^ n1660 ;
  assign n26795 = n26794 ^ n26793 ^ n4229 ;
  assign n26796 = n9619 ^ n9242 ^ 1'b0 ;
  assign n26797 = n19880 | n26796 ;
  assign n26798 = ~n11190 & n17966 ;
  assign n26799 = ~n24507 & n26798 ;
  assign n26800 = n1745 & ~n17571 ;
  assign n26801 = ( n17827 & ~n20373 ) | ( n17827 & n26800 ) | ( ~n20373 & n26800 ) ;
  assign n26802 = n3442 & n4497 ;
  assign n26803 = n26802 ^ n15676 ^ n6977 ;
  assign n26804 = n26233 ^ n19767 ^ n4950 ;
  assign n26805 = n8343 | n15789 ;
  assign n26806 = ~n7040 & n26805 ;
  assign n26807 = n26806 ^ n25561 ^ n372 ;
  assign n26808 = n1937 | n15304 ;
  assign n26809 = n15221 & ~n26808 ;
  assign n26810 = n16771 & n25520 ;
  assign n26812 = ~n4618 & n17769 ;
  assign n26813 = n8519 | n26812 ;
  assign n26811 = n4527 & ~n11960 ;
  assign n26814 = n26813 ^ n26811 ^ 1'b0 ;
  assign n26815 = ( n4226 & n4669 ) | ( n4226 & ~n5059 ) | ( n4669 & ~n5059 ) ;
  assign n26816 = ~n900 & n4434 ;
  assign n26817 = ( n140 & n26815 ) | ( n140 & n26816 ) | ( n26815 & n26816 ) ;
  assign n26818 = n4806 & ~n8092 ;
  assign n26819 = ~n26817 & n26818 ;
  assign n26820 = n24071 ^ n2110 ^ 1'b0 ;
  assign n26821 = n2789 & n26820 ;
  assign n26822 = n10420 ^ n5569 ^ 1'b0 ;
  assign n26823 = ~n12628 & n26822 ;
  assign n26824 = ( n8729 & ~n21884 ) | ( n8729 & n22368 ) | ( ~n21884 & n22368 ) ;
  assign n26825 = n21886 ^ n11211 ^ 1'b0 ;
  assign n26826 = n3674 | n8160 ;
  assign n26827 = ( ~n1184 & n18065 ) | ( ~n1184 & n26826 ) | ( n18065 & n26826 ) ;
  assign n26828 = ~n3072 & n10154 ;
  assign n26829 = ~n10154 & n26828 ;
  assign n26830 = n1519 | n26829 ;
  assign n26831 = n26830 ^ n17619 ^ 1'b0 ;
  assign n26832 = n26831 ^ n24743 ^ n13693 ;
  assign n26833 = n13112 | n26832 ;
  assign n26834 = n14697 | n26833 ;
  assign n26835 = n8406 ^ n3247 ^ 1'b0 ;
  assign n26836 = ~n1449 & n26835 ;
  assign n26837 = n11560 | n26836 ;
  assign n26838 = n23621 ^ n22476 ^ 1'b0 ;
  assign n26839 = n17908 ^ n8272 ^ 1'b0 ;
  assign n26840 = ( n982 & n26838 ) | ( n982 & n26839 ) | ( n26838 & n26839 ) ;
  assign n26841 = n9168 | n13391 ;
  assign n26842 = n12965 | n26841 ;
  assign n26843 = n270 | n2200 ;
  assign n26844 = n6258 | n26843 ;
  assign n26845 = n18218 ^ n17290 ^ n3447 ;
  assign n26846 = ~n6813 & n18733 ;
  assign n26847 = ~n2931 & n26846 ;
  assign n26848 = ~n15414 & n24208 ;
  assign n26849 = n26848 ^ n24481 ^ 1'b0 ;
  assign n26850 = ~n10556 & n16362 ;
  assign n26851 = n7201 ^ n6087 ^ 1'b0 ;
  assign n26852 = n7022 & ~n26851 ;
  assign n26853 = n252 & n1876 ;
  assign n26854 = n12268 & n26853 ;
  assign n26855 = n8648 ^ n206 ^ 1'b0 ;
  assign n26856 = n26854 | n26855 ;
  assign n26857 = n10539 | n21724 ;
  assign n26858 = ~n21468 & n22257 ;
  assign n26859 = n5223 & n26858 ;
  assign n26860 = ( n285 & n2971 ) | ( n285 & ~n26859 ) | ( n2971 & ~n26859 ) ;
  assign n26861 = n9845 | n10476 ;
  assign n26862 = n2586 | n7658 ;
  assign n26863 = n701 & n20112 ;
  assign n26864 = n26863 ^ n1713 ^ 1'b0 ;
  assign n26865 = ~n14573 & n26864 ;
  assign n26866 = n24405 ^ n20873 ^ 1'b0 ;
  assign n26867 = n17076 | n26866 ;
  assign n26868 = ~n18252 & n24494 ;
  assign n26869 = ~n5814 & n26868 ;
  assign n26870 = n6423 & ~n22130 ;
  assign n26871 = n20454 & n26870 ;
  assign n26872 = n13645 ^ n10797 ^ 1'b0 ;
  assign n26873 = n16121 | n26872 ;
  assign n26874 = x11 & n3582 ;
  assign n26875 = n2422 & n26874 ;
  assign n26876 = n26873 & n26875 ;
  assign n26877 = n20413 | n24646 ;
  assign n26878 = n14240 ^ n13128 ^ n12203 ;
  assign n26879 = n7910 ^ n6349 ^ n5155 ;
  assign n26880 = n4598 & ~n5840 ;
  assign n26881 = ~n23467 & n26880 ;
  assign n26882 = n20335 ^ n191 ^ 1'b0 ;
  assign n26883 = n4045 | n26882 ;
  assign n26884 = n9017 ^ n5812 ^ 1'b0 ;
  assign n26885 = n4197 & ~n26884 ;
  assign n26886 = n3466 & ~n4857 ;
  assign n26888 = ( ~n5726 & n10464 ) | ( ~n5726 & n19395 ) | ( n10464 & n19395 ) ;
  assign n26887 = ~n18355 & n18649 ;
  assign n26889 = n26888 ^ n26887 ^ 1'b0 ;
  assign n26890 = n22177 ^ n8929 ^ 1'b0 ;
  assign n26891 = n8201 | n26890 ;
  assign n26892 = n26891 ^ n14143 ^ 1'b0 ;
  assign n26893 = n6275 ^ x49 ^ 1'b0 ;
  assign n26894 = ( ~n13904 & n25306 ) | ( ~n13904 & n26893 ) | ( n25306 & n26893 ) ;
  assign n26895 = ~n6935 & n16470 ;
  assign n26896 = n12990 ^ n3157 ^ 1'b0 ;
  assign n26897 = n992 ^ n314 ^ 1'b0 ;
  assign n26898 = n1200 & ~n26897 ;
  assign n26899 = n4841 & ~n18324 ;
  assign n26900 = ( n1888 & ~n3545 ) | ( n1888 & n14387 ) | ( ~n3545 & n14387 ) ;
  assign n26901 = ~n5123 & n26900 ;
  assign n26902 = n10867 & ~n15542 ;
  assign n26903 = n26902 ^ n18350 ^ 1'b0 ;
  assign n26904 = n5900 & ~n13620 ;
  assign n26907 = n6325 & n12295 ;
  assign n26906 = n3618 & n15863 ;
  assign n26905 = ( n824 & ~n7475 ) | ( n824 & n17117 ) | ( ~n7475 & n17117 ) ;
  assign n26908 = n26907 ^ n26906 ^ n26905 ;
  assign n26909 = n19465 ^ n16611 ^ 1'b0 ;
  assign n26910 = ( ~n6552 & n18004 ) | ( ~n6552 & n25088 ) | ( n18004 & n25088 ) ;
  assign n26911 = ( n5611 & n13653 ) | ( n5611 & ~n26605 ) | ( n13653 & ~n26605 ) ;
  assign n26912 = n24504 | n26911 ;
  assign n26913 = ~n1892 & n14452 ;
  assign n26914 = n2785 & n21009 ;
  assign n26915 = ~n1093 & n26914 ;
  assign n26916 = n5995 | n26915 ;
  assign n26917 = n10112 & ~n26916 ;
  assign n26918 = n3638 & ~n4929 ;
  assign n26919 = n3263 ^ n2437 ^ 1'b0 ;
  assign n26920 = n10588 | n26919 ;
  assign n26921 = n8503 ^ n1373 ^ 1'b0 ;
  assign n26922 = n2647 & ~n26921 ;
  assign n26923 = n26922 ^ n8346 ^ 1'b0 ;
  assign n26924 = n12299 ^ x45 ^ 1'b0 ;
  assign n26925 = ( n4620 & ~n22725 ) | ( n4620 & n26924 ) | ( ~n22725 & n26924 ) ;
  assign n26926 = ( n6310 & n21160 ) | ( n6310 & n21949 ) | ( n21160 & n21949 ) ;
  assign n26932 = n8097 & ~n8599 ;
  assign n26927 = n6886 & ~n11412 ;
  assign n26928 = n26927 ^ n7625 ^ 1'b0 ;
  assign n26929 = n5915 | n26928 ;
  assign n26930 = n26929 ^ n18145 ^ 1'b0 ;
  assign n26931 = n5463 & ~n26930 ;
  assign n26933 = n26932 ^ n26931 ^ n25916 ;
  assign n26934 = n9520 ^ n8828 ^ 1'b0 ;
  assign n26935 = n25716 & ~n26934 ;
  assign n26936 = n9933 ^ n7328 ^ 1'b0 ;
  assign n26937 = ~n6744 & n17581 ;
  assign n26938 = ~n9039 & n26937 ;
  assign n26939 = n17314 ^ n6247 ^ n3567 ;
  assign n26940 = n15577 & n26939 ;
  assign n26941 = n22742 ^ n20184 ^ n17142 ;
  assign n26942 = n4641 ^ n3855 ^ 1'b0 ;
  assign n26943 = n26942 ^ n23628 ^ n1956 ;
  assign n26944 = n5175 | n8944 ;
  assign n26945 = n16853 | n26944 ;
  assign n26946 = n3552 & n21065 ;
  assign n26947 = n26946 ^ n24119 ^ 1'b0 ;
  assign n26948 = n26947 ^ n15724 ^ 1'b0 ;
  assign n26949 = ( n6981 & n26945 ) | ( n6981 & n26948 ) | ( n26945 & n26948 ) ;
  assign n26950 = n15734 ^ n12809 ^ 1'b0 ;
  assign n26951 = ~n10700 & n26950 ;
  assign n26952 = n17591 ^ n1858 ^ 1'b0 ;
  assign n26953 = ~n12225 & n26952 ;
  assign n26954 = ~n4570 & n11084 ;
  assign n26955 = ~n21985 & n26954 ;
  assign n26956 = n26955 ^ n17517 ^ 1'b0 ;
  assign n26957 = n7481 ^ n6461 ^ 1'b0 ;
  assign n26958 = n5352 & n26957 ;
  assign n26959 = n26958 ^ n824 ^ 1'b0 ;
  assign n26960 = n26959 ^ n10925 ^ 1'b0 ;
  assign n26963 = n2897 & ~n5566 ;
  assign n26964 = ~n828 & n26963 ;
  assign n26961 = n3263 | n5649 ;
  assign n26962 = n26961 ^ n7077 ^ 1'b0 ;
  assign n26965 = n26964 ^ n26962 ^ n18927 ;
  assign n26966 = n14585 ^ n2366 ^ 1'b0 ;
  assign n26967 = n26966 ^ n26858 ^ x78 ;
  assign n26968 = n25814 ^ n8815 ^ 1'b0 ;
  assign n26969 = n26968 ^ n20884 ^ n1483 ;
  assign n26970 = n9488 ^ n9262 ^ 1'b0 ;
  assign n26971 = ~n17775 & n26970 ;
  assign n26972 = n2308 & n4175 ;
  assign n26973 = n3968 & n8127 ;
  assign n26974 = n25849 ^ n21805 ^ 1'b0 ;
  assign n26975 = ~n13700 & n15817 ;
  assign n26976 = n9982 & ~n26975 ;
  assign n26977 = n732 & n13993 ;
  assign n26978 = n26977 ^ n1927 ^ 1'b0 ;
  assign n26979 = ( n2426 & ~n6345 ) | ( n2426 & n26978 ) | ( ~n6345 & n26978 ) ;
  assign n26980 = n19770 & n26979 ;
  assign n26981 = n15440 ^ n9464 ^ n2789 ;
  assign n26982 = ~n16733 & n26981 ;
  assign n26983 = ~n6126 & n6906 ;
  assign n26984 = n20910 | n26293 ;
  assign n26985 = n26984 ^ n25862 ^ 1'b0 ;
  assign n26986 = n25421 | n26819 ;
  assign n26987 = n26986 ^ n14618 ^ 1'b0 ;
  assign n26988 = n4625 & ~n19313 ;
  assign n26989 = n6249 & ~n26988 ;
  assign n26990 = n936 & n9963 ;
  assign n26991 = n26990 ^ n173 ^ 1'b0 ;
  assign n26992 = n6430 | n23504 ;
  assign n26993 = n13819 | n23505 ;
  assign n26994 = n23429 ^ n6798 ^ n3163 ;
  assign n26995 = ~n2459 & n6583 ;
  assign n26996 = n26995 ^ n2432 ^ 1'b0 ;
  assign n26997 = n26996 ^ n4592 ^ 1'b0 ;
  assign n26998 = n6916 ^ n5885 ^ 1'b0 ;
  assign n26999 = n23586 | n26998 ;
  assign n27000 = n26999 ^ n8777 ^ 1'b0 ;
  assign n27001 = n20979 & ~n27000 ;
  assign n27002 = n4261 & ~n14694 ;
  assign n27003 = n27002 ^ n1280 ^ 1'b0 ;
  assign n27004 = n17767 ^ n9888 ^ 1'b0 ;
  assign n27005 = n5813 ^ n2647 ^ 1'b0 ;
  assign n27006 = n136 & ~n3257 ;
  assign n27007 = n16227 ^ n10723 ^ 1'b0 ;
  assign n27008 = n7304 & ~n27007 ;
  assign n27009 = ( ~n7618 & n13414 ) | ( ~n7618 & n20118 ) | ( n13414 & n20118 ) ;
  assign n27010 = ( n3697 & n6347 ) | ( n3697 & n25650 ) | ( n6347 & n25650 ) ;
  assign n27011 = n14341 ^ n1408 ^ 1'b0 ;
  assign n27012 = n445 & n2254 ;
  assign n27013 = n27011 & n27012 ;
  assign n27014 = n17643 & ~n19213 ;
  assign n27015 = n27013 & n27014 ;
  assign n27016 = ( n12062 & ~n20325 ) | ( n12062 & n27015 ) | ( ~n20325 & n27015 ) ;
  assign n27017 = n6903 ^ n5663 ^ 1'b0 ;
  assign n27018 = n14781 | n27017 ;
  assign n27019 = n24640 | n27018 ;
  assign n27020 = n10131 ^ n5613 ^ 1'b0 ;
  assign n27021 = ~n27019 & n27020 ;
  assign n27022 = n2381 & n12555 ;
  assign n27023 = ~n630 & n27022 ;
  assign n27024 = n6398 & ~n22987 ;
  assign n27025 = n1831 & n4038 ;
  assign n27026 = n2089 & ~n3657 ;
  assign n27027 = n27025 & n27026 ;
  assign n27028 = n17420 ^ n800 ^ 1'b0 ;
  assign n27029 = n3012 | n27028 ;
  assign n27030 = n14787 | n27029 ;
  assign n27031 = n27030 ^ n6186 ^ n3389 ;
  assign n27032 = ~n2870 & n12913 ;
  assign n27033 = n13631 & n27032 ;
  assign n27034 = n27033 ^ n25627 ^ 1'b0 ;
  assign n27035 = ( x41 & n27031 ) | ( x41 & ~n27034 ) | ( n27031 & ~n27034 ) ;
  assign n27036 = n21964 ^ x101 ^ 1'b0 ;
  assign n27037 = ( ~n15747 & n22235 ) | ( ~n15747 & n27036 ) | ( n22235 & n27036 ) ;
  assign n27038 = n7473 ^ n2452 ^ 1'b0 ;
  assign n27039 = n20313 | n27038 ;
  assign n27040 = n27039 ^ n4387 ^ n3022 ;
  assign n27041 = n20847 ^ n3185 ^ 1'b0 ;
  assign n27042 = n27040 | n27041 ;
  assign n27043 = ( n9575 & n14594 ) | ( n9575 & n27042 ) | ( n14594 & n27042 ) ;
  assign n27044 = ~n14164 & n21488 ;
  assign n27045 = n11142 & ~n12678 ;
  assign n27046 = n27045 ^ n18253 ^ 1'b0 ;
  assign n27047 = ~n15301 & n16638 ;
  assign n27048 = n2303 & n3012 ;
  assign n27049 = n27048 ^ n3345 ^ 1'b0 ;
  assign n27050 = n10672 & ~n18320 ;
  assign n27051 = n6137 & n27050 ;
  assign n27052 = ( n6454 & ~n15226 ) | ( n6454 & n20986 ) | ( ~n15226 & n20986 ) ;
  assign n27053 = ( n6821 & ~n17811 ) | ( n6821 & n27052 ) | ( ~n17811 & n27052 ) ;
  assign n27054 = n27053 ^ n7953 ^ 1'b0 ;
  assign n27055 = ( ~n4945 & n21503 ) | ( ~n4945 & n25288 ) | ( n21503 & n25288 ) ;
  assign n27056 = n1382 & ~n22569 ;
  assign n27057 = ( n4866 & n8466 ) | ( n4866 & n27056 ) | ( n8466 & n27056 ) ;
  assign n27058 = x49 & n8965 ;
  assign n27059 = ~n12321 & n27058 ;
  assign n27060 = n12877 & n13292 ;
  assign n27061 = ~n23500 & n27060 ;
  assign n27062 = n6409 & ~n22846 ;
  assign n27063 = n27062 ^ n325 ^ 1'b0 ;
  assign n27064 = n11996 ^ n7727 ^ 1'b0 ;
  assign n27065 = n17870 | n27064 ;
  assign n27066 = n27065 ^ n7848 ^ 1'b0 ;
  assign n27067 = n11409 | n27019 ;
  assign n27068 = ( n8031 & ~n21807 ) | ( n8031 & n24245 ) | ( ~n21807 & n24245 ) ;
  assign n27070 = n13195 ^ n4012 ^ n3888 ;
  assign n27071 = n20392 ^ n16535 ^ 1'b0 ;
  assign n27072 = n27070 & ~n27071 ;
  assign n27073 = n915 & n13008 ;
  assign n27074 = ~n27072 & n27073 ;
  assign n27069 = n1994 & n3581 ;
  assign n27075 = n27074 ^ n27069 ^ 1'b0 ;
  assign n27077 = n4498 ^ n2323 ^ n2285 ;
  assign n27078 = ~n4926 & n27077 ;
  assign n27076 = ~n20713 & n22533 ;
  assign n27079 = n27078 ^ n27076 ^ 1'b0 ;
  assign n27080 = n3329 | n17468 ;
  assign n27081 = n9693 & ~n17449 ;
  assign n27082 = n27081 ^ n608 ^ 1'b0 ;
  assign n27083 = n27082 ^ n2904 ^ 1'b0 ;
  assign n27084 = n8056 | n27083 ;
  assign n27085 = n20209 ^ n3703 ^ n302 ;
  assign n27086 = n16291 & n27085 ;
  assign n27087 = n1839 & n27086 ;
  assign n27088 = ( n1728 & n2723 ) | ( n1728 & ~n24244 ) | ( n2723 & ~n24244 ) ;
  assign n27089 = n11872 ^ n8447 ^ n6121 ;
  assign n27090 = ( n3561 & n3806 ) | ( n3561 & ~n5317 ) | ( n3806 & ~n5317 ) ;
  assign n27091 = n21168 | n27090 ;
  assign n27092 = n27091 ^ n11770 ^ 1'b0 ;
  assign n27093 = ( n3807 & n4802 ) | ( n3807 & n19618 ) | ( n4802 & n19618 ) ;
  assign n27094 = n16652 & n19873 ;
  assign n27096 = ( ~n2209 & n4945 ) | ( ~n2209 & n14314 ) | ( n4945 & n14314 ) ;
  assign n27097 = n3766 ^ n509 ^ 1'b0 ;
  assign n27098 = n27096 & n27097 ;
  assign n27095 = n1854 & ~n2923 ;
  assign n27099 = n27098 ^ n27095 ^ 1'b0 ;
  assign n27101 = n5743 | n8558 ;
  assign n27100 = n11987 & n17495 ;
  assign n27102 = n27101 ^ n27100 ^ 1'b0 ;
  assign n27103 = n21288 | n22308 ;
  assign n27104 = n27103 ^ n10888 ^ 1'b0 ;
  assign n27106 = n6127 | n15106 ;
  assign n27107 = n281 & ~n27106 ;
  assign n27108 = n27107 ^ n17067 ^ 1'b0 ;
  assign n27105 = x89 & n10433 ;
  assign n27109 = n27108 ^ n27105 ^ 1'b0 ;
  assign n27110 = n10713 & n11805 ;
  assign n27111 = n8453 & n27110 ;
  assign n27112 = ( n9110 & ~n16243 ) | ( n9110 & n27111 ) | ( ~n16243 & n27111 ) ;
  assign n27113 = ( ~n247 & n6196 ) | ( ~n247 & n14311 ) | ( n6196 & n14311 ) ;
  assign n27114 = ( n10388 & ~n20700 ) | ( n10388 & n27113 ) | ( ~n20700 & n27113 ) ;
  assign n27115 = ~n3162 & n5257 ;
  assign n27116 = n27115 ^ n4387 ^ 1'b0 ;
  assign n27117 = ~n14709 & n27116 ;
  assign n27118 = x104 & ~n1596 ;
  assign n27119 = n27118 ^ n11868 ^ n4149 ;
  assign n27120 = n3832 & n27119 ;
  assign n27121 = ~n20411 & n24881 ;
  assign n27122 = n13552 & n27121 ;
  assign n27123 = n21242 & ~n25766 ;
  assign n27124 = n27123 ^ n5771 ^ 1'b0 ;
  assign n27125 = n4527 ^ n4321 ^ n234 ;
  assign n27126 = ( n12950 & n17982 ) | ( n12950 & ~n27125 ) | ( n17982 & ~n27125 ) ;
  assign n27127 = n13807 & n15319 ;
  assign n27128 = ~n1224 & n24440 ;
  assign n27129 = n27128 ^ n15291 ^ n7474 ;
  assign n27130 = ~n11949 & n14575 ;
  assign n27131 = n4919 ^ n1939 ^ 1'b0 ;
  assign n27132 = n13914 & n27131 ;
  assign n27133 = n22033 ^ n14143 ^ 1'b0 ;
  assign n27134 = n13434 | n27133 ;
  assign n27135 = n27134 ^ n19788 ^ 1'b0 ;
  assign n27136 = n14094 & n27135 ;
  assign n27138 = ~n3381 & n8869 ;
  assign n27139 = n4223 & n27138 ;
  assign n27137 = n2421 & n25238 ;
  assign n27140 = n27139 ^ n27137 ^ 1'b0 ;
  assign n27141 = n17780 ^ n2889 ^ 1'b0 ;
  assign n27142 = ~n15631 & n15821 ;
  assign n27143 = n27141 & n27142 ;
  assign n27144 = n1503 & ~n27143 ;
  assign n27146 = n12361 ^ n1396 ^ 1'b0 ;
  assign n27147 = n10972 | n27146 ;
  assign n27145 = n5513 | n18008 ;
  assign n27148 = n27147 ^ n27145 ^ n13248 ;
  assign n27149 = n2353 & n17641 ;
  assign n27150 = n6806 ^ n5517 ^ n2796 ;
  assign n27151 = ~n3723 & n27150 ;
  assign n27152 = x103 & ~n9472 ;
  assign n27153 = n3158 & n14393 ;
  assign n27154 = ~n7292 & n27153 ;
  assign n27155 = n3636 | n11748 ;
  assign n27156 = n18571 | n27155 ;
  assign n27157 = ~n15195 & n22942 ;
  assign n27158 = n27157 ^ n9175 ^ 1'b0 ;
  assign n27159 = n6632 ^ n5005 ^ 1'b0 ;
  assign n27160 = n27159 ^ n20192 ^ n210 ;
  assign n27161 = n27160 ^ n5475 ^ 1'b0 ;
  assign n27162 = n13512 & ~n27161 ;
  assign n27163 = n8468 & ~n20324 ;
  assign n27164 = ( n9675 & n16685 ) | ( n9675 & ~n27163 ) | ( n16685 & ~n27163 ) ;
  assign n27165 = n8007 & ~n8744 ;
  assign n27166 = n15614 & ~n27165 ;
  assign n27167 = n7200 ^ n7108 ^ 1'b0 ;
  assign n27168 = n8759 ^ n2323 ^ 1'b0 ;
  assign n27169 = n8446 | n27168 ;
  assign n27170 = n2598 & ~n6440 ;
  assign n27171 = ~n14314 & n27170 ;
  assign n27172 = n5490 & n7861 ;
  assign n27173 = n14528 & n27172 ;
  assign n27174 = ~n3716 & n10186 ;
  assign n27175 = n1723 & ~n9504 ;
  assign n27176 = n6851 ^ n3951 ^ 1'b0 ;
  assign n27177 = n27175 | n27176 ;
  assign n27178 = n5973 & n23943 ;
  assign n27179 = ~n12970 & n27178 ;
  assign n27180 = n6862 | n25529 ;
  assign n27181 = ~n3296 & n10066 ;
  assign n27182 = ~n20441 & n24363 ;
  assign n27183 = n16408 ^ n2737 ^ n690 ;
  assign n27184 = n27183 ^ n10212 ^ 1'b0 ;
  assign n27187 = n7949 & n8708 ;
  assign n27188 = n27187 ^ n8853 ^ 1'b0 ;
  assign n27189 = n11181 & ~n27188 ;
  assign n27190 = ~n11362 & n27189 ;
  assign n27191 = n19221 | n27190 ;
  assign n27185 = x56 & ~n8126 ;
  assign n27186 = ~n25666 & n27185 ;
  assign n27192 = n27191 ^ n27186 ^ 1'b0 ;
  assign n27193 = n24146 ^ n2542 ^ 1'b0 ;
  assign n27194 = n14755 & ~n27193 ;
  assign n27195 = n14240 & n25295 ;
  assign n27196 = n27195 ^ n4143 ^ 1'b0 ;
  assign n27197 = n11098 ^ n8741 ^ 1'b0 ;
  assign n27198 = n27196 | n27197 ;
  assign n27199 = ~n1563 & n7895 ;
  assign n27200 = n27199 ^ n11316 ^ 1'b0 ;
  assign n27201 = n27200 ^ n644 ^ 1'b0 ;
  assign n27202 = ( n17449 & ~n21564 ) | ( n17449 & n22918 ) | ( ~n21564 & n22918 ) ;
  assign n27203 = n18958 ^ n4717 ^ n3856 ;
  assign n27204 = n20054 & ~n27203 ;
  assign n27205 = n27204 ^ n15536 ^ 1'b0 ;
  assign n27206 = n9528 | n23610 ;
  assign n27207 = n27206 ^ n3293 ^ 1'b0 ;
  assign n27208 = ( n14251 & ~n24232 ) | ( n14251 & n27207 ) | ( ~n24232 & n27207 ) ;
  assign n27209 = n470 | n20343 ;
  assign n27210 = ( ~n1851 & n27208 ) | ( ~n1851 & n27209 ) | ( n27208 & n27209 ) ;
  assign n27211 = n24567 ^ n7641 ^ n4117 ;
  assign n27212 = n27211 ^ n3274 ^ 1'b0 ;
  assign n27213 = n7254 ^ n4994 ^ 1'b0 ;
  assign n27214 = n1184 & n27213 ;
  assign n27215 = n9316 & n27214 ;
  assign n27216 = n26521 ^ n18496 ^ n12062 ;
  assign n27217 = n1588 & ~n8848 ;
  assign n27218 = n27217 ^ n12564 ^ 1'b0 ;
  assign n27219 = n27216 & ~n27218 ;
  assign n27220 = n7762 ^ n881 ^ 1'b0 ;
  assign n27221 = ~n18735 & n19170 ;
  assign n27222 = n8253 & ~n21738 ;
  assign n27223 = n7950 ^ n7813 ^ 1'b0 ;
  assign n27224 = ~n11425 & n13128 ;
  assign n27225 = n27224 ^ n1733 ^ 1'b0 ;
  assign n27226 = ( n1280 & n27223 ) | ( n1280 & n27225 ) | ( n27223 & n27225 ) ;
  assign n27227 = ( ~n3279 & n5774 ) | ( ~n3279 & n17641 ) | ( n5774 & n17641 ) ;
  assign n27228 = n1362 | n27227 ;
  assign n27230 = n10576 ^ n1152 ^ 1'b0 ;
  assign n27231 = n8102 & ~n27230 ;
  assign n27232 = n27231 ^ n3908 ^ 1'b0 ;
  assign n27233 = n27232 ^ n24882 ^ n9153 ;
  assign n27229 = n2743 & ~n12386 ;
  assign n27234 = n27233 ^ n27229 ^ 1'b0 ;
  assign n27236 = n3472 & ~n15373 ;
  assign n27237 = ~n6424 & n27236 ;
  assign n27235 = n5599 & n12987 ;
  assign n27238 = n27237 ^ n27235 ^ 1'b0 ;
  assign n27239 = n27238 ^ n6741 ^ 1'b0 ;
  assign n27240 = n5163 ^ n2167 ^ 1'b0 ;
  assign n27241 = n10348 ^ x5 ^ 1'b0 ;
  assign n27242 = n27240 & n27241 ;
  assign n27243 = ~n4200 & n8634 ;
  assign n27244 = n27243 ^ n17557 ^ n15943 ;
  assign n27245 = n15254 ^ n10030 ^ 1'b0 ;
  assign n27246 = ( n4236 & ~n5940 ) | ( n4236 & n26642 ) | ( ~n5940 & n26642 ) ;
  assign n27247 = n21009 ^ n17791 ^ n16381 ;
  assign n27248 = n1365 & n25880 ;
  assign n27249 = n27248 ^ n12414 ^ 1'b0 ;
  assign n27250 = n26058 ^ n11232 ^ 1'b0 ;
  assign n27251 = n9432 ^ n2395 ^ 1'b0 ;
  assign n27252 = n27250 | n27251 ;
  assign n27253 = n2296 | n11391 ;
  assign n27254 = n27253 ^ n13188 ^ n2420 ;
  assign n27255 = n4351 ^ n1584 ^ 1'b0 ;
  assign n27256 = n9933 | n27255 ;
  assign n27257 = n27254 | n27256 ;
  assign n27258 = n19784 ^ n10021 ^ 1'b0 ;
  assign n27259 = n23709 & n27258 ;
  assign n27260 = n5483 & n13232 ;
  assign n27261 = n10536 & n27260 ;
  assign n27262 = n17233 & n17557 ;
  assign n27263 = n27262 ^ n9107 ^ 1'b0 ;
  assign n27264 = n7650 & n19728 ;
  assign n27265 = ~n27263 & n27264 ;
  assign n27266 = n25110 ^ n14778 ^ 1'b0 ;
  assign n27267 = n6342 & ~n27266 ;
  assign n27268 = n1373 | n17372 ;
  assign n27269 = n27267 | n27268 ;
  assign n27270 = n8805 & ~n15106 ;
  assign n27271 = n27270 ^ n11430 ^ n10532 ;
  assign n27272 = n16457 ^ n9251 ^ n4250 ;
  assign n27273 = n6890 | n25910 ;
  assign n27274 = n432 & n11074 ;
  assign n27275 = n18053 & n27274 ;
  assign n27277 = n5686 & ~n6347 ;
  assign n27278 = n27277 ^ n16622 ^ 1'b0 ;
  assign n27276 = n5742 & n5966 ;
  assign n27279 = n27278 ^ n27276 ^ 1'b0 ;
  assign n27280 = ~n4697 & n27279 ;
  assign n27281 = n27280 ^ n10155 ^ 1'b0 ;
  assign n27282 = n7337 & ~n11425 ;
  assign n27283 = n7023 & n27282 ;
  assign n27284 = n27283 ^ n13615 ^ 1'b0 ;
  assign n27285 = n3666 | n27284 ;
  assign n27286 = ~n1049 & n1829 ;
  assign n27287 = n27286 ^ n4995 ^ 1'b0 ;
  assign n27288 = n17450 ^ n7364 ^ n746 ;
  assign n27289 = n6507 ^ n5389 ^ 1'b0 ;
  assign n27290 = n12306 & ~n27289 ;
  assign n27291 = n12312 ^ n12208 ^ n6629 ;
  assign n27292 = n27290 & n27291 ;
  assign n27293 = n19084 ^ n16224 ^ n9835 ;
  assign n27294 = n6304 | n20555 ;
  assign n27295 = n1266 | n27294 ;
  assign n27296 = n9927 ^ n5583 ^ 1'b0 ;
  assign n27297 = n21874 & ~n27296 ;
  assign n27298 = n27297 ^ n23041 ^ 1'b0 ;
  assign n27299 = n27298 ^ n2276 ^ 1'b0 ;
  assign n27300 = ( n1994 & n27295 ) | ( n1994 & n27299 ) | ( n27295 & n27299 ) ;
  assign n27301 = n21457 ^ n14587 ^ 1'b0 ;
  assign n27302 = ( n6474 & n10706 ) | ( n6474 & n12638 ) | ( n10706 & n12638 ) ;
  assign n27303 = n775 & n13207 ;
  assign n27304 = ~n4224 & n27303 ;
  assign n27305 = ~n27302 & n27304 ;
  assign n27306 = n9478 ^ n5568 ^ n1996 ;
  assign n27307 = n27306 ^ n7975 ^ 1'b0 ;
  assign n27308 = n24008 ^ n15187 ^ 1'b0 ;
  assign n27309 = n18370 & ~n27308 ;
  assign n27310 = n22493 ^ n9013 ^ 1'b0 ;
  assign n27311 = n17994 ^ n14553 ^ 1'b0 ;
  assign n27312 = n3395 & n20112 ;
  assign n27313 = x93 & n24663 ;
  assign n27314 = n11432 & n27313 ;
  assign n27315 = ~n4917 & n27314 ;
  assign n27316 = n27315 ^ n3777 ^ 1'b0 ;
  assign n27317 = n8721 & ~n17051 ;
  assign n27318 = ( ~n3106 & n22026 ) | ( ~n3106 & n27317 ) | ( n22026 & n27317 ) ;
  assign n27319 = ~n4075 & n7932 ;
  assign n27320 = n3621 & n27319 ;
  assign n27321 = ~n23394 & n27320 ;
  assign n27322 = n10912 ^ n9234 ^ 1'b0 ;
  assign n27323 = n13188 | n15491 ;
  assign n27324 = n21729 | n27323 ;
  assign n27325 = n27324 ^ n3284 ^ 1'b0 ;
  assign n27326 = n18980 & ~n27325 ;
  assign n27327 = n27326 ^ n15360 ^ 1'b0 ;
  assign n27328 = ~n7051 & n9748 ;
  assign n27329 = n27328 ^ n12100 ^ 1'b0 ;
  assign n27330 = n15889 | n18771 ;
  assign n27331 = n27330 ^ n9638 ^ 1'b0 ;
  assign n27332 = ~n15237 & n23491 ;
  assign n27333 = n27332 ^ n21864 ^ 1'b0 ;
  assign n27334 = n5202 ^ n4665 ^ 1'b0 ;
  assign n27335 = n27334 ^ n27082 ^ n6274 ;
  assign n27336 = n18588 | n27335 ;
  assign n27337 = ( n7116 & n17587 ) | ( n7116 & n25411 ) | ( n17587 & n25411 ) ;
  assign n27338 = ( n6537 & ~n8601 ) | ( n6537 & n23354 ) | ( ~n8601 & n23354 ) ;
  assign n27339 = n11333 ^ n11136 ^ n9546 ;
  assign n27340 = n8660 & ~n27339 ;
  assign n27341 = n2665 & n27340 ;
  assign n27342 = n9406 & ~n21891 ;
  assign n27343 = n27342 ^ n7091 ^ 1'b0 ;
  assign n27344 = n14914 ^ n302 ^ 1'b0 ;
  assign n27345 = n3393 | n27344 ;
  assign n27346 = n13153 ^ n5168 ^ n3851 ;
  assign n27347 = n27346 ^ n19702 ^ 1'b0 ;
  assign n27348 = n8146 ^ n5438 ^ 1'b0 ;
  assign n27349 = ~n20667 & n27348 ;
  assign n27350 = n7675 | n20457 ;
  assign n27351 = n788 & n27350 ;
  assign n27352 = n20683 & n27351 ;
  assign n27353 = n7104 ^ n2075 ^ n154 ;
  assign n27354 = n25905 ^ n25687 ^ n1131 ;
  assign n27355 = ~n608 & n2855 ;
  assign n27356 = n11806 & n27355 ;
  assign n27357 = ( ~n14570 & n25880 ) | ( ~n14570 & n27356 ) | ( n25880 & n27356 ) ;
  assign n27358 = ( n7307 & n20745 ) | ( n7307 & n27357 ) | ( n20745 & n27357 ) ;
  assign n27359 = n7723 ^ n358 ^ 1'b0 ;
  assign n27360 = n5139 | n27359 ;
  assign n27361 = n12981 & n27360 ;
  assign n27362 = n15445 ^ n2000 ^ 1'b0 ;
  assign n27363 = n5163 ^ n2423 ^ 1'b0 ;
  assign n27364 = n12478 ^ n6326 ^ 1'b0 ;
  assign n27365 = n27363 & ~n27364 ;
  assign n27366 = n9606 | n13626 ;
  assign n27367 = n27366 ^ n1271 ^ 1'b0 ;
  assign n27368 = n354 & n4610 ;
  assign n27369 = n3852 & n27368 ;
  assign n27370 = x13 & ~n12995 ;
  assign n27371 = n27370 ^ n22852 ^ 1'b0 ;
  assign n27372 = n26270 & n27371 ;
  assign n27373 = n16384 ^ n15469 ^ n13488 ;
  assign n27374 = ~n2879 & n4217 ;
  assign n27375 = n22659 & n27374 ;
  assign n27376 = n23812 ^ n6594 ^ 1'b0 ;
  assign n27377 = n15632 ^ n6365 ^ 1'b0 ;
  assign n27378 = ( n7700 & ~n7780 ) | ( n7700 & n9464 ) | ( ~n7780 & n9464 ) ;
  assign n27379 = ~n11308 & n24889 ;
  assign n27380 = n27379 ^ n14196 ^ 1'b0 ;
  assign n27381 = ( n358 & ~n746 ) | ( n358 & n8708 ) | ( ~n746 & n8708 ) ;
  assign n27382 = ~n3144 & n27381 ;
  assign n27383 = n12849 ^ n8814 ^ n2921 ;
  assign n27384 = n2992 & n6750 ;
  assign n27385 = n20075 | n27384 ;
  assign n27386 = n27383 | n27385 ;
  assign n27387 = n1310 | n18319 ;
  assign n27388 = n23171 & ~n27387 ;
  assign n27389 = ( n12109 & ~n24469 ) | ( n12109 & n27139 ) | ( ~n24469 & n27139 ) ;
  assign n27390 = n5088 & ~n12862 ;
  assign n27392 = n14321 | n20970 ;
  assign n27391 = n24479 ^ n3514 ^ 1'b0 ;
  assign n27393 = n27392 ^ n27391 ^ n6382 ;
  assign n27394 = ( n20360 & n27390 ) | ( n20360 & n27393 ) | ( n27390 & n27393 ) ;
  assign n27395 = n11553 ^ n9656 ^ n1186 ;
  assign n27396 = ~n8738 & n14148 ;
  assign n27397 = n24994 ^ n10967 ^ n5378 ;
  assign n27398 = ~n7158 & n27397 ;
  assign n27399 = n15580 | n17745 ;
  assign n27400 = ~n8049 & n12859 ;
  assign n27401 = n27400 ^ n9573 ^ 1'b0 ;
  assign n27402 = n27401 ^ n5548 ^ 1'b0 ;
  assign n27403 = n17209 ^ n13729 ^ n965 ;
  assign n27404 = n11416 ^ n7004 ^ 1'b0 ;
  assign n27405 = n15242 & n18599 ;
  assign n27406 = n27405 ^ n13004 ^ 1'b0 ;
  assign n27407 = n27406 ^ n2173 ^ 1'b0 ;
  assign n27408 = n5868 & ~n19392 ;
  assign n27409 = n15927 & ~n16241 ;
  assign n27410 = n469 & ~n25060 ;
  assign n27411 = n11274 ^ n10575 ^ 1'b0 ;
  assign n27412 = n7824 ^ n3827 ^ 1'b0 ;
  assign n27413 = n2038 & ~n27412 ;
  assign n27414 = n11539 | n18288 ;
  assign n27415 = n3180 & ~n27414 ;
  assign n27416 = ( n4776 & ~n14495 ) | ( n4776 & n19405 ) | ( ~n14495 & n19405 ) ;
  assign n27417 = ( n14697 & ~n18925 ) | ( n14697 & n27416 ) | ( ~n18925 & n27416 ) ;
  assign n27418 = ( n2874 & n17091 ) | ( n2874 & n17144 ) | ( n17091 & n17144 ) ;
  assign n27419 = n2251 & n14066 ;
  assign n27420 = n27419 ^ n10271 ^ 1'b0 ;
  assign n27421 = n4123 | n27420 ;
  assign n27422 = n3726 & n11210 ;
  assign n27423 = n6913 & ~n17310 ;
  assign n27424 = n27423 ^ n20801 ^ 1'b0 ;
  assign n27425 = n5185 & n12314 ;
  assign n27426 = n20250 ^ n15884 ^ 1'b0 ;
  assign n27427 = ~n19198 & n23775 ;
  assign n27428 = n27427 ^ n1150 ^ 1'b0 ;
  assign n27429 = n11887 | n27428 ;
  assign n27430 = ~n1770 & n5838 ;
  assign n27431 = n27430 ^ n15073 ^ 1'b0 ;
  assign n27432 = ~n14100 & n27431 ;
  assign n27433 = n27432 ^ n10663 ^ 1'b0 ;
  assign n27434 = ( ~n17536 & n17843 ) | ( ~n17536 & n22524 ) | ( n17843 & n22524 ) ;
  assign n27435 = n27433 | n27434 ;
  assign n27436 = ( n18369 & n27429 ) | ( n18369 & ~n27435 ) | ( n27429 & ~n27435 ) ;
  assign n27437 = ( n5149 & n13901 ) | ( n5149 & n20643 ) | ( n13901 & n20643 ) ;
  assign n27438 = n432 | n12306 ;
  assign n27439 = ( n8129 & ~n23487 ) | ( n8129 & n27438 ) | ( ~n23487 & n27438 ) ;
  assign n27440 = n6083 & n18592 ;
  assign n27441 = n23938 & n27440 ;
  assign n27442 = n20026 ^ n2186 ^ 1'b0 ;
  assign n27443 = n1049 | n27442 ;
  assign n27444 = n14317 | n26281 ;
  assign n27445 = ( n3382 & n3634 ) | ( n3382 & ~n11757 ) | ( n3634 & ~n11757 ) ;
  assign n27446 = n7032 | n22795 ;
  assign n27447 = n27445 & ~n27446 ;
  assign n27448 = n23570 ^ n11875 ^ n9201 ;
  assign n27449 = n27448 ^ n22106 ^ n18139 ;
  assign n27450 = ~n15878 & n27449 ;
  assign n27451 = n3461 & n19376 ;
  assign n27452 = n27451 ^ n5767 ^ n1653 ;
  assign n27453 = ( n11485 & ~n20341 ) | ( n11485 & n27452 ) | ( ~n20341 & n27452 ) ;
  assign n27454 = n10344 ^ n870 ^ 1'b0 ;
  assign n27455 = ~n5089 & n27454 ;
  assign n27456 = n27455 ^ n22667 ^ 1'b0 ;
  assign n27457 = ~n14280 & n16299 ;
  assign n27458 = n27457 ^ n10489 ^ 1'b0 ;
  assign n27459 = n15162 | n23660 ;
  assign n27460 = n21359 ^ n5453 ^ 1'b0 ;
  assign n27461 = n25012 & ~n27460 ;
  assign n27462 = n26659 & n27461 ;
  assign n27463 = n27462 ^ n9192 ^ 1'b0 ;
  assign n27465 = n16217 & n22344 ;
  assign n27466 = n6935 & n27465 ;
  assign n27464 = ~n11165 & n21089 ;
  assign n27467 = n27466 ^ n27464 ^ 1'b0 ;
  assign n27468 = ( ~n735 & n4180 ) | ( ~n735 & n27467 ) | ( n4180 & n27467 ) ;
  assign n27469 = n27468 ^ n10962 ^ 1'b0 ;
  assign n27471 = ~n4279 & n7060 ;
  assign n27472 = n5045 & n27471 ;
  assign n27470 = n10362 & ~n16482 ;
  assign n27473 = n27472 ^ n27470 ^ 1'b0 ;
  assign n27474 = n9303 | n11755 ;
  assign n27475 = n6966 | n9197 ;
  assign n27476 = ( ~n270 & n4020 ) | ( ~n270 & n7839 ) | ( n4020 & n7839 ) ;
  assign n27477 = ( n16884 & n27475 ) | ( n16884 & ~n27476 ) | ( n27475 & ~n27476 ) ;
  assign n27478 = n3809 & n3988 ;
  assign n27479 = n16687 ^ n892 ^ 1'b0 ;
  assign n27480 = n9651 ^ n8079 ^ n325 ;
  assign n27481 = n27480 ^ n22375 ^ n2189 ;
  assign n27482 = ~n2989 & n27481 ;
  assign n27483 = n9846 ^ n4478 ^ n4428 ;
  assign n27484 = n15246 ^ n15195 ^ 1'b0 ;
  assign n27485 = n27483 | n27484 ;
  assign n27486 = n1307 & ~n27485 ;
  assign n27487 = n3478 & n27486 ;
  assign n27488 = ~n12619 & n16685 ;
  assign n27489 = n6317 & n27488 ;
  assign n27490 = n1660 & n19001 ;
  assign n27491 = n5238 & n27490 ;
  assign n27492 = n15059 ^ n2452 ^ 1'b0 ;
  assign n27493 = n27492 ^ n19481 ^ 1'b0 ;
  assign n27494 = n27491 & ~n27493 ;
  assign n27495 = ( n3438 & n14087 ) | ( n3438 & ~n27494 ) | ( n14087 & ~n27494 ) ;
  assign n27496 = n13853 ^ n9255 ^ 1'b0 ;
  assign n27497 = n23349 ^ n16028 ^ n6412 ;
  assign n27498 = n12151 ^ n802 ^ 1'b0 ;
  assign n27499 = n27498 ^ n17965 ^ n11934 ;
  assign n27500 = n11428 ^ n6232 ^ 1'b0 ;
  assign n27501 = n13732 ^ n6228 ^ 1'b0 ;
  assign n27502 = n2331 ^ n148 ^ 1'b0 ;
  assign n27503 = n27501 & n27502 ;
  assign n27504 = n15125 ^ n9049 ^ 1'b0 ;
  assign n27505 = n796 & ~n6761 ;
  assign n27506 = ~n27504 & n27505 ;
  assign n27507 = ~n6043 & n16344 ;
  assign n27508 = ~n5137 & n27507 ;
  assign n27509 = n17009 & ~n27508 ;
  assign n27510 = ~n2839 & n11823 ;
  assign n27511 = n18051 ^ n5574 ^ n3195 ;
  assign n27512 = n27510 & n27511 ;
  assign n27513 = n27512 ^ n7233 ^ 1'b0 ;
  assign n27514 = ( n5609 & ~n24551 ) | ( n5609 & n27513 ) | ( ~n24551 & n27513 ) ;
  assign n27515 = n27514 ^ n5327 ^ 1'b0 ;
  assign n27516 = n8773 ^ n740 ^ x10 ;
  assign n27517 = ~n23918 & n23997 ;
  assign n27518 = n7571 ^ n1138 ^ 1'b0 ;
  assign n27519 = ~n27517 & n27518 ;
  assign n27520 = ( n7718 & ~n16948 ) | ( n7718 & n27519 ) | ( ~n16948 & n27519 ) ;
  assign n27521 = n11695 ^ n4186 ^ n892 ;
  assign n27522 = n10745 & n12221 ;
  assign n27523 = n27522 ^ n3923 ^ 1'b0 ;
  assign n27524 = ~n3320 & n24479 ;
  assign n27525 = n26200 & n27524 ;
  assign n27526 = ( ~n1257 & n7482 ) | ( ~n1257 & n17127 ) | ( n7482 & n17127 ) ;
  assign n27527 = n27526 ^ n22790 ^ 1'b0 ;
  assign n27528 = ~n4964 & n14417 ;
  assign n27529 = ~n27527 & n27528 ;
  assign n27530 = ~n6896 & n7774 ;
  assign n27531 = n23704 ^ n4227 ^ 1'b0 ;
  assign n27532 = n10652 & n15551 ;
  assign n27533 = ( n6838 & n20216 ) | ( n6838 & n20926 ) | ( n20216 & n20926 ) ;
  assign n27537 = n19682 ^ n9956 ^ n8826 ;
  assign n27534 = n9497 & n9527 ;
  assign n27535 = ( n2460 & n7108 ) | ( n2460 & ~n27534 ) | ( n7108 & ~n27534 ) ;
  assign n27536 = ( ~n637 & n13677 ) | ( ~n637 & n27535 ) | ( n13677 & n27535 ) ;
  assign n27538 = n27537 ^ n27536 ^ n25716 ;
  assign n27539 = n15779 ^ n221 ^ 1'b0 ;
  assign n27540 = n3961 & n12577 ;
  assign n27541 = n27540 ^ n10061 ^ 1'b0 ;
  assign n27542 = ~n2844 & n12644 ;
  assign n27543 = n11037 & n27542 ;
  assign n27544 = n9259 | n27543 ;
  assign n27545 = n27544 ^ n4170 ^ 1'b0 ;
  assign n27547 = n1586 | n7931 ;
  assign n27546 = ~n4495 & n19943 ;
  assign n27548 = n27547 ^ n27546 ^ n21537 ;
  assign n27549 = n13318 ^ n7775 ^ 1'b0 ;
  assign n27550 = ( n1113 & n9555 ) | ( n1113 & ~n27549 ) | ( n9555 & ~n27549 ) ;
  assign n27551 = ( n933 & n5788 ) | ( n933 & n11946 ) | ( n5788 & n11946 ) ;
  assign n27552 = n10304 ^ n3090 ^ n960 ;
  assign n27553 = ( n11236 & n27551 ) | ( n11236 & ~n27552 ) | ( n27551 & ~n27552 ) ;
  assign n27555 = ( n2796 & n3584 ) | ( n2796 & n14769 ) | ( n3584 & n14769 ) ;
  assign n27554 = n8096 & n10826 ;
  assign n27556 = n27555 ^ n27554 ^ 1'b0 ;
  assign n27557 = n27556 ^ n1300 ^ 1'b0 ;
  assign n27558 = ~n2462 & n10032 ;
  assign n27559 = n20966 & n27558 ;
  assign n27560 = n14094 ^ n13821 ^ n4069 ;
  assign n27561 = n27559 | n27560 ;
  assign n27562 = n25627 ^ n18540 ^ n9795 ;
  assign n27563 = n14698 & ~n17388 ;
  assign n27564 = n27562 & n27563 ;
  assign n27565 = ~n6290 & n21175 ;
  assign n27566 = ~n3829 & n27565 ;
  assign n27567 = n8527 ^ x11 ^ 1'b0 ;
  assign n27568 = n4255 | n27567 ;
  assign n27569 = n2248 | n12440 ;
  assign n27570 = n23288 ^ n5090 ^ 1'b0 ;
  assign n27571 = n27569 | n27570 ;
  assign n27572 = n8453 ^ n5855 ^ n3088 ;
  assign n27575 = ~n593 & n9483 ;
  assign n27576 = n27575 ^ n4798 ^ 1'b0 ;
  assign n27573 = n21874 ^ n13684 ^ 1'b0 ;
  assign n27574 = n641 | n27573 ;
  assign n27577 = n27576 ^ n27574 ^ 1'b0 ;
  assign n27578 = n2609 & n9593 ;
  assign n27579 = n27578 ^ n12120 ^ 1'b0 ;
  assign n27580 = n7034 & ~n8982 ;
  assign n27581 = n27580 ^ n11478 ^ 1'b0 ;
  assign n27582 = n27581 ^ n2717 ^ 1'b0 ;
  assign n27583 = n13699 & n27582 ;
  assign n27584 = n24163 ^ n6505 ^ 1'b0 ;
  assign n27585 = n3049 & ~n27584 ;
  assign n27586 = ~n6905 & n9193 ;
  assign n27587 = n27586 ^ n1994 ^ 1'b0 ;
  assign n27588 = ( ~n6946 & n25452 ) | ( ~n6946 & n26579 ) | ( n25452 & n26579 ) ;
  assign n27589 = n19947 & ~n21937 ;
  assign n27590 = ~n12464 & n27589 ;
  assign n27591 = n2440 & n27590 ;
  assign n27592 = n2937 | n10100 ;
  assign n27593 = ~n10958 & n16790 ;
  assign n27594 = n4983 & n27593 ;
  assign n27595 = ~n15611 & n27594 ;
  assign n27596 = n27595 ^ n1431 ^ 1'b0 ;
  assign n27597 = ~n27592 & n27596 ;
  assign n27598 = n7788 | n23495 ;
  assign n27599 = n820 & ~n27598 ;
  assign n27600 = n21884 ^ n5246 ^ 1'b0 ;
  assign n27601 = n11269 & ~n27600 ;
  assign n27602 = n6640 ^ n1863 ^ 1'b0 ;
  assign n27603 = n3824 & n4378 ;
  assign n27604 = ~n6233 & n27603 ;
  assign n27605 = n6203 & ~n27604 ;
  assign n27606 = ~n27602 & n27605 ;
  assign n27607 = n9059 ^ n6867 ^ 1'b0 ;
  assign n27608 = n13814 ^ n13085 ^ 1'b0 ;
  assign n27609 = n389 & n10864 ;
  assign n27610 = ~n1648 & n27609 ;
  assign n27611 = n3334 & ~n27610 ;
  assign n27612 = n27611 ^ n1795 ^ 1'b0 ;
  assign n27613 = n27612 ^ n9729 ^ 1'b0 ;
  assign n27614 = ~n27608 & n27613 ;
  assign n27615 = n1199 | n16621 ;
  assign n27616 = n1441 & ~n8188 ;
  assign n27617 = n27616 ^ n2321 ^ 1'b0 ;
  assign n27618 = n9150 ^ n2303 ^ 1'b0 ;
  assign n27619 = ~n27617 & n27618 ;
  assign n27620 = n27619 ^ n25102 ^ n4911 ;
  assign n27621 = n24574 ^ n7439 ^ 1'b0 ;
  assign n27622 = n979 | n12297 ;
  assign n27623 = ~n6036 & n10468 ;
  assign n27624 = n27623 ^ n7868 ^ 1'b0 ;
  assign n27630 = ( n6456 & n19224 ) | ( n6456 & ~n27255 ) | ( n19224 & ~n27255 ) ;
  assign n27625 = ~n6999 & n22037 ;
  assign n27626 = n27625 ^ n2189 ^ 1'b0 ;
  assign n27627 = x29 & n3894 ;
  assign n27628 = n27626 & n27627 ;
  assign n27629 = n21359 | n27628 ;
  assign n27631 = n27630 ^ n27629 ^ 1'b0 ;
  assign n27633 = n726 & ~n3997 ;
  assign n27634 = n27633 ^ n7624 ^ n5246 ;
  assign n27632 = ~n1820 & n9379 ;
  assign n27635 = n27634 ^ n27632 ^ 1'b0 ;
  assign n27636 = ( n1924 & ~n5262 ) | ( n1924 & n15044 ) | ( ~n5262 & n15044 ) ;
  assign n27637 = n27636 ^ n1489 ^ 1'b0 ;
  assign n27640 = n5201 & n5804 ;
  assign n27638 = n13273 ^ n7297 ^ n4119 ;
  assign n27639 = n1761 & ~n27638 ;
  assign n27641 = n27640 ^ n27639 ^ n11435 ;
  assign n27642 = n18812 & n27641 ;
  assign n27643 = n2290 & n27642 ;
  assign n27644 = n9492 ^ n9306 ^ 1'b0 ;
  assign n27645 = ( n980 & n4511 ) | ( n980 & ~n7514 ) | ( n4511 & ~n7514 ) ;
  assign n27646 = n12799 ^ n10420 ^ n800 ;
  assign n27647 = ( n22201 & n26445 ) | ( n22201 & ~n27646 ) | ( n26445 & ~n27646 ) ;
  assign n27648 = n2726 & ~n3359 ;
  assign n27649 = n850 | n1779 ;
  assign n27650 = n18512 & n27649 ;
  assign n27651 = n4113 & ~n27650 ;
  assign n27652 = n7021 & ~n9542 ;
  assign n27653 = n27652 ^ n21224 ^ 1'b0 ;
  assign n27654 = ( ~n1995 & n7612 ) | ( ~n1995 & n22114 ) | ( n7612 & n22114 ) ;
  assign n27655 = n14332 ^ n9903 ^ 1'b0 ;
  assign n27656 = n7232 & ~n27655 ;
  assign n27657 = n27656 ^ n3312 ^ 1'b0 ;
  assign n27658 = ~n27654 & n27657 ;
  assign n27659 = n16117 ^ n7189 ^ 1'b0 ;
  assign n27660 = n21064 | n27659 ;
  assign n27661 = n9431 & ~n27660 ;
  assign n27662 = n27661 ^ n18688 ^ 1'b0 ;
  assign n27663 = n17033 ^ n13449 ^ 1'b0 ;
  assign n27664 = n1505 & ~n27663 ;
  assign n27665 = n18219 ^ n3902 ^ 1'b0 ;
  assign n27666 = n27665 ^ n11772 ^ n9682 ;
  assign n27667 = n13502 & n18484 ;
  assign n27668 = ~n5257 & n27667 ;
  assign n27669 = n8757 & ~n13302 ;
  assign n27670 = ~n8689 & n27669 ;
  assign n27671 = n27670 ^ n23305 ^ 1'b0 ;
  assign n27672 = n13819 & n14541 ;
  assign n27673 = n26126 ^ n1062 ^ 1'b0 ;
  assign n27674 = n6339 | n27673 ;
  assign n27675 = n27674 ^ n19270 ^ 1'b0 ;
  assign n27676 = n10045 & ~n18427 ;
  assign n27677 = ~n8680 & n27676 ;
  assign n27678 = n4569 ^ n3600 ^ 1'b0 ;
  assign n27679 = n4978 & ~n8952 ;
  assign n27680 = n27679 ^ n10729 ^ 1'b0 ;
  assign n27681 = n8097 & ~n8799 ;
  assign n27682 = n27681 ^ n2449 ^ 1'b0 ;
  assign n27683 = ( ~n10699 & n15779 ) | ( ~n10699 & n18161 ) | ( n15779 & n18161 ) ;
  assign n27684 = ~n12396 & n24932 ;
  assign n27685 = n14534 | n27684 ;
  assign n27686 = n9668 ^ n6623 ^ 1'b0 ;
  assign n27687 = ~n2772 & n27686 ;
  assign n27688 = n27078 ^ n18580 ^ n5821 ;
  assign n27689 = n27688 ^ n10492 ^ n6220 ;
  assign n27690 = ~n5676 & n25807 ;
  assign n27691 = n1858 ^ n1518 ^ 1'b0 ;
  assign n27692 = n3227 | n27691 ;
  assign n27693 = n14387 | n26620 ;
  assign n27694 = n1740 & n10630 ;
  assign n27695 = ( n2161 & n5193 ) | ( n2161 & n5955 ) | ( n5193 & n5955 ) ;
  assign n27699 = n8079 ^ n1874 ^ 1'b0 ;
  assign n27700 = n10010 & ~n27699 ;
  assign n27696 = n1481 | n4068 ;
  assign n27697 = n27696 ^ n2849 ^ 1'b0 ;
  assign n27698 = n5229 & n27697 ;
  assign n27701 = n27700 ^ n27698 ^ 1'b0 ;
  assign n27702 = ~n21105 & n27070 ;
  assign n27703 = n2926 | n5613 ;
  assign n27704 = n1733 & n27703 ;
  assign n27705 = n27704 ^ n21402 ^ n15995 ;
  assign n27706 = n13042 ^ n2307 ^ 1'b0 ;
  assign n27707 = n9749 | n19287 ;
  assign n27708 = n27707 ^ n15683 ^ 1'b0 ;
  assign n27709 = n5589 | n20444 ;
  assign n27710 = n4235 | n27709 ;
  assign n27711 = n14416 ^ n3227 ^ 1'b0 ;
  assign n27712 = ~n4265 & n6907 ;
  assign n27713 = n5759 & ~n23262 ;
  assign n27714 = ~n27712 & n27713 ;
  assign n27715 = n9512 | n27714 ;
  assign n27716 = n27715 ^ n1195 ^ 1'b0 ;
  assign n27717 = n1848 ^ n876 ^ n708 ;
  assign n27718 = n21057 & n27717 ;
  assign n27719 = ( n9349 & n9845 ) | ( n9349 & n26480 ) | ( n9845 & n26480 ) ;
  assign n27720 = n5828 & ~n10875 ;
  assign n27721 = n27720 ^ n9736 ^ 1'b0 ;
  assign n27722 = ( ~n9646 & n15193 ) | ( ~n9646 & n27721 ) | ( n15193 & n27721 ) ;
  assign n27727 = ~n1374 & n8425 ;
  assign n27728 = n27727 ^ n7822 ^ 1'b0 ;
  assign n27724 = n293 & n1915 ;
  assign n27725 = n27724 ^ n2992 ^ 1'b0 ;
  assign n27726 = n27725 ^ n15036 ^ n13242 ;
  assign n27729 = n27728 ^ n27726 ^ n3289 ;
  assign n27723 = ~n8374 & n21577 ;
  assign n27730 = n27729 ^ n27723 ^ 1'b0 ;
  assign n27731 = ( n8702 & ~n15762 ) | ( n8702 & n20939 ) | ( ~n15762 & n20939 ) ;
  assign n27732 = n11433 & ~n13752 ;
  assign n27733 = n27732 ^ n20128 ^ 1'b0 ;
  assign n27734 = n10338 ^ n10222 ^ 1'b0 ;
  assign n27735 = n22160 | n27734 ;
  assign n27736 = n2743 & ~n12454 ;
  assign n27737 = ~n8078 & n27736 ;
  assign n27738 = ~n4489 & n27737 ;
  assign n27739 = ~n6651 & n14845 ;
  assign n27740 = n3538 & n27739 ;
  assign n27741 = n8240 | n23616 ;
  assign n27742 = n19778 & ~n27741 ;
  assign n27744 = n20706 ^ n13002 ^ n4813 ;
  assign n27743 = n12377 & n17628 ;
  assign n27745 = n27744 ^ n27743 ^ n1709 ;
  assign n27746 = n3828 & ~n20208 ;
  assign n27747 = n25627 | n27746 ;
  assign n27748 = n3361 | n27747 ;
  assign n27749 = n6166 | n27748 ;
  assign n27750 = n14737 ^ n13832 ^ n7253 ;
  assign n27751 = n16190 | n27750 ;
  assign n27752 = n14290 | n27751 ;
  assign n27753 = ~n9084 & n9598 ;
  assign n27754 = ~n20665 & n27753 ;
  assign n27755 = n7497 ^ n4954 ^ 1'b0 ;
  assign n27756 = ( n3866 & ~n27754 ) | ( n3866 & n27755 ) | ( ~n27754 & n27755 ) ;
  assign n27757 = n16247 | n24341 ;
  assign n27758 = n7451 | n7462 ;
  assign n27759 = n24618 & ~n27758 ;
  assign n27760 = n6201 ^ n3726 ^ 1'b0 ;
  assign n27761 = ~n12529 & n27760 ;
  assign n27762 = ~n1555 & n1787 ;
  assign n27763 = n27762 ^ n3756 ^ 1'b0 ;
  assign n27764 = n7540 | n27763 ;
  assign n27765 = ( n12699 & n14541 ) | ( n12699 & n20548 ) | ( n14541 & n20548 ) ;
  assign n27766 = n16539 ^ n15869 ^ 1'b0 ;
  assign n27767 = n5335 & n12277 ;
  assign n27768 = n3521 ^ x3 ^ 1'b0 ;
  assign n27769 = ~n22569 & n27768 ;
  assign n27770 = n14143 & n27769 ;
  assign n27771 = ~n16213 & n20100 ;
  assign n27772 = ~n1971 & n27771 ;
  assign n27773 = n7011 & n21240 ;
  assign n27774 = n26542 | n27318 ;
  assign n27775 = n27774 ^ n21198 ^ 1'b0 ;
  assign n27776 = n19347 ^ n10756 ^ 1'b0 ;
  assign n27777 = n7514 & n27776 ;
  assign n27778 = n2528 & n20354 ;
  assign n27779 = n8708 & ~n10340 ;
  assign n27780 = n11790 & n27779 ;
  assign n27781 = n27780 ^ n12809 ^ n9679 ;
  assign n27782 = ~n2231 & n2470 ;
  assign n27783 = ( n3871 & ~n5139 ) | ( n3871 & n27782 ) | ( ~n5139 & n27782 ) ;
  assign n27784 = ( n8395 & ~n15248 ) | ( n8395 & n24199 ) | ( ~n15248 & n24199 ) ;
  assign n27785 = n17129 & ~n20817 ;
  assign n27786 = n27785 ^ n11406 ^ 1'b0 ;
  assign n27787 = ( n4104 & n4757 ) | ( n4104 & n7063 ) | ( n4757 & n7063 ) ;
  assign n27788 = ( n362 & ~n8255 ) | ( n362 & n27787 ) | ( ~n8255 & n27787 ) ;
  assign n27789 = n27788 ^ n22401 ^ 1'b0 ;
  assign n27790 = n15468 ^ n1899 ^ 1'b0 ;
  assign n27791 = ~n7412 & n12965 ;
  assign n27792 = n27791 ^ n6346 ^ 1'b0 ;
  assign n27793 = n25428 & n25830 ;
  assign n27794 = ~n4761 & n27793 ;
  assign n27795 = n19688 | n25893 ;
  assign n27796 = n4632 | n27795 ;
  assign n27797 = n1554 & ~n7706 ;
  assign n27798 = ( ~n1531 & n11791 ) | ( ~n1531 & n27508 ) | ( n11791 & n27508 ) ;
  assign n27799 = ( ~n5953 & n27691 ) | ( ~n5953 & n27798 ) | ( n27691 & n27798 ) ;
  assign n27800 = n4472 ^ x22 ^ 1'b0 ;
  assign n27801 = n20239 ^ n3045 ^ 1'b0 ;
  assign n27802 = ~n173 & n824 ;
  assign n27803 = ~n2038 & n27802 ;
  assign n27804 = ~n9064 & n27803 ;
  assign n27805 = n27804 ^ n22253 ^ n5357 ;
  assign n27806 = ~n4510 & n10076 ;
  assign n27807 = ~n10076 & n27806 ;
  assign n27808 = n19396 ^ n17311 ^ 1'b0 ;
  assign n27809 = ~n27807 & n27808 ;
  assign n27810 = n8560 ^ n2308 ^ 1'b0 ;
  assign n27811 = n22093 ^ n12307 ^ 1'b0 ;
  assign n27812 = ( ~n8891 & n13148 ) | ( ~n8891 & n19596 ) | ( n13148 & n19596 ) ;
  assign n27813 = ( n5616 & n11136 ) | ( n5616 & n20454 ) | ( n11136 & n20454 ) ;
  assign n27814 = n12923 ^ n7821 ^ 1'b0 ;
  assign n27815 = n7522 | n27594 ;
  assign n27816 = n27815 ^ n6318 ^ 1'b0 ;
  assign n27817 = ~n704 & n1850 ;
  assign n27818 = n27817 ^ n10169 ^ 1'b0 ;
  assign n27819 = n27818 ^ n12061 ^ 1'b0 ;
  assign n27820 = n3063 & n27819 ;
  assign n27821 = ( n2258 & n27816 ) | ( n2258 & ~n27820 ) | ( n27816 & ~n27820 ) ;
  assign n27825 = n7368 ^ n6581 ^ 1'b0 ;
  assign n27826 = ~n20235 & n27825 ;
  assign n27822 = n9875 ^ n5103 ^ 1'b0 ;
  assign n27823 = n8144 & ~n27822 ;
  assign n27824 = n2836 & n27823 ;
  assign n27827 = n27826 ^ n27824 ^ 1'b0 ;
  assign n27828 = n17480 & ~n22464 ;
  assign n27829 = ~n10771 & n27828 ;
  assign n27830 = n10468 & ~n11004 ;
  assign n27831 = n11625 & n27830 ;
  assign n27832 = n4546 | n21200 ;
  assign n27833 = n27832 ^ n14347 ^ 1'b0 ;
  assign n27834 = ( n7182 & n9685 ) | ( n7182 & n19005 ) | ( n9685 & n19005 ) ;
  assign n27835 = n7099 | n27834 ;
  assign n27836 = ( ~n211 & n8321 ) | ( ~n211 & n20084 ) | ( n8321 & n20084 ) ;
  assign n27837 = ( n3016 & n5138 ) | ( n3016 & n10584 ) | ( n5138 & n10584 ) ;
  assign n27838 = n27837 ^ n22866 ^ n1317 ;
  assign n27839 = n5236 ^ n3575 ^ 1'b0 ;
  assign n27840 = n27839 ^ n6522 ^ n915 ;
  assign n27841 = ( n9043 & n20455 ) | ( n9043 & n27634 ) | ( n20455 & n27634 ) ;
  assign n27842 = ( n6166 & ~n7928 ) | ( n6166 & n27841 ) | ( ~n7928 & n27841 ) ;
  assign n27843 = n18125 & ~n18654 ;
  assign n27844 = n1236 & n27843 ;
  assign n27845 = n13871 ^ n4071 ^ 1'b0 ;
  assign n27846 = ~n18993 & n20510 ;
  assign n27847 = n6934 | n27846 ;
  assign n27848 = n27845 & ~n27847 ;
  assign n27849 = n21004 ^ n12930 ^ 1'b0 ;
  assign n27850 = n3606 & ~n8976 ;
  assign n27851 = n3714 & ~n27850 ;
  assign n27852 = n27851 ^ n4420 ^ 1'b0 ;
  assign n27853 = n21181 ^ n1400 ^ 1'b0 ;
  assign n27854 = n12020 ^ n6539 ^ n2092 ;
  assign n27855 = n20441 & ~n27854 ;
  assign n27856 = n853 & ~n17015 ;
  assign n27857 = n27855 | n27856 ;
  assign n27858 = n12945 | n27857 ;
  assign n27859 = n15738 & n27858 ;
  assign n27860 = ( n1100 & n27853 ) | ( n1100 & n27859 ) | ( n27853 & n27859 ) ;
  assign n27861 = n7581 ^ n5951 ^ n1025 ;
  assign n27862 = n18683 ^ n12122 ^ n1129 ;
  assign n27863 = n27862 ^ n1027 ^ n491 ;
  assign n27864 = n2712 & ~n23268 ;
  assign n27865 = ~n11179 & n27864 ;
  assign n27866 = n1125 & n9373 ;
  assign n27867 = n22284 & n27866 ;
  assign n27868 = n14817 | n27867 ;
  assign n27869 = n27868 ^ n14249 ^ 1'b0 ;
  assign n27870 = n1591 & ~n13046 ;
  assign n27871 = n24065 ^ n4109 ^ 1'b0 ;
  assign n27872 = n2383 & ~n11399 ;
  assign n27873 = n6687 & ~n8022 ;
  assign n27874 = n6497 & n27873 ;
  assign n27875 = n23023 & n27874 ;
  assign n27876 = n19334 ^ n8864 ^ n1295 ;
  assign n27877 = n8145 ^ n5635 ^ x113 ;
  assign n27878 = n3319 | n3666 ;
  assign n27879 = n27878 ^ n21284 ^ 1'b0 ;
  assign n27880 = n23985 ^ n11586 ^ n10768 ;
  assign n27881 = n14115 ^ n9116 ^ 1'b0 ;
  assign n27882 = n27880 & n27881 ;
  assign n27883 = ~n5669 & n20048 ;
  assign n27884 = n22732 ^ n4236 ^ 1'b0 ;
  assign n27885 = ( n4155 & n4331 ) | ( n4155 & ~n8126 ) | ( n4331 & ~n8126 ) ;
  assign n27886 = ~n5753 & n27885 ;
  assign n27887 = ~n27884 & n27886 ;
  assign n27888 = n15384 & n25773 ;
  assign n27889 = ~n14921 & n15070 ;
  assign n27890 = n13203 ^ n1311 ^ n1136 ;
  assign n27891 = n11632 ^ n10908 ^ 1'b0 ;
  assign n27892 = n13112 & ~n27891 ;
  assign n27893 = n23750 ^ n3826 ^ 1'b0 ;
  assign n27894 = n3828 | n27893 ;
  assign n27895 = n27894 ^ n1106 ^ 1'b0 ;
  assign n27896 = n27895 ^ n17248 ^ 1'b0 ;
  assign n27897 = n1322 & ~n1358 ;
  assign n27898 = ~n8209 & n27897 ;
  assign n27899 = ~n3611 & n7392 ;
  assign n27900 = n27898 & n27899 ;
  assign n27901 = n13602 ^ n8891 ^ 1'b0 ;
  assign n27902 = n1915 & ~n21018 ;
  assign n27903 = n2430 & n11720 ;
  assign n27904 = ~n21184 & n27903 ;
  assign n27905 = ( n530 & ~n1611 ) | ( n530 & n12979 ) | ( ~n1611 & n12979 ) ;
  assign n27906 = n9775 ^ n855 ^ 1'b0 ;
  assign n27907 = ~n5782 & n12279 ;
  assign n27908 = n27907 ^ n19693 ^ 1'b0 ;
  assign n27909 = n27908 ^ n24805 ^ 1'b0 ;
  assign n27910 = n9200 | n25883 ;
  assign n27911 = n11450 | n27910 ;
  assign n27912 = n25420 ^ n7158 ^ 1'b0 ;
  assign n27913 = ~n13721 & n27912 ;
  assign n27914 = n6183 | n23428 ;
  assign n27915 = n767 & ~n27914 ;
  assign n27916 = ~n11151 & n19617 ;
  assign n27917 = n24146 ^ n6752 ^ x90 ;
  assign n27918 = n26429 ^ n23746 ^ n10665 ;
  assign n27919 = ( n6614 & n16565 ) | ( n6614 & ~n27918 ) | ( n16565 & ~n27918 ) ;
  assign n27921 = n27633 ^ n2745 ^ 1'b0 ;
  assign n27920 = n9760 | n13268 ;
  assign n27922 = n27921 ^ n27920 ^ 1'b0 ;
  assign n27923 = n27922 ^ n8719 ^ 1'b0 ;
  assign n27924 = ( n3011 & ~n19170 ) | ( n3011 & n27923 ) | ( ~n19170 & n27923 ) ;
  assign n27925 = n18104 & ~n27924 ;
  assign n27926 = ~n14462 & n27925 ;
  assign n27927 = n13778 ^ n4940 ^ 1'b0 ;
  assign n27928 = n19192 & ~n27927 ;
  assign n27929 = n25332 ^ n15475 ^ 1'b0 ;
  assign n27930 = n15228 & n27929 ;
  assign n27931 = n20413 ^ n9512 ^ 1'b0 ;
  assign n27932 = n10388 & n14957 ;
  assign n27933 = n16983 ^ n1205 ^ 1'b0 ;
  assign n27934 = n3218 & ~n27933 ;
  assign n27938 = n7094 & ~n9114 ;
  assign n27939 = ~n17945 & n27938 ;
  assign n27937 = n20469 ^ n11515 ^ n1725 ;
  assign n27940 = n27939 ^ n27937 ^ n8236 ;
  assign n27935 = ~n5421 & n11540 ;
  assign n27936 = ~n420 & n27935 ;
  assign n27941 = n27940 ^ n27936 ^ n17220 ;
  assign n27943 = n24532 ^ n15296 ^ 1'b0 ;
  assign n27942 = ( ~n6092 & n14079 ) | ( ~n6092 & n21944 ) | ( n14079 & n21944 ) ;
  assign n27944 = n27943 ^ n27942 ^ n22079 ;
  assign n27945 = n25786 ^ n744 ^ 1'b0 ;
  assign n27946 = n10540 & ~n27945 ;
  assign n27947 = ( n23837 & n24888 ) | ( n23837 & ~n27946 ) | ( n24888 & ~n27946 ) ;
  assign n27948 = n5372 & n8845 ;
  assign n27949 = ( ~n4802 & n23460 ) | ( ~n4802 & n27948 ) | ( n23460 & n27948 ) ;
  assign n27950 = n27949 ^ n2650 ^ n2106 ;
  assign n27951 = n27950 ^ n19052 ^ 1'b0 ;
  assign n27952 = ( ~n377 & n10390 ) | ( ~n377 & n14257 ) | ( n10390 & n14257 ) ;
  assign n27953 = n5552 | n27952 ;
  assign n27954 = n17530 & ~n27953 ;
  assign n27955 = ~n504 & n9835 ;
  assign n27956 = n25343 ^ n19372 ^ n234 ;
  assign n27957 = n27955 & ~n27956 ;
  assign n27958 = n17102 ^ n7768 ^ 1'b0 ;
  assign n27959 = n27957 & n27958 ;
  assign n27960 = n3034 & ~n11493 ;
  assign n27961 = n972 & n27960 ;
  assign n27962 = n5384 & n8101 ;
  assign n27963 = n27961 & n27962 ;
  assign n27964 = n5425 | n14528 ;
  assign n27965 = n802 ^ n232 ^ 1'b0 ;
  assign n27966 = n9089 & n27965 ;
  assign n27967 = ~n7053 & n27966 ;
  assign n27968 = n434 | n5046 ;
  assign n27969 = n20251 & ~n27968 ;
  assign n27970 = ( n5147 & ~n11418 ) | ( n5147 & n27969 ) | ( ~n11418 & n27969 ) ;
  assign n27971 = ~n2406 & n4020 ;
  assign n27972 = n27971 ^ n2573 ^ 1'b0 ;
  assign n27973 = ~n14201 & n27972 ;
  assign n27974 = n4224 & n27973 ;
  assign n27975 = ( n22511 & n26299 ) | ( n22511 & ~n27974 ) | ( n26299 & ~n27974 ) ;
  assign n27976 = n23869 ^ n11389 ^ 1'b0 ;
  assign n27977 = ~n12053 & n12410 ;
  assign n27978 = n7989 & n27977 ;
  assign n27979 = n20478 ^ n755 ^ 1'b0 ;
  assign n27980 = ~n15471 & n27979 ;
  assign n27981 = n9075 & ~n16370 ;
  assign n27982 = n12235 & n20582 ;
  assign n27983 = n22462 ^ n3815 ^ 1'b0 ;
  assign n27984 = n27982 | n27983 ;
  assign n27985 = n24973 ^ x92 ^ 1'b0 ;
  assign n27986 = n3211 | n27985 ;
  assign n27987 = ( n11296 & n15001 ) | ( n11296 & n25591 ) | ( n15001 & n25591 ) ;
  assign n27988 = n25558 ^ n11193 ^ n10429 ;
  assign n27989 = n22590 ^ n11186 ^ 1'b0 ;
  assign n27991 = ~n9461 & n17179 ;
  assign n27992 = ~n17179 & n27991 ;
  assign n27990 = n975 & ~n2693 ;
  assign n27993 = n27992 ^ n27990 ^ 1'b0 ;
  assign n27994 = n726 & ~n2767 ;
  assign n27995 = ~n726 & n27994 ;
  assign n27996 = n12131 | n27995 ;
  assign n27997 = n27995 & ~n27996 ;
  assign n27998 = n1898 | n5630 ;
  assign n27999 = n1898 & ~n27998 ;
  assign n28000 = n27999 ^ n3905 ^ 1'b0 ;
  assign n28001 = n27997 | n28000 ;
  assign n28002 = ( n2040 & ~n11115 ) | ( n2040 & n28001 ) | ( ~n11115 & n28001 ) ;
  assign n28003 = ~n10085 & n28002 ;
  assign n28004 = ~n27993 & n28003 ;
  assign n28005 = n28004 ^ n22348 ^ n15901 ;
  assign n28006 = n15723 | n28005 ;
  assign n28007 = n16015 ^ n13133 ^ 1'b0 ;
  assign n28008 = n20575 ^ n11150 ^ 1'b0 ;
  assign n28009 = ~n8524 & n16831 ;
  assign n28010 = n28009 ^ n897 ^ 1'b0 ;
  assign n28011 = n10851 & n13851 ;
  assign n28012 = n6137 & n28011 ;
  assign n28013 = n6158 & n28012 ;
  assign n28014 = n13838 | n27653 ;
  assign n28015 = n26874 | n28014 ;
  assign n28016 = n7656 | n15141 ;
  assign n28017 = n28016 ^ n14893 ^ 1'b0 ;
  assign n28018 = n28017 ^ n20555 ^ 1'b0 ;
  assign n28022 = n4541 | n22268 ;
  assign n28023 = n28022 ^ n5400 ^ 1'b0 ;
  assign n28024 = n28023 ^ n2247 ^ 1'b0 ;
  assign n28025 = n6772 & ~n28024 ;
  assign n28019 = ( n7192 & n7794 ) | ( n7192 & ~n9985 ) | ( n7794 & ~n9985 ) ;
  assign n28020 = n28019 ^ n14060 ^ 1'b0 ;
  assign n28021 = n28020 ^ n3231 ^ n1819 ;
  assign n28026 = n28025 ^ n28021 ^ n19392 ;
  assign n28027 = ( x21 & ~n3888 ) | ( x21 & n26738 ) | ( ~n3888 & n26738 ) ;
  assign n28028 = n28027 ^ n17056 ^ 1'b0 ;
  assign n28031 = ~n19312 & n20854 ;
  assign n28029 = n2401 ^ n593 ^ 1'b0 ;
  assign n28030 = n15625 | n28029 ;
  assign n28032 = n28031 ^ n28030 ^ 1'b0 ;
  assign n28033 = n14507 ^ n10639 ^ n4815 ;
  assign n28034 = n28033 ^ n13652 ^ n2167 ;
  assign n28035 = ( ~n8548 & n14902 ) | ( ~n8548 & n28034 ) | ( n14902 & n28034 ) ;
  assign n28036 = n26841 ^ n14677 ^ 1'b0 ;
  assign n28037 = n28035 | n28036 ;
  assign n28038 = ~n20154 & n27077 ;
  assign n28039 = n20852 ^ n14943 ^ 1'b0 ;
  assign n28040 = n1012 & ~n18177 ;
  assign n28041 = n11821 ^ n11513 ^ n5555 ;
  assign n28042 = ( n5854 & ~n10281 ) | ( n5854 & n28041 ) | ( ~n10281 & n28041 ) ;
  assign n28043 = n8826 & ~n8988 ;
  assign n28044 = n13168 | n17627 ;
  assign n28045 = n28044 ^ n20352 ^ 1'b0 ;
  assign n28046 = n22416 ^ n17664 ^ n6227 ;
  assign n28047 = n18158 ^ n2072 ^ 1'b0 ;
  assign n28048 = ~n15420 & n28047 ;
  assign n28049 = n16597 ^ n7892 ^ 1'b0 ;
  assign n28050 = n5469 & ~n28049 ;
  assign n28051 = ( ~n2934 & n14201 ) | ( ~n2934 & n24726 ) | ( n14201 & n24726 ) ;
  assign n28052 = n9766 & ~n10317 ;
  assign n28053 = n28051 & n28052 ;
  assign n28054 = n15549 ^ n2411 ^ n1094 ;
  assign n28055 = n28054 ^ n23512 ^ n3886 ;
  assign n28056 = n9306 ^ n6070 ^ 1'b0 ;
  assign n28057 = n17090 ^ n16212 ^ x29 ;
  assign n28060 = ( ~n5603 & n8312 ) | ( ~n5603 & n12418 ) | ( n8312 & n12418 ) ;
  assign n28058 = n4380 & n24503 ;
  assign n28059 = n28058 ^ n27592 ^ 1'b0 ;
  assign n28061 = n28060 ^ n28059 ^ n2085 ;
  assign n28062 = n19558 ^ n9380 ^ 1'b0 ;
  assign n28063 = n14180 & ~n24792 ;
  assign n28064 = n7658 ^ n6840 ^ 1'b0 ;
  assign n28065 = n20306 & ~n28064 ;
  assign n28066 = n8601 ^ n1867 ^ 1'b0 ;
  assign n28067 = ( n895 & ~n2510 ) | ( n895 & n4937 ) | ( ~n2510 & n4937 ) ;
  assign n28068 = n6010 & ~n9562 ;
  assign n28069 = n28068 ^ n18644 ^ 1'b0 ;
  assign n28070 = ~n2272 & n5369 ;
  assign n28071 = ~n10118 & n28070 ;
  assign n28072 = n28071 ^ n9113 ^ n3744 ;
  assign n28073 = ( n28067 & n28069 ) | ( n28067 & n28072 ) | ( n28069 & n28072 ) ;
  assign n28074 = ( n2833 & ~n5416 ) | ( n2833 & n8574 ) | ( ~n5416 & n8574 ) ;
  assign n28075 = ~n8436 & n28074 ;
  assign n28076 = n28075 ^ n13233 ^ 1'b0 ;
  assign n28077 = ~n8705 & n28076 ;
  assign n28078 = ~n28073 & n28077 ;
  assign n28079 = n21088 & ~n25101 ;
  assign n28080 = n28079 ^ n4103 ^ 1'b0 ;
  assign n28081 = n24507 ^ n10883 ^ 1'b0 ;
  assign n28082 = n9215 ^ n3661 ^ 1'b0 ;
  assign n28083 = n28081 & n28082 ;
  assign n28084 = n15140 ^ n6447 ^ n4499 ;
  assign n28085 = n28083 & ~n28084 ;
  assign n28086 = n25697 ^ n18333 ^ n8212 ;
  assign n28087 = ( n10660 & n17185 ) | ( n10660 & n20650 ) | ( n17185 & n20650 ) ;
  assign n28088 = n28087 ^ n3316 ^ 1'b0 ;
  assign n28089 = n28088 ^ n20732 ^ n17311 ;
  assign n28091 = n7351 ^ n1700 ^ 1'b0 ;
  assign n28090 = n7844 ^ n1986 ^ 1'b0 ;
  assign n28092 = n28091 ^ n28090 ^ n2364 ;
  assign n28093 = n5370 | n14095 ;
  assign n28094 = n28093 ^ n8700 ^ 1'b0 ;
  assign n28095 = n13615 ^ n3389 ^ 1'b0 ;
  assign n28096 = n9004 & n22031 ;
  assign n28097 = ~n2143 & n28096 ;
  assign n28098 = n11415 & ~n28097 ;
  assign n28099 = n15440 & n28098 ;
  assign n28100 = n28099 ^ n13983 ^ 1'b0 ;
  assign n28101 = n839 & n17451 ;
  assign n28102 = ( ~n18756 & n22754 ) | ( ~n18756 & n28101 ) | ( n22754 & n28101 ) ;
  assign n28104 = ~n3873 & n12557 ;
  assign n28105 = ~n5533 & n28104 ;
  assign n28103 = ( n316 & ~n9021 ) | ( n316 & n17789 ) | ( ~n9021 & n17789 ) ;
  assign n28106 = n28105 ^ n28103 ^ n22299 ;
  assign n28107 = n17483 ^ n12110 ^ x108 ;
  assign n28108 = n2554 & n28107 ;
  assign n28109 = n28108 ^ n20034 ^ n389 ;
  assign n28110 = n9522 | n13779 ;
  assign n28111 = n28110 ^ n27884 ^ 1'b0 ;
  assign n28112 = n27320 ^ n16804 ^ 1'b0 ;
  assign n28113 = n3611 | n9659 ;
  assign n28114 = n667 & ~n28113 ;
  assign n28115 = ( n1420 & n13310 ) | ( n1420 & ~n28114 ) | ( n13310 & ~n28114 ) ;
  assign n28117 = n7377 & ~n8569 ;
  assign n28118 = n20097 ^ n3113 ^ 1'b0 ;
  assign n28119 = ~n28117 & n28118 ;
  assign n28116 = n20038 ^ n12445 ^ 1'b0 ;
  assign n28120 = n28119 ^ n28116 ^ n14064 ;
  assign n28121 = n28120 ^ n11065 ^ 1'b0 ;
  assign n28122 = n28115 & n28121 ;
  assign n28123 = n5997 & n6445 ;
  assign n28124 = n28123 ^ n11312 ^ 1'b0 ;
  assign n28125 = n19087 | n27891 ;
  assign n28126 = n8345 ^ n4231 ^ 1'b0 ;
  assign n28127 = ~n2976 & n19185 ;
  assign n28128 = ~n1212 & n28127 ;
  assign n28129 = ~n14711 & n22590 ;
  assign n28130 = ( n15907 & ~n19196 ) | ( n15907 & n20614 ) | ( ~n19196 & n20614 ) ;
  assign n28131 = ( n7540 & n10807 ) | ( n7540 & ~n22994 ) | ( n10807 & ~n22994 ) ;
  assign n28133 = ~n8645 & n14185 ;
  assign n28134 = n28133 ^ n5531 ^ 1'b0 ;
  assign n28132 = n13547 & n25090 ;
  assign n28135 = n28134 ^ n28132 ^ 1'b0 ;
  assign n28136 = ~n13409 & n16769 ;
  assign n28137 = n19705 ^ n8552 ^ 1'b0 ;
  assign n28138 = ~n22647 & n28137 ;
  assign n28139 = n9619 | n22978 ;
  assign n28140 = n15614 ^ n10148 ^ 1'b0 ;
  assign n28141 = n1250 & n6294 ;
  assign n28142 = n28141 ^ n13932 ^ n5759 ;
  assign n28143 = n6445 | n23878 ;
  assign n28144 = n28143 ^ n9638 ^ 1'b0 ;
  assign n28145 = n28144 ^ n16033 ^ n8321 ;
  assign n28146 = n795 | n14838 ;
  assign n28147 = n28146 ^ n6142 ^ 1'b0 ;
  assign n28148 = n3816 & ~n4608 ;
  assign n28149 = n20442 & n28148 ;
  assign n28150 = n11198 ^ n163 ^ 1'b0 ;
  assign n28151 = ~n27855 & n28150 ;
  assign n28152 = n8351 ^ n374 ^ 1'b0 ;
  assign n28153 = n13120 ^ n5881 ^ 1'b0 ;
  assign n28154 = n17407 | n28153 ;
  assign n28155 = n12974 & ~n16669 ;
  assign n28156 = n28155 ^ n7021 ^ n3879 ;
  assign n28157 = n16926 ^ n9858 ^ 1'b0 ;
  assign n28158 = ( n2715 & n11409 ) | ( n2715 & ~n28157 ) | ( n11409 & ~n28157 ) ;
  assign n28159 = n14338 | n24239 ;
  assign n28160 = n24724 ^ n18746 ^ x68 ;
  assign n28161 = ~n16162 & n25015 ;
  assign n28162 = n28160 & n28161 ;
  assign n28163 = n6111 & ~n7137 ;
  assign n28164 = n28069 ^ n424 ^ 1'b0 ;
  assign n28165 = x1 & n28164 ;
  assign n28166 = n4929 & n7171 ;
  assign n28167 = n28166 ^ n11480 ^ 1'b0 ;
  assign n28168 = n28165 & n28167 ;
  assign n28169 = n18490 ^ n1546 ^ 1'b0 ;
  assign n28170 = ~n18223 & n28169 ;
  assign n28171 = ~n827 & n28170 ;
  assign n28172 = ~n218 & n28171 ;
  assign n28173 = n10860 ^ n445 ^ 1'b0 ;
  assign n28174 = ( n3777 & n12408 ) | ( n3777 & ~n28173 ) | ( n12408 & ~n28173 ) ;
  assign n28175 = n28174 ^ n10323 ^ 1'b0 ;
  assign n28176 = n20080 ^ n14941 ^ n12815 ;
  assign n28177 = n21385 ^ n17165 ^ 1'b0 ;
  assign n28178 = n12949 | n24785 ;
  assign n28179 = n28178 ^ n24442 ^ n6422 ;
  assign n28180 = n7311 & ~n12961 ;
  assign n28181 = ~n1990 & n28180 ;
  assign n28182 = n15636 ^ n2942 ^ 1'b0 ;
  assign n28183 = n13541 ^ n5973 ^ 1'b0 ;
  assign n28184 = n18965 & ~n28183 ;
  assign n28185 = n7056 | n9786 ;
  assign n28186 = n28184 | n28185 ;
  assign n28187 = n28186 ^ n1365 ^ 1'b0 ;
  assign n28188 = n2239 ^ n941 ^ 1'b0 ;
  assign n28189 = n6601 & ~n28188 ;
  assign n28190 = n309 & n28189 ;
  assign n28191 = n28190 ^ n9075 ^ 1'b0 ;
  assign n28192 = n10369 ^ n5752 ^ n4996 ;
  assign n28193 = n28192 ^ n5890 ^ 1'b0 ;
  assign n28194 = n9793 & ~n28193 ;
  assign n28195 = ( n967 & n3442 ) | ( n967 & ~n24883 ) | ( n3442 & ~n24883 ) ;
  assign n28196 = ( n15499 & n19812 ) | ( n15499 & n28195 ) | ( n19812 & n28195 ) ;
  assign n28197 = n1067 & ~n17152 ;
  assign n28198 = n28197 ^ n3803 ^ n2241 ;
  assign n28199 = ( n210 & n8321 ) | ( n210 & n19943 ) | ( n8321 & n19943 ) ;
  assign n28200 = n9733 ^ n8101 ^ 1'b0 ;
  assign n28201 = n24386 & ~n28200 ;
  assign n28202 = n21982 & n28201 ;
  assign n28203 = n2921 & n28202 ;
  assign n28204 = n14923 & n21302 ;
  assign n28205 = n23028 | n23236 ;
  assign n28206 = n28204 & ~n28205 ;
  assign n28207 = n10850 ^ n4085 ^ 1'b0 ;
  assign n28208 = ~n1743 & n2648 ;
  assign n28209 = n3406 | n28208 ;
  assign n28210 = n18262 & ~n28209 ;
  assign n28211 = n21066 | n28210 ;
  assign n28212 = n28207 & ~n28211 ;
  assign n28213 = n8539 & n27559 ;
  assign n28214 = n28213 ^ n15319 ^ n14039 ;
  assign n28215 = n10114 & ~n13880 ;
  assign n28216 = ( n4688 & n25615 ) | ( n4688 & n28215 ) | ( n25615 & n28215 ) ;
  assign n28217 = n795 | n4614 ;
  assign n28218 = n28217 ^ n3010 ^ 1'b0 ;
  assign n28219 = ( n10840 & n16208 ) | ( n10840 & ~n28218 ) | ( n16208 & ~n28218 ) ;
  assign n28220 = n20661 & ~n22593 ;
  assign n28221 = n28220 ^ n19904 ^ n11206 ;
  assign n28222 = n19211 & ~n28221 ;
  assign n28223 = n25115 | n26766 ;
  assign n28224 = ~x92 & n5187 ;
  assign n28225 = ~n7058 & n24056 ;
  assign n28226 = n15049 & n28225 ;
  assign n28227 = n10103 & n18145 ;
  assign n28228 = n5920 & ~n10527 ;
  assign n28229 = n16418 & n28228 ;
  assign n28230 = n18704 & n28229 ;
  assign n28231 = ( n14820 & n19142 ) | ( n14820 & ~n20661 ) | ( n19142 & ~n20661 ) ;
  assign n28232 = n24928 ^ n20510 ^ 1'b0 ;
  assign n28233 = n1826 & n28232 ;
  assign n28234 = ( n1522 & n5612 ) | ( n1522 & ~n6809 ) | ( n5612 & ~n6809 ) ;
  assign n28235 = ~n8865 & n28234 ;
  assign n28236 = n28235 ^ n20119 ^ 1'b0 ;
  assign n28237 = n28233 & n28236 ;
  assign n28239 = n8204 ^ n7420 ^ n3169 ;
  assign n28238 = ( ~n1477 & n4123 ) | ( ~n1477 & n25306 ) | ( n4123 & n25306 ) ;
  assign n28240 = n28239 ^ n28238 ^ n13114 ;
  assign n28241 = n15452 ^ n9990 ^ n1690 ;
  assign n28242 = n15969 & ~n28241 ;
  assign n28243 = n23381 ^ n2389 ^ 1'b0 ;
  assign n28244 = n28243 ^ n27636 ^ n26843 ;
  assign n28245 = n21143 | n28244 ;
  assign n28246 = n28245 ^ n7302 ^ 1'b0 ;
  assign n28247 = n2957 | n6830 ;
  assign n28248 = n28247 ^ n5191 ^ 1'b0 ;
  assign n28249 = n9807 | n28248 ;
  assign n28250 = n28249 ^ n9126 ^ 1'b0 ;
  assign n28251 = ( ~n5301 & n9304 ) | ( ~n5301 & n17047 ) | ( n9304 & n17047 ) ;
  assign n28252 = ( n3707 & ~n21686 ) | ( n3707 & n28251 ) | ( ~n21686 & n28251 ) ;
  assign n28253 = ~n4789 & n26749 ;
  assign n28254 = ~n28252 & n28253 ;
  assign n28255 = n25365 ^ n18549 ^ 1'b0 ;
  assign n28256 = n21987 ^ n4057 ^ x31 ;
  assign n28257 = n5956 & n28256 ;
  assign n28258 = ( ~n2239 & n6088 ) | ( ~n2239 & n17501 ) | ( n6088 & n17501 ) ;
  assign n28259 = n28258 ^ n13650 ^ n8937 ;
  assign n28260 = n1485 | n3281 ;
  assign n28261 = n5314 & ~n28260 ;
  assign n28262 = n14659 & n28261 ;
  assign n28263 = n28262 ^ n22393 ^ n9380 ;
  assign n28264 = n19959 ^ n7094 ^ n3828 ;
  assign n28265 = n18002 ^ n3968 ^ 1'b0 ;
  assign n28266 = n11784 ^ n2181 ^ 1'b0 ;
  assign n28267 = n10122 & n28266 ;
  assign n28268 = n4090 & n4220 ;
  assign n28269 = n10775 ^ n8987 ^ 1'b0 ;
  assign n28270 = n1697 | n18425 ;
  assign n28271 = n25145 & ~n28270 ;
  assign n28272 = n365 | n9147 ;
  assign n28273 = n28272 ^ n3244 ^ n2917 ;
  assign n28274 = n4498 | n9603 ;
  assign n28275 = n28274 ^ n22130 ^ n9569 ;
  assign n28276 = n18190 ^ n6986 ^ n5807 ;
  assign n28277 = n28276 ^ n4349 ^ n2845 ;
  assign n28278 = n4593 & n9771 ;
  assign n28279 = n28278 ^ n7726 ^ 1'b0 ;
  assign n28280 = n28279 ^ n5098 ^ 1'b0 ;
  assign n28281 = n7425 ^ n1068 ^ 1'b0 ;
  assign n28282 = ( n8130 & ~n10875 ) | ( n8130 & n24942 ) | ( ~n10875 & n24942 ) ;
  assign n28283 = n8871 & ~n28282 ;
  assign n28284 = ~n2219 & n16581 ;
  assign n28285 = n4289 ^ n3482 ^ 1'b0 ;
  assign n28286 = n12295 ^ n5840 ^ 1'b0 ;
  assign n28287 = ( n8204 & ~n27952 ) | ( n8204 & n28286 ) | ( ~n27952 & n28286 ) ;
  assign n28288 = n15744 & n16599 ;
  assign n28289 = n26482 ^ n7550 ^ 1'b0 ;
  assign n28290 = n8551 | n11688 ;
  assign n28291 = n9556 & n28290 ;
  assign n28292 = n14945 & n28291 ;
  assign n28293 = ~n2619 & n2945 ;
  assign n28294 = n3815 & n28293 ;
  assign n28295 = ( ~x29 & n19659 ) | ( ~x29 & n20345 ) | ( n19659 & n20345 ) ;
  assign n28296 = n28295 ^ n6619 ^ n4397 ;
  assign n28297 = n13464 ^ n12747 ^ 1'b0 ;
  assign n28298 = ( n28294 & n28296 ) | ( n28294 & ~n28297 ) | ( n28296 & ~n28297 ) ;
  assign n28299 = n2275 | n28298 ;
  assign n28300 = n28299 ^ n4746 ^ 1'b0 ;
  assign n28301 = n8299 & n15220 ;
  assign n28302 = n3072 & n28301 ;
  assign n28303 = n7707 & n24861 ;
  assign n28304 = ~n356 & n28303 ;
  assign n28305 = n17891 ^ n10991 ^ n798 ;
  assign n28306 = ( n5009 & ~n11143 ) | ( n5009 & n14826 ) | ( ~n11143 & n14826 ) ;
  assign n28307 = n9787 ^ n8643 ^ 1'b0 ;
  assign n28308 = n20427 ^ n4055 ^ n3211 ;
  assign n28309 = n3621 ^ n2216 ^ 1'b0 ;
  assign n28311 = n21105 ^ n6483 ^ 1'b0 ;
  assign n28310 = n2872 & n15980 ;
  assign n28312 = n28311 ^ n28310 ^ 1'b0 ;
  assign n28313 = n21167 ^ n4186 ^ 1'b0 ;
  assign n28314 = n17554 & ~n28313 ;
  assign n28315 = n23824 ^ n3834 ^ 1'b0 ;
  assign n28316 = ~n3779 & n28315 ;
  assign n28317 = n2806 & n28316 ;
  assign n28318 = n19234 ^ n2827 ^ 1'b0 ;
  assign n28319 = n10262 | n28318 ;
  assign n28322 = ~n2976 & n6085 ;
  assign n28323 = n28322 ^ n9406 ^ 1'b0 ;
  assign n28320 = n1489 ^ n904 ^ 1'b0 ;
  assign n28321 = n3345 | n28320 ;
  assign n28324 = n28323 ^ n28321 ^ n14196 ;
  assign n28325 = ( ~n12419 & n15650 ) | ( ~n12419 & n28324 ) | ( n15650 & n28324 ) ;
  assign n28326 = n28325 ^ n9607 ^ 1'b0 ;
  assign n28327 = ( n2036 & n3119 ) | ( n2036 & ~n5911 ) | ( n3119 & ~n5911 ) ;
  assign n28328 = n8521 & n28327 ;
  assign n28329 = n10431 & n28328 ;
  assign n28330 = n28329 ^ n18842 ^ 1'b0 ;
  assign n28331 = ( n1147 & ~n2437 ) | ( n1147 & n23746 ) | ( ~n2437 & n23746 ) ;
  assign n28332 = n13807 ^ n4029 ^ 1'b0 ;
  assign n28333 = ~n19465 & n28332 ;
  assign n28334 = ( n9105 & ~n28331 ) | ( n9105 & n28333 ) | ( ~n28331 & n28333 ) ;
  assign n28335 = n10956 & ~n14836 ;
  assign n28336 = n28335 ^ n15768 ^ 1'b0 ;
  assign n28337 = ( n10659 & ~n15089 ) | ( n10659 & n17484 ) | ( ~n15089 & n17484 ) ;
  assign n28338 = n13936 & ~n14900 ;
  assign n28339 = n28338 ^ n10960 ^ 1'b0 ;
  assign n28340 = n17129 ^ n15836 ^ 1'b0 ;
  assign n28341 = n1942 | n28340 ;
  assign n28342 = n11791 | n28341 ;
  assign n28346 = n12558 ^ n1415 ^ 1'b0 ;
  assign n28347 = n15596 | n28346 ;
  assign n28343 = n5817 & ~n8729 ;
  assign n28344 = ~n1068 & n9938 ;
  assign n28345 = ~n28343 & n28344 ;
  assign n28348 = n28347 ^ n28345 ^ n25754 ;
  assign n28349 = n23660 ^ n17407 ^ 1'b0 ;
  assign n28350 = n26929 ^ n7248 ^ n4515 ;
  assign n28351 = ( ~n6661 & n25878 ) | ( ~n6661 & n28350 ) | ( n25878 & n28350 ) ;
  assign n28352 = n15705 ^ n14363 ^ n5873 ;
  assign n28353 = ~n2961 & n22189 ;
  assign n28354 = n1031 & ~n27873 ;
  assign n28355 = ~n28353 & n28354 ;
  assign n28356 = ( ~n1750 & n2293 ) | ( ~n1750 & n8808 ) | ( n2293 & n8808 ) ;
  assign n28357 = n17236 | n28356 ;
  assign n28358 = n19511 & ~n28357 ;
  assign n28359 = n11274 | n28358 ;
  assign n28360 = n28359 ^ n20086 ^ 1'b0 ;
  assign n28361 = n27401 ^ n3059 ^ 1'b0 ;
  assign n28362 = n12644 & n28361 ;
  assign n28363 = n4868 ^ n4267 ^ 1'b0 ;
  assign n28364 = ~n10597 & n28363 ;
  assign n28365 = n12913 ^ n9507 ^ 1'b0 ;
  assign n28366 = n1365 & ~n28365 ;
  assign n28367 = n6356 & n25851 ;
  assign n28368 = n19151 & ~n28367 ;
  assign n28369 = n28368 ^ n2559 ^ 1'b0 ;
  assign n28370 = n20319 ^ n8105 ^ 1'b0 ;
  assign n28371 = ( ~n203 & n749 ) | ( ~n203 & n1529 ) | ( n749 & n1529 ) ;
  assign n28372 = n28371 ^ n14451 ^ 1'b0 ;
  assign n28373 = ( n248 & ~n12870 ) | ( n248 & n28372 ) | ( ~n12870 & n28372 ) ;
  assign n28374 = n23749 ^ n21671 ^ n449 ;
  assign n28375 = n9016 & ~n11468 ;
  assign n28376 = n6112 & n14353 ;
  assign n28377 = n8945 & ~n17569 ;
  assign n28378 = ~n5658 & n28377 ;
  assign n28381 = n14115 & n17077 ;
  assign n28382 = ~n19018 & n28381 ;
  assign n28379 = n22208 ^ n2906 ^ n1055 ;
  assign n28380 = n4343 & ~n28379 ;
  assign n28383 = n28382 ^ n28380 ^ 1'b0 ;
  assign n28384 = ( n10687 & ~n22537 ) | ( n10687 & n28383 ) | ( ~n22537 & n28383 ) ;
  assign n28385 = n15529 ^ n10370 ^ n6483 ;
  assign n28386 = n28385 ^ n7994 ^ 1'b0 ;
  assign n28387 = n3246 & ~n24201 ;
  assign n28388 = n23286 ^ n16497 ^ n10266 ;
  assign n28389 = ( n5000 & n10398 ) | ( n5000 & n18676 ) | ( n10398 & n18676 ) ;
  assign n28390 = n27345 ^ n16226 ^ 1'b0 ;
  assign n28391 = n28389 | n28390 ;
  assign n28392 = n8355 & n24300 ;
  assign n28393 = ~x73 & n28392 ;
  assign n28394 = n11616 ^ n9668 ^ 1'b0 ;
  assign n28395 = n8958 ^ n8363 ^ 1'b0 ;
  assign n28396 = n4431 | n28395 ;
  assign n28397 = n5914 | n14606 ;
  assign n28398 = n11236 & ~n28397 ;
  assign n28399 = n28398 ^ n25748 ^ 1'b0 ;
  assign n28400 = n3762 | n5195 ;
  assign n28401 = n28400 ^ n9327 ^ 1'b0 ;
  assign n28402 = ( n9679 & ~n24402 ) | ( n9679 & n28401 ) | ( ~n24402 & n28401 ) ;
  assign n28403 = ( n965 & n9482 ) | ( n965 & n18949 ) | ( n9482 & n18949 ) ;
  assign n28404 = ( n5349 & n8689 ) | ( n5349 & n10943 ) | ( n8689 & n10943 ) ;
  assign n28405 = n28404 ^ n6036 ^ 1'b0 ;
  assign n28406 = n19563 | n24241 ;
  assign n28407 = n15615 | n28406 ;
  assign n28408 = n16360 & n26201 ;
  assign n28409 = n11261 ^ n10584 ^ 1'b0 ;
  assign n28410 = n491 | n1118 ;
  assign n28411 = n8271 | n28410 ;
  assign n28412 = n13660 & n28411 ;
  assign n28413 = n1499 & n28412 ;
  assign n28414 = n27150 ^ n15837 ^ 1'b0 ;
  assign n28415 = n6982 | n28414 ;
  assign n28416 = n28413 & ~n28415 ;
  assign n28417 = n15789 ^ n6543 ^ 1'b0 ;
  assign n28418 = n16090 ^ n6131 ^ 1'b0 ;
  assign n28419 = ~n18453 & n27885 ;
  assign n28420 = n28419 ^ n1418 ^ 1'b0 ;
  assign n28421 = n25330 ^ n6326 ^ n6035 ;
  assign n28422 = ( ~n1539 & n24520 ) | ( ~n1539 & n28421 ) | ( n24520 & n28421 ) ;
  assign n28423 = n24498 ^ n4264 ^ n3141 ;
  assign n28424 = n17460 ^ n3023 ^ n1427 ;
  assign n28425 = n11630 | n21412 ;
  assign n28426 = n5870 | n28425 ;
  assign n28427 = n24040 ^ n20949 ^ 1'b0 ;
  assign n28428 = n14143 ^ n1123 ^ 1'b0 ;
  assign n28429 = n26234 & n28428 ;
  assign n28430 = ~n5691 & n28429 ;
  assign n28431 = ~n2189 & n28430 ;
  assign n28432 = n8161 ^ n847 ^ 1'b0 ;
  assign n28433 = n12728 & ~n28432 ;
  assign n28434 = n6300 ^ n3316 ^ 1'b0 ;
  assign n28435 = n25517 & n28434 ;
  assign n28436 = n21721 & n28435 ;
  assign n28437 = n21982 & n28436 ;
  assign y0 = x2 ;
  assign y1 = x16 ;
  assign y2 = x17 ;
  assign y3 = x23 ;
  assign y4 = x31 ;
  assign y5 = x35 ;
  assign y6 = x36 ;
  assign y7 = x39 ;
  assign y8 = x48 ;
  assign y9 = x53 ;
  assign y10 = x56 ;
  assign y11 = x61 ;
  assign y12 = x63 ;
  assign y13 = x64 ;
  assign y14 = x65 ;
  assign y15 = x66 ;
  assign y16 = x69 ;
  assign y17 = x79 ;
  assign y18 = x82 ;
  assign y19 = x92 ;
  assign y20 = x93 ;
  assign y21 = x103 ;
  assign y22 = x104 ;
  assign y23 = x105 ;
  assign y24 = x114 ;
  assign y25 = x117 ;
  assign y26 = x124 ;
  assign y27 = n129 ;
  assign y28 = ~n131 ;
  assign y29 = ~1'b0 ;
  assign y30 = ~1'b0 ;
  assign y31 = ~n134 ;
  assign y32 = ~n136 ;
  assign y33 = ~n138 ;
  assign y34 = n139 ;
  assign y35 = ~n143 ;
  assign y36 = ~1'b0 ;
  assign y37 = ~1'b0 ;
  assign y38 = ~n146 ;
  assign y39 = n148 ;
  assign y40 = ~n153 ;
  assign y41 = ~n157 ;
  assign y42 = n162 ;
  assign y43 = ~n163 ;
  assign y44 = ~n167 ;
  assign y45 = n168 ;
  assign y46 = n170 ;
  assign y47 = ~1'b0 ;
  assign y48 = ~n180 ;
  assign y49 = n181 ;
  assign y50 = ~n182 ;
  assign y51 = n184 ;
  assign y52 = ~n189 ;
  assign y53 = ~1'b0 ;
  assign y54 = ~n190 ;
  assign y55 = n191 ;
  assign y56 = n193 ;
  assign y57 = ~1'b0 ;
  assign y58 = ~n196 ;
  assign y59 = n197 ;
  assign y60 = n199 ;
  assign y61 = ~1'b0 ;
  assign y62 = n206 ;
  assign y63 = ~n209 ;
  assign y64 = ~n211 ;
  assign y65 = ~n216 ;
  assign y66 = ~n220 ;
  assign y67 = n222 ;
  assign y68 = ~n223 ;
  assign y69 = ~n227 ;
  assign y70 = ~1'b0 ;
  assign y71 = ~n229 ;
  assign y72 = n232 ;
  assign y73 = n234 ;
  assign y74 = ~n238 ;
  assign y75 = n243 ;
  assign y76 = n246 ;
  assign y77 = ~1'b0 ;
  assign y78 = n250 ;
  assign y79 = ~n260 ;
  assign y80 = ~1'b0 ;
  assign y81 = n265 ;
  assign y82 = ~n267 ;
  assign y83 = ~1'b0 ;
  assign y84 = ~1'b0 ;
  assign y85 = n272 ;
  assign y86 = n278 ;
  assign y87 = ~1'b0 ;
  assign y88 = ~n279 ;
  assign y89 = n286 ;
  assign y90 = ~1'b0 ;
  assign y91 = ~n288 ;
  assign y92 = n289 ;
  assign y93 = n290 ;
  assign y94 = ~n293 ;
  assign y95 = ~n296 ;
  assign y96 = ~n300 ;
  assign y97 = ~n303 ;
  assign y98 = ~1'b0 ;
  assign y99 = ~n305 ;
  assign y100 = n309 ;
  assign y101 = n310 ;
  assign y102 = n312 ;
  assign y103 = ~n319 ;
  assign y104 = n320 ;
  assign y105 = ~n325 ;
  assign y106 = n328 ;
  assign y107 = ~n331 ;
  assign y108 = n332 ;
  assign y109 = n334 ;
  assign y110 = n335 ;
  assign y111 = ~n341 ;
  assign y112 = ~1'b0 ;
  assign y113 = n354 ;
  assign y114 = ~n358 ;
  assign y115 = ~1'b0 ;
  assign y116 = ~n360 ;
  assign y117 = n363 ;
  assign y118 = n366 ;
  assign y119 = ~1'b0 ;
  assign y120 = n367 ;
  assign y121 = ~n379 ;
  assign y122 = n381 ;
  assign y123 = ~n384 ;
  assign y124 = ~n386 ;
  assign y125 = ~n391 ;
  assign y126 = ~n393 ;
  assign y127 = n402 ;
  assign y128 = n404 ;
  assign y129 = ~n406 ;
  assign y130 = ~n410 ;
  assign y131 = ~n415 ;
  assign y132 = ~n416 ;
  assign y133 = n419 ;
  assign y134 = ~1'b0 ;
  assign y135 = n424 ;
  assign y136 = ~n425 ;
  assign y137 = ~1'b0 ;
  assign y138 = n431 ;
  assign y139 = n432 ;
  assign y140 = n433 ;
  assign y141 = ~n434 ;
  assign y142 = ~1'b0 ;
  assign y143 = n442 ;
  assign y144 = n444 ;
  assign y145 = n448 ;
  assign y146 = ~n451 ;
  assign y147 = n453 ;
  assign y148 = ~n462 ;
  assign y149 = n463 ;
  assign y150 = n471 ;
  assign y151 = ~n480 ;
  assign y152 = ~n482 ;
  assign y153 = n487 ;
  assign y154 = ~n489 ;
  assign y155 = ~n491 ;
  assign y156 = ~n494 ;
  assign y157 = n496 ;
  assign y158 = ~1'b0 ;
  assign y159 = n499 ;
  assign y160 = n501 ;
  assign y161 = ~n504 ;
  assign y162 = ~n508 ;
  assign y163 = ~n509 ;
  assign y164 = n511 ;
  assign y165 = ~n515 ;
  assign y166 = n520 ;
  assign y167 = n521 ;
  assign y168 = ~1'b0 ;
  assign y169 = n529 ;
  assign y170 = ~n531 ;
  assign y171 = ~n535 ;
  assign y172 = n537 ;
  assign y173 = n543 ;
  assign y174 = ~n548 ;
  assign y175 = n553 ;
  assign y176 = ~n555 ;
  assign y177 = ~n557 ;
  assign y178 = n562 ;
  assign y179 = n565 ;
  assign y180 = ~1'b0 ;
  assign y181 = ~n568 ;
  assign y182 = ~n285 ;
  assign y183 = ~n569 ;
  assign y184 = ~n572 ;
  assign y185 = ~n579 ;
  assign y186 = n580 ;
  assign y187 = ~n584 ;
  assign y188 = n585 ;
  assign y189 = n586 ;
  assign y190 = n587 ;
  assign y191 = ~n593 ;
  assign y192 = n599 ;
  assign y193 = ~n613 ;
  assign y194 = n622 ;
  assign y195 = ~n624 ;
  assign y196 = ~x49 ;
  assign y197 = n625 ;
  assign y198 = ~1'b0 ;
  assign y199 = ~n630 ;
  assign y200 = ~n631 ;
  assign y201 = n634 ;
  assign y202 = ~1'b0 ;
  assign y203 = ~1'b0 ;
  assign y204 = n644 ;
  assign y205 = ~n646 ;
  assign y206 = ~n652 ;
  assign y207 = n653 ;
  assign y208 = ~n654 ;
  assign y209 = ~n660 ;
  assign y210 = ~n664 ;
  assign y211 = n670 ;
  assign y212 = n673 ;
  assign y213 = ~n685 ;
  assign y214 = ~1'b0 ;
  assign y215 = n688 ;
  assign y216 = ~n690 ;
  assign y217 = ~n693 ;
  assign y218 = ~n694 ;
  assign y219 = ~1'b0 ;
  assign y220 = n697 ;
  assign y221 = ~n700 ;
  assign y222 = n701 ;
  assign y223 = n293 ;
  assign y224 = n709 ;
  assign y225 = ~n711 ;
  assign y226 = ~1'b0 ;
  assign y227 = ~1'b0 ;
  assign y228 = n712 ;
  assign y229 = n714 ;
  assign y230 = ~n719 ;
  assign y231 = ~1'b0 ;
  assign y232 = ~n726 ;
  assign y233 = ~n727 ;
  assign y234 = ~n729 ;
  assign y235 = n732 ;
  assign y236 = ~1'b0 ;
  assign y237 = n739 ;
  assign y238 = n744 ;
  assign y239 = n746 ;
  assign y240 = ~n747 ;
  assign y241 = ~n751 ;
  assign y242 = n753 ;
  assign y243 = n763 ;
  assign y244 = n770 ;
  assign y245 = n773 ;
  assign y246 = ~1'b0 ;
  assign y247 = ~n778 ;
  assign y248 = ~n782 ;
  assign y249 = ~1'b0 ;
  assign y250 = ~1'b0 ;
  assign y251 = ~n148 ;
  assign y252 = ~n785 ;
  assign y253 = ~1'b0 ;
  assign y254 = ~1'b0 ;
  assign y255 = n786 ;
  assign y256 = n788 ;
  assign y257 = ~1'b0 ;
  assign y258 = n790 ;
  assign y259 = n793 ;
  assign y260 = ~n794 ;
  assign y261 = ~n795 ;
  assign y262 = n796 ;
  assign y263 = n799 ;
  assign y264 = ~1'b0 ;
  assign y265 = ~n801 ;
  assign y266 = ~1'b0 ;
  assign y267 = ~n803 ;
  assign y268 = ~n316 ;
  assign y269 = n805 ;
  assign y270 = ~n808 ;
  assign y271 = ~1'b0 ;
  assign y272 = n809 ;
  assign y273 = ~1'b0 ;
  assign y274 = ~n812 ;
  assign y275 = n823 ;
  assign y276 = ~n827 ;
  assign y277 = ~n832 ;
  assign y278 = n834 ;
  assign y279 = ~n841 ;
  assign y280 = ~1'b0 ;
  assign y281 = ~n844 ;
  assign y282 = ~n845 ;
  assign y283 = ~n847 ;
  assign y284 = n848 ;
  assign y285 = n857 ;
  assign y286 = ~n859 ;
  assign y287 = ~n860 ;
  assign y288 = n870 ;
  assign y289 = n872 ;
  assign y290 = n877 ;
  assign y291 = ~n879 ;
  assign y292 = n882 ;
  assign y293 = ~n836 ;
  assign y294 = ~n885 ;
  assign y295 = n887 ;
  assign y296 = ~n901 ;
  assign y297 = ~n904 ;
  assign y298 = ~n906 ;
  assign y299 = ~n909 ;
  assign y300 = ~n914 ;
  assign y301 = ~n923 ;
  assign y302 = n928 ;
  assign y303 = n934 ;
  assign y304 = n936 ;
  assign y305 = n937 ;
  assign y306 = ~n947 ;
  assign y307 = ~n953 ;
  assign y308 = n954 ;
  assign y309 = ~1'b0 ;
  assign y310 = ~1'b0 ;
  assign y311 = n960 ;
  assign y312 = ~n970 ;
  assign y313 = ~n986 ;
  assign y314 = ~n1002 ;
  assign y315 = ~1'b0 ;
  assign y316 = n1004 ;
  assign y317 = ~1'b0 ;
  assign y318 = ~n1011 ;
  assign y319 = ~n1015 ;
  assign y320 = ~n1017 ;
  assign y321 = ~1'b0 ;
  assign y322 = ~1'b0 ;
  assign y323 = n1018 ;
  assign y324 = n1031 ;
  assign y325 = n1033 ;
  assign y326 = n1036 ;
  assign y327 = n1039 ;
  assign y328 = n1042 ;
  assign y329 = n1047 ;
  assign y330 = ~n1055 ;
  assign y331 = ~1'b0 ;
  assign y332 = n1060 ;
  assign y333 = ~n1064 ;
  assign y334 = n1065 ;
  assign y335 = ~n1068 ;
  assign y336 = ~n1074 ;
  assign y337 = n1078 ;
  assign y338 = ~n1079 ;
  assign y339 = ~n1080 ;
  assign y340 = n1083 ;
  assign y341 = ~1'b0 ;
  assign y342 = ~n1086 ;
  assign y343 = n1090 ;
  assign y344 = n1098 ;
  assign y345 = ~1'b0 ;
  assign y346 = ~n1099 ;
  assign y347 = ~n1104 ;
  assign y348 = n1114 ;
  assign y349 = n1121 ;
  assign y350 = n1124 ;
  assign y351 = ~n1127 ;
  assign y352 = n1131 ;
  assign y353 = ~n1133 ;
  assign y354 = n1138 ;
  assign y355 = ~n1143 ;
  assign y356 = ~n1146 ;
  assign y357 = ~1'b0 ;
  assign y358 = n824 ;
  assign y359 = ~n1153 ;
  assign y360 = ~n744 ;
  assign y361 = n1157 ;
  assign y362 = ~1'b0 ;
  assign y363 = n1167 ;
  assign y364 = n1179 ;
  assign y365 = n1181 ;
  assign y366 = n1184 ;
  assign y367 = ~n1185 ;
  assign y368 = ~1'b0 ;
  assign y369 = ~n1188 ;
  assign y370 = ~1'b0 ;
  assign y371 = n1194 ;
  assign y372 = ~n1198 ;
  assign y373 = ~1'b0 ;
  assign y374 = n1199 ;
  assign y375 = ~1'b0 ;
  assign y376 = n1201 ;
  assign y377 = n1207 ;
  assign y378 = ~1'b0 ;
  assign y379 = ~n1211 ;
  assign y380 = n1221 ;
  assign y381 = ~n1224 ;
  assign y382 = n1227 ;
  assign y383 = ~n1234 ;
  assign y384 = n1236 ;
  assign y385 = ~1'b0 ;
  assign y386 = ~1'b0 ;
  assign y387 = ~n1253 ;
  assign y388 = n1257 ;
  assign y389 = n1259 ;
  assign y390 = n1268 ;
  assign y391 = ~n1271 ;
  assign y392 = n1274 ;
  assign y393 = n1281 ;
  assign y394 = n1288 ;
  assign y395 = ~1'b0 ;
  assign y396 = n1291 ;
  assign y397 = ~n1292 ;
  assign y398 = ~1'b0 ;
  assign y399 = ~n1297 ;
  assign y400 = ~n1299 ;
  assign y401 = ~1'b0 ;
  assign y402 = ~n1302 ;
  assign y403 = n1305 ;
  assign y404 = n1309 ;
  assign y405 = ~1'b0 ;
  assign y406 = ~n1314 ;
  assign y407 = ~n1316 ;
  assign y408 = ~1'b0 ;
  assign y409 = n1318 ;
  assign y410 = ~1'b0 ;
  assign y411 = ~n1320 ;
  assign y412 = n1322 ;
  assign y413 = ~1'b0 ;
  assign y414 = ~n1332 ;
  assign y415 = ~1'b0 ;
  assign y416 = ~1'b0 ;
  assign y417 = ~n1335 ;
  assign y418 = ~n1338 ;
  assign y419 = ~n1341 ;
  assign y420 = n1343 ;
  assign y421 = ~1'b0 ;
  assign y422 = ~n1349 ;
  assign y423 = n1351 ;
  assign y424 = ~n1363 ;
  assign y425 = n1365 ;
  assign y426 = ~n1368 ;
  assign y427 = ~n1374 ;
  assign y428 = n1376 ;
  assign y429 = ~n1381 ;
  assign y430 = ~1'b0 ;
  assign y431 = ~n1383 ;
  assign y432 = n1384 ;
  assign y433 = ~n1392 ;
  assign y434 = ~1'b0 ;
  assign y435 = ~1'b0 ;
  assign y436 = ~1'b0 ;
  assign y437 = n1394 ;
  assign y438 = ~1'b0 ;
  assign y439 = n1396 ;
  assign y440 = ~n1403 ;
  assign y441 = ~n1410 ;
  assign y442 = ~n1418 ;
  assign y443 = n1420 ;
  assign y444 = ~n1428 ;
  assign y445 = ~n1433 ;
  assign y446 = ~n1434 ;
  assign y447 = n1435 ;
  assign y448 = ~1'b0 ;
  assign y449 = 1'b0 ;
  assign y450 = n1440 ;
  assign y451 = n1441 ;
  assign y452 = n251 ;
  assign y453 = ~1'b0 ;
  assign y454 = ~x78 ;
  assign y455 = ~1'b0 ;
  assign y456 = ~1'b0 ;
  assign y457 = n1442 ;
  assign y458 = ~1'b0 ;
  assign y459 = ~n795 ;
  assign y460 = ~1'b0 ;
  assign y461 = n1448 ;
  assign y462 = ~1'b0 ;
  assign y463 = ~1'b0 ;
  assign y464 = ~n1449 ;
  assign y465 = ~n1462 ;
  assign y466 = n1465 ;
  assign y467 = n1467 ;
  assign y468 = ~1'b0 ;
  assign y469 = ~n1472 ;
  assign y470 = ~n1476 ;
  assign y471 = n1480 ;
  assign y472 = ~n1481 ;
  assign y473 = ~1'b0 ;
  assign y474 = ~n1485 ;
  assign y475 = n1489 ;
  assign y476 = ~1'b0 ;
  assign y477 = ~1'b0 ;
  assign y478 = n1491 ;
  assign y479 = ~n1496 ;
  assign y480 = n1497 ;
  assign y481 = n1498 ;
  assign y482 = ~1'b0 ;
  assign y483 = ~n1503 ;
  assign y484 = n1506 ;
  assign y485 = n1507 ;
  assign y486 = ~n1513 ;
  assign y487 = n1515 ;
  assign y488 = ~1'b0 ;
  assign y489 = ~1'b0 ;
  assign y490 = n1518 ;
  assign y491 = ~n1519 ;
  assign y492 = ~1'b0 ;
  assign y493 = ~n1524 ;
  assign y494 = ~1'b0 ;
  assign y495 = n968 ;
  assign y496 = n1525 ;
  assign y497 = ~1'b0 ;
  assign y498 = ~n1527 ;
  assign y499 = n1528 ;
  assign y500 = ~1'b0 ;
  assign y501 = ~n1529 ;
  assign y502 = n1535 ;
  assign y503 = n1537 ;
  assign y504 = n1543 ;
  assign y505 = ~1'b0 ;
  assign y506 = ~n1554 ;
  assign y507 = ~n1555 ;
  assign y508 = ~n1561 ;
  assign y509 = ~n1571 ;
  assign y510 = ~n1573 ;
  assign y511 = ~n1577 ;
  assign y512 = ~1'b0 ;
  assign y513 = ~n1589 ;
  assign y514 = ~n1596 ;
  assign y515 = ~n1600 ;
  assign y516 = ~n411 ;
  assign y517 = n1602 ;
  assign y518 = ~n1603 ;
  assign y519 = n1605 ;
  assign y520 = n1612 ;
  assign y521 = ~1'b0 ;
  assign y522 = n1613 ;
  assign y523 = ~n1614 ;
  assign y524 = ~1'b0 ;
  assign y525 = n1617 ;
  assign y526 = n1618 ;
  assign y527 = ~1'b0 ;
  assign y528 = n1619 ;
  assign y529 = ~n1622 ;
  assign y530 = n1626 ;
  assign y531 = ~n1629 ;
  assign y532 = ~1'b0 ;
  assign y533 = ~n1632 ;
  assign y534 = ~n1634 ;
  assign y535 = ~1'b0 ;
  assign y536 = n1636 ;
  assign y537 = ~1'b0 ;
  assign y538 = ~n1639 ;
  assign y539 = n1642 ;
  assign y540 = n1645 ;
  assign y541 = n1652 ;
  assign y542 = ~1'b0 ;
  assign y543 = ~1'b0 ;
  assign y544 = n1656 ;
  assign y545 = n1657 ;
  assign y546 = n1376 ;
  assign y547 = ~n1658 ;
  assign y548 = ~n1664 ;
  assign y549 = ~n1667 ;
  assign y550 = ~1'b0 ;
  assign y551 = ~n1671 ;
  assign y552 = ~n1673 ;
  assign y553 = n1678 ;
  assign y554 = ~n1679 ;
  assign y555 = x103 ;
  assign y556 = n1680 ;
  assign y557 = ~x123 ;
  assign y558 = ~1'b0 ;
  assign y559 = n1685 ;
  assign y560 = n1689 ;
  assign y561 = ~n1690 ;
  assign y562 = ~n1692 ;
  assign y563 = n1696 ;
  assign y564 = ~1'b0 ;
  assign y565 = ~1'b0 ;
  assign y566 = ~n1697 ;
  assign y567 = n1702 ;
  assign y568 = ~n1703 ;
  assign y569 = n1542 ;
  assign y570 = ~n1704 ;
  assign y571 = ~1'b0 ;
  assign y572 = ~n1710 ;
  assign y573 = ~n1713 ;
  assign y574 = ~n1718 ;
  assign y575 = ~n1726 ;
  assign y576 = ~n1727 ;
  assign y577 = n1731 ;
  assign y578 = n1732 ;
  assign y579 = ~n1739 ;
  assign y580 = n1740 ;
  assign y581 = n1752 ;
  assign y582 = ~n1758 ;
  assign y583 = n1759 ;
  assign y584 = ~n1767 ;
  assign y585 = ~1'b0 ;
  assign y586 = n1772 ;
  assign y587 = ~n1773 ;
  assign y588 = ~n1781 ;
  assign y589 = ~n1788 ;
  assign y590 = ~n1791 ;
  assign y591 = n1794 ;
  assign y592 = ~n1795 ;
  assign y593 = ~1'b0 ;
  assign y594 = 1'b0 ;
  assign y595 = n1797 ;
  assign y596 = n1802 ;
  assign y597 = ~n1806 ;
  assign y598 = ~n1818 ;
  assign y599 = ~n1820 ;
  assign y600 = ~n1828 ;
  assign y601 = n1829 ;
  assign y602 = ~n1832 ;
  assign y603 = ~n1834 ;
  assign y604 = n1836 ;
  assign y605 = n1837 ;
  assign y606 = n1842 ;
  assign y607 = n1848 ;
  assign y608 = n1850 ;
  assign y609 = n1855 ;
  assign y610 = n1860 ;
  assign y611 = ~n1861 ;
  assign y612 = ~1'b0 ;
  assign y613 = n1863 ;
  assign y614 = ~1'b0 ;
  assign y615 = ~1'b0 ;
  assign y616 = n1873 ;
  assign y617 = ~n1878 ;
  assign y618 = ~1'b0 ;
  assign y619 = ~n1884 ;
  assign y620 = ~n1515 ;
  assign y621 = ~n1890 ;
  assign y622 = ~n1892 ;
  assign y623 = ~1'b0 ;
  assign y624 = ~1'b0 ;
  assign y625 = ~n1895 ;
  assign y626 = ~n1900 ;
  assign y627 = ~n1906 ;
  assign y628 = ~n1910 ;
  assign y629 = n1917 ;
  assign y630 = ~n1919 ;
  assign y631 = 1'b0 ;
  assign y632 = 1'b0 ;
  assign y633 = ~n1920 ;
  assign y634 = ~1'b0 ;
  assign y635 = ~n1925 ;
  assign y636 = ~n1928 ;
  assign y637 = n1930 ;
  assign y638 = ~1'b0 ;
  assign y639 = ~n1938 ;
  assign y640 = n1939 ;
  assign y641 = n1943 ;
  assign y642 = ~n1953 ;
  assign y643 = ~1'b0 ;
  assign y644 = ~1'b0 ;
  assign y645 = ~n1959 ;
  assign y646 = n1962 ;
  assign y647 = ~n1974 ;
  assign y648 = ~1'b0 ;
  assign y649 = ~n1979 ;
  assign y650 = ~n1981 ;
  assign y651 = ~n992 ;
  assign y652 = n1983 ;
  assign y653 = n1984 ;
  assign y654 = n1988 ;
  assign y655 = ~n1993 ;
  assign y656 = ~n1162 ;
  assign y657 = n1996 ;
  assign y658 = n2007 ;
  assign y659 = n2008 ;
  assign y660 = ~n2009 ;
  assign y661 = ~n2011 ;
  assign y662 = ~n2017 ;
  assign y663 = n2026 ;
  assign y664 = ~1'b0 ;
  assign y665 = n2032 ;
  assign y666 = n2040 ;
  assign y667 = ~n2041 ;
  assign y668 = ~n2046 ;
  assign y669 = n2047 ;
  assign y670 = n1929 ;
  assign y671 = ~1'b0 ;
  assign y672 = n2048 ;
  assign y673 = n2054 ;
  assign y674 = ~n2059 ;
  assign y675 = n2060 ;
  assign y676 = ~n2062 ;
  assign y677 = ~1'b0 ;
  assign y678 = ~1'b0 ;
  assign y679 = n2063 ;
  assign y680 = n2064 ;
  assign y681 = ~n2066 ;
  assign y682 = ~n2069 ;
  assign y683 = n2070 ;
  assign y684 = ~n2074 ;
  assign y685 = ~n2078 ;
  assign y686 = ~n2084 ;
  assign y687 = ~n2086 ;
  assign y688 = ~n2097 ;
  assign y689 = ~1'b0 ;
  assign y690 = ~n2101 ;
  assign y691 = n2108 ;
  assign y692 = ~n2110 ;
  assign y693 = n2115 ;
  assign y694 = ~n2120 ;
  assign y695 = ~n2124 ;
  assign y696 = ~n2129 ;
  assign y697 = ~1'b0 ;
  assign y698 = ~1'b0 ;
  assign y699 = n2130 ;
  assign y700 = ~n2131 ;
  assign y701 = ~n2134 ;
  assign y702 = ~n2138 ;
  assign y703 = ~1'b0 ;
  assign y704 = ~1'b0 ;
  assign y705 = ~n2139 ;
  assign y706 = n2148 ;
  assign y707 = ~1'b0 ;
  assign y708 = ~1'b0 ;
  assign y709 = n2151 ;
  assign y710 = n2159 ;
  assign y711 = ~n2167 ;
  assign y712 = ~n2176 ;
  assign y713 = ~1'b0 ;
  assign y714 = ~n2179 ;
  assign y715 = ~n2181 ;
  assign y716 = ~n2183 ;
  assign y717 = n2187 ;
  assign y718 = n2195 ;
  assign y719 = n2197 ;
  assign y720 = n2201 ;
  assign y721 = ~n2202 ;
  assign y722 = ~1'b0 ;
  assign y723 = n2213 ;
  assign y724 = ~1'b0 ;
  assign y725 = ~1'b0 ;
  assign y726 = n2215 ;
  assign y727 = ~n2217 ;
  assign y728 = ~1'b0 ;
  assign y729 = ~n2218 ;
  assign y730 = n2219 ;
  assign y731 = ~n2222 ;
  assign y732 = ~n2228 ;
  assign y733 = ~n2231 ;
  assign y734 = ~n2235 ;
  assign y735 = n2239 ;
  assign y736 = ~n2243 ;
  assign y737 = ~n2256 ;
  assign y738 = n2267 ;
  assign y739 = n2269 ;
  assign y740 = ~1'b0 ;
  assign y741 = ~n2275 ;
  assign y742 = ~n2276 ;
  assign y743 = n2280 ;
  assign y744 = ~n2282 ;
  assign y745 = ~1'b0 ;
  assign y746 = n2283 ;
  assign y747 = ~n2285 ;
  assign y748 = ~n2286 ;
  assign y749 = ~n2288 ;
  assign y750 = ~n2310 ;
  assign y751 = n2320 ;
  assign y752 = ~1'b0 ;
  assign y753 = n2321 ;
  assign y754 = ~1'b0 ;
  assign y755 = ~n2324 ;
  assign y756 = n2326 ;
  assign y757 = n2332 ;
  assign y758 = ~n2340 ;
  assign y759 = ~n2347 ;
  assign y760 = ~n2359 ;
  assign y761 = n2368 ;
  assign y762 = n2372 ;
  assign y763 = ~n2374 ;
  assign y764 = ~1'b0 ;
  assign y765 = ~n2375 ;
  assign y766 = ~1'b0 ;
  assign y767 = n2381 ;
  assign y768 = n2387 ;
  assign y769 = n2388 ;
  assign y770 = ~n2389 ;
  assign y771 = ~n2393 ;
  assign y772 = ~1'b0 ;
  assign y773 = n2395 ;
  assign y774 = n2399 ;
  assign y775 = ~n2404 ;
  assign y776 = ~n2406 ;
  assign y777 = n2408 ;
  assign y778 = ~n2413 ;
  assign y779 = n2415 ;
  assign y780 = n2416 ;
  assign y781 = ~1'b0 ;
  assign y782 = ~n2427 ;
  assign y783 = ~n2438 ;
  assign y784 = ~n1150 ;
  assign y785 = n2441 ;
  assign y786 = n2444 ;
  assign y787 = ~1'b0 ;
  assign y788 = ~1'b0 ;
  assign y789 = ~n2447 ;
  assign y790 = x107 ;
  assign y791 = n2448 ;
  assign y792 = ~1'b0 ;
  assign y793 = n2450 ;
  assign y794 = n2455 ;
  assign y795 = ~1'b0 ;
  assign y796 = ~n2462 ;
  assign y797 = ~n2470 ;
  assign y798 = n2471 ;
  assign y799 = ~n2477 ;
  assign y800 = ~n2478 ;
  assign y801 = ~n2479 ;
  assign y802 = ~n2486 ;
  assign y803 = ~1'b0 ;
  assign y804 = n2487 ;
  assign y805 = n2488 ;
  assign y806 = n2492 ;
  assign y807 = ~n2494 ;
  assign y808 = ~1'b0 ;
  assign y809 = ~1'b0 ;
  assign y810 = n2499 ;
  assign y811 = n2500 ;
  assign y812 = ~1'b0 ;
  assign y813 = n2501 ;
  assign y814 = n1104 ;
  assign y815 = n2506 ;
  assign y816 = n2508 ;
  assign y817 = n2511 ;
  assign y818 = ~1'b0 ;
  assign y819 = n2514 ;
  assign y820 = ~1'b0 ;
  assign y821 = n2516 ;
  assign y822 = ~1'b0 ;
  assign y823 = ~1'b0 ;
  assign y824 = ~1'b0 ;
  assign y825 = n2526 ;
  assign y826 = n2527 ;
  assign y827 = n2536 ;
  assign y828 = ~1'b0 ;
  assign y829 = n2422 ;
  assign y830 = ~1'b0 ;
  assign y831 = n2542 ;
  assign y832 = ~n2544 ;
  assign y833 = ~n2547 ;
  assign y834 = ~n2551 ;
  assign y835 = ~n2563 ;
  assign y836 = n2566 ;
  assign y837 = ~1'b0 ;
  assign y838 = ~n2574 ;
  assign y839 = ~1'b0 ;
  assign y840 = n2577 ;
  assign y841 = ~1'b0 ;
  assign y842 = ~1'b0 ;
  assign y843 = ~n2580 ;
  assign y844 = n2582 ;
  assign y845 = n2584 ;
  assign y846 = ~1'b0 ;
  assign y847 = n2589 ;
  assign y848 = ~n2590 ;
  assign y849 = ~1'b0 ;
  assign y850 = ~1'b0 ;
  assign y851 = ~n2592 ;
  assign y852 = n2593 ;
  assign y853 = ~n2066 ;
  assign y854 = ~n2595 ;
  assign y855 = ~n2596 ;
  assign y856 = ~n2597 ;
  assign y857 = n2598 ;
  assign y858 = ~1'b0 ;
  assign y859 = ~1'b0 ;
  assign y860 = n2609 ;
  assign y861 = n2611 ;
  assign y862 = ~n2612 ;
  assign y863 = n2614 ;
  assign y864 = ~1'b0 ;
  assign y865 = ~n2616 ;
  assign y866 = ~n2619 ;
  assign y867 = ~1'b0 ;
  assign y868 = n1470 ;
  assign y869 = n2630 ;
  assign y870 = n2633 ;
  assign y871 = ~n2648 ;
  assign y872 = ~1'b0 ;
  assign y873 = ~n2655 ;
  assign y874 = ~n2660 ;
  assign y875 = n2661 ;
  assign y876 = ~n2664 ;
  assign y877 = ~n2670 ;
  assign y878 = ~n2677 ;
  assign y879 = ~1'b0 ;
  assign y880 = n2685 ;
  assign y881 = ~n2686 ;
  assign y882 = ~n2687 ;
  assign y883 = n2692 ;
  assign y884 = ~n2693 ;
  assign y885 = ~n2700 ;
  assign y886 = ~1'b0 ;
  assign y887 = ~n2709 ;
  assign y888 = ~n2716 ;
  assign y889 = ~1'b0 ;
  assign y890 = ~n2717 ;
  assign y891 = ~n2731 ;
  assign y892 = n2734 ;
  assign y893 = ~n2736 ;
  assign y894 = ~n2737 ;
  assign y895 = ~n2741 ;
  assign y896 = n2743 ;
  assign y897 = n2745 ;
  assign y898 = n2750 ;
  assign y899 = ~1'b0 ;
  assign y900 = n2751 ;
  assign y901 = ~n2755 ;
  assign y902 = ~1'b0 ;
  assign y903 = ~1'b0 ;
  assign y904 = ~n2758 ;
  assign y905 = ~n2759 ;
  assign y906 = ~1'b0 ;
  assign y907 = ~1'b0 ;
  assign y908 = ~1'b0 ;
  assign y909 = ~n2761 ;
  assign y910 = ~1'b0 ;
  assign y911 = ~1'b0 ;
  assign y912 = ~n579 ;
  assign y913 = ~n2771 ;
  assign y914 = n2779 ;
  assign y915 = ~n2781 ;
  assign y916 = ~n2782 ;
  assign y917 = n2783 ;
  assign y918 = n2798 ;
  assign y919 = n2799 ;
  assign y920 = ~n2801 ;
  assign y921 = n2804 ;
  assign y922 = ~n2817 ;
  assign y923 = n2819 ;
  assign y924 = n2820 ;
  assign y925 = n2822 ;
  assign y926 = ~1'b0 ;
  assign y927 = ~n2827 ;
  assign y928 = n2836 ;
  assign y929 = ~n2844 ;
  assign y930 = n2846 ;
  assign y931 = n2849 ;
  assign y932 = ~n2854 ;
  assign y933 = n2856 ;
  assign y934 = n2859 ;
  assign y935 = ~n2862 ;
  assign y936 = n2865 ;
  assign y937 = n2872 ;
  assign y938 = ~n2873 ;
  assign y939 = n2880 ;
  assign y940 = ~n2888 ;
  assign y941 = ~n2890 ;
  assign y942 = n2891 ;
  assign y943 = n2895 ;
  assign y944 = ~n2896 ;
  assign y945 = ~1'b0 ;
  assign y946 = n2898 ;
  assign y947 = ~n2900 ;
  assign y948 = ~n2904 ;
  assign y949 = n2907 ;
  assign y950 = ~1'b0 ;
  assign y951 = ~n2909 ;
  assign y952 = ~1'b0 ;
  assign y953 = ~1'b0 ;
  assign y954 = n2912 ;
  assign y955 = n2915 ;
  assign y956 = ~n2926 ;
  assign y957 = n2928 ;
  assign y958 = ~n2929 ;
  assign y959 = ~n2935 ;
  assign y960 = n2939 ;
  assign y961 = n2940 ;
  assign y962 = ~n2942 ;
  assign y963 = ~n2944 ;
  assign y964 = ~1'b0 ;
  assign y965 = ~n2946 ;
  assign y966 = ~1'b0 ;
  assign y967 = ~1'b0 ;
  assign y968 = n2956 ;
  assign y969 = ~1'b0 ;
  assign y970 = ~n2961 ;
  assign y971 = ~1'b0 ;
  assign y972 = ~n2969 ;
  assign y973 = ~1'b0 ;
  assign y974 = ~n2972 ;
  assign y975 = ~n2974 ;
  assign y976 = n2981 ;
  assign y977 = n2984 ;
  assign y978 = n2989 ;
  assign y979 = ~n2991 ;
  assign y980 = n2993 ;
  assign y981 = ~1'b0 ;
  assign y982 = n2995 ;
  assign y983 = ~1'b0 ;
  assign y984 = ~n3002 ;
  assign y985 = n3007 ;
  assign y986 = ~n3010 ;
  assign y987 = n3011 ;
  assign y988 = n3012 ;
  assign y989 = ~1'b0 ;
  assign y990 = ~1'b0 ;
  assign y991 = ~n3013 ;
  assign y992 = n3020 ;
  assign y993 = ~n3025 ;
  assign y994 = ~n3029 ;
  assign y995 = n3032 ;
  assign y996 = n3033 ;
  assign y997 = n1715 ;
  assign y998 = ~1'b0 ;
  assign y999 = ~1'b0 ;
  assign y1000 = n3035 ;
  assign y1001 = n3043 ;
  assign y1002 = ~n3044 ;
  assign y1003 = ~1'b0 ;
  assign y1004 = n3047 ;
  assign y1005 = n3049 ;
  assign y1006 = ~1'b0 ;
  assign y1007 = n3053 ;
  assign y1008 = ~1'b0 ;
  assign y1009 = ~1'b0 ;
  assign y1010 = n3054 ;
  assign y1011 = n3056 ;
  assign y1012 = n3059 ;
  assign y1013 = ~n3060 ;
  assign y1014 = n3062 ;
  assign y1015 = n3066 ;
  assign y1016 = ~1'b0 ;
  assign y1017 = n3068 ;
  assign y1018 = n3070 ;
  assign y1019 = n3076 ;
  assign y1020 = ~n2107 ;
  assign y1021 = n3084 ;
  assign y1022 = n3091 ;
  assign y1023 = ~n3092 ;
  assign y1024 = ~1'b0 ;
  assign y1025 = n3100 ;
  assign y1026 = ~n3114 ;
  assign y1027 = ~n3118 ;
  assign y1028 = ~1'b0 ;
  assign y1029 = n3119 ;
  assign y1030 = n3126 ;
  assign y1031 = ~n3127 ;
  assign y1032 = n3128 ;
  assign y1033 = ~n3129 ;
  assign y1034 = n3136 ;
  assign y1035 = ~1'b0 ;
  assign y1036 = ~n3139 ;
  assign y1037 = ~1'b0 ;
  assign y1038 = n3140 ;
  assign y1039 = ~n3141 ;
  assign y1040 = ~1'b0 ;
  assign y1041 = ~n3142 ;
  assign y1042 = n3149 ;
  assign y1043 = ~1'b0 ;
  assign y1044 = ~n3150 ;
  assign y1045 = ~1'b0 ;
  assign y1046 = n3155 ;
  assign y1047 = ~1'b0 ;
  assign y1048 = ~1'b0 ;
  assign y1049 = n3158 ;
  assign y1050 = n3159 ;
  assign y1051 = ~n3166 ;
  assign y1052 = n3171 ;
  assign y1053 = ~n3173 ;
  assign y1054 = ~n3176 ;
  assign y1055 = ~n3178 ;
  assign y1056 = ~1'b0 ;
  assign y1057 = n3181 ;
  assign y1058 = n3184 ;
  assign y1059 = ~n3185 ;
  assign y1060 = ~n3186 ;
  assign y1061 = ~n3191 ;
  assign y1062 = ~n3192 ;
  assign y1063 = ~n3196 ;
  assign y1064 = n3198 ;
  assign y1065 = n3203 ;
  assign y1066 = ~1'b0 ;
  assign y1067 = n3205 ;
  assign y1068 = ~n3215 ;
  assign y1069 = ~n3219 ;
  assign y1070 = ~n3224 ;
  assign y1071 = ~n3230 ;
  assign y1072 = ~n3232 ;
  assign y1073 = ~n3234 ;
  assign y1074 = ~1'b0 ;
  assign y1075 = ~1'b0 ;
  assign y1076 = n3236 ;
  assign y1077 = ~n3237 ;
  assign y1078 = n3238 ;
  assign y1079 = ~n3239 ;
  assign y1080 = n3241 ;
  assign y1081 = ~n3248 ;
  assign y1082 = n3254 ;
  assign y1083 = ~n3258 ;
  assign y1084 = ~n3263 ;
  assign y1085 = ~n3264 ;
  assign y1086 = ~n3275 ;
  assign y1087 = ~n3276 ;
  assign y1088 = ~n3281 ;
  assign y1089 = ~n3282 ;
  assign y1090 = ~1'b0 ;
  assign y1091 = ~n3284 ;
  assign y1092 = n3289 ;
  assign y1093 = ~1'b0 ;
  assign y1094 = ~n3294 ;
  assign y1095 = ~1'b0 ;
  assign y1096 = n1487 ;
  assign y1097 = n3298 ;
  assign y1098 = n3300 ;
  assign y1099 = ~1'b0 ;
  assign y1100 = n3302 ;
  assign y1101 = ~n3305 ;
  assign y1102 = n3308 ;
  assign y1103 = n2653 ;
  assign y1104 = ~1'b0 ;
  assign y1105 = n3312 ;
  assign y1106 = 1'b0 ;
  assign y1107 = ~n3314 ;
  assign y1108 = ~n3315 ;
  assign y1109 = n3317 ;
  assign y1110 = ~n3318 ;
  assign y1111 = ~n3320 ;
  assign y1112 = ~n3329 ;
  assign y1113 = n3334 ;
  assign y1114 = n3335 ;
  assign y1115 = n3338 ;
  assign y1116 = ~1'b0 ;
  assign y1117 = ~n3340 ;
  assign y1118 = ~n3348 ;
  assign y1119 = ~1'b0 ;
  assign y1120 = ~n3353 ;
  assign y1121 = ~n853 ;
  assign y1122 = n3362 ;
  assign y1123 = ~n3364 ;
  assign y1124 = ~n3367 ;
  assign y1125 = ~n3373 ;
  assign y1126 = ~1'b0 ;
  assign y1127 = ~n3390 ;
  assign y1128 = ~1'b0 ;
  assign y1129 = n3392 ;
  assign y1130 = n3398 ;
  assign y1131 = ~1'b0 ;
  assign y1132 = ~n3399 ;
  assign y1133 = ~n3401 ;
  assign y1134 = ~1'b0 ;
  assign y1135 = ~n3404 ;
  assign y1136 = ~n3406 ;
  assign y1137 = ~n3413 ;
  assign y1138 = ~1'b0 ;
  assign y1139 = ~n3416 ;
  assign y1140 = ~1'b0 ;
  assign y1141 = n3417 ;
  assign y1142 = n3421 ;
  assign y1143 = ~n3430 ;
  assign y1144 = ~n3433 ;
  assign y1145 = n1257 ;
  assign y1146 = ~n3441 ;
  assign y1147 = ~n3446 ;
  assign y1148 = ~n3449 ;
  assign y1149 = ~n3452 ;
  assign y1150 = ~1'b0 ;
  assign y1151 = ~n3455 ;
  assign y1152 = n3459 ;
  assign y1153 = ~1'b0 ;
  assign y1154 = ~n3465 ;
  assign y1155 = n3466 ;
  assign y1156 = ~n3467 ;
  assign y1157 = ~1'b0 ;
  assign y1158 = ~1'b0 ;
  assign y1159 = ~n3469 ;
  assign y1160 = ~n3470 ;
  assign y1161 = ~n3471 ;
  assign y1162 = n3474 ;
  assign y1163 = n3478 ;
  assign y1164 = n3479 ;
  assign y1165 = ~1'b0 ;
  assign y1166 = n3483 ;
  assign y1167 = ~n3488 ;
  assign y1168 = ~n3493 ;
  assign y1169 = n3494 ;
  assign y1170 = n3496 ;
  assign y1171 = ~n3501 ;
  assign y1172 = ~n3504 ;
  assign y1173 = ~n3509 ;
  assign y1174 = ~n3514 ;
  assign y1175 = n3515 ;
  assign y1176 = ~n3517 ;
  assign y1177 = ~n3519 ;
  assign y1178 = n3524 ;
  assign y1179 = n3526 ;
  assign y1180 = ~n3528 ;
  assign y1181 = ~n3530 ;
  assign y1182 = ~1'b0 ;
  assign y1183 = ~n3541 ;
  assign y1184 = ~n3543 ;
  assign y1185 = ~n3546 ;
  assign y1186 = n3548 ;
  assign y1187 = n3551 ;
  assign y1188 = ~n3552 ;
  assign y1189 = ~n3560 ;
  assign y1190 = ~n3561 ;
  assign y1191 = ~n3570 ;
  assign y1192 = ~n3575 ;
  assign y1193 = ~n3578 ;
  assign y1194 = ~n3587 ;
  assign y1195 = n3594 ;
  assign y1196 = n3597 ;
  assign y1197 = ~n3598 ;
  assign y1198 = ~n3599 ;
  assign y1199 = n3608 ;
  assign y1200 = ~n3611 ;
  assign y1201 = ~n3612 ;
  assign y1202 = n3614 ;
  assign y1203 = ~n3615 ;
  assign y1204 = ~n3621 ;
  assign y1205 = ~n3622 ;
  assign y1206 = n1448 ;
  assign y1207 = ~n3626 ;
  assign y1208 = ~n3629 ;
  assign y1209 = ~1'b0 ;
  assign y1210 = ~n3649 ;
  assign y1211 = ~n3652 ;
  assign y1212 = ~n3654 ;
  assign y1213 = ~n3657 ;
  assign y1214 = n3658 ;
  assign y1215 = ~n3659 ;
  assign y1216 = n3664 ;
  assign y1217 = ~n3666 ;
  assign y1218 = n3669 ;
  assign y1219 = ~1'b0 ;
  assign y1220 = ~n3671 ;
  assign y1221 = ~1'b0 ;
  assign y1222 = n3673 ;
  assign y1223 = n3316 ;
  assign y1224 = n3676 ;
  assign y1225 = ~1'b0 ;
  assign y1226 = n3677 ;
  assign y1227 = n3681 ;
  assign y1228 = n3695 ;
  assign y1229 = n3696 ;
  assign y1230 = n1491 ;
  assign y1231 = ~n3704 ;
  assign y1232 = n3706 ;
  assign y1233 = ~n3711 ;
  assign y1234 = ~n3713 ;
  assign y1235 = n3714 ;
  assign y1236 = ~n3720 ;
  assign y1237 = n3723 ;
  assign y1238 = n3726 ;
  assign y1239 = ~n3730 ;
  assign y1240 = n3731 ;
  assign y1241 = ~1'b0 ;
  assign y1242 = 1'b0 ;
  assign y1243 = ~1'b0 ;
  assign y1244 = ~n3732 ;
  assign y1245 = ~n3737 ;
  assign y1246 = ~n3743 ;
  assign y1247 = ~1'b0 ;
  assign y1248 = ~1'b0 ;
  assign y1249 = ~n3748 ;
  assign y1250 = ~n3755 ;
  assign y1251 = ~n3760 ;
  assign y1252 = n3762 ;
  assign y1253 = n3766 ;
  assign y1254 = ~n3769 ;
  assign y1255 = n3770 ;
  assign y1256 = n3771 ;
  assign y1257 = n3772 ;
  assign y1258 = ~1'b0 ;
  assign y1259 = n3778 ;
  assign y1260 = ~n3779 ;
  assign y1261 = n1305 ;
  assign y1262 = ~1'b0 ;
  assign y1263 = n3780 ;
  assign y1264 = ~1'b0 ;
  assign y1265 = ~1'b0 ;
  assign y1266 = n3781 ;
  assign y1267 = n3783 ;
  assign y1268 = ~1'b0 ;
  assign y1269 = ~1'b0 ;
  assign y1270 = ~1'b0 ;
  assign y1271 = ~n3784 ;
  assign y1272 = ~n3811 ;
  assign y1273 = ~1'b0 ;
  assign y1274 = ~1'b0 ;
  assign y1275 = ~n3814 ;
  assign y1276 = ~1'b0 ;
  assign y1277 = ~n3815 ;
  assign y1278 = ~n3820 ;
  assign y1279 = ~1'b0 ;
  assign y1280 = n3823 ;
  assign y1281 = n3824 ;
  assign y1282 = n402 ;
  assign y1283 = ~n3826 ;
  assign y1284 = 1'b0 ;
  assign y1285 = ~n3828 ;
  assign y1286 = ~n3836 ;
  assign y1287 = ~1'b0 ;
  assign y1288 = ~1'b0 ;
  assign y1289 = ~n3838 ;
  assign y1290 = n3840 ;
  assign y1291 = n3842 ;
  assign y1292 = ~1'b0 ;
  assign y1293 = n3847 ;
  assign y1294 = ~n3676 ;
  assign y1295 = ~n3848 ;
  assign y1296 = ~1'b0 ;
  assign y1297 = ~1'b0 ;
  assign y1298 = ~n3851 ;
  assign y1299 = ~n3853 ;
  assign y1300 = ~n3855 ;
  assign y1301 = ~1'b0 ;
  assign y1302 = n3863 ;
  assign y1303 = ~n3876 ;
  assign y1304 = ~n477 ;
  assign y1305 = ~n3883 ;
  assign y1306 = ~n3886 ;
  assign y1307 = ~n3888 ;
  assign y1308 = ~n3892 ;
  assign y1309 = n3894 ;
  assign y1310 = ~n1748 ;
  assign y1311 = n3896 ;
  assign y1312 = n3902 ;
  assign y1313 = ~n3905 ;
  assign y1314 = ~1'b0 ;
  assign y1315 = ~n2933 ;
  assign y1316 = ~n3908 ;
  assign y1317 = n3912 ;
  assign y1318 = n3916 ;
  assign y1319 = n3919 ;
  assign y1320 = n3920 ;
  assign y1321 = n3931 ;
  assign y1322 = ~1'b0 ;
  assign y1323 = ~n3934 ;
  assign y1324 = ~1'b0 ;
  assign y1325 = n3935 ;
  assign y1326 = n3941 ;
  assign y1327 = ~1'b0 ;
  assign y1328 = n3942 ;
  assign y1329 = n3943 ;
  assign y1330 = n2592 ;
  assign y1331 = n3946 ;
  assign y1332 = ~n3947 ;
  assign y1333 = ~n3955 ;
  assign y1334 = ~n3960 ;
  assign y1335 = n3962 ;
  assign y1336 = n3973 ;
  assign y1337 = ~n3987 ;
  assign y1338 = n3988 ;
  assign y1339 = ~1'b0 ;
  assign y1340 = ~n3989 ;
  assign y1341 = ~n3993 ;
  assign y1342 = n3994 ;
  assign y1343 = ~n3995 ;
  assign y1344 = ~n3997 ;
  assign y1345 = n4006 ;
  assign y1346 = ~1'b0 ;
  assign y1347 = n4009 ;
  assign y1348 = ~n4010 ;
  assign y1349 = ~n4015 ;
  assign y1350 = ~n4021 ;
  assign y1351 = ~n4031 ;
  assign y1352 = n4042 ;
  assign y1353 = ~n4046 ;
  assign y1354 = ~n4050 ;
  assign y1355 = ~n4052 ;
  assign y1356 = ~1'b0 ;
  assign y1357 = n4065 ;
  assign y1358 = ~n4066 ;
  assign y1359 = ~n4067 ;
  assign y1360 = n4074 ;
  assign y1361 = ~1'b0 ;
  assign y1362 = n4079 ;
  assign y1363 = ~n4084 ;
  assign y1364 = ~n4086 ;
  assign y1365 = ~n4087 ;
  assign y1366 = ~1'b0 ;
  assign y1367 = n3836 ;
  assign y1368 = n4088 ;
  assign y1369 = n4090 ;
  assign y1370 = n4097 ;
  assign y1371 = n4110 ;
  assign y1372 = n4111 ;
  assign y1373 = ~n4112 ;
  assign y1374 = ~1'b0 ;
  assign y1375 = n4119 ;
  assign y1376 = ~n4121 ;
  assign y1377 = ~n4122 ;
  assign y1378 = n4123 ;
  assign y1379 = n4125 ;
  assign y1380 = ~n4128 ;
  assign y1381 = ~n4130 ;
  assign y1382 = ~n4131 ;
  assign y1383 = ~n4133 ;
  assign y1384 = n4134 ;
  assign y1385 = n4137 ;
  assign y1386 = ~n4149 ;
  assign y1387 = n4156 ;
  assign y1388 = ~n4163 ;
  assign y1389 = 1'b0 ;
  assign y1390 = ~1'b0 ;
  assign y1391 = n4167 ;
  assign y1392 = ~1'b0 ;
  assign y1393 = n4172 ;
  assign y1394 = ~n4174 ;
  assign y1395 = ~1'b0 ;
  assign y1396 = ~n4175 ;
  assign y1397 = ~n4179 ;
  assign y1398 = ~1'b0 ;
  assign y1399 = ~n4181 ;
  assign y1400 = ~n4185 ;
  assign y1401 = n4188 ;
  assign y1402 = ~n4193 ;
  assign y1403 = n4195 ;
  assign y1404 = ~n4201 ;
  assign y1405 = n4204 ;
  assign y1406 = ~1'b0 ;
  assign y1407 = n4208 ;
  assign y1408 = n2552 ;
  assign y1409 = n4216 ;
  assign y1410 = ~1'b0 ;
  assign y1411 = n4217 ;
  assign y1412 = ~n4221 ;
  assign y1413 = ~n4226 ;
  assign y1414 = ~1'b0 ;
  assign y1415 = n4231 ;
  assign y1416 = ~n4238 ;
  assign y1417 = ~n4239 ;
  assign y1418 = n4247 ;
  assign y1419 = ~1'b0 ;
  assign y1420 = ~n4253 ;
  assign y1421 = ~n4257 ;
  assign y1422 = ~1'b0 ;
  assign y1423 = n4261 ;
  assign y1424 = n4284 ;
  assign y1425 = ~n4288 ;
  assign y1426 = n4292 ;
  assign y1427 = ~n4296 ;
  assign y1428 = n4298 ;
  assign y1429 = n4303 ;
  assign y1430 = ~n4306 ;
  assign y1431 = n4308 ;
  assign y1432 = ~n4324 ;
  assign y1433 = n4328 ;
  assign y1434 = ~1'b0 ;
  assign y1435 = n4330 ;
  assign y1436 = n4334 ;
  assign y1437 = n4337 ;
  assign y1438 = 1'b0 ;
  assign y1439 = n4338 ;
  assign y1440 = n4343 ;
  assign y1441 = n4350 ;
  assign y1442 = n3035 ;
  assign y1443 = ~1'b0 ;
  assign y1444 = n4354 ;
  assign y1445 = ~n4355 ;
  assign y1446 = ~1'b0 ;
  assign y1447 = ~1'b0 ;
  assign y1448 = n4358 ;
  assign y1449 = ~1'b0 ;
  assign y1450 = n4360 ;
  assign y1451 = ~n4361 ;
  assign y1452 = n4370 ;
  assign y1453 = ~n4372 ;
  assign y1454 = ~n4373 ;
  assign y1455 = ~1'b0 ;
  assign y1456 = n4378 ;
  assign y1457 = n4380 ;
  assign y1458 = n4382 ;
  assign y1459 = n4383 ;
  assign y1460 = ~1'b0 ;
  assign y1461 = ~n4384 ;
  assign y1462 = ~n4388 ;
  assign y1463 = ~1'b0 ;
  assign y1464 = n4389 ;
  assign y1465 = ~n4404 ;
  assign y1466 = ~n4094 ;
  assign y1467 = ~1'b0 ;
  assign y1468 = ~n4411 ;
  assign y1469 = n4413 ;
  assign y1470 = n4414 ;
  assign y1471 = ~n4415 ;
  assign y1472 = n4417 ;
  assign y1473 = ~n4422 ;
  assign y1474 = ~n4426 ;
  assign y1475 = n4428 ;
  assign y1476 = ~n4430 ;
  assign y1477 = ~1'b0 ;
  assign y1478 = ~n4434 ;
  assign y1479 = ~n4441 ;
  assign y1480 = ~1'b0 ;
  assign y1481 = n4443 ;
  assign y1482 = ~n4446 ;
  assign y1483 = n4447 ;
  assign y1484 = ~1'b0 ;
  assign y1485 = n4449 ;
  assign y1486 = ~n4450 ;
  assign y1487 = n4452 ;
  assign y1488 = ~n4455 ;
  assign y1489 = n4461 ;
  assign y1490 = ~n4465 ;
  assign y1491 = ~1'b0 ;
  assign y1492 = ~n4468 ;
  assign y1493 = n4476 ;
  assign y1494 = ~1'b0 ;
  assign y1495 = n4478 ;
  assign y1496 = n4479 ;
  assign y1497 = ~n4480 ;
  assign y1498 = ~1'b0 ;
  assign y1499 = ~n4482 ;
  assign y1500 = ~n4483 ;
  assign y1501 = ~n4484 ;
  assign y1502 = n4487 ;
  assign y1503 = ~n4490 ;
  assign y1504 = n1854 ;
  assign y1505 = ~1'b0 ;
  assign y1506 = ~n4494 ;
  assign y1507 = n4497 ;
  assign y1508 = ~n4498 ;
  assign y1509 = ~1'b0 ;
  assign y1510 = ~n4499 ;
  assign y1511 = n4501 ;
  assign y1512 = ~n4504 ;
  assign y1513 = ~n4510 ;
  assign y1514 = n4512 ;
  assign y1515 = n4513 ;
  assign y1516 = n4517 ;
  assign y1517 = n4519 ;
  assign y1518 = ~n4524 ;
  assign y1519 = n4525 ;
  assign y1520 = n4526 ;
  assign y1521 = n4527 ;
  assign y1522 = n4542 ;
  assign y1523 = ~1'b0 ;
  assign y1524 = ~n4543 ;
  assign y1525 = ~n4544 ;
  assign y1526 = ~n4552 ;
  assign y1527 = ~n4553 ;
  assign y1528 = n4555 ;
  assign y1529 = ~n4557 ;
  assign y1530 = ~1'b0 ;
  assign y1531 = ~1'b0 ;
  assign y1532 = n4559 ;
  assign y1533 = ~1'b0 ;
  assign y1534 = ~n4562 ;
  assign y1535 = ~n2930 ;
  assign y1536 = n4572 ;
  assign y1537 = ~n4576 ;
  assign y1538 = n4580 ;
  assign y1539 = n4588 ;
  assign y1540 = ~n4590 ;
  assign y1541 = n4594 ;
  assign y1542 = n4598 ;
  assign y1543 = ~n4600 ;
  assign y1544 = n4608 ;
  assign y1545 = ~1'b0 ;
  assign y1546 = ~n4612 ;
  assign y1547 = ~n4615 ;
  assign y1548 = n4625 ;
  assign y1549 = ~1'b0 ;
  assign y1550 = ~n4644 ;
  assign y1551 = n4647 ;
  assign y1552 = n4649 ;
  assign y1553 = ~1'b0 ;
  assign y1554 = ~n4650 ;
  assign y1555 = ~n4653 ;
  assign y1556 = ~n4657 ;
  assign y1557 = n4660 ;
  assign y1558 = ~n4661 ;
  assign y1559 = ~n4662 ;
  assign y1560 = ~1'b0 ;
  assign y1561 = n3044 ;
  assign y1562 = ~n4671 ;
  assign y1563 = n4673 ;
  assign y1564 = n4679 ;
  assign y1565 = n4680 ;
  assign y1566 = ~1'b0 ;
  assign y1567 = n4681 ;
  assign y1568 = ~n4687 ;
  assign y1569 = ~n4696 ;
  assign y1570 = ~n4697 ;
  assign y1571 = n4700 ;
  assign y1572 = ~n4704 ;
  assign y1573 = n4707 ;
  assign y1574 = ~n4710 ;
  assign y1575 = ~1'b0 ;
  assign y1576 = ~n4713 ;
  assign y1577 = n4714 ;
  assign y1578 = ~n4716 ;
  assign y1579 = ~1'b0 ;
  assign y1580 = n4718 ;
  assign y1581 = n4720 ;
  assign y1582 = n4724 ;
  assign y1583 = ~n4726 ;
  assign y1584 = ~1'b0 ;
  assign y1585 = n4728 ;
  assign y1586 = n4733 ;
  assign y1587 = ~n4741 ;
  assign y1588 = ~1'b0 ;
  assign y1589 = n4743 ;
  assign y1590 = ~1'b0 ;
  assign y1591 = ~1'b0 ;
  assign y1592 = ~n4745 ;
  assign y1593 = ~n4748 ;
  assign y1594 = ~n4754 ;
  assign y1595 = n4756 ;
  assign y1596 = ~n4757 ;
  assign y1597 = n4762 ;
  assign y1598 = n4768 ;
  assign y1599 = n4770 ;
  assign y1600 = n4772 ;
  assign y1601 = ~n4777 ;
  assign y1602 = n4778 ;
  assign y1603 = ~n2748 ;
  assign y1604 = n4783 ;
  assign y1605 = n4785 ;
  assign y1606 = ~n4789 ;
  assign y1607 = ~n4790 ;
  assign y1608 = ~1'b0 ;
  assign y1609 = ~n4794 ;
  assign y1610 = n4797 ;
  assign y1611 = ~n4801 ;
  assign y1612 = ~n4803 ;
  assign y1613 = ~n4808 ;
  assign y1614 = n4810 ;
  assign y1615 = ~1'b0 ;
  assign y1616 = ~n4811 ;
  assign y1617 = ~n4819 ;
  assign y1618 = n4822 ;
  assign y1619 = ~n4828 ;
  assign y1620 = ~n4832 ;
  assign y1621 = ~n4835 ;
  assign y1622 = ~1'b0 ;
  assign y1623 = ~n4843 ;
  assign y1624 = n4849 ;
  assign y1625 = ~n4850 ;
  assign y1626 = ~n4852 ;
  assign y1627 = ~n4859 ;
  assign y1628 = ~n4860 ;
  assign y1629 = ~1'b0 ;
  assign y1630 = ~n4861 ;
  assign y1631 = ~1'b0 ;
  assign y1632 = ~n4868 ;
  assign y1633 = ~n4875 ;
  assign y1634 = ~1'b0 ;
  assign y1635 = ~n4882 ;
  assign y1636 = ~n4884 ;
  assign y1637 = n4889 ;
  assign y1638 = n4896 ;
  assign y1639 = ~n4899 ;
  assign y1640 = n4901 ;
  assign y1641 = ~n4906 ;
  assign y1642 = n4909 ;
  assign y1643 = n4913 ;
  assign y1644 = n4216 ;
  assign y1645 = ~n4914 ;
  assign y1646 = ~1'b0 ;
  assign y1647 = ~n4916 ;
  assign y1648 = ~n4924 ;
  assign y1649 = ~n4925 ;
  assign y1650 = n1842 ;
  assign y1651 = ~1'b0 ;
  assign y1652 = ~n4933 ;
  assign y1653 = ~n4934 ;
  assign y1654 = ~n4938 ;
  assign y1655 = ~n4939 ;
  assign y1656 = ~1'b0 ;
  assign y1657 = ~n4941 ;
  assign y1658 = 1'b0 ;
  assign y1659 = ~n4943 ;
  assign y1660 = ~n4948 ;
  assign y1661 = ~n4954 ;
  assign y1662 = ~n4958 ;
  assign y1663 = n4961 ;
  assign y1664 = ~n4964 ;
  assign y1665 = n4966 ;
  assign y1666 = ~n4967 ;
  assign y1667 = ~n1203 ;
  assign y1668 = n4975 ;
  assign y1669 = n4978 ;
  assign y1670 = ~n4979 ;
  assign y1671 = ~n4983 ;
  assign y1672 = ~n4986 ;
  assign y1673 = n4988 ;
  assign y1674 = n4989 ;
  assign y1675 = ~n4993 ;
  assign y1676 = ~n4994 ;
  assign y1677 = n4997 ;
  assign y1678 = n3503 ;
  assign y1679 = n4999 ;
  assign y1680 = n5002 ;
  assign y1681 = n5003 ;
  assign y1682 = ~1'b0 ;
  assign y1683 = ~n5011 ;
  assign y1684 = ~n5012 ;
  assign y1685 = n5018 ;
  assign y1686 = n5022 ;
  assign y1687 = ~n5026 ;
  assign y1688 = n5037 ;
  assign y1689 = n5038 ;
  assign y1690 = n5040 ;
  assign y1691 = ~n5041 ;
  assign y1692 = n5044 ;
  assign y1693 = ~1'b0 ;
  assign y1694 = ~n5045 ;
  assign y1695 = n5048 ;
  assign y1696 = ~1'b0 ;
  assign y1697 = n5051 ;
  assign y1698 = ~n5053 ;
  assign y1699 = n5054 ;
  assign y1700 = ~n5056 ;
  assign y1701 = ~n5057 ;
  assign y1702 = n5061 ;
  assign y1703 = ~1'b0 ;
  assign y1704 = n5065 ;
  assign y1705 = n5066 ;
  assign y1706 = ~1'b0 ;
  assign y1707 = ~1'b0 ;
  assign y1708 = n5068 ;
  assign y1709 = n5070 ;
  assign y1710 = n5076 ;
  assign y1711 = ~1'b0 ;
  assign y1712 = ~n5081 ;
  assign y1713 = ~n5087 ;
  assign y1714 = ~n5089 ;
  assign y1715 = ~n5090 ;
  assign y1716 = ~n5104 ;
  assign y1717 = n5108 ;
  assign y1718 = ~n5112 ;
  assign y1719 = ~n5113 ;
  assign y1720 = ~1'b0 ;
  assign y1721 = n5116 ;
  assign y1722 = n5125 ;
  assign y1723 = n5131 ;
  assign y1724 = ~n5134 ;
  assign y1725 = n5145 ;
  assign y1726 = ~1'b0 ;
  assign y1727 = ~n5154 ;
  assign y1728 = ~n5156 ;
  assign y1729 = n5158 ;
  assign y1730 = ~1'b0 ;
  assign y1731 = n5160 ;
  assign y1732 = ~n5161 ;
  assign y1733 = ~1'b0 ;
  assign y1734 = ~n5165 ;
  assign y1735 = ~n2538 ;
  assign y1736 = ~1'b0 ;
  assign y1737 = n5167 ;
  assign y1738 = ~n5170 ;
  assign y1739 = ~n5172 ;
  assign y1740 = ~n5176 ;
  assign y1741 = ~n5178 ;
  assign y1742 = ~n5180 ;
  assign y1743 = ~1'b0 ;
  assign y1744 = n5192 ;
  assign y1745 = ~n5196 ;
  assign y1746 = ~1'b0 ;
  assign y1747 = ~1'b0 ;
  assign y1748 = n5198 ;
  assign y1749 = n5199 ;
  assign y1750 = n5202 ;
  assign y1751 = ~n4586 ;
  assign y1752 = ~n5208 ;
  assign y1753 = n5210 ;
  assign y1754 = ~1'b0 ;
  assign y1755 = n5213 ;
  assign y1756 = ~n5224 ;
  assign y1757 = n5225 ;
  assign y1758 = n5227 ;
  assign y1759 = ~n5231 ;
  assign y1760 = ~n5233 ;
  assign y1761 = ~n5234 ;
  assign y1762 = ~n5235 ;
  assign y1763 = ~n5236 ;
  assign y1764 = ~n5237 ;
  assign y1765 = n5242 ;
  assign y1766 = ~n5243 ;
  assign y1767 = n5246 ;
  assign y1768 = ~n5256 ;
  assign y1769 = ~n5264 ;
  assign y1770 = ~n5270 ;
  assign y1771 = ~1'b0 ;
  assign y1772 = ~n5272 ;
  assign y1773 = ~n5279 ;
  assign y1774 = ~n5281 ;
  assign y1775 = n5283 ;
  assign y1776 = n5285 ;
  assign y1777 = n5286 ;
  assign y1778 = ~n5287 ;
  assign y1779 = n5293 ;
  assign y1780 = ~1'b0 ;
  assign y1781 = ~1'b0 ;
  assign y1782 = n5294 ;
  assign y1783 = n5300 ;
  assign y1784 = ~n5303 ;
  assign y1785 = ~1'b0 ;
  assign y1786 = ~n5305 ;
  assign y1787 = ~n5308 ;
  assign y1788 = ~1'b0 ;
  assign y1789 = ~n5313 ;
  assign y1790 = n5314 ;
  assign y1791 = n5315 ;
  assign y1792 = ~n5316 ;
  assign y1793 = ~n377 ;
  assign y1794 = ~n5320 ;
  assign y1795 = n5323 ;
  assign y1796 = ~n5327 ;
  assign y1797 = ~n5328 ;
  assign y1798 = ~n5329 ;
  assign y1799 = ~n5331 ;
  assign y1800 = n5332 ;
  assign y1801 = n3726 ;
  assign y1802 = n5333 ;
  assign y1803 = ~1'b0 ;
  assign y1804 = n5347 ;
  assign y1805 = ~n5354 ;
  assign y1806 = ~n5360 ;
  assign y1807 = ~n5366 ;
  assign y1808 = ~n5370 ;
  assign y1809 = ~n5372 ;
  assign y1810 = n5378 ;
  assign y1811 = n5384 ;
  assign y1812 = ~n5387 ;
  assign y1813 = n5393 ;
  assign y1814 = n5394 ;
  assign y1815 = ~n5399 ;
  assign y1816 = n5403 ;
  assign y1817 = ~n5404 ;
  assign y1818 = ~n5406 ;
  assign y1819 = ~n5414 ;
  assign y1820 = n5419 ;
  assign y1821 = n5422 ;
  assign y1822 = ~1'b0 ;
  assign y1823 = ~1'b0 ;
  assign y1824 = ~n5423 ;
  assign y1825 = ~n5426 ;
  assign y1826 = ~1'b0 ;
  assign y1827 = ~n5436 ;
  assign y1828 = ~n5439 ;
  assign y1829 = ~n1712 ;
  assign y1830 = ~1'b0 ;
  assign y1831 = ~n5442 ;
  assign y1832 = n5443 ;
  assign y1833 = n5448 ;
  assign y1834 = n5453 ;
  assign y1835 = ~1'b0 ;
  assign y1836 = ~n5457 ;
  assign y1837 = n5458 ;
  assign y1838 = n5459 ;
  assign y1839 = n5462 ;
  assign y1840 = ~n5471 ;
  assign y1841 = ~n5475 ;
  assign y1842 = ~1'b0 ;
  assign y1843 = n5478 ;
  assign y1844 = ~n5482 ;
  assign y1845 = ~1'b0 ;
  assign y1846 = ~n5487 ;
  assign y1847 = ~n5488 ;
  assign y1848 = ~1'b0 ;
  assign y1849 = ~n5493 ;
  assign y1850 = n5501 ;
  assign y1851 = ~n5504 ;
  assign y1852 = ~1'b0 ;
  assign y1853 = ~n5506 ;
  assign y1854 = ~n5513 ;
  assign y1855 = ~1'b0 ;
  assign y1856 = n5514 ;
  assign y1857 = ~n5519 ;
  assign y1858 = n5520 ;
  assign y1859 = ~n5522 ;
  assign y1860 = ~n5530 ;
  assign y1861 = ~n5532 ;
  assign y1862 = n5533 ;
  assign y1863 = ~n5536 ;
  assign y1864 = n5538 ;
  assign y1865 = ~n3611 ;
  assign y1866 = n5539 ;
  assign y1867 = ~n5540 ;
  assign y1868 = n5543 ;
  assign y1869 = ~1'b0 ;
  assign y1870 = ~n5544 ;
  assign y1871 = ~n5550 ;
  assign y1872 = ~n5552 ;
  assign y1873 = ~n5557 ;
  assign y1874 = ~1'b0 ;
  assign y1875 = 1'b0 ;
  assign y1876 = ~1'b0 ;
  assign y1877 = ~1'b0 ;
  assign y1878 = ~1'b0 ;
  assign y1879 = ~n5558 ;
  assign y1880 = ~n1196 ;
  assign y1881 = ~n2499 ;
  assign y1882 = n5561 ;
  assign y1883 = ~n5566 ;
  assign y1884 = ~n5570 ;
  assign y1885 = ~1'b0 ;
  assign y1886 = n5574 ;
  assign y1887 = ~n5575 ;
  assign y1888 = ~n5576 ;
  assign y1889 = n5578 ;
  assign y1890 = ~n5580 ;
  assign y1891 = ~n2361 ;
  assign y1892 = ~n5582 ;
  assign y1893 = n5585 ;
  assign y1894 = ~n432 ;
  assign y1895 = ~1'b0 ;
  assign y1896 = n5586 ;
  assign y1897 = n3581 ;
  assign y1898 = ~n5587 ;
  assign y1899 = ~1'b0 ;
  assign y1900 = n5588 ;
  assign y1901 = ~1'b0 ;
  assign y1902 = n5589 ;
  assign y1903 = ~n5591 ;
  assign y1904 = n5597 ;
  assign y1905 = ~n5598 ;
  assign y1906 = n5599 ;
  assign y1907 = n5611 ;
  assign y1908 = ~n5612 ;
  assign y1909 = ~n5615 ;
  assign y1910 = ~1'b0 ;
  assign y1911 = ~n5619 ;
  assign y1912 = n5620 ;
  assign y1913 = ~n5621 ;
  assign y1914 = n5627 ;
  assign y1915 = ~n5631 ;
  assign y1916 = ~n5632 ;
  assign y1917 = ~n2019 ;
  assign y1918 = n5637 ;
  assign y1919 = ~n5641 ;
  assign y1920 = n5642 ;
  assign y1921 = ~n5649 ;
  assign y1922 = n5650 ;
  assign y1923 = ~1'b0 ;
  assign y1924 = ~1'b0 ;
  assign y1925 = ~n5652 ;
  assign y1926 = ~n5654 ;
  assign y1927 = ~1'b0 ;
  assign y1928 = n5655 ;
  assign y1929 = n5659 ;
  assign y1930 = n5660 ;
  assign y1931 = n5661 ;
  assign y1932 = ~n5662 ;
  assign y1933 = n5663 ;
  assign y1934 = ~n5666 ;
  assign y1935 = n5677 ;
  assign y1936 = ~n5683 ;
  assign y1937 = ~n1928 ;
  assign y1938 = ~1'b0 ;
  assign y1939 = ~n5684 ;
  assign y1940 = n5685 ;
  assign y1941 = ~n5689 ;
  assign y1942 = ~n5690 ;
  assign y1943 = ~n5691 ;
  assign y1944 = ~n5692 ;
  assign y1945 = ~n5694 ;
  assign y1946 = n5700 ;
  assign y1947 = n5702 ;
  assign y1948 = ~1'b0 ;
  assign y1949 = n5706 ;
  assign y1950 = ~n5714 ;
  assign y1951 = n5716 ;
  assign y1952 = n5721 ;
  assign y1953 = ~1'b0 ;
  assign y1954 = n5726 ;
  assign y1955 = ~n5728 ;
  assign y1956 = n5735 ;
  assign y1957 = n5737 ;
  assign y1958 = ~n5738 ;
  assign y1959 = ~n5741 ;
  assign y1960 = ~1'b0 ;
  assign y1961 = n5742 ;
  assign y1962 = n5745 ;
  assign y1963 = n5746 ;
  assign y1964 = n5747 ;
  assign y1965 = ~n5750 ;
  assign y1966 = ~1'b0 ;
  assign y1967 = ~n5753 ;
  assign y1968 = n5756 ;
  assign y1969 = n5758 ;
  assign y1970 = ~1'b0 ;
  assign y1971 = ~n5765 ;
  assign y1972 = ~1'b0 ;
  assign y1973 = ~n5769 ;
  assign y1974 = n5772 ;
  assign y1975 = ~n5775 ;
  assign y1976 = ~1'b0 ;
  assign y1977 = ~n5776 ;
  assign y1978 = ~1'b0 ;
  assign y1979 = ~n5777 ;
  assign y1980 = n5781 ;
  assign y1981 = ~1'b0 ;
  assign y1982 = n5785 ;
  assign y1983 = ~1'b0 ;
  assign y1984 = ~n5791 ;
  assign y1985 = ~n5794 ;
  assign y1986 = n5800 ;
  assign y1987 = n5801 ;
  assign y1988 = n5804 ;
  assign y1989 = n5808 ;
  assign y1990 = ~1'b0 ;
  assign y1991 = n5809 ;
  assign y1992 = ~n5810 ;
  assign y1993 = n5813 ;
  assign y1994 = ~n5815 ;
  assign y1995 = n5818 ;
  assign y1996 = ~n5819 ;
  assign y1997 = ~1'b0 ;
  assign y1998 = ~n5821 ;
  assign y1999 = ~n1770 ;
  assign y2000 = ~n5826 ;
  assign y2001 = ~n5827 ;
  assign y2002 = n5829 ;
  assign y2003 = ~1'b0 ;
  assign y2004 = n5834 ;
  assign y2005 = n5836 ;
  assign y2006 = n5837 ;
  assign y2007 = ~1'b0 ;
  assign y2008 = n5838 ;
  assign y2009 = n5839 ;
  assign y2010 = ~n5844 ;
  assign y2011 = n5858 ;
  assign y2012 = ~1'b0 ;
  assign y2013 = ~n5859 ;
  assign y2014 = ~1'b0 ;
  assign y2015 = ~n5861 ;
  assign y2016 = 1'b0 ;
  assign y2017 = ~1'b0 ;
  assign y2018 = n5867 ;
  assign y2019 = n5871 ;
  assign y2020 = ~n5872 ;
  assign y2021 = ~1'b0 ;
  assign y2022 = n5878 ;
  assign y2023 = n5880 ;
  assign y2024 = n5881 ;
  assign y2025 = ~n5882 ;
  assign y2026 = ~n5884 ;
  assign y2027 = ~n5885 ;
  assign y2028 = ~1'b0 ;
  assign y2029 = n5689 ;
  assign y2030 = ~n5888 ;
  assign y2031 = ~n5890 ;
  assign y2032 = ~1'b0 ;
  assign y2033 = ~1'b0 ;
  assign y2034 = ~1'b0 ;
  assign y2035 = ~n5893 ;
  assign y2036 = n5895 ;
  assign y2037 = ~1'b0 ;
  assign y2038 = n5897 ;
  assign y2039 = ~n5909 ;
  assign y2040 = ~n5912 ;
  assign y2041 = ~n5914 ;
  assign y2042 = ~n5916 ;
  assign y2043 = n5918 ;
  assign y2044 = n5920 ;
  assign y2045 = n3329 ;
  assign y2046 = ~1'b0 ;
  assign y2047 = ~1'b0 ;
  assign y2048 = n5926 ;
  assign y2049 = n4927 ;
  assign y2050 = n5928 ;
  assign y2051 = ~1'b0 ;
  assign y2052 = n5930 ;
  assign y2053 = ~1'b0 ;
  assign y2054 = ~n5931 ;
  assign y2055 = ~n5937 ;
  assign y2056 = ~n5944 ;
  assign y2057 = ~1'b0 ;
  assign y2058 = ~1'b0 ;
  assign y2059 = ~1'b0 ;
  assign y2060 = ~n5947 ;
  assign y2061 = n5948 ;
  assign y2062 = n5954 ;
  assign y2063 = n746 ;
  assign y2064 = ~n5958 ;
  assign y2065 = n5959 ;
  assign y2066 = n5961 ;
  assign y2067 = ~n5965 ;
  assign y2068 = n5966 ;
  assign y2069 = ~1'b0 ;
  assign y2070 = ~n5974 ;
  assign y2071 = ~n5984 ;
  assign y2072 = ~n5986 ;
  assign y2073 = n5988 ;
  assign y2074 = n5992 ;
  assign y2075 = ~n5995 ;
  assign y2076 = 1'b0 ;
  assign y2077 = n6001 ;
  assign y2078 = ~1'b0 ;
  assign y2079 = n6014 ;
  assign y2080 = n6015 ;
  assign y2081 = ~n6019 ;
  assign y2082 = ~n6021 ;
  assign y2083 = n6023 ;
  assign y2084 = ~n6024 ;
  assign y2085 = ~1'b0 ;
  assign y2086 = ~n6026 ;
  assign y2087 = ~n6030 ;
  assign y2088 = ~1'b0 ;
  assign y2089 = ~n6035 ;
  assign y2090 = ~n6038 ;
  assign y2091 = n6039 ;
  assign y2092 = n6040 ;
  assign y2093 = ~n6042 ;
  assign y2094 = ~n6044 ;
  assign y2095 = ~n726 ;
  assign y2096 = n5851 ;
  assign y2097 = ~n6047 ;
  assign y2098 = ~1'b0 ;
  assign y2099 = ~n6049 ;
  assign y2100 = ~n6050 ;
  assign y2101 = ~n6051 ;
  assign y2102 = ~n6052 ;
  assign y2103 = ~n6056 ;
  assign y2104 = ~n6061 ;
  assign y2105 = ~n6063 ;
  assign y2106 = ~n6066 ;
  assign y2107 = n6068 ;
  assign y2108 = n6083 ;
  assign y2109 = n6085 ;
  assign y2110 = n6090 ;
  assign y2111 = 1'b0 ;
  assign y2112 = ~n6096 ;
  assign y2113 = n6105 ;
  assign y2114 = ~1'b0 ;
  assign y2115 = ~1'b0 ;
  assign y2116 = n6110 ;
  assign y2117 = ~1'b0 ;
  assign y2118 = ~n6111 ;
  assign y2119 = ~n5589 ;
  assign y2120 = ~n6124 ;
  assign y2121 = ~n6130 ;
  assign y2122 = ~1'b0 ;
  assign y2123 = ~1'b0 ;
  assign y2124 = ~n6132 ;
  assign y2125 = n6133 ;
  assign y2126 = n4341 ;
  assign y2127 = n6134 ;
  assign y2128 = ~1'b0 ;
  assign y2129 = ~n6145 ;
  assign y2130 = n6147 ;
  assign y2131 = n6150 ;
  assign y2132 = ~1'b0 ;
  assign y2133 = ~n6152 ;
  assign y2134 = ~n6154 ;
  assign y2135 = ~1'b0 ;
  assign y2136 = ~n6160 ;
  assign y2137 = n6161 ;
  assign y2138 = n6165 ;
  assign y2139 = ~1'b0 ;
  assign y2140 = ~1'b0 ;
  assign y2141 = n6167 ;
  assign y2142 = ~n6170 ;
  assign y2143 = ~n6172 ;
  assign y2144 = ~1'b0 ;
  assign y2145 = n6173 ;
  assign y2146 = ~n6180 ;
  assign y2147 = ~n6182 ;
  assign y2148 = ~n6183 ;
  assign y2149 = n6186 ;
  assign y2150 = ~n6189 ;
  assign y2151 = ~n6191 ;
  assign y2152 = ~n6197 ;
  assign y2153 = ~1'b0 ;
  assign y2154 = ~1'b0 ;
  assign y2155 = n6200 ;
  assign y2156 = n6203 ;
  assign y2157 = n6207 ;
  assign y2158 = ~n6222 ;
  assign y2159 = ~n6230 ;
  assign y2160 = n6235 ;
  assign y2161 = n6236 ;
  assign y2162 = n6245 ;
  assign y2163 = n6250 ;
  assign y2164 = n6255 ;
  assign y2165 = n6262 ;
  assign y2166 = n6264 ;
  assign y2167 = ~1'b0 ;
  assign y2168 = ~1'b0 ;
  assign y2169 = ~n6267 ;
  assign y2170 = ~n6275 ;
  assign y2171 = n6276 ;
  assign y2172 = ~n1023 ;
  assign y2173 = n6282 ;
  assign y2174 = ~1'b0 ;
  assign y2175 = ~1'b0 ;
  assign y2176 = ~1'b0 ;
  assign y2177 = ~n6284 ;
  assign y2178 = ~1'b0 ;
  assign y2179 = ~n6298 ;
  assign y2180 = n6305 ;
  assign y2181 = ~1'b0 ;
  assign y2182 = n6306 ;
  assign y2183 = n6309 ;
  assign y2184 = n6310 ;
  assign y2185 = ~n6313 ;
  assign y2186 = ~1'b0 ;
  assign y2187 = n6318 ;
  assign y2188 = ~n6320 ;
  assign y2189 = ~1'b0 ;
  assign y2190 = ~n6322 ;
  assign y2191 = ~n6326 ;
  assign y2192 = ~n6336 ;
  assign y2193 = n6337 ;
  assign y2194 = n1125 ;
  assign y2195 = ~n6341 ;
  assign y2196 = n6342 ;
  assign y2197 = n6348 ;
  assign y2198 = n6351 ;
  assign y2199 = ~1'b0 ;
  assign y2200 = ~n6355 ;
  assign y2201 = n6357 ;
  assign y2202 = n6360 ;
  assign y2203 = ~n6366 ;
  assign y2204 = ~n6372 ;
  assign y2205 = ~n6373 ;
  assign y2206 = n6374 ;
  assign y2207 = n6378 ;
  assign y2208 = n6383 ;
  assign y2209 = ~n6387 ;
  assign y2210 = 1'b0 ;
  assign y2211 = ~n6392 ;
  assign y2212 = ~n6393 ;
  assign y2213 = ~n6395 ;
  assign y2214 = n6398 ;
  assign y2215 = ~n6400 ;
  assign y2216 = ~n6401 ;
  assign y2217 = n6404 ;
  assign y2218 = n6410 ;
  assign y2219 = n6423 ;
  assign y2220 = ~1'b0 ;
  assign y2221 = n6427 ;
  assign y2222 = ~n6428 ;
  assign y2223 = ~n6430 ;
  assign y2224 = n6435 ;
  assign y2225 = ~1'b0 ;
  assign y2226 = n6436 ;
  assign y2227 = n6437 ;
  assign y2228 = ~n1633 ;
  assign y2229 = n6445 ;
  assign y2230 = n6446 ;
  assign y2231 = ~n6449 ;
  assign y2232 = ~1'b0 ;
  assign y2233 = n6451 ;
  assign y2234 = n6452 ;
  assign y2235 = ~n6456 ;
  assign y2236 = ~n6459 ;
  assign y2237 = n6460 ;
  assign y2238 = ~n6461 ;
  assign y2239 = n6467 ;
  assign y2240 = ~n6479 ;
  assign y2241 = ~n6480 ;
  assign y2242 = n436 ;
  assign y2243 = n6481 ;
  assign y2244 = ~n6485 ;
  assign y2245 = ~n6488 ;
  assign y2246 = n3610 ;
  assign y2247 = ~1'b0 ;
  assign y2248 = ~1'b0 ;
  assign y2249 = ~n6489 ;
  assign y2250 = ~1'b0 ;
  assign y2251 = n6491 ;
  assign y2252 = ~n6492 ;
  assign y2253 = ~1'b0 ;
  assign y2254 = ~n6493 ;
  assign y2255 = n6494 ;
  assign y2256 = n6503 ;
  assign y2257 = n6506 ;
  assign y2258 = ~n593 ;
  assign y2259 = ~n6513 ;
  assign y2260 = n6515 ;
  assign y2261 = ~1'b0 ;
  assign y2262 = n6517 ;
  assign y2263 = n6519 ;
  assign y2264 = ~1'b0 ;
  assign y2265 = ~n6520 ;
  assign y2266 = n6521 ;
  assign y2267 = ~1'b0 ;
  assign y2268 = n6527 ;
  assign y2269 = ~n6531 ;
  assign y2270 = ~n6535 ;
  assign y2271 = n6536 ;
  assign y2272 = ~n6538 ;
  assign y2273 = ~n6541 ;
  assign y2274 = ~n6543 ;
  assign y2275 = n6550 ;
  assign y2276 = n6552 ;
  assign y2277 = ~n5789 ;
  assign y2278 = ~1'b0 ;
  assign y2279 = ~n6553 ;
  assign y2280 = n6557 ;
  assign y2281 = ~n6564 ;
  assign y2282 = n6568 ;
  assign y2283 = ~1'b0 ;
  assign y2284 = ~n6571 ;
  assign y2285 = ~n6573 ;
  assign y2286 = ~1'b0 ;
  assign y2287 = ~n6576 ;
  assign y2288 = ~n6578 ;
  assign y2289 = n6589 ;
  assign y2290 = ~n6596 ;
  assign y2291 = n6609 ;
  assign y2292 = ~n6610 ;
  assign y2293 = ~1'b0 ;
  assign y2294 = n6611 ;
  assign y2295 = n6612 ;
  assign y2296 = ~n6623 ;
  assign y2297 = ~1'b0 ;
  assign y2298 = n6627 ;
  assign y2299 = n6632 ;
  assign y2300 = ~n6634 ;
  assign y2301 = ~n6635 ;
  assign y2302 = ~1'b0 ;
  assign y2303 = ~n6638 ;
  assign y2304 = n6641 ;
  assign y2305 = n6643 ;
  assign y2306 = ~1'b0 ;
  assign y2307 = n6645 ;
  assign y2308 = ~n6651 ;
  assign y2309 = ~n6654 ;
  assign y2310 = n6656 ;
  assign y2311 = n6660 ;
  assign y2312 = ~n6664 ;
  assign y2313 = ~n6667 ;
  assign y2314 = ~1'b0 ;
  assign y2315 = ~n6670 ;
  assign y2316 = ~n6672 ;
  assign y2317 = n6680 ;
  assign y2318 = n2038 ;
  assign y2319 = n6681 ;
  assign y2320 = ~n6685 ;
  assign y2321 = n6686 ;
  assign y2322 = n6690 ;
  assign y2323 = n6691 ;
  assign y2324 = ~n6693 ;
  assign y2325 = n6697 ;
  assign y2326 = ~n6698 ;
  assign y2327 = ~n6699 ;
  assign y2328 = ~n6701 ;
  assign y2329 = n6703 ;
  assign y2330 = ~1'b0 ;
  assign y2331 = n6709 ;
  assign y2332 = ~n6711 ;
  assign y2333 = ~n6712 ;
  assign y2334 = ~1'b0 ;
  assign y2335 = 1'b0 ;
  assign y2336 = ~n6715 ;
  assign y2337 = n6716 ;
  assign y2338 = ~1'b0 ;
  assign y2339 = ~n6723 ;
  assign y2340 = n6725 ;
  assign y2341 = n6726 ;
  assign y2342 = ~1'b0 ;
  assign y2343 = ~n6732 ;
  assign y2344 = ~n6733 ;
  assign y2345 = ~n6741 ;
  assign y2346 = n6749 ;
  assign y2347 = n6751 ;
  assign y2348 = n6752 ;
  assign y2349 = n6753 ;
  assign y2350 = ~n6754 ;
  assign y2351 = ~n6760 ;
  assign y2352 = ~1'b0 ;
  assign y2353 = ~n6764 ;
  assign y2354 = n6766 ;
  assign y2355 = ~n6768 ;
  assign y2356 = ~n6769 ;
  assign y2357 = n6776 ;
  assign y2358 = ~1'b0 ;
  assign y2359 = ~1'b0 ;
  assign y2360 = n6782 ;
  assign y2361 = n6784 ;
  assign y2362 = n6787 ;
  assign y2363 = ~n6789 ;
  assign y2364 = ~1'b0 ;
  assign y2365 = n6791 ;
  assign y2366 = n6792 ;
  assign y2367 = n6793 ;
  assign y2368 = ~1'b0 ;
  assign y2369 = ~n6799 ;
  assign y2370 = ~n6800 ;
  assign y2371 = n6801 ;
  assign y2372 = ~n6806 ;
  assign y2373 = n6811 ;
  assign y2374 = n6812 ;
  assign y2375 = ~n6813 ;
  assign y2376 = ~1'b0 ;
  assign y2377 = ~n6814 ;
  assign y2378 = ~n6816 ;
  assign y2379 = ~1'b0 ;
  assign y2380 = n6820 ;
  assign y2381 = ~1'b0 ;
  assign y2382 = ~n6829 ;
  assign y2383 = ~n6830 ;
  assign y2384 = n6840 ;
  assign y2385 = ~n6843 ;
  assign y2386 = n6845 ;
  assign y2387 = ~n6846 ;
  assign y2388 = ~n6848 ;
  assign y2389 = n6851 ;
  assign y2390 = ~1'b0 ;
  assign y2391 = n6859 ;
  assign y2392 = n6865 ;
  assign y2393 = ~n6868 ;
  assign y2394 = ~1'b0 ;
  assign y2395 = ~1'b0 ;
  assign y2396 = ~n6870 ;
  assign y2397 = ~1'b0 ;
  assign y2398 = ~n6876 ;
  assign y2399 = n6881 ;
  assign y2400 = ~1'b0 ;
  assign y2401 = n6882 ;
  assign y2402 = n6888 ;
  assign y2403 = ~1'b0 ;
  assign y2404 = n6891 ;
  assign y2405 = ~n6893 ;
  assign y2406 = n6894 ;
  assign y2407 = ~n6897 ;
  assign y2408 = ~1'b0 ;
  assign y2409 = n6906 ;
  assign y2410 = ~n6909 ;
  assign y2411 = n6913 ;
  assign y2412 = n6916 ;
  assign y2413 = ~n6917 ;
  assign y2414 = n6918 ;
  assign y2415 = ~n6920 ;
  assign y2416 = ~1'b0 ;
  assign y2417 = n6921 ;
  assign y2418 = ~1'b0 ;
  assign y2419 = ~n6925 ;
  assign y2420 = ~n6934 ;
  assign y2421 = ~n6935 ;
  assign y2422 = n4158 ;
  assign y2423 = n6938 ;
  assign y2424 = ~n6939 ;
  assign y2425 = ~n6945 ;
  assign y2426 = ~n6949 ;
  assign y2427 = ~1'b0 ;
  assign y2428 = n6952 ;
  assign y2429 = ~n6958 ;
  assign y2430 = ~n6960 ;
  assign y2431 = n6967 ;
  assign y2432 = ~n6968 ;
  assign y2433 = n6972 ;
  assign y2434 = ~n6973 ;
  assign y2435 = ~n6976 ;
  assign y2436 = ~n6982 ;
  assign y2437 = n6984 ;
  assign y2438 = ~1'b0 ;
  assign y2439 = n6988 ;
  assign y2440 = ~1'b0 ;
  assign y2441 = ~n6993 ;
  assign y2442 = ~n6999 ;
  assign y2443 = ~n7002 ;
  assign y2444 = ~1'b0 ;
  assign y2445 = ~1'b0 ;
  assign y2446 = n7009 ;
  assign y2447 = n7013 ;
  assign y2448 = ~n7017 ;
  assign y2449 = ~n7018 ;
  assign y2450 = ~1'b0 ;
  assign y2451 = n7019 ;
  assign y2452 = ~n7025 ;
  assign y2453 = n7029 ;
  assign y2454 = ~n7031 ;
  assign y2455 = ~n7033 ;
  assign y2456 = ~n7040 ;
  assign y2457 = n7043 ;
  assign y2458 = ~1'b0 ;
  assign y2459 = ~1'b0 ;
  assign y2460 = ~n7045 ;
  assign y2461 = ~1'b0 ;
  assign y2462 = ~n7047 ;
  assign y2463 = n7052 ;
  assign y2464 = n7055 ;
  assign y2465 = 1'b0 ;
  assign y2466 = ~1'b0 ;
  assign y2467 = ~n7058 ;
  assign y2468 = n7062 ;
  assign y2469 = ~n7066 ;
  assign y2470 = n7067 ;
  assign y2471 = n7084 ;
  assign y2472 = n7085 ;
  assign y2473 = ~n7088 ;
  assign y2474 = ~n7093 ;
  assign y2475 = n7099 ;
  assign y2476 = ~1'b0 ;
  assign y2477 = ~n7101 ;
  assign y2478 = ~1'b0 ;
  assign y2479 = ~1'b0 ;
  assign y2480 = n7105 ;
  assign y2481 = ~1'b0 ;
  assign y2482 = ~1'b0 ;
  assign y2483 = 1'b0 ;
  assign y2484 = n7114 ;
  assign y2485 = n7123 ;
  assign y2486 = ~n7128 ;
  assign y2487 = ~n5352 ;
  assign y2488 = ~n7131 ;
  assign y2489 = n250 ;
  assign y2490 = ~n7139 ;
  assign y2491 = n7143 ;
  assign y2492 = n7146 ;
  assign y2493 = n7148 ;
  assign y2494 = n7150 ;
  assign y2495 = n2246 ;
  assign y2496 = ~n7156 ;
  assign y2497 = ~1'b0 ;
  assign y2498 = ~n1748 ;
  assign y2499 = ~1'b0 ;
  assign y2500 = n7158 ;
  assign y2501 = ~n3946 ;
  assign y2502 = ~n2641 ;
  assign y2503 = ~n7168 ;
  assign y2504 = n7171 ;
  assign y2505 = ~1'b0 ;
  assign y2506 = ~n7173 ;
  assign y2507 = n7174 ;
  assign y2508 = n7175 ;
  assign y2509 = n7177 ;
  assign y2510 = ~1'b0 ;
  assign y2511 = ~1'b0 ;
  assign y2512 = ~1'b0 ;
  assign y2513 = n7180 ;
  assign y2514 = n7183 ;
  assign y2515 = n7184 ;
  assign y2516 = n7186 ;
  assign y2517 = ~n7191 ;
  assign y2518 = ~1'b0 ;
  assign y2519 = n7192 ;
  assign y2520 = ~n7193 ;
  assign y2521 = ~n7199 ;
  assign y2522 = ~n7204 ;
  assign y2523 = ~1'b0 ;
  assign y2524 = ~n7206 ;
  assign y2525 = ~n7210 ;
  assign y2526 = ~1'b0 ;
  assign y2527 = n7211 ;
  assign y2528 = n7212 ;
  assign y2529 = ~1'b0 ;
  assign y2530 = 1'b0 ;
  assign y2531 = n7213 ;
  assign y2532 = n7214 ;
  assign y2533 = ~1'b0 ;
  assign y2534 = n7217 ;
  assign y2535 = ~1'b0 ;
  assign y2536 = ~n7224 ;
  assign y2537 = ~1'b0 ;
  assign y2538 = n7225 ;
  assign y2539 = ~1'b0 ;
  assign y2540 = n7231 ;
  assign y2541 = n7235 ;
  assign y2542 = ~n7247 ;
  assign y2543 = ~n7249 ;
  assign y2544 = n7251 ;
  assign y2545 = ~1'b0 ;
  assign y2546 = ~1'b0 ;
  assign y2547 = ~n7260 ;
  assign y2548 = ~n7261 ;
  assign y2549 = ~1'b0 ;
  assign y2550 = ~n7263 ;
  assign y2551 = ~n7272 ;
  assign y2552 = n7274 ;
  assign y2553 = ~n7283 ;
  assign y2554 = ~n7301 ;
  assign y2555 = ~1'b0 ;
  assign y2556 = n7303 ;
  assign y2557 = ~1'b0 ;
  assign y2558 = ~n7307 ;
  assign y2559 = ~n7310 ;
  assign y2560 = n7311 ;
  assign y2561 = ~n7313 ;
  assign y2562 = ~n7314 ;
  assign y2563 = n7321 ;
  assign y2564 = ~1'b0 ;
  assign y2565 = n7323 ;
  assign y2566 = ~n7328 ;
  assign y2567 = 1'b0 ;
  assign y2568 = n7329 ;
  assign y2569 = n7334 ;
  assign y2570 = n7338 ;
  assign y2571 = ~1'b0 ;
  assign y2572 = ~n7340 ;
  assign y2573 = n1715 ;
  assign y2574 = n7341 ;
  assign y2575 = ~1'b0 ;
  assign y2576 = ~n7342 ;
  assign y2577 = ~n7343 ;
  assign y2578 = n7344 ;
  assign y2579 = ~n7346 ;
  assign y2580 = ~1'b0 ;
  assign y2581 = n7349 ;
  assign y2582 = ~n7350 ;
  assign y2583 = n181 ;
  assign y2584 = ~n7351 ;
  assign y2585 = n7359 ;
  assign y2586 = ~n7360 ;
  assign y2587 = ~n7366 ;
  assign y2588 = n7368 ;
  assign y2589 = n7372 ;
  assign y2590 = n7376 ;
  assign y2591 = ~n7379 ;
  assign y2592 = n7387 ;
  assign y2593 = ~n7389 ;
  assign y2594 = ~n7396 ;
  assign y2595 = n7397 ;
  assign y2596 = ~n7402 ;
  assign y2597 = n7404 ;
  assign y2598 = n7406 ;
  assign y2599 = ~n7408 ;
  assign y2600 = ~n7409 ;
  assign y2601 = ~n7410 ;
  assign y2602 = ~1'b0 ;
  assign y2603 = ~1'b0 ;
  assign y2604 = ~n7412 ;
  assign y2605 = ~n7424 ;
  assign y2606 = n7425 ;
  assign y2607 = ~1'b0 ;
  assign y2608 = ~n7434 ;
  assign y2609 = ~n7451 ;
  assign y2610 = ~1'b0 ;
  assign y2611 = ~n7453 ;
  assign y2612 = n7457 ;
  assign y2613 = ~n7460 ;
  assign y2614 = n7463 ;
  assign y2615 = n7464 ;
  assign y2616 = ~n7471 ;
  assign y2617 = ~n7473 ;
  assign y2618 = ~1'b0 ;
  assign y2619 = n7484 ;
  assign y2620 = n7485 ;
  assign y2621 = n7489 ;
  assign y2622 = ~n7493 ;
  assign y2623 = ~n7494 ;
  assign y2624 = ~n7499 ;
  assign y2625 = ~1'b0 ;
  assign y2626 = n7513 ;
  assign y2627 = ~n7517 ;
  assign y2628 = ~n7524 ;
  assign y2629 = n7528 ;
  assign y2630 = n7532 ;
  assign y2631 = n7538 ;
  assign y2632 = ~n7541 ;
  assign y2633 = ~1'b0 ;
  assign y2634 = ~n7553 ;
  assign y2635 = ~n7558 ;
  assign y2636 = ~n7562 ;
  assign y2637 = ~1'b0 ;
  assign y2638 = n7566 ;
  assign y2639 = ~1'b0 ;
  assign y2640 = n7567 ;
  assign y2641 = ~n7572 ;
  assign y2642 = ~1'b0 ;
  assign y2643 = n7573 ;
  assign y2644 = ~n7574 ;
  assign y2645 = n7575 ;
  assign y2646 = ~1'b0 ;
  assign y2647 = ~1'b0 ;
  assign y2648 = n7578 ;
  assign y2649 = ~n7580 ;
  assign y2650 = n7589 ;
  assign y2651 = ~n7595 ;
  assign y2652 = n7596 ;
  assign y2653 = n7602 ;
  assign y2654 = ~n7604 ;
  assign y2655 = ~n7607 ;
  assign y2656 = n7616 ;
  assign y2657 = ~n7620 ;
  assign y2658 = n7622 ;
  assign y2659 = ~n7629 ;
  assign y2660 = n7632 ;
  assign y2661 = n7636 ;
  assign y2662 = ~1'b0 ;
  assign y2663 = n7641 ;
  assign y2664 = ~n7642 ;
  assign y2665 = n7644 ;
  assign y2666 = ~n7646 ;
  assign y2667 = ~1'b0 ;
  assign y2668 = n7648 ;
  assign y2669 = n7652 ;
  assign y2670 = ~n7654 ;
  assign y2671 = ~n7655 ;
  assign y2672 = ~n7659 ;
  assign y2673 = ~n7663 ;
  assign y2674 = n7665 ;
  assign y2675 = ~n7668 ;
  assign y2676 = ~1'b0 ;
  assign y2677 = ~n7669 ;
  assign y2678 = ~n7671 ;
  assign y2679 = ~1'b0 ;
  assign y2680 = ~n7672 ;
  assign y2681 = n7674 ;
  assign y2682 = ~n7675 ;
  assign y2683 = n7679 ;
  assign y2684 = ~n7682 ;
  assign y2685 = 1'b0 ;
  assign y2686 = n7685 ;
  assign y2687 = ~1'b0 ;
  assign y2688 = ~1'b0 ;
  assign y2689 = ~n7686 ;
  assign y2690 = n7687 ;
  assign y2691 = n7694 ;
  assign y2692 = n7696 ;
  assign y2693 = n7697 ;
  assign y2694 = ~1'b0 ;
  assign y2695 = ~n7703 ;
  assign y2696 = n7274 ;
  assign y2697 = 1'b0 ;
  assign y2698 = ~1'b0 ;
  assign y2699 = ~1'b0 ;
  assign y2700 = n4193 ;
  assign y2701 = n7707 ;
  assign y2702 = ~n7708 ;
  assign y2703 = ~n7713 ;
  assign y2704 = n7719 ;
  assign y2705 = n7724 ;
  assign y2706 = n7727 ;
  assign y2707 = ~n7729 ;
  assign y2708 = ~1'b0 ;
  assign y2709 = n7730 ;
  assign y2710 = ~n3566 ;
  assign y2711 = ~n7734 ;
  assign y2712 = n7736 ;
  assign y2713 = n7740 ;
  assign y2714 = ~n7741 ;
  assign y2715 = ~1'b0 ;
  assign y2716 = ~n7742 ;
  assign y2717 = n7745 ;
  assign y2718 = ~n3241 ;
  assign y2719 = ~1'b0 ;
  assign y2720 = 1'b0 ;
  assign y2721 = ~n7748 ;
  assign y2722 = ~1'b0 ;
  assign y2723 = ~n7754 ;
  assign y2724 = n7762 ;
  assign y2725 = n7765 ;
  assign y2726 = ~n7767 ;
  assign y2727 = ~n7768 ;
  assign y2728 = n7774 ;
  assign y2729 = ~n7777 ;
  assign y2730 = ~n7778 ;
  assign y2731 = ~n7791 ;
  assign y2732 = ~1'b0 ;
  assign y2733 = n7795 ;
  assign y2734 = ~n7798 ;
  assign y2735 = n7800 ;
  assign y2736 = ~1'b0 ;
  assign y2737 = ~n7804 ;
  assign y2738 = n7805 ;
  assign y2739 = ~n7808 ;
  assign y2740 = n7811 ;
  assign y2741 = ~n7813 ;
  assign y2742 = n7815 ;
  assign y2743 = ~n7816 ;
  assign y2744 = n7818 ;
  assign y2745 = n7824 ;
  assign y2746 = ~n7831 ;
  assign y2747 = ~n7832 ;
  assign y2748 = n7833 ;
  assign y2749 = n7838 ;
  assign y2750 = ~n7841 ;
  assign y2751 = ~n7842 ;
  assign y2752 = n7846 ;
  assign y2753 = ~1'b0 ;
  assign y2754 = n7850 ;
  assign y2755 = ~n7856 ;
  assign y2756 = n7860 ;
  assign y2757 = n7861 ;
  assign y2758 = ~1'b0 ;
  assign y2759 = ~n7867 ;
  assign y2760 = ~n7869 ;
  assign y2761 = ~n7870 ;
  assign y2762 = ~n7873 ;
  assign y2763 = ~1'b0 ;
  assign y2764 = ~1'b0 ;
  assign y2765 = ~1'b0 ;
  assign y2766 = n7874 ;
  assign y2767 = ~n7884 ;
  assign y2768 = n7886 ;
  assign y2769 = ~n7887 ;
  assign y2770 = ~n7898 ;
  assign y2771 = ~1'b0 ;
  assign y2772 = n7908 ;
  assign y2773 = n7912 ;
  assign y2774 = ~n7914 ;
  assign y2775 = ~1'b0 ;
  assign y2776 = n7915 ;
  assign y2777 = n7917 ;
  assign y2778 = ~1'b0 ;
  assign y2779 = ~n7919 ;
  assign y2780 = ~1'b0 ;
  assign y2781 = n7927 ;
  assign y2782 = ~n7930 ;
  assign y2783 = ~n7931 ;
  assign y2784 = ~n7935 ;
  assign y2785 = ~n5387 ;
  assign y2786 = ~1'b0 ;
  assign y2787 = n7937 ;
  assign y2788 = ~n7943 ;
  assign y2789 = ~1'b0 ;
  assign y2790 = ~n7947 ;
  assign y2791 = n7950 ;
  assign y2792 = ~1'b0 ;
  assign y2793 = n7954 ;
  assign y2794 = n7955 ;
  assign y2795 = n7957 ;
  assign y2796 = n7963 ;
  assign y2797 = n7968 ;
  assign y2798 = ~n7970 ;
  assign y2799 = ~n7971 ;
  assign y2800 = n7975 ;
  assign y2801 = n1433 ;
  assign y2802 = ~1'b0 ;
  assign y2803 = ~n7979 ;
  assign y2804 = ~n7981 ;
  assign y2805 = ~1'b0 ;
  assign y2806 = n7984 ;
  assign y2807 = ~n7986 ;
  assign y2808 = n7987 ;
  assign y2809 = ~n7990 ;
  assign y2810 = ~n7999 ;
  assign y2811 = ~n8001 ;
  assign y2812 = n8005 ;
  assign y2813 = ~n8006 ;
  assign y2814 = ~1'b0 ;
  assign y2815 = n8010 ;
  assign y2816 = ~n8012 ;
  assign y2817 = ~n8014 ;
  assign y2818 = ~n8019 ;
  assign y2819 = ~n1349 ;
  assign y2820 = ~n8020 ;
  assign y2821 = n8023 ;
  assign y2822 = n8024 ;
  assign y2823 = ~n8030 ;
  assign y2824 = ~1'b0 ;
  assign y2825 = n8032 ;
  assign y2826 = n8039 ;
  assign y2827 = n4483 ;
  assign y2828 = ~n3168 ;
  assign y2829 = ~n8041 ;
  assign y2830 = ~1'b0 ;
  assign y2831 = ~1'b0 ;
  assign y2832 = n7221 ;
  assign y2833 = ~n8043 ;
  assign y2834 = n8045 ;
  assign y2835 = ~n8049 ;
  assign y2836 = ~n8050 ;
  assign y2837 = ~1'b0 ;
  assign y2838 = n8054 ;
  assign y2839 = n8058 ;
  assign y2840 = n8061 ;
  assign y2841 = ~1'b0 ;
  assign y2842 = ~1'b0 ;
  assign y2843 = ~n8062 ;
  assign y2844 = ~n8066 ;
  assign y2845 = ~n8073 ;
  assign y2846 = ~1'b0 ;
  assign y2847 = ~1'b0 ;
  assign y2848 = ~n8076 ;
  assign y2849 = n8079 ;
  assign y2850 = n8081 ;
  assign y2851 = ~n8088 ;
  assign y2852 = ~n8092 ;
  assign y2853 = ~1'b0 ;
  assign y2854 = n8096 ;
  assign y2855 = ~n8106 ;
  assign y2856 = ~1'b0 ;
  assign y2857 = n8110 ;
  assign y2858 = ~n8111 ;
  assign y2859 = ~n8113 ;
  assign y2860 = ~1'b0 ;
  assign y2861 = ~1'b0 ;
  assign y2862 = n8120 ;
  assign y2863 = ~n8122 ;
  assign y2864 = n4815 ;
  assign y2865 = ~1'b0 ;
  assign y2866 = ~1'b0 ;
  assign y2867 = n8137 ;
  assign y2868 = ~n8138 ;
  assign y2869 = ~n8142 ;
  assign y2870 = ~1'b0 ;
  assign y2871 = ~n8143 ;
  assign y2872 = ~n8146 ;
  assign y2873 = n8147 ;
  assign y2874 = ~1'b0 ;
  assign y2875 = ~n8149 ;
  assign y2876 = ~n8150 ;
  assign y2877 = n8154 ;
  assign y2878 = n8157 ;
  assign y2879 = n8167 ;
  assign y2880 = ~n8173 ;
  assign y2881 = ~n8066 ;
  assign y2882 = n8176 ;
  assign y2883 = ~n8178 ;
  assign y2884 = ~1'b0 ;
  assign y2885 = ~1'b0 ;
  assign y2886 = ~n7774 ;
  assign y2887 = ~1'b0 ;
  assign y2888 = ~1'b0 ;
  assign y2889 = ~1'b0 ;
  assign y2890 = n8182 ;
  assign y2891 = n8183 ;
  assign y2892 = n8184 ;
  assign y2893 = n8187 ;
  assign y2894 = ~n8188 ;
  assign y2895 = ~n8190 ;
  assign y2896 = n8197 ;
  assign y2897 = n8202 ;
  assign y2898 = ~n8207 ;
  assign y2899 = 1'b0 ;
  assign y2900 = ~1'b0 ;
  assign y2901 = ~n8214 ;
  assign y2902 = n8219 ;
  assign y2903 = n8221 ;
  assign y2904 = ~n8222 ;
  assign y2905 = ~n8225 ;
  assign y2906 = ~1'b0 ;
  assign y2907 = ~n8227 ;
  assign y2908 = ~n8233 ;
  assign y2909 = n8234 ;
  assign y2910 = ~n8239 ;
  assign y2911 = ~1'b0 ;
  assign y2912 = ~n8243 ;
  assign y2913 = n8245 ;
  assign y2914 = n8246 ;
  assign y2915 = n8248 ;
  assign y2916 = 1'b0 ;
  assign y2917 = n8250 ;
  assign y2918 = ~n8252 ;
  assign y2919 = n8260 ;
  assign y2920 = ~1'b0 ;
  assign y2921 = n8261 ;
  assign y2922 = ~n8262 ;
  assign y2923 = ~1'b0 ;
  assign y2924 = ~n8265 ;
  assign y2925 = ~n8268 ;
  assign y2926 = n8271 ;
  assign y2927 = n8276 ;
  assign y2928 = n6908 ;
  assign y2929 = ~1'b0 ;
  assign y2930 = n8281 ;
  assign y2931 = n8282 ;
  assign y2932 = ~1'b0 ;
  assign y2933 = ~1'b0 ;
  assign y2934 = ~n8286 ;
  assign y2935 = n8287 ;
  assign y2936 = ~n8288 ;
  assign y2937 = ~n8292 ;
  assign y2938 = 1'b0 ;
  assign y2939 = n8295 ;
  assign y2940 = ~n8296 ;
  assign y2941 = ~n8300 ;
  assign y2942 = ~n8304 ;
  assign y2943 = ~n8305 ;
  assign y2944 = ~1'b0 ;
  assign y2945 = n8306 ;
  assign y2946 = n8307 ;
  assign y2947 = ~n8308 ;
  assign y2948 = ~n8312 ;
  assign y2949 = ~1'b0 ;
  assign y2950 = ~n8314 ;
  assign y2951 = ~1'b0 ;
  assign y2952 = n8316 ;
  assign y2953 = ~n8323 ;
  assign y2954 = n8331 ;
  assign y2955 = n8338 ;
  assign y2956 = n8340 ;
  assign y2957 = ~1'b0 ;
  assign y2958 = ~1'b0 ;
  assign y2959 = ~n8341 ;
  assign y2960 = ~1'b0 ;
  assign y2961 = n8355 ;
  assign y2962 = n8358 ;
  assign y2963 = n8359 ;
  assign y2964 = ~n8365 ;
  assign y2965 = n8368 ;
  assign y2966 = ~n8375 ;
  assign y2967 = ~n8385 ;
  assign y2968 = n8387 ;
  assign y2969 = ~1'b0 ;
  assign y2970 = n8390 ;
  assign y2971 = ~n8394 ;
  assign y2972 = n8396 ;
  assign y2973 = ~1'b0 ;
  assign y2974 = ~1'b0 ;
  assign y2975 = ~1'b0 ;
  assign y2976 = n8400 ;
  assign y2977 = ~1'b0 ;
  assign y2978 = n8402 ;
  assign y2979 = n8404 ;
  assign y2980 = n8408 ;
  assign y2981 = ~n8409 ;
  assign y2982 = ~1'b0 ;
  assign y2983 = ~n8412 ;
  assign y2984 = ~n8414 ;
  assign y2985 = ~n8415 ;
  assign y2986 = n8424 ;
  assign y2987 = n8425 ;
  assign y2988 = n8426 ;
  assign y2989 = ~1'b0 ;
  assign y2990 = n8427 ;
  assign y2991 = ~n8430 ;
  assign y2992 = ~n8431 ;
  assign y2993 = n8432 ;
  assign y2994 = ~n8436 ;
  assign y2995 = n8439 ;
  assign y2996 = n3482 ;
  assign y2997 = n8442 ;
  assign y2998 = ~1'b0 ;
  assign y2999 = ~1'b0 ;
  assign y3000 = ~1'b0 ;
  assign y3001 = ~n8443 ;
  assign y3002 = ~n8448 ;
  assign y3003 = ~1'b0 ;
  assign y3004 = ~n8452 ;
  assign y3005 = ~n8453 ;
  assign y3006 = ~n8455 ;
  assign y3007 = ~n8457 ;
  assign y3008 = ~1'b0 ;
  assign y3009 = ~n8463 ;
  assign y3010 = ~n8469 ;
  assign y3011 = ~1'b0 ;
  assign y3012 = n8473 ;
  assign y3013 = ~n8476 ;
  assign y3014 = n8477 ;
  assign y3015 = ~1'b0 ;
  assign y3016 = ~n8479 ;
  assign y3017 = n8484 ;
  assign y3018 = n8485 ;
  assign y3019 = n8488 ;
  assign y3020 = ~n8494 ;
  assign y3021 = n5784 ;
  assign y3022 = ~n8497 ;
  assign y3023 = n8501 ;
  assign y3024 = n8515 ;
  assign y3025 = n8520 ;
  assign y3026 = n8184 ;
  assign y3027 = n8521 ;
  assign y3028 = ~n8525 ;
  assign y3029 = ~1'b0 ;
  assign y3030 = ~n8526 ;
  assign y3031 = ~n8527 ;
  assign y3032 = ~n8531 ;
  assign y3033 = n8541 ;
  assign y3034 = n8547 ;
  assign y3035 = ~n8551 ;
  assign y3036 = ~1'b0 ;
  assign y3037 = ~1'b0 ;
  assign y3038 = n8555 ;
  assign y3039 = ~n8556 ;
  assign y3040 = n8560 ;
  assign y3041 = ~n8568 ;
  assign y3042 = ~1'b0 ;
  assign y3043 = ~1'b0 ;
  assign y3044 = ~1'b0 ;
  assign y3045 = ~1'b0 ;
  assign y3046 = ~1'b0 ;
  assign y3047 = ~n8571 ;
  assign y3048 = ~n8577 ;
  assign y3049 = n8586 ;
  assign y3050 = n8587 ;
  assign y3051 = ~n8589 ;
  assign y3052 = ~n8591 ;
  assign y3053 = n8593 ;
  assign y3054 = ~n8598 ;
  assign y3055 = ~1'b0 ;
  assign y3056 = n8601 ;
  assign y3057 = n8605 ;
  assign y3058 = ~1'b0 ;
  assign y3059 = ~n8608 ;
  assign y3060 = ~n8613 ;
  assign y3061 = n8614 ;
  assign y3062 = ~1'b0 ;
  assign y3063 = n8615 ;
  assign y3064 = ~n1205 ;
  assign y3065 = n8618 ;
  assign y3066 = ~1'b0 ;
  assign y3067 = ~1'b0 ;
  assign y3068 = ~n8619 ;
  assign y3069 = ~1'b0 ;
  assign y3070 = ~n8621 ;
  assign y3071 = ~1'b0 ;
  assign y3072 = ~n8625 ;
  assign y3073 = ~1'b0 ;
  assign y3074 = ~n8631 ;
  assign y3075 = ~n8633 ;
  assign y3076 = n8634 ;
  assign y3077 = n8635 ;
  assign y3078 = ~1'b0 ;
  assign y3079 = ~1'b0 ;
  assign y3080 = ~n8636 ;
  assign y3081 = ~n8641 ;
  assign y3082 = ~n8647 ;
  assign y3083 = ~n8652 ;
  assign y3084 = n8656 ;
  assign y3085 = ~n8657 ;
  assign y3086 = n8660 ;
  assign y3087 = ~n8663 ;
  assign y3088 = n8676 ;
  assign y3089 = ~1'b0 ;
  assign y3090 = ~n8679 ;
  assign y3091 = n8682 ;
  assign y3092 = n8684 ;
  assign y3093 = n8688 ;
  assign y3094 = ~n8689 ;
  assign y3095 = ~n8691 ;
  assign y3096 = ~1'b0 ;
  assign y3097 = ~n8697 ;
  assign y3098 = ~n8701 ;
  assign y3099 = n8704 ;
  assign y3100 = ~n8705 ;
  assign y3101 = ~n8719 ;
  assign y3102 = ~1'b0 ;
  assign y3103 = ~n8722 ;
  assign y3104 = n8729 ;
  assign y3105 = ~1'b0 ;
  assign y3106 = n627 ;
  assign y3107 = ~n8730 ;
  assign y3108 = n8732 ;
  assign y3109 = ~n8741 ;
  assign y3110 = ~1'b0 ;
  assign y3111 = n8742 ;
  assign y3112 = ~n3408 ;
  assign y3113 = ~n8750 ;
  assign y3114 = n8751 ;
  assign y3115 = n8754 ;
  assign y3116 = n8757 ;
  assign y3117 = ~n8759 ;
  assign y3118 = ~n8765 ;
  assign y3119 = ~n8766 ;
  assign y3120 = ~n8767 ;
  assign y3121 = n8774 ;
  assign y3122 = ~1'b0 ;
  assign y3123 = n8777 ;
  assign y3124 = ~n8781 ;
  assign y3125 = ~1'b0 ;
  assign y3126 = ~n8784 ;
  assign y3127 = n8787 ;
  assign y3128 = ~n8791 ;
  assign y3129 = ~1'b0 ;
  assign y3130 = ~1'b0 ;
  assign y3131 = ~1'b0 ;
  assign y3132 = ~1'b0 ;
  assign y3133 = ~n8794 ;
  assign y3134 = ~n6838 ;
  assign y3135 = ~n8799 ;
  assign y3136 = ~n8811 ;
  assign y3137 = ~n8814 ;
  assign y3138 = ~n8815 ;
  assign y3139 = n8821 ;
  assign y3140 = ~n8827 ;
  assign y3141 = n8828 ;
  assign y3142 = n8677 ;
  assign y3143 = n8835 ;
  assign y3144 = ~1'b0 ;
  assign y3145 = ~n5000 ;
  assign y3146 = n8836 ;
  assign y3147 = ~n8837 ;
  assign y3148 = ~1'b0 ;
  assign y3149 = n8838 ;
  assign y3150 = n8844 ;
  assign y3151 = ~1'b0 ;
  assign y3152 = n8847 ;
  assign y3153 = ~n8850 ;
  assign y3154 = ~1'b0 ;
  assign y3155 = n8855 ;
  assign y3156 = n8857 ;
  assign y3157 = n8858 ;
  assign y3158 = ~n8859 ;
  assign y3159 = ~n8865 ;
  assign y3160 = ~n8871 ;
  assign y3161 = n8872 ;
  assign y3162 = n8875 ;
  assign y3163 = ~1'b0 ;
  assign y3164 = ~1'b0 ;
  assign y3165 = ~n6336 ;
  assign y3166 = n8878 ;
  assign y3167 = n8880 ;
  assign y3168 = ~n8887 ;
  assign y3169 = n8888 ;
  assign y3170 = ~1'b0 ;
  assign y3171 = ~n8894 ;
  assign y3172 = n8896 ;
  assign y3173 = ~n8897 ;
  assign y3174 = ~n8904 ;
  assign y3175 = n8905 ;
  assign y3176 = ~1'b0 ;
  assign y3177 = ~n8911 ;
  assign y3178 = n8913 ;
  assign y3179 = n6110 ;
  assign y3180 = n8918 ;
  assign y3181 = ~n3636 ;
  assign y3182 = n8919 ;
  assign y3183 = ~n5963 ;
  assign y3184 = n8921 ;
  assign y3185 = ~1'b0 ;
  assign y3186 = ~1'b0 ;
  assign y3187 = ~1'b0 ;
  assign y3188 = n8923 ;
  assign y3189 = ~n8926 ;
  assign y3190 = ~n8927 ;
  assign y3191 = ~n8944 ;
  assign y3192 = ~n7996 ;
  assign y3193 = ~1'b0 ;
  assign y3194 = n8945 ;
  assign y3195 = n8947 ;
  assign y3196 = n8949 ;
  assign y3197 = n8951 ;
  assign y3198 = ~n8953 ;
  assign y3199 = ~n8957 ;
  assign y3200 = ~1'b0 ;
  assign y3201 = n8958 ;
  assign y3202 = ~n8963 ;
  assign y3203 = n8965 ;
  assign y3204 = ~n8972 ;
  assign y3205 = n8976 ;
  assign y3206 = ~1'b0 ;
  assign y3207 = n8979 ;
  assign y3208 = ~1'b0 ;
  assign y3209 = ~n8982 ;
  assign y3210 = ~n8987 ;
  assign y3211 = ~n8990 ;
  assign y3212 = n5955 ;
  assign y3213 = n8994 ;
  assign y3214 = ~1'b0 ;
  assign y3215 = n4147 ;
  assign y3216 = n8996 ;
  assign y3217 = ~n8998 ;
  assign y3218 = ~n9000 ;
  assign y3219 = ~1'b0 ;
  assign y3220 = ~n9002 ;
  assign y3221 = n9007 ;
  assign y3222 = ~n9017 ;
  assign y3223 = ~1'b0 ;
  assign y3224 = n9018 ;
  assign y3225 = ~n9019 ;
  assign y3226 = ~1'b0 ;
  assign y3227 = n9026 ;
  assign y3228 = n9027 ;
  assign y3229 = n9029 ;
  assign y3230 = ~n9031 ;
  assign y3231 = ~n9034 ;
  assign y3232 = ~n9041 ;
  assign y3233 = ~n9044 ;
  assign y3234 = ~n9045 ;
  assign y3235 = n9047 ;
  assign y3236 = ~n9048 ;
  assign y3237 = ~1'b0 ;
  assign y3238 = ~1'b0 ;
  assign y3239 = ~n9050 ;
  assign y3240 = ~n9057 ;
  assign y3241 = ~n9059 ;
  assign y3242 = ~1'b0 ;
  assign y3243 = ~n9060 ;
  assign y3244 = n9063 ;
  assign y3245 = n9065 ;
  assign y3246 = n9072 ;
  assign y3247 = ~1'b0 ;
  assign y3248 = n9075 ;
  assign y3249 = ~n9076 ;
  assign y3250 = n9077 ;
  assign y3251 = n9078 ;
  assign y3252 = n9081 ;
  assign y3253 = n9083 ;
  assign y3254 = ~n9084 ;
  assign y3255 = ~n9087 ;
  assign y3256 = ~n9090 ;
  assign y3257 = ~1'b0 ;
  assign y3258 = n9091 ;
  assign y3259 = ~n9094 ;
  assign y3260 = n9097 ;
  assign y3261 = ~n9106 ;
  assign y3262 = n9109 ;
  assign y3263 = ~n9111 ;
  assign y3264 = n9116 ;
  assign y3265 = ~1'b0 ;
  assign y3266 = n9117 ;
  assign y3267 = ~n9123 ;
  assign y3268 = ~1'b0 ;
  assign y3269 = ~1'b0 ;
  assign y3270 = ~n9125 ;
  assign y3271 = ~n9126 ;
  assign y3272 = ~n9129 ;
  assign y3273 = ~n9130 ;
  assign y3274 = ~1'b0 ;
  assign y3275 = n9138 ;
  assign y3276 = ~n9142 ;
  assign y3277 = ~n9149 ;
  assign y3278 = ~n9154 ;
  assign y3279 = ~1'b0 ;
  assign y3280 = ~n9155 ;
  assign y3281 = ~n9159 ;
  assign y3282 = ~n9160 ;
  assign y3283 = n9165 ;
  assign y3284 = n9171 ;
  assign y3285 = n9174 ;
  assign y3286 = n9193 ;
  assign y3287 = ~1'b0 ;
  assign y3288 = ~n9195 ;
  assign y3289 = n9196 ;
  assign y3290 = ~1'b0 ;
  assign y3291 = n9197 ;
  assign y3292 = n9198 ;
  assign y3293 = ~n9200 ;
  assign y3294 = ~n9204 ;
  assign y3295 = ~1'b0 ;
  assign y3296 = ~1'b0 ;
  assign y3297 = ~n9208 ;
  assign y3298 = ~n9209 ;
  assign y3299 = ~n9210 ;
  assign y3300 = ~n9212 ;
  assign y3301 = n5575 ;
  assign y3302 = ~n9213 ;
  assign y3303 = ~1'b0 ;
  assign y3304 = ~n9215 ;
  assign y3305 = n9218 ;
  assign y3306 = ~n9220 ;
  assign y3307 = ~n9222 ;
  assign y3308 = ~n9227 ;
  assign y3309 = ~1'b0 ;
  assign y3310 = ~n9230 ;
  assign y3311 = ~n9234 ;
  assign y3312 = n9240 ;
  assign y3313 = n9242 ;
  assign y3314 = ~n9247 ;
  assign y3315 = ~n9249 ;
  assign y3316 = ~1'b0 ;
  assign y3317 = n9252 ;
  assign y3318 = ~n9254 ;
  assign y3319 = ~n9259 ;
  assign y3320 = ~n9260 ;
  assign y3321 = ~n9264 ;
  assign y3322 = ~1'b0 ;
  assign y3323 = ~n9266 ;
  assign y3324 = ~n9267 ;
  assign y3325 = n9268 ;
  assign y3326 = ~1'b0 ;
  assign y3327 = ~1'b0 ;
  assign y3328 = n9270 ;
  assign y3329 = ~1'b0 ;
  assign y3330 = n9277 ;
  assign y3331 = n9280 ;
  assign y3332 = n9284 ;
  assign y3333 = ~1'b0 ;
  assign y3334 = ~n9285 ;
  assign y3335 = ~n9286 ;
  assign y3336 = n9289 ;
  assign y3337 = n214 ;
  assign y3338 = ~n9293 ;
  assign y3339 = ~1'b0 ;
  assign y3340 = ~1'b0 ;
  assign y3341 = ~1'b0 ;
  assign y3342 = ~n9298 ;
  assign y3343 = n9300 ;
  assign y3344 = n9311 ;
  assign y3345 = n9312 ;
  assign y3346 = ~n9313 ;
  assign y3347 = n853 ;
  assign y3348 = ~n9314 ;
  assign y3349 = 1'b0 ;
  assign y3350 = n265 ;
  assign y3351 = ~n9315 ;
  assign y3352 = ~n9319 ;
  assign y3353 = ~n9324 ;
  assign y3354 = ~1'b0 ;
  assign y3355 = ~1'b0 ;
  assign y3356 = ~1'b0 ;
  assign y3357 = ~n9325 ;
  assign y3358 = n9328 ;
  assign y3359 = ~n9330 ;
  assign y3360 = ~1'b0 ;
  assign y3361 = ~n9336 ;
  assign y3362 = ~1'b0 ;
  assign y3363 = n9337 ;
  assign y3364 = ~n9340 ;
  assign y3365 = ~n9342 ;
  assign y3366 = ~n9345 ;
  assign y3367 = ~n9347 ;
  assign y3368 = ~n7201 ;
  assign y3369 = n9348 ;
  assign y3370 = n5578 ;
  assign y3371 = ~1'b0 ;
  assign y3372 = n9352 ;
  assign y3373 = ~n9356 ;
  assign y3374 = n9359 ;
  assign y3375 = ~1'b0 ;
  assign y3376 = n9362 ;
  assign y3377 = ~1'b0 ;
  assign y3378 = ~n9367 ;
  assign y3379 = n9371 ;
  assign y3380 = ~n9372 ;
  assign y3381 = ~1'b0 ;
  assign y3382 = ~n9374 ;
  assign y3383 = ~n9377 ;
  assign y3384 = n9382 ;
  assign y3385 = ~n9386 ;
  assign y3386 = n9388 ;
  assign y3387 = ~n9395 ;
  assign y3388 = ~1'b0 ;
  assign y3389 = n9397 ;
  assign y3390 = n9398 ;
  assign y3391 = ~n9399 ;
  assign y3392 = ~n9400 ;
  assign y3393 = ~1'b0 ;
  assign y3394 = ~n9404 ;
  assign y3395 = n9405 ;
  assign y3396 = n9414 ;
  assign y3397 = n9422 ;
  assign y3398 = n9431 ;
  assign y3399 = n9433 ;
  assign y3400 = ~n9438 ;
  assign y3401 = n9440 ;
  assign y3402 = n9443 ;
  assign y3403 = n9449 ;
  assign y3404 = ~1'b0 ;
  assign y3405 = ~n9450 ;
  assign y3406 = ~n9454 ;
  assign y3407 = ~n9461 ;
  assign y3408 = n9470 ;
  assign y3409 = n9474 ;
  assign y3410 = ~1'b0 ;
  assign y3411 = ~n9485 ;
  assign y3412 = ~n9488 ;
  assign y3413 = ~1'b0 ;
  assign y3414 = ~n9490 ;
  assign y3415 = ~n9494 ;
  assign y3416 = ~1'b0 ;
  assign y3417 = ~n9497 ;
  assign y3418 = n9505 ;
  assign y3419 = ~n9512 ;
  assign y3420 = ~1'b0 ;
  assign y3421 = n9514 ;
  assign y3422 = ~n9518 ;
  assign y3423 = n9519 ;
  assign y3424 = ~n9521 ;
  assign y3425 = ~n9528 ;
  assign y3426 = n9538 ;
  assign y3427 = n9540 ;
  assign y3428 = ~n9542 ;
  assign y3429 = n9545 ;
  assign y3430 = n9552 ;
  assign y3431 = n9556 ;
  assign y3432 = n9565 ;
  assign y3433 = ~1'b0 ;
  assign y3434 = n9566 ;
  assign y3435 = n9570 ;
  assign y3436 = ~n9572 ;
  assign y3437 = ~n9577 ;
  assign y3438 = n9581 ;
  assign y3439 = ~1'b0 ;
  assign y3440 = ~n9583 ;
  assign y3441 = n9585 ;
  assign y3442 = ~n9587 ;
  assign y3443 = n9588 ;
  assign y3444 = ~1'b0 ;
  assign y3445 = ~n9589 ;
  assign y3446 = n9590 ;
  assign y3447 = ~n9596 ;
  assign y3448 = n9600 ;
  assign y3449 = ~n9603 ;
  assign y3450 = ~n9606 ;
  assign y3451 = n9607 ;
  assign y3452 = n9610 ;
  assign y3453 = ~n9613 ;
  assign y3454 = ~n9614 ;
  assign y3455 = n9618 ;
  assign y3456 = n9622 ;
  assign y3457 = n9625 ;
  assign y3458 = ~n9626 ;
  assign y3459 = ~n9634 ;
  assign y3460 = n9635 ;
  assign y3461 = n9639 ;
  assign y3462 = ~n9640 ;
  assign y3463 = n9641 ;
  assign y3464 = ~n9643 ;
  assign y3465 = ~n9644 ;
  assign y3466 = n9647 ;
  assign y3467 = ~n9653 ;
  assign y3468 = ~1'b0 ;
  assign y3469 = ~n9655 ;
  assign y3470 = ~1'b0 ;
  assign y3471 = n9657 ;
  assign y3472 = ~n9659 ;
  assign y3473 = ~1'b0 ;
  assign y3474 = n9664 ;
  assign y3475 = ~n9667 ;
  assign y3476 = ~n9670 ;
  assign y3477 = ~n9685 ;
  assign y3478 = ~1'b0 ;
  assign y3479 = ~n9687 ;
  assign y3480 = ~n9691 ;
  assign y3481 = ~n9692 ;
  assign y3482 = ~1'b0 ;
  assign y3483 = n9693 ;
  assign y3484 = ~n3729 ;
  assign y3485 = n9695 ;
  assign y3486 = ~n9696 ;
  assign y3487 = ~n9699 ;
  assign y3488 = n9701 ;
  assign y3489 = ~n9708 ;
  assign y3490 = ~n9714 ;
  assign y3491 = ~n9716 ;
  assign y3492 = ~n9717 ;
  assign y3493 = n9719 ;
  assign y3494 = n9721 ;
  assign y3495 = ~n9723 ;
  assign y3496 = ~n9726 ;
  assign y3497 = ~1'b0 ;
  assign y3498 = ~1'b0 ;
  assign y3499 = ~n9727 ;
  assign y3500 = ~n9729 ;
  assign y3501 = ~n9733 ;
  assign y3502 = ~n9734 ;
  assign y3503 = ~n9738 ;
  assign y3504 = ~n9740 ;
  assign y3505 = ~n9742 ;
  assign y3506 = ~n9745 ;
  assign y3507 = n9748 ;
  assign y3508 = ~1'b0 ;
  assign y3509 = ~1'b0 ;
  assign y3510 = ~n9749 ;
  assign y3511 = ~n9751 ;
  assign y3512 = n9753 ;
  assign y3513 = ~n9756 ;
  assign y3514 = n9763 ;
  assign y3515 = n9766 ;
  assign y3516 = n9768 ;
  assign y3517 = ~n2296 ;
  assign y3518 = n368 ;
  assign y3519 = n9771 ;
  assign y3520 = ~n9776 ;
  assign y3521 = ~n9778 ;
  assign y3522 = 1'b0 ;
  assign y3523 = n9783 ;
  assign y3524 = ~n9786 ;
  assign y3525 = n9790 ;
  assign y3526 = ~n9799 ;
  assign y3527 = n9805 ;
  assign y3528 = n9806 ;
  assign y3529 = ~n2695 ;
  assign y3530 = ~1'b0 ;
  assign y3531 = ~n9807 ;
  assign y3532 = n9810 ;
  assign y3533 = n9813 ;
  assign y3534 = ~1'b0 ;
  assign y3535 = n9824 ;
  assign y3536 = ~1'b0 ;
  assign y3537 = ~1'b0 ;
  assign y3538 = n9825 ;
  assign y3539 = n9826 ;
  assign y3540 = ~1'b0 ;
  assign y3541 = ~1'b0 ;
  assign y3542 = n9827 ;
  assign y3543 = ~n9828 ;
  assign y3544 = ~1'b0 ;
  assign y3545 = ~n9836 ;
  assign y3546 = n9837 ;
  assign y3547 = ~n9844 ;
  assign y3548 = ~n9851 ;
  assign y3549 = ~1'b0 ;
  assign y3550 = ~n9852 ;
  assign y3551 = ~n9853 ;
  assign y3552 = ~n9854 ;
  assign y3553 = n9856 ;
  assign y3554 = ~n9869 ;
  assign y3555 = ~1'b0 ;
  assign y3556 = n5269 ;
  assign y3557 = ~1'b0 ;
  assign y3558 = x13 ;
  assign y3559 = n9871 ;
  assign y3560 = ~n9874 ;
  assign y3561 = ~1'b0 ;
  assign y3562 = ~n9879 ;
  assign y3563 = ~1'b0 ;
  assign y3564 = ~n4550 ;
  assign y3565 = ~1'b0 ;
  assign y3566 = ~1'b0 ;
  assign y3567 = n9880 ;
  assign y3568 = n6872 ;
  assign y3569 = n9884 ;
  assign y3570 = n9888 ;
  assign y3571 = ~n6249 ;
  assign y3572 = n9891 ;
  assign y3573 = n9895 ;
  assign y3574 = ~n9896 ;
  assign y3575 = ~1'b0 ;
  assign y3576 = ~1'b0 ;
  assign y3577 = n9898 ;
  assign y3578 = ~n9900 ;
  assign y3579 = n9902 ;
  assign y3580 = ~n9906 ;
  assign y3581 = ~1'b0 ;
  assign y3582 = ~n9908 ;
  assign y3583 = n9909 ;
  assign y3584 = n9916 ;
  assign y3585 = ~n9918 ;
  assign y3586 = ~n9920 ;
  assign y3587 = ~n471 ;
  assign y3588 = ~1'b0 ;
  assign y3589 = ~n9924 ;
  assign y3590 = ~n9927 ;
  assign y3591 = n9932 ;
  assign y3592 = ~1'b0 ;
  assign y3593 = ~n9933 ;
  assign y3594 = n9936 ;
  assign y3595 = ~1'b0 ;
  assign y3596 = n9938 ;
  assign y3597 = n9939 ;
  assign y3598 = ~n9942 ;
  assign y3599 = ~n9947 ;
  assign y3600 = ~n9951 ;
  assign y3601 = ~1'b0 ;
  assign y3602 = ~1'b0 ;
  assign y3603 = n9964 ;
  assign y3604 = n9965 ;
  assign y3605 = ~n9968 ;
  assign y3606 = ~n9971 ;
  assign y3607 = ~n3610 ;
  assign y3608 = n9975 ;
  assign y3609 = n9978 ;
  assign y3610 = ~n9980 ;
  assign y3611 = n9985 ;
  assign y3612 = n9986 ;
  assign y3613 = n9988 ;
  assign y3614 = n9990 ;
  assign y3615 = ~n9996 ;
  assign y3616 = ~1'b0 ;
  assign y3617 = n9998 ;
  assign y3618 = n10000 ;
  assign y3619 = ~n10002 ;
  assign y3620 = n10009 ;
  assign y3621 = n10018 ;
  assign y3622 = ~1'b0 ;
  assign y3623 = ~n10021 ;
  assign y3624 = n10026 ;
  assign y3625 = ~1'b0 ;
  assign y3626 = ~1'b0 ;
  assign y3627 = n10028 ;
  assign y3628 = n10033 ;
  assign y3629 = n10045 ;
  assign y3630 = ~1'b0 ;
  assign y3631 = ~n10046 ;
  assign y3632 = n10054 ;
  assign y3633 = ~1'b0 ;
  assign y3634 = ~n10056 ;
  assign y3635 = n10059 ;
  assign y3636 = ~n10063 ;
  assign y3637 = ~n10065 ;
  assign y3638 = n10068 ;
  assign y3639 = ~n10069 ;
  assign y3640 = ~1'b0 ;
  assign y3641 = ~n10073 ;
  assign y3642 = ~n10074 ;
  assign y3643 = ~1'b0 ;
  assign y3644 = ~n10078 ;
  assign y3645 = n10081 ;
  assign y3646 = ~n10083 ;
  assign y3647 = ~n10085 ;
  assign y3648 = n10086 ;
  assign y3649 = ~n10088 ;
  assign y3650 = n10090 ;
  assign y3651 = n10092 ;
  assign y3652 = n10093 ;
  assign y3653 = n10097 ;
  assign y3654 = ~1'b0 ;
  assign y3655 = ~n10098 ;
  assign y3656 = ~1'b0 ;
  assign y3657 = ~n10099 ;
  assign y3658 = ~n10100 ;
  assign y3659 = ~1'b0 ;
  assign y3660 = ~1'b0 ;
  assign y3661 = n10102 ;
  assign y3662 = n10103 ;
  assign y3663 = ~1'b0 ;
  assign y3664 = ~n10105 ;
  assign y3665 = ~1'b0 ;
  assign y3666 = ~n10109 ;
  assign y3667 = ~n10115 ;
  assign y3668 = n10120 ;
  assign y3669 = n10122 ;
  assign y3670 = n10127 ;
  assign y3671 = ~n10128 ;
  assign y3672 = ~n10137 ;
  assign y3673 = ~n10140 ;
  assign y3674 = ~1'b0 ;
  assign y3675 = ~n10143 ;
  assign y3676 = ~1'b0 ;
  assign y3677 = ~1'b0 ;
  assign y3678 = ~n10147 ;
  assign y3679 = n10149 ;
  assign y3680 = n10153 ;
  assign y3681 = n10161 ;
  assign y3682 = n10164 ;
  assign y3683 = n10167 ;
  assign y3684 = n10174 ;
  assign y3685 = ~1'b0 ;
  assign y3686 = ~n10176 ;
  assign y3687 = ~n10179 ;
  assign y3688 = n10181 ;
  assign y3689 = ~n10183 ;
  assign y3690 = n10186 ;
  assign y3691 = n10188 ;
  assign y3692 = n10191 ;
  assign y3693 = ~1'b0 ;
  assign y3694 = ~n10193 ;
  assign y3695 = n10195 ;
  assign y3696 = ~n10201 ;
  assign y3697 = n10204 ;
  assign y3698 = n10207 ;
  assign y3699 = ~1'b0 ;
  assign y3700 = ~n10216 ;
  assign y3701 = ~n10217 ;
  assign y3702 = ~n10227 ;
  assign y3703 = n4329 ;
  assign y3704 = n903 ;
  assign y3705 = n10229 ;
  assign y3706 = n10230 ;
  assign y3707 = ~n10234 ;
  assign y3708 = n10235 ;
  assign y3709 = ~n10242 ;
  assign y3710 = n10244 ;
  assign y3711 = ~n10248 ;
  assign y3712 = n10254 ;
  assign y3713 = n10263 ;
  assign y3714 = ~n10265 ;
  assign y3715 = ~n10269 ;
  assign y3716 = ~1'b0 ;
  assign y3717 = ~n10276 ;
  assign y3718 = ~n10281 ;
  assign y3719 = 1'b0 ;
  assign y3720 = n10287 ;
  assign y3721 = n10288 ;
  assign y3722 = ~1'b0 ;
  assign y3723 = n10289 ;
  assign y3724 = n10293 ;
  assign y3725 = ~n10294 ;
  assign y3726 = ~1'b0 ;
  assign y3727 = n10295 ;
  assign y3728 = n10297 ;
  assign y3729 = ~1'b0 ;
  assign y3730 = ~1'b0 ;
  assign y3731 = ~n10298 ;
  assign y3732 = ~n10302 ;
  assign y3733 = ~n10307 ;
  assign y3734 = ~n10310 ;
  assign y3735 = n6914 ;
  assign y3736 = n10313 ;
  assign y3737 = ~n10315 ;
  assign y3738 = n10318 ;
  assign y3739 = n10331 ;
  assign y3740 = n10337 ;
  assign y3741 = ~1'b0 ;
  assign y3742 = ~n10338 ;
  assign y3743 = n10339 ;
  assign y3744 = n10342 ;
  assign y3745 = ~n10344 ;
  assign y3746 = ~n10345 ;
  assign y3747 = n10346 ;
  assign y3748 = ~n10347 ;
  assign y3749 = n10348 ;
  assign y3750 = ~n10349 ;
  assign y3751 = n10351 ;
  assign y3752 = n10354 ;
  assign y3753 = ~1'b0 ;
  assign y3754 = ~n10356 ;
  assign y3755 = n10357 ;
  assign y3756 = n10364 ;
  assign y3757 = ~n10366 ;
  assign y3758 = ~n10374 ;
  assign y3759 = ~n10375 ;
  assign y3760 = ~n10380 ;
  assign y3761 = ~1'b0 ;
  assign y3762 = ~n10382 ;
  assign y3763 = n10384 ;
  assign y3764 = ~n10386 ;
  assign y3765 = ~1'b0 ;
  assign y3766 = ~n10391 ;
  assign y3767 = n10394 ;
  assign y3768 = ~n10396 ;
  assign y3769 = n10399 ;
  assign y3770 = ~n10401 ;
  assign y3771 = ~n10403 ;
  assign y3772 = ~1'b0 ;
  assign y3773 = ~n10409 ;
  assign y3774 = n10412 ;
  assign y3775 = n10416 ;
  assign y3776 = n10420 ;
  assign y3777 = n10421 ;
  assign y3778 = n10425 ;
  assign y3779 = ~1'b0 ;
  assign y3780 = ~n10428 ;
  assign y3781 = n10433 ;
  assign y3782 = ~n10434 ;
  assign y3783 = ~n10438 ;
  assign y3784 = n10441 ;
  assign y3785 = n10443 ;
  assign y3786 = ~1'b0 ;
  assign y3787 = n10448 ;
  assign y3788 = ~n10451 ;
  assign y3789 = ~n10455 ;
  assign y3790 = ~n10456 ;
  assign y3791 = ~n1188 ;
  assign y3792 = ~1'b0 ;
  assign y3793 = ~n10457 ;
  assign y3794 = n10458 ;
  assign y3795 = ~n10459 ;
  assign y3796 = n10461 ;
  assign y3797 = ~n10465 ;
  assign y3798 = n10468 ;
  assign y3799 = ~n10469 ;
  assign y3800 = n10470 ;
  assign y3801 = ~1'b0 ;
  assign y3802 = n10472 ;
  assign y3803 = n10475 ;
  assign y3804 = ~n10480 ;
  assign y3805 = ~n10481 ;
  assign y3806 = n10482 ;
  assign y3807 = ~n8952 ;
  assign y3808 = 1'b0 ;
  assign y3809 = ~1'b0 ;
  assign y3810 = ~n10485 ;
  assign y3811 = ~n7622 ;
  assign y3812 = n10487 ;
  assign y3813 = n10491 ;
  assign y3814 = ~1'b0 ;
  assign y3815 = n10495 ;
  assign y3816 = n10496 ;
  assign y3817 = 1'b0 ;
  assign y3818 = ~1'b0 ;
  assign y3819 = n10509 ;
  assign y3820 = n10511 ;
  assign y3821 = ~n10512 ;
  assign y3822 = 1'b0 ;
  assign y3823 = ~1'b0 ;
  assign y3824 = ~n10513 ;
  assign y3825 = ~n10515 ;
  assign y3826 = ~1'b0 ;
  assign y3827 = ~1'b0 ;
  assign y3828 = n10517 ;
  assign y3829 = ~n10518 ;
  assign y3830 = 1'b0 ;
  assign y3831 = n10521 ;
  assign y3832 = ~n10530 ;
  assign y3833 = ~n10546 ;
  assign y3834 = ~n10550 ;
  assign y3835 = ~1'b0 ;
  assign y3836 = ~n10552 ;
  assign y3837 = n10561 ;
  assign y3838 = ~1'b0 ;
  assign y3839 = n10564 ;
  assign y3840 = ~n7023 ;
  assign y3841 = ~1'b0 ;
  assign y3842 = 1'b0 ;
  assign y3843 = ~n4416 ;
  assign y3844 = n10566 ;
  assign y3845 = n10571 ;
  assign y3846 = n10572 ;
  assign y3847 = n10578 ;
  assign y3848 = n10584 ;
  assign y3849 = n10586 ;
  assign y3850 = ~n10587 ;
  assign y3851 = n10594 ;
  assign y3852 = ~n10596 ;
  assign y3853 = ~1'b0 ;
  assign y3854 = n10597 ;
  assign y3855 = ~n10598 ;
  assign y3856 = ~n10601 ;
  assign y3857 = ~1'b0 ;
  assign y3858 = ~1'b0 ;
  assign y3859 = ~n10604 ;
  assign y3860 = ~1'b0 ;
  assign y3861 = ~n10607 ;
  assign y3862 = n10612 ;
  assign y3863 = n10615 ;
  assign y3864 = ~n10617 ;
  assign y3865 = ~1'b0 ;
  assign y3866 = ~n10624 ;
  assign y3867 = ~n10632 ;
  assign y3868 = n10634 ;
  assign y3869 = n10635 ;
  assign y3870 = ~1'b0 ;
  assign y3871 = ~n3012 ;
  assign y3872 = n10637 ;
  assign y3873 = n10641 ;
  assign y3874 = ~n10644 ;
  assign y3875 = ~1'b0 ;
  assign y3876 = ~n10648 ;
  assign y3877 = ~n10651 ;
  assign y3878 = n5880 ;
  assign y3879 = ~1'b0 ;
  assign y3880 = ~n10653 ;
  assign y3881 = ~n10655 ;
  assign y3882 = ~n10661 ;
  assign y3883 = ~n10664 ;
  assign y3884 = n10670 ;
  assign y3885 = n10672 ;
  assign y3886 = ~1'b0 ;
  assign y3887 = ~1'b0 ;
  assign y3888 = ~1'b0 ;
  assign y3889 = ~n10676 ;
  assign y3890 = ~n10679 ;
  assign y3891 = n10681 ;
  assign y3892 = ~1'b0 ;
  assign y3893 = ~n10685 ;
  assign y3894 = ~1'b0 ;
  assign y3895 = ~n10687 ;
  assign y3896 = n10690 ;
  assign y3897 = ~n10694 ;
  assign y3898 = ~1'b0 ;
  assign y3899 = ~1'b0 ;
  assign y3900 = n10696 ;
  assign y3901 = ~n10701 ;
  assign y3902 = ~1'b0 ;
  assign y3903 = ~n10703 ;
  assign y3904 = ~n10718 ;
  assign y3905 = ~n10722 ;
  assign y3906 = ~n10725 ;
  assign y3907 = ~n10727 ;
  assign y3908 = 1'b0 ;
  assign y3909 = ~1'b0 ;
  assign y3910 = n10736 ;
  assign y3911 = ~n10741 ;
  assign y3912 = ~1'b0 ;
  assign y3913 = ~n10742 ;
  assign y3914 = ~n10746 ;
  assign y3915 = ~1'b0 ;
  assign y3916 = n10750 ;
  assign y3917 = ~n10758 ;
  assign y3918 = ~n10759 ;
  assign y3919 = n10760 ;
  assign y3920 = n4719 ;
  assign y3921 = n10767 ;
  assign y3922 = n10773 ;
  assign y3923 = n10782 ;
  assign y3924 = ~n10785 ;
  assign y3925 = ~1'b0 ;
  assign y3926 = ~n10791 ;
  assign y3927 = ~n10796 ;
  assign y3928 = ~n8272 ;
  assign y3929 = ~n10799 ;
  assign y3930 = ~n10802 ;
  assign y3931 = n10806 ;
  assign y3932 = n10808 ;
  assign y3933 = ~n10811 ;
  assign y3934 = n10817 ;
  assign y3935 = ~1'b0 ;
  assign y3936 = ~n10820 ;
  assign y3937 = ~1'b0 ;
  assign y3938 = n10821 ;
  assign y3939 = ~n10823 ;
  assign y3940 = n10827 ;
  assign y3941 = n10829 ;
  assign y3942 = ~1'b0 ;
  assign y3943 = ~1'b0 ;
  assign y3944 = ~1'b0 ;
  assign y3945 = ~n10832 ;
  assign y3946 = ~1'b0 ;
  assign y3947 = ~n10845 ;
  assign y3948 = ~1'b0 ;
  assign y3949 = n10851 ;
  assign y3950 = n10852 ;
  assign y3951 = ~1'b0 ;
  assign y3952 = ~1'b0 ;
  assign y3953 = n10853 ;
  assign y3954 = n10856 ;
  assign y3955 = ~n10858 ;
  assign y3956 = ~1'b0 ;
  assign y3957 = n10859 ;
  assign y3958 = ~n10863 ;
  assign y3959 = ~n10870 ;
  assign y3960 = n10871 ;
  assign y3961 = ~1'b0 ;
  assign y3962 = ~1'b0 ;
  assign y3963 = n1867 ;
  assign y3964 = n10878 ;
  assign y3965 = ~n10880 ;
  assign y3966 = ~1'b0 ;
  assign y3967 = n10882 ;
  assign y3968 = n10891 ;
  assign y3969 = ~n10892 ;
  assign y3970 = ~n10893 ;
  assign y3971 = n10894 ;
  assign y3972 = ~n10896 ;
  assign y3973 = ~1'b0 ;
  assign y3974 = n10897 ;
  assign y3975 = n10898 ;
  assign y3976 = n10901 ;
  assign y3977 = n10907 ;
  assign y3978 = ~n10909 ;
  assign y3979 = n10916 ;
  assign y3980 = n10918 ;
  assign y3981 = n10921 ;
  assign y3982 = n10924 ;
  assign y3983 = n10925 ;
  assign y3984 = ~1'b0 ;
  assign y3985 = n3796 ;
  assign y3986 = n10928 ;
  assign y3987 = ~n10931 ;
  assign y3988 = n10932 ;
  assign y3989 = ~n10935 ;
  assign y3990 = ~n10938 ;
  assign y3991 = n10940 ;
  assign y3992 = n10945 ;
  assign y3993 = ~n10946 ;
  assign y3994 = ~n10947 ;
  assign y3995 = ~n10952 ;
  assign y3996 = n10954 ;
  assign y3997 = ~1'b0 ;
  assign y3998 = x3 ;
  assign y3999 = n10956 ;
  assign y4000 = n10961 ;
  assign y4001 = ~1'b0 ;
  assign y4002 = ~n10962 ;
  assign y4003 = ~1'b0 ;
  assign y4004 = ~n10963 ;
  assign y4005 = ~n10966 ;
  assign y4006 = ~1'b0 ;
  assign y4007 = n10967 ;
  assign y4008 = ~1'b0 ;
  assign y4009 = ~n10973 ;
  assign y4010 = ~1'b0 ;
  assign y4011 = n10977 ;
  assign y4012 = n10981 ;
  assign y4013 = ~n10984 ;
  assign y4014 = n10985 ;
  assign y4015 = n10988 ;
  assign y4016 = ~n10990 ;
  assign y4017 = ~1'b0 ;
  assign y4018 = 1'b0 ;
  assign y4019 = n10995 ;
  assign y4020 = ~n10999 ;
  assign y4021 = n11000 ;
  assign y4022 = ~1'b0 ;
  assign y4023 = ~n10665 ;
  assign y4024 = n11002 ;
  assign y4025 = n11012 ;
  assign y4026 = ~n11013 ;
  assign y4027 = n11016 ;
  assign y4028 = n11030 ;
  assign y4029 = n11034 ;
  assign y4030 = ~n11038 ;
  assign y4031 = ~n11044 ;
  assign y4032 = n11054 ;
  assign y4033 = ~1'b0 ;
  assign y4034 = ~n11061 ;
  assign y4035 = n11062 ;
  assign y4036 = n11065 ;
  assign y4037 = ~n11068 ;
  assign y4038 = ~n11075 ;
  assign y4039 = ~n11076 ;
  assign y4040 = ~n11079 ;
  assign y4041 = n11088 ;
  assign y4042 = n11090 ;
  assign y4043 = ~1'b0 ;
  assign y4044 = ~1'b0 ;
  assign y4045 = n11092 ;
  assign y4046 = n11096 ;
  assign y4047 = ~n11103 ;
  assign y4048 = ~1'b0 ;
  assign y4049 = ~1'b0 ;
  assign y4050 = ~n11104 ;
  assign y4051 = n11110 ;
  assign y4052 = n11112 ;
  assign y4053 = ~1'b0 ;
  assign y4054 = ~n11114 ;
  assign y4055 = ~n11121 ;
  assign y4056 = n11124 ;
  assign y4057 = n11125 ;
  assign y4058 = ~1'b0 ;
  assign y4059 = ~n11127 ;
  assign y4060 = ~n11128 ;
  assign y4061 = n11131 ;
  assign y4062 = ~n11134 ;
  assign y4063 = ~1'b0 ;
  assign y4064 = ~n11138 ;
  assign y4065 = n11139 ;
  assign y4066 = n11140 ;
  assign y4067 = ~1'b0 ;
  assign y4068 = ~n11141 ;
  assign y4069 = n11142 ;
  assign y4070 = n11150 ;
  assign y4071 = n7663 ;
  assign y4072 = n11162 ;
  assign y4073 = n11171 ;
  assign y4074 = ~n11173 ;
  assign y4075 = ~n11174 ;
  assign y4076 = n11181 ;
  assign y4077 = n11183 ;
  assign y4078 = ~n11184 ;
  assign y4079 = ~1'b0 ;
  assign y4080 = n11192 ;
  assign y4081 = n11196 ;
  assign y4082 = ~n11199 ;
  assign y4083 = ~n11201 ;
  assign y4084 = n11202 ;
  assign y4085 = ~n11208 ;
  assign y4086 = n1914 ;
  assign y4087 = ~1'b0 ;
  assign y4088 = ~n11210 ;
  assign y4089 = ~1'b0 ;
  assign y4090 = ~n11213 ;
  assign y4091 = ~1'b0 ;
  assign y4092 = ~n11217 ;
  assign y4093 = ~n11218 ;
  assign y4094 = ~n11223 ;
  assign y4095 = n11225 ;
  assign y4096 = n11227 ;
  assign y4097 = ~n11240 ;
  assign y4098 = ~n11244 ;
  assign y4099 = n11246 ;
  assign y4100 = n11247 ;
  assign y4101 = ~1'b0 ;
  assign y4102 = ~n11250 ;
  assign y4103 = ~1'b0 ;
  assign y4104 = ~n11251 ;
  assign y4105 = ~n11252 ;
  assign y4106 = n11255 ;
  assign y4107 = n11258 ;
  assign y4108 = ~n11260 ;
  assign y4109 = ~1'b0 ;
  assign y4110 = n11263 ;
  assign y4111 = n11264 ;
  assign y4112 = ~n11267 ;
  assign y4113 = ~n11268 ;
  assign y4114 = n11271 ;
  assign y4115 = ~n11274 ;
  assign y4116 = ~n11277 ;
  assign y4117 = n11280 ;
  assign y4118 = 1'b0 ;
  assign y4119 = n11284 ;
  assign y4120 = ~n11286 ;
  assign y4121 = n11289 ;
  assign y4122 = n11298 ;
  assign y4123 = n11299 ;
  assign y4124 = ~1'b0 ;
  assign y4125 = ~n11308 ;
  assign y4126 = n11313 ;
  assign y4127 = n11314 ;
  assign y4128 = n11315 ;
  assign y4129 = n11317 ;
  assign y4130 = ~n11318 ;
  assign y4131 = n11320 ;
  assign y4132 = ~1'b0 ;
  assign y4133 = n7685 ;
  assign y4134 = 1'b0 ;
  assign y4135 = n11325 ;
  assign y4136 = ~n11331 ;
  assign y4137 = ~n11334 ;
  assign y4138 = ~1'b0 ;
  assign y4139 = n11336 ;
  assign y4140 = n11337 ;
  assign y4141 = ~n11350 ;
  assign y4142 = n11354 ;
  assign y4143 = ~n325 ;
  assign y4144 = ~n11358 ;
  assign y4145 = n11359 ;
  assign y4146 = ~n11366 ;
  assign y4147 = n11372 ;
  assign y4148 = n4054 ;
  assign y4149 = n11373 ;
  assign y4150 = n201 ;
  assign y4151 = ~n11377 ;
  assign y4152 = ~1'b0 ;
  assign y4153 = ~1'b0 ;
  assign y4154 = ~1'b0 ;
  assign y4155 = n11378 ;
  assign y4156 = ~n11385 ;
  assign y4157 = ~1'b0 ;
  assign y4158 = ~n11390 ;
  assign y4159 = ~1'b0 ;
  assign y4160 = ~n11402 ;
  assign y4161 = ~n11403 ;
  assign y4162 = n11404 ;
  assign y4163 = n11407 ;
  assign y4164 = n11415 ;
  assign y4165 = ~n11417 ;
  assign y4166 = ~1'b0 ;
  assign y4167 = ~1'b0 ;
  assign y4168 = n6444 ;
  assign y4169 = ~n11421 ;
  assign y4170 = ~n11425 ;
  assign y4171 = n11426 ;
  assign y4172 = n11427 ;
  assign y4173 = ~n11428 ;
  assign y4174 = ~n11437 ;
  assign y4175 = n11439 ;
  assign y4176 = ~n11445 ;
  assign y4177 = ~n11453 ;
  assign y4178 = n11476 ;
  assign y4179 = ~n11480 ;
  assign y4180 = ~1'b0 ;
  assign y4181 = n11483 ;
  assign y4182 = ~1'b0 ;
  assign y4183 = ~n11486 ;
  assign y4184 = ~n11487 ;
  assign y4185 = 1'b0 ;
  assign y4186 = ~n11490 ;
  assign y4187 = ~n11492 ;
  assign y4188 = ~1'b0 ;
  assign y4189 = ~n11493 ;
  assign y4190 = ~n11502 ;
  assign y4191 = n11503 ;
  assign y4192 = n11506 ;
  assign y4193 = ~n11508 ;
  assign y4194 = n11511 ;
  assign y4195 = ~n11512 ;
  assign y4196 = n11513 ;
  assign y4197 = n11515 ;
  assign y4198 = ~n11517 ;
  assign y4199 = ~n11518 ;
  assign y4200 = n11519 ;
  assign y4201 = n11522 ;
  assign y4202 = n11526 ;
  assign y4203 = n11529 ;
  assign y4204 = n11535 ;
  assign y4205 = n11540 ;
  assign y4206 = ~n9324 ;
  assign y4207 = ~n11544 ;
  assign y4208 = ~n11545 ;
  assign y4209 = n11548 ;
  assign y4210 = n11552 ;
  assign y4211 = n11555 ;
  assign y4212 = ~n11559 ;
  assign y4213 = n11568 ;
  assign y4214 = n11571 ;
  assign y4215 = ~n11574 ;
  assign y4216 = ~1'b0 ;
  assign y4217 = ~n11577 ;
  assign y4218 = ~n11578 ;
  assign y4219 = ~1'b0 ;
  assign y4220 = ~1'b0 ;
  assign y4221 = n11580 ;
  assign y4222 = n11582 ;
  assign y4223 = n11585 ;
  assign y4224 = ~n11587 ;
  assign y4225 = ~n11588 ;
  assign y4226 = ~n7221 ;
  assign y4227 = ~1'b0 ;
  assign y4228 = ~n11594 ;
  assign y4229 = ~1'b0 ;
  assign y4230 = n11597 ;
  assign y4231 = ~n6017 ;
  assign y4232 = ~n11599 ;
  assign y4233 = ~1'b0 ;
  assign y4234 = n11602 ;
  assign y4235 = ~n11603 ;
  assign y4236 = ~n11606 ;
  assign y4237 = ~n11607 ;
  assign y4238 = n11610 ;
  assign y4239 = ~n11612 ;
  assign y4240 = n11613 ;
  assign y4241 = ~1'b0 ;
  assign y4242 = n11615 ;
  assign y4243 = ~n11620 ;
  assign y4244 = ~1'b0 ;
  assign y4245 = ~1'b0 ;
  assign y4246 = ~1'b0 ;
  assign y4247 = ~n11622 ;
  assign y4248 = n11628 ;
  assign y4249 = ~n11632 ;
  assign y4250 = ~n11633 ;
  assign y4251 = ~n11634 ;
  assign y4252 = ~n11635 ;
  assign y4253 = n11636 ;
  assign y4254 = ~1'b0 ;
  assign y4255 = ~1'b0 ;
  assign y4256 = ~n11639 ;
  assign y4257 = ~1'b0 ;
  assign y4258 = n11641 ;
  assign y4259 = ~n11642 ;
  assign y4260 = ~n11644 ;
  assign y4261 = ~1'b0 ;
  assign y4262 = n11649 ;
  assign y4263 = ~n11652 ;
  assign y4264 = ~n11655 ;
  assign y4265 = ~n11656 ;
  assign y4266 = n11661 ;
  assign y4267 = ~1'b0 ;
  assign y4268 = ~1'b0 ;
  assign y4269 = n11662 ;
  assign y4270 = ~n11663 ;
  assign y4271 = ~n11669 ;
  assign y4272 = n11681 ;
  assign y4273 = n11686 ;
  assign y4274 = n11687 ;
  assign y4275 = ~n11690 ;
  assign y4276 = ~n11697 ;
  assign y4277 = ~n11701 ;
  assign y4278 = ~n11702 ;
  assign y4279 = n11704 ;
  assign y4280 = n11710 ;
  assign y4281 = ~n11711 ;
  assign y4282 = n11712 ;
  assign y4283 = ~1'b0 ;
  assign y4284 = ~1'b0 ;
  assign y4285 = ~n374 ;
  assign y4286 = ~n11714 ;
  assign y4287 = n11716 ;
  assign y4288 = n11720 ;
  assign y4289 = ~n11725 ;
  assign y4290 = n11729 ;
  assign y4291 = ~1'b0 ;
  assign y4292 = ~n7824 ;
  assign y4293 = n11735 ;
  assign y4294 = n11738 ;
  assign y4295 = ~1'b0 ;
  assign y4296 = ~n11739 ;
  assign y4297 = n9703 ;
  assign y4298 = ~1'b0 ;
  assign y4299 = n11742 ;
  assign y4300 = n11746 ;
  assign y4301 = ~n11749 ;
  assign y4302 = n11752 ;
  assign y4303 = ~n11753 ;
  assign y4304 = n11757 ;
  assign y4305 = ~1'b0 ;
  assign y4306 = ~n11762 ;
  assign y4307 = ~n11767 ;
  assign y4308 = ~1'b0 ;
  assign y4309 = n11771 ;
  assign y4310 = ~1'b0 ;
  assign y4311 = ~1'b0 ;
  assign y4312 = ~n11773 ;
  assign y4313 = n11775 ;
  assign y4314 = ~n11777 ;
  assign y4315 = n11781 ;
  assign y4316 = 1'b0 ;
  assign y4317 = n11784 ;
  assign y4318 = n11785 ;
  assign y4319 = n11791 ;
  assign y4320 = ~n11801 ;
  assign y4321 = ~1'b0 ;
  assign y4322 = ~n11630 ;
  assign y4323 = ~n11803 ;
  assign y4324 = ~1'b0 ;
  assign y4325 = ~1'b0 ;
  assign y4326 = ~1'b0 ;
  assign y4327 = ~1'b0 ;
  assign y4328 = ~n11804 ;
  assign y4329 = ~n11806 ;
  assign y4330 = ~n11807 ;
  assign y4331 = ~n11811 ;
  assign y4332 = n11812 ;
  assign y4333 = ~n11813 ;
  assign y4334 = n11814 ;
  assign y4335 = n11817 ;
  assign y4336 = ~1'b0 ;
  assign y4337 = ~n11820 ;
  assign y4338 = ~n11824 ;
  assign y4339 = ~n11827 ;
  assign y4340 = ~1'b0 ;
  assign y4341 = ~1'b0 ;
  assign y4342 = ~n11828 ;
  assign y4343 = ~n11829 ;
  assign y4344 = ~n11831 ;
  assign y4345 = n11834 ;
  assign y4346 = n11835 ;
  assign y4347 = n11838 ;
  assign y4348 = ~1'b0 ;
  assign y4349 = ~1'b0 ;
  assign y4350 = n11839 ;
  assign y4351 = ~n11844 ;
  assign y4352 = n11846 ;
  assign y4353 = ~n11847 ;
  assign y4354 = n11855 ;
  assign y4355 = 1'b0 ;
  assign y4356 = 1'b0 ;
  assign y4357 = ~1'b0 ;
  assign y4358 = n11863 ;
  assign y4359 = n11865 ;
  assign y4360 = ~1'b0 ;
  assign y4361 = ~n3011 ;
  assign y4362 = n11866 ;
  assign y4363 = ~1'b0 ;
  assign y4364 = n11867 ;
  assign y4365 = n11868 ;
  assign y4366 = ~n11874 ;
  assign y4367 = n6560 ;
  assign y4368 = ~n11876 ;
  assign y4369 = n11878 ;
  assign y4370 = ~1'b0 ;
  assign y4371 = ~1'b0 ;
  assign y4372 = ~1'b0 ;
  assign y4373 = ~1'b0 ;
  assign y4374 = ~1'b0 ;
  assign y4375 = ~1'b0 ;
  assign y4376 = ~n11885 ;
  assign y4377 = n11886 ;
  assign y4378 = n11889 ;
  assign y4379 = ~1'b0 ;
  assign y4380 = ~n11891 ;
  assign y4381 = n11893 ;
  assign y4382 = ~1'b0 ;
  assign y4383 = n7837 ;
  assign y4384 = ~1'b0 ;
  assign y4385 = n11901 ;
  assign y4386 = n11907 ;
  assign y4387 = ~n11913 ;
  assign y4388 = n11916 ;
  assign y4389 = ~n11917 ;
  assign y4390 = ~n11919 ;
  assign y4391 = n11922 ;
  assign y4392 = ~n11928 ;
  assign y4393 = n11933 ;
  assign y4394 = n11939 ;
  assign y4395 = ~n11940 ;
  assign y4396 = ~n11949 ;
  assign y4397 = ~n11952 ;
  assign y4398 = n11955 ;
  assign y4399 = ~1'b0 ;
  assign y4400 = ~n11957 ;
  assign y4401 = ~1'b0 ;
  assign y4402 = ~n11963 ;
  assign y4403 = n11964 ;
  assign y4404 = ~n11966 ;
  assign y4405 = ~n11969 ;
  assign y4406 = n11972 ;
  assign y4407 = ~n11976 ;
  assign y4408 = n11977 ;
  assign y4409 = ~n11982 ;
  assign y4410 = ~n11985 ;
  assign y4411 = n11987 ;
  assign y4412 = ~n11988 ;
  assign y4413 = n11991 ;
  assign y4414 = ~1'b0 ;
  assign y4415 = n216 ;
  assign y4416 = n11992 ;
  assign y4417 = n11993 ;
  assign y4418 = n11997 ;
  assign y4419 = n11999 ;
  assign y4420 = n12002 ;
  assign y4421 = ~n12005 ;
  assign y4422 = n12008 ;
  assign y4423 = ~1'b0 ;
  assign y4424 = ~n12010 ;
  assign y4425 = n12013 ;
  assign y4426 = ~1'b0 ;
  assign y4427 = n12014 ;
  assign y4428 = n12021 ;
  assign y4429 = ~n12022 ;
  assign y4430 = ~n12025 ;
  assign y4431 = ~n12029 ;
  assign y4432 = n12036 ;
  assign y4433 = ~1'b0 ;
  assign y4434 = ~n9016 ;
  assign y4435 = n12038 ;
  assign y4436 = ~1'b0 ;
  assign y4437 = n12040 ;
  assign y4438 = n12041 ;
  assign y4439 = ~n12044 ;
  assign y4440 = n12048 ;
  assign y4441 = ~n12053 ;
  assign y4442 = n12057 ;
  assign y4443 = ~n12061 ;
  assign y4444 = ~n12064 ;
  assign y4445 = n12065 ;
  assign y4446 = n12066 ;
  assign y4447 = ~n12069 ;
  assign y4448 = ~n12072 ;
  assign y4449 = n12073 ;
  assign y4450 = ~1'b0 ;
  assign y4451 = ~n12075 ;
  assign y4452 = ~n12077 ;
  assign y4453 = n12078 ;
  assign y4454 = n12082 ;
  assign y4455 = n12087 ;
  assign y4456 = ~1'b0 ;
  assign y4457 = n12090 ;
  assign y4458 = n12091 ;
  assign y4459 = n12100 ;
  assign y4460 = n12102 ;
  assign y4461 = n12105 ;
  assign y4462 = ~n12106 ;
  assign y4463 = ~n12113 ;
  assign y4464 = n10841 ;
  assign y4465 = n12114 ;
  assign y4466 = ~n12116 ;
  assign y4467 = n12124 ;
  assign y4468 = n12125 ;
  assign y4469 = ~n12129 ;
  assign y4470 = n12132 ;
  assign y4471 = n12134 ;
  assign y4472 = n12135 ;
  assign y4473 = n12138 ;
  assign y4474 = n12140 ;
  assign y4475 = n12141 ;
  assign y4476 = n12146 ;
  assign y4477 = ~1'b0 ;
  assign y4478 = ~1'b0 ;
  assign y4479 = n12147 ;
  assign y4480 = ~n12149 ;
  assign y4481 = ~1'b0 ;
  assign y4482 = ~n12150 ;
  assign y4483 = n12152 ;
  assign y4484 = ~1'b0 ;
  assign y4485 = ~n12155 ;
  assign y4486 = ~1'b0 ;
  assign y4487 = n12162 ;
  assign y4488 = ~n12164 ;
  assign y4489 = ~n12165 ;
  assign y4490 = n12167 ;
  assign y4491 = n12172 ;
  assign y4492 = n12176 ;
  assign y4493 = ~n12178 ;
  assign y4494 = ~1'b0 ;
  assign y4495 = ~n12180 ;
  assign y4496 = ~n12181 ;
  assign y4497 = ~n12183 ;
  assign y4498 = ~1'b0 ;
  assign y4499 = ~n12186 ;
  assign y4500 = ~1'b0 ;
  assign y4501 = n12196 ;
  assign y4502 = ~1'b0 ;
  assign y4503 = n12197 ;
  assign y4504 = ~n12198 ;
  assign y4505 = n12201 ;
  assign y4506 = n12204 ;
  assign y4507 = n12205 ;
  assign y4508 = n12206 ;
  assign y4509 = ~1'b0 ;
  assign y4510 = ~n12207 ;
  assign y4511 = ~n12211 ;
  assign y4512 = ~1'b0 ;
  assign y4513 = n12221 ;
  assign y4514 = ~n6038 ;
  assign y4515 = ~1'b0 ;
  assign y4516 = n12225 ;
  assign y4517 = ~1'b0 ;
  assign y4518 = ~n12230 ;
  assign y4519 = ~n12231 ;
  assign y4520 = n12236 ;
  assign y4521 = ~n12238 ;
  assign y4522 = ~n12239 ;
  assign y4523 = ~n12246 ;
  assign y4524 = ~n12253 ;
  assign y4525 = ~1'b0 ;
  assign y4526 = ~1'b0 ;
  assign y4527 = ~n12254 ;
  assign y4528 = ~1'b0 ;
  assign y4529 = ~n12256 ;
  assign y4530 = ~n12257 ;
  assign y4531 = ~1'b0 ;
  assign y4532 = ~n12259 ;
  assign y4533 = ~1'b0 ;
  assign y4534 = n12261 ;
  assign y4535 = ~1'b0 ;
  assign y4536 = ~n12262 ;
  assign y4537 = ~n12263 ;
  assign y4538 = ~n12265 ;
  assign y4539 = ~1'b0 ;
  assign y4540 = n12267 ;
  assign y4541 = ~n12268 ;
  assign y4542 = n12269 ;
  assign y4543 = n12271 ;
  assign y4544 = ~1'b0 ;
  assign y4545 = ~n12273 ;
  assign y4546 = ~n4414 ;
  assign y4547 = n12274 ;
  assign y4548 = ~1'b0 ;
  assign y4549 = n12275 ;
  assign y4550 = ~1'b0 ;
  assign y4551 = n12277 ;
  assign y4552 = n12279 ;
  assign y4553 = n12281 ;
  assign y4554 = n12283 ;
  assign y4555 = ~n12284 ;
  assign y4556 = ~n12286 ;
  assign y4557 = ~1'b0 ;
  assign y4558 = ~n12288 ;
  assign y4559 = n12289 ;
  assign y4560 = n12291 ;
  assign y4561 = ~1'b0 ;
  assign y4562 = ~n12293 ;
  assign y4563 = ~n12296 ;
  assign y4564 = n12301 ;
  assign y4565 = ~n10423 ;
  assign y4566 = n3186 ;
  assign y4567 = ~n12303 ;
  assign y4568 = ~1'b0 ;
  assign y4569 = n12309 ;
  assign y4570 = n12319 ;
  assign y4571 = ~1'b0 ;
  assign y4572 = ~n12323 ;
  assign y4573 = ~n12326 ;
  assign y4574 = ~1'b0 ;
  assign y4575 = ~n12330 ;
  assign y4576 = n6003 ;
  assign y4577 = ~n12331 ;
  assign y4578 = n10931 ;
  assign y4579 = ~n12335 ;
  assign y4580 = ~n12347 ;
  assign y4581 = n12348 ;
  assign y4582 = n12350 ;
  assign y4583 = ~1'b0 ;
  assign y4584 = ~n12352 ;
  assign y4585 = ~n12353 ;
  assign y4586 = ~n12358 ;
  assign y4587 = n12360 ;
  assign y4588 = ~1'b0 ;
  assign y4589 = ~n12369 ;
  assign y4590 = ~n7554 ;
  assign y4591 = n12374 ;
  assign y4592 = ~1'b0 ;
  assign y4593 = n12377 ;
  assign y4594 = n12381 ;
  assign y4595 = ~1'b0 ;
  assign y4596 = n12382 ;
  assign y4597 = ~1'b0 ;
  assign y4598 = n6787 ;
  assign y4599 = n12384 ;
  assign y4600 = ~n12389 ;
  assign y4601 = ~1'b0 ;
  assign y4602 = ~1'b0 ;
  assign y4603 = ~1'b0 ;
  assign y4604 = n12393 ;
  assign y4605 = n12394 ;
  assign y4606 = n12398 ;
  assign y4607 = ~n12401 ;
  assign y4608 = n12406 ;
  assign y4609 = ~1'b0 ;
  assign y4610 = ~1'b0 ;
  assign y4611 = ~n12411 ;
  assign y4612 = n12412 ;
  assign y4613 = n12421 ;
  assign y4614 = ~1'b0 ;
  assign y4615 = n12423 ;
  assign y4616 = ~n12424 ;
  assign y4617 = ~n3762 ;
  assign y4618 = ~n12427 ;
  assign y4619 = ~n12433 ;
  assign y4620 = ~n12435 ;
  assign y4621 = ~n12440 ;
  assign y4622 = ~1'b0 ;
  assign y4623 = ~1'b0 ;
  assign y4624 = n12445 ;
  assign y4625 = n12446 ;
  assign y4626 = ~n12447 ;
  assign y4627 = ~1'b0 ;
  assign y4628 = n12448 ;
  assign y4629 = ~n12452 ;
  assign y4630 = ~n12456 ;
  assign y4631 = ~1'b0 ;
  assign y4632 = ~1'b0 ;
  assign y4633 = n12460 ;
  assign y4634 = ~n12465 ;
  assign y4635 = ~1'b0 ;
  assign y4636 = n12475 ;
  assign y4637 = ~n12480 ;
  assign y4638 = 1'b0 ;
  assign y4639 = ~n12481 ;
  assign y4640 = ~n12483 ;
  assign y4641 = n12486 ;
  assign y4642 = ~1'b0 ;
  assign y4643 = ~n12490 ;
  assign y4644 = ~n12492 ;
  assign y4645 = ~1'b0 ;
  assign y4646 = n12495 ;
  assign y4647 = n12496 ;
  assign y4648 = ~n12497 ;
  assign y4649 = ~n12500 ;
  assign y4650 = n10131 ;
  assign y4651 = ~n12501 ;
  assign y4652 = n12504 ;
  assign y4653 = n12510 ;
  assign y4654 = ~1'b0 ;
  assign y4655 = n4045 ;
  assign y4656 = ~n12511 ;
  assign y4657 = ~n12515 ;
  assign y4658 = n12522 ;
  assign y4659 = ~n12524 ;
  assign y4660 = ~n12525 ;
  assign y4661 = ~1'b0 ;
  assign y4662 = ~n12527 ;
  assign y4663 = ~n12528 ;
  assign y4664 = ~1'b0 ;
  assign y4665 = ~1'b0 ;
  assign y4666 = n12530 ;
  assign y4667 = ~n12531 ;
  assign y4668 = n12532 ;
  assign y4669 = n12536 ;
  assign y4670 = ~n12539 ;
  assign y4671 = ~n12545 ;
  assign y4672 = ~1'b0 ;
  assign y4673 = ~1'b0 ;
  assign y4674 = ~n8716 ;
  assign y4675 = ~n12549 ;
  assign y4676 = ~n12558 ;
  assign y4677 = n12564 ;
  assign y4678 = ~n12566 ;
  assign y4679 = ~n4601 ;
  assign y4680 = n12569 ;
  assign y4681 = ~1'b0 ;
  assign y4682 = ~1'b0 ;
  assign y4683 = n12570 ;
  assign y4684 = ~n12572 ;
  assign y4685 = ~n12574 ;
  assign y4686 = n12577 ;
  assign y4687 = n12580 ;
  assign y4688 = n12583 ;
  assign y4689 = ~n12585 ;
  assign y4690 = n12587 ;
  assign y4691 = n12597 ;
  assign y4692 = n12599 ;
  assign y4693 = ~1'b0 ;
  assign y4694 = n12600 ;
  assign y4695 = n12602 ;
  assign y4696 = n12605 ;
  assign y4697 = ~n12607 ;
  assign y4698 = ~1'b0 ;
  assign y4699 = n12612 ;
  assign y4700 = ~1'b0 ;
  assign y4701 = ~1'b0 ;
  assign y4702 = n12615 ;
  assign y4703 = ~n12616 ;
  assign y4704 = n12617 ;
  assign y4705 = ~n12624 ;
  assign y4706 = n12631 ;
  assign y4707 = ~1'b0 ;
  assign y4708 = n1127 ;
  assign y4709 = n12634 ;
  assign y4710 = ~1'b0 ;
  assign y4711 = ~1'b0 ;
  assign y4712 = n12639 ;
  assign y4713 = n12640 ;
  assign y4714 = ~n12643 ;
  assign y4715 = n12648 ;
  assign y4716 = ~n12652 ;
  assign y4717 = n12654 ;
  assign y4718 = n12656 ;
  assign y4719 = ~n12659 ;
  assign y4720 = n12660 ;
  assign y4721 = ~n12669 ;
  assign y4722 = n12670 ;
  assign y4723 = ~n12675 ;
  assign y4724 = ~1'b0 ;
  assign y4725 = ~1'b0 ;
  assign y4726 = ~n12679 ;
  assign y4727 = ~n12685 ;
  assign y4728 = n12690 ;
  assign y4729 = n12691 ;
  assign y4730 = n12694 ;
  assign y4731 = ~1'b0 ;
  assign y4732 = ~n12695 ;
  assign y4733 = ~n12697 ;
  assign y4734 = n12705 ;
  assign y4735 = ~n12706 ;
  assign y4736 = ~x100 ;
  assign y4737 = n12708 ;
  assign y4738 = n12709 ;
  assign y4739 = n12710 ;
  assign y4740 = ~n12715 ;
  assign y4741 = ~1'b0 ;
  assign y4742 = n12723 ;
  assign y4743 = n4929 ;
  assign y4744 = ~n12728 ;
  assign y4745 = n12731 ;
  assign y4746 = ~n12733 ;
  assign y4747 = n12735 ;
  assign y4748 = n12739 ;
  assign y4749 = n12740 ;
  assign y4750 = n12746 ;
  assign y4751 = ~1'b0 ;
  assign y4752 = ~n12749 ;
  assign y4753 = ~1'b0 ;
  assign y4754 = n12752 ;
  assign y4755 = ~n12762 ;
  assign y4756 = ~n12764 ;
  assign y4757 = n12766 ;
  assign y4758 = ~n12769 ;
  assign y4759 = n12775 ;
  assign y4760 = ~n12777 ;
  assign y4761 = ~1'b0 ;
  assign y4762 = ~n12780 ;
  assign y4763 = n12783 ;
  assign y4764 = ~1'b0 ;
  assign y4765 = ~n12784 ;
  assign y4766 = ~n4432 ;
  assign y4767 = ~1'b0 ;
  assign y4768 = n12787 ;
  assign y4769 = n12792 ;
  assign y4770 = ~n12793 ;
  assign y4771 = ~1'b0 ;
  assign y4772 = ~n12795 ;
  assign y4773 = ~n12799 ;
  assign y4774 = ~n8138 ;
  assign y4775 = ~1'b0 ;
  assign y4776 = ~n12802 ;
  assign y4777 = ~n12811 ;
  assign y4778 = n12817 ;
  assign y4779 = ~n12820 ;
  assign y4780 = ~n12823 ;
  assign y4781 = ~n12825 ;
  assign y4782 = n153 ;
  assign y4783 = ~1'b0 ;
  assign y4784 = ~1'b0 ;
  assign y4785 = n12828 ;
  assign y4786 = ~n12833 ;
  assign y4787 = ~n12837 ;
  assign y4788 = n12840 ;
  assign y4789 = ~n12841 ;
  assign y4790 = ~n12843 ;
  assign y4791 = ~1'b0 ;
  assign y4792 = ~1'b0 ;
  assign y4793 = n12845 ;
  assign y4794 = ~n12849 ;
  assign y4795 = ~n12853 ;
  assign y4796 = n12859 ;
  assign y4797 = ~1'b0 ;
  assign y4798 = n12860 ;
  assign y4799 = ~n12864 ;
  assign y4800 = n12879 ;
  assign y4801 = ~1'b0 ;
  assign y4802 = ~n12884 ;
  assign y4803 = n12886 ;
  assign y4804 = ~n12889 ;
  assign y4805 = n12895 ;
  assign y4806 = ~1'b0 ;
  assign y4807 = ~n3887 ;
  assign y4808 = n12899 ;
  assign y4809 = ~n12910 ;
  assign y4810 = n12913 ;
  assign y4811 = ~n12919 ;
  assign y4812 = ~1'b0 ;
  assign y4813 = n12921 ;
  assign y4814 = ~1'b0 ;
  assign y4815 = n12926 ;
  assign y4816 = ~n12927 ;
  assign y4817 = n12928 ;
  assign y4818 = ~1'b0 ;
  assign y4819 = n12930 ;
  assign y4820 = ~n12934 ;
  assign y4821 = ~n11616 ;
  assign y4822 = n12935 ;
  assign y4823 = ~1'b0 ;
  assign y4824 = ~1'b0 ;
  assign y4825 = ~1'b0 ;
  assign y4826 = ~n12936 ;
  assign y4827 = n12940 ;
  assign y4828 = ~n12941 ;
  assign y4829 = ~n12949 ;
  assign y4830 = n12951 ;
  assign y4831 = ~1'b0 ;
  assign y4832 = ~n12952 ;
  assign y4833 = n12955 ;
  assign y4834 = ~n12957 ;
  assign y4835 = ~n12960 ;
  assign y4836 = ~n12962 ;
  assign y4837 = ~n12966 ;
  assign y4838 = ~1'b0 ;
  assign y4839 = ~1'b0 ;
  assign y4840 = ~n12973 ;
  assign y4841 = ~n12976 ;
  assign y4842 = n12978 ;
  assign y4843 = ~n12979 ;
  assign y4844 = ~1'b0 ;
  assign y4845 = ~n2772 ;
  assign y4846 = n12983 ;
  assign y4847 = ~n12984 ;
  assign y4848 = ~n12986 ;
  assign y4849 = n12987 ;
  assign y4850 = ~n12989 ;
  assign y4851 = ~1'b0 ;
  assign y4852 = ~1'b0 ;
  assign y4853 = ~1'b0 ;
  assign y4854 = n12994 ;
  assign y4855 = ~n12995 ;
  assign y4856 = ~1'b0 ;
  assign y4857 = ~n12997 ;
  assign y4858 = n13001 ;
  assign y4859 = n13005 ;
  assign y4860 = ~n13010 ;
  assign y4861 = n13012 ;
  assign y4862 = n13016 ;
  assign y4863 = n13017 ;
  assign y4864 = ~1'b0 ;
  assign y4865 = ~n13018 ;
  assign y4866 = ~n13021 ;
  assign y4867 = ~n13023 ;
  assign y4868 = n13026 ;
  assign y4869 = n13028 ;
  assign y4870 = ~n13031 ;
  assign y4871 = ~1'b0 ;
  assign y4872 = 1'b0 ;
  assign y4873 = ~n13036 ;
  assign y4874 = n13038 ;
  assign y4875 = n13043 ;
  assign y4876 = n13044 ;
  assign y4877 = ~n13048 ;
  assign y4878 = ~n13051 ;
  assign y4879 = n13056 ;
  assign y4880 = ~n13057 ;
  assign y4881 = ~n13062 ;
  assign y4882 = ~n13063 ;
  assign y4883 = ~n13064 ;
  assign y4884 = n13067 ;
  assign y4885 = ~n13068 ;
  assign y4886 = n13070 ;
  assign y4887 = ~n13071 ;
  assign y4888 = ~n13076 ;
  assign y4889 = n13079 ;
  assign y4890 = ~n13083 ;
  assign y4891 = ~n778 ;
  assign y4892 = n13084 ;
  assign y4893 = ~n5821 ;
  assign y4894 = n13087 ;
  assign y4895 = ~n13089 ;
  assign y4896 = ~n13091 ;
  assign y4897 = ~n13092 ;
  assign y4898 = ~n13094 ;
  assign y4899 = n13095 ;
  assign y4900 = ~n13100 ;
  assign y4901 = n13104 ;
  assign y4902 = ~n13109 ;
  assign y4903 = n13116 ;
  assign y4904 = ~1'b0 ;
  assign y4905 = n13125 ;
  assign y4906 = ~1'b0 ;
  assign y4907 = n13131 ;
  assign y4908 = ~1'b0 ;
  assign y4909 = ~n13135 ;
  assign y4910 = ~n13139 ;
  assign y4911 = n13144 ;
  assign y4912 = ~1'b0 ;
  assign y4913 = n13150 ;
  assign y4914 = n13151 ;
  assign y4915 = ~n13154 ;
  assign y4916 = n13155 ;
  assign y4917 = ~1'b0 ;
  assign y4918 = n13157 ;
  assign y4919 = ~1'b0 ;
  assign y4920 = ~n13159 ;
  assign y4921 = ~n13164 ;
  assign y4922 = ~n13166 ;
  assign y4923 = ~n13169 ;
  assign y4924 = n13171 ;
  assign y4925 = ~n13175 ;
  assign y4926 = ~n13176 ;
  assign y4927 = n13182 ;
  assign y4928 = n13184 ;
  assign y4929 = ~n13189 ;
  assign y4930 = ~n13191 ;
  assign y4931 = ~1'b0 ;
  assign y4932 = ~n13192 ;
  assign y4933 = ~n13193 ;
  assign y4934 = ~n13196 ;
  assign y4935 = n13200 ;
  assign y4936 = ~1'b0 ;
  assign y4937 = ~n13204 ;
  assign y4938 = n13206 ;
  assign y4939 = ~n13208 ;
  assign y4940 = ~1'b0 ;
  assign y4941 = ~n13211 ;
  assign y4942 = n13217 ;
  assign y4943 = ~n13222 ;
  assign y4944 = ~1'b0 ;
  assign y4945 = ~n13228 ;
  assign y4946 = n13231 ;
  assign y4947 = n13232 ;
  assign y4948 = ~1'b0 ;
  assign y4949 = ~n13239 ;
  assign y4950 = ~n13240 ;
  assign y4951 = ~n13241 ;
  assign y4952 = ~n13242 ;
  assign y4953 = ~n3941 ;
  assign y4954 = ~1'b0 ;
  assign y4955 = n13251 ;
  assign y4956 = n13252 ;
  assign y4957 = n13253 ;
  assign y4958 = n13255 ;
  assign y4959 = n13260 ;
  assign y4960 = ~n13262 ;
  assign y4961 = n13267 ;
  assign y4962 = n13269 ;
  assign y4963 = ~1'b0 ;
  assign y4964 = n13274 ;
  assign y4965 = ~n13279 ;
  assign y4966 = n13283 ;
  assign y4967 = n13287 ;
  assign y4968 = n13292 ;
  assign y4969 = ~n13293 ;
  assign y4970 = n13297 ;
  assign y4971 = n13298 ;
  assign y4972 = ~n13299 ;
  assign y4973 = n13300 ;
  assign y4974 = ~n13303 ;
  assign y4975 = n13304 ;
  assign y4976 = n8550 ;
  assign y4977 = n13312 ;
  assign y4978 = n13315 ;
  assign y4979 = ~1'b0 ;
  assign y4980 = n13317 ;
  assign y4981 = ~n13321 ;
  assign y4982 = ~n13324 ;
  assign y4983 = n13326 ;
  assign y4984 = ~n13327 ;
  assign y4985 = ~n13329 ;
  assign y4986 = n13330 ;
  assign y4987 = ~n13342 ;
  assign y4988 = ~n13344 ;
  assign y4989 = n13347 ;
  assign y4990 = ~1'b0 ;
  assign y4991 = ~1'b0 ;
  assign y4992 = ~n13355 ;
  assign y4993 = ~1'b0 ;
  assign y4994 = ~n13358 ;
  assign y4995 = ~n13363 ;
  assign y4996 = ~n13366 ;
  assign y4997 = ~1'b0 ;
  assign y4998 = n13372 ;
  assign y4999 = n13376 ;
  assign y5000 = ~1'b0 ;
  assign y5001 = n13379 ;
  assign y5002 = ~n13382 ;
  assign y5003 = n13383 ;
  assign y5004 = ~n13384 ;
  assign y5005 = ~1'b0 ;
  assign y5006 = ~n13386 ;
  assign y5007 = ~n13392 ;
  assign y5008 = ~1'b0 ;
  assign y5009 = ~n13394 ;
  assign y5010 = ~1'b0 ;
  assign y5011 = ~1'b0 ;
  assign y5012 = ~n13396 ;
  assign y5013 = ~n13397 ;
  assign y5014 = ~n13399 ;
  assign y5015 = n13403 ;
  assign y5016 = ~n13408 ;
  assign y5017 = n13419 ;
  assign y5018 = ~n13420 ;
  assign y5019 = n13421 ;
  assign y5020 = ~n13423 ;
  assign y5021 = ~n13427 ;
  assign y5022 = ~n13429 ;
  assign y5023 = ~n7333 ;
  assign y5024 = ~n13436 ;
  assign y5025 = ~n9259 ;
  assign y5026 = ~1'b0 ;
  assign y5027 = ~n13443 ;
  assign y5028 = ~n13445 ;
  assign y5029 = ~1'b0 ;
  assign y5030 = ~n13448 ;
  assign y5031 = ~n13449 ;
  assign y5032 = n13450 ;
  assign y5033 = n13453 ;
  assign y5034 = n13456 ;
  assign y5035 = ~n13458 ;
  assign y5036 = n13461 ;
  assign y5037 = ~n13463 ;
  assign y5038 = n13466 ;
  assign y5039 = n13468 ;
  assign y5040 = ~1'b0 ;
  assign y5041 = ~1'b0 ;
  assign y5042 = 1'b0 ;
  assign y5043 = ~1'b0 ;
  assign y5044 = ~n13479 ;
  assign y5045 = ~n13483 ;
  assign y5046 = n13486 ;
  assign y5047 = ~1'b0 ;
  assign y5048 = ~n13492 ;
  assign y5049 = ~n13495 ;
  assign y5050 = n13501 ;
  assign y5051 = ~n13507 ;
  assign y5052 = n13512 ;
  assign y5053 = ~n13523 ;
  assign y5054 = ~1'b0 ;
  assign y5055 = ~1'b0 ;
  assign y5056 = ~n13527 ;
  assign y5057 = n13530 ;
  assign y5058 = n13534 ;
  assign y5059 = ~n13537 ;
  assign y5060 = n13538 ;
  assign y5061 = n13546 ;
  assign y5062 = n6808 ;
  assign y5063 = ~1'b0 ;
  assign y5064 = n13547 ;
  assign y5065 = n13548 ;
  assign y5066 = ~n13550 ;
  assign y5067 = ~n13555 ;
  assign y5068 = ~1'b0 ;
  assign y5069 = ~n13558 ;
  assign y5070 = ~n13563 ;
  assign y5071 = ~n13570 ;
  assign y5072 = n13574 ;
  assign y5073 = n13578 ;
  assign y5074 = ~n13579 ;
  assign y5075 = n13580 ;
  assign y5076 = n13588 ;
  assign y5077 = ~n13589 ;
  assign y5078 = ~1'b0 ;
  assign y5079 = ~1'b0 ;
  assign y5080 = n13591 ;
  assign y5081 = n13593 ;
  assign y5082 = n13595 ;
  assign y5083 = n13596 ;
  assign y5084 = n4607 ;
  assign y5085 = n13198 ;
  assign y5086 = n13597 ;
  assign y5087 = ~n13598 ;
  assign y5088 = n13599 ;
  assign y5089 = ~n13602 ;
  assign y5090 = ~1'b0 ;
  assign y5091 = ~n13603 ;
  assign y5092 = ~n13608 ;
  assign y5093 = ~n13610 ;
  assign y5094 = ~n13613 ;
  assign y5095 = n13617 ;
  assign y5096 = n13622 ;
  assign y5097 = ~n13624 ;
  assign y5098 = n13629 ;
  assign y5099 = ~n13634 ;
  assign y5100 = n13635 ;
  assign y5101 = n13636 ;
  assign y5102 = ~n13637 ;
  assign y5103 = ~1'b0 ;
  assign y5104 = ~1'b0 ;
  assign y5105 = ~n13640 ;
  assign y5106 = n13644 ;
  assign y5107 = n13646 ;
  assign y5108 = ~1'b0 ;
  assign y5109 = ~1'b0 ;
  assign y5110 = n13647 ;
  assign y5111 = n13649 ;
  assign y5112 = ~n13655 ;
  assign y5113 = n13661 ;
  assign y5114 = ~n13668 ;
  assign y5115 = ~1'b0 ;
  assign y5116 = n13673 ;
  assign y5117 = n13675 ;
  assign y5118 = ~n13676 ;
  assign y5119 = ~n13678 ;
  assign y5120 = ~1'b0 ;
  assign y5121 = n11103 ;
  assign y5122 = ~1'b0 ;
  assign y5123 = n13680 ;
  assign y5124 = n13682 ;
  assign y5125 = ~1'b0 ;
  assign y5126 = ~1'b0 ;
  assign y5127 = n13686 ;
  assign y5128 = n13688 ;
  assign y5129 = n9385 ;
  assign y5130 = ~1'b0 ;
  assign y5131 = n13689 ;
  assign y5132 = n13690 ;
  assign y5133 = ~n13695 ;
  assign y5134 = n13698 ;
  assign y5135 = ~n13706 ;
  assign y5136 = ~1'b0 ;
  assign y5137 = ~1'b0 ;
  assign y5138 = ~n13536 ;
  assign y5139 = ~n13708 ;
  assign y5140 = ~n13712 ;
  assign y5141 = ~1'b0 ;
  assign y5142 = ~1'b0 ;
  assign y5143 = n3068 ;
  assign y5144 = ~1'b0 ;
  assign y5145 = n13713 ;
  assign y5146 = ~n13716 ;
  assign y5147 = n13726 ;
  assign y5148 = ~1'b0 ;
  assign y5149 = ~n11487 ;
  assign y5150 = ~n13731 ;
  assign y5151 = ~n13735 ;
  assign y5152 = ~n13737 ;
  assign y5153 = ~n13743 ;
  assign y5154 = n13744 ;
  assign y5155 = ~n13747 ;
  assign y5156 = ~n13752 ;
  assign y5157 = n13753 ;
  assign y5158 = n13760 ;
  assign y5159 = n6433 ;
  assign y5160 = ~n13764 ;
  assign y5161 = ~n13766 ;
  assign y5162 = ~1'b0 ;
  assign y5163 = ~1'b0 ;
  assign y5164 = n13772 ;
  assign y5165 = n10080 ;
  assign y5166 = ~1'b0 ;
  assign y5167 = n13773 ;
  assign y5168 = n13774 ;
  assign y5169 = ~1'b0 ;
  assign y5170 = n13778 ;
  assign y5171 = ~1'b0 ;
  assign y5172 = ~n13779 ;
  assign y5173 = ~n13780 ;
  assign y5174 = ~n13783 ;
  assign y5175 = n13784 ;
  assign y5176 = n13786 ;
  assign y5177 = ~n13789 ;
  assign y5178 = ~n13791 ;
  assign y5179 = ~n13792 ;
  assign y5180 = ~n13797 ;
  assign y5181 = ~n13802 ;
  assign y5182 = ~n13804 ;
  assign y5183 = ~n13806 ;
  assign y5184 = n13809 ;
  assign y5185 = n13810 ;
  assign y5186 = n4448 ;
  assign y5187 = ~1'b0 ;
  assign y5188 = n13812 ;
  assign y5189 = ~n13814 ;
  assign y5190 = ~n13815 ;
  assign y5191 = ~n13816 ;
  assign y5192 = ~n13825 ;
  assign y5193 = ~1'b0 ;
  assign y5194 = n13826 ;
  assign y5195 = ~1'b0 ;
  assign y5196 = ~n13832 ;
  assign y5197 = ~n13833 ;
  assign y5198 = ~n13837 ;
  assign y5199 = ~1'b0 ;
  assign y5200 = ~1'b0 ;
  assign y5201 = ~n13840 ;
  assign y5202 = n13846 ;
  assign y5203 = ~n13849 ;
  assign y5204 = ~1'b0 ;
  assign y5205 = n13855 ;
  assign y5206 = n13861 ;
  assign y5207 = n13864 ;
  assign y5208 = ~n13866 ;
  assign y5209 = ~n13867 ;
  assign y5210 = ~n13874 ;
  assign y5211 = ~n13875 ;
  assign y5212 = n13876 ;
  assign y5213 = ~1'b0 ;
  assign y5214 = ~1'b0 ;
  assign y5215 = ~n13879 ;
  assign y5216 = ~1'b0 ;
  assign y5217 = ~n13887 ;
  assign y5218 = ~n13890 ;
  assign y5219 = ~n13899 ;
  assign y5220 = ~1'b0 ;
  assign y5221 = ~1'b0 ;
  assign y5222 = ~1'b0 ;
  assign y5223 = n13900 ;
  assign y5224 = n13906 ;
  assign y5225 = ~n3753 ;
  assign y5226 = ~1'b0 ;
  assign y5227 = ~n13907 ;
  assign y5228 = ~n13913 ;
  assign y5229 = n13915 ;
  assign y5230 = ~n13918 ;
  assign y5231 = ~1'b0 ;
  assign y5232 = n13919 ;
  assign y5233 = ~1'b0 ;
  assign y5234 = ~n13920 ;
  assign y5235 = n13921 ;
  assign y5236 = ~n13923 ;
  assign y5237 = ~1'b0 ;
  assign y5238 = ~n13925 ;
  assign y5239 = ~n13927 ;
  assign y5240 = n13928 ;
  assign y5241 = n13929 ;
  assign y5242 = n13930 ;
  assign y5243 = n13931 ;
  assign y5244 = n13934 ;
  assign y5245 = ~1'b0 ;
  assign y5246 = n13936 ;
  assign y5247 = 1'b0 ;
  assign y5248 = ~1'b0 ;
  assign y5249 = n13937 ;
  assign y5250 = ~n7784 ;
  assign y5251 = n13939 ;
  assign y5252 = n13941 ;
  assign y5253 = ~1'b0 ;
  assign y5254 = ~n13942 ;
  assign y5255 = ~n13948 ;
  assign y5256 = ~n13955 ;
  assign y5257 = n13956 ;
  assign y5258 = ~n13959 ;
  assign y5259 = n13968 ;
  assign y5260 = ~n13976 ;
  assign y5261 = ~n13978 ;
  assign y5262 = ~n13979 ;
  assign y5263 = ~n13980 ;
  assign y5264 = ~n13981 ;
  assign y5265 = ~n13983 ;
  assign y5266 = n13988 ;
  assign y5267 = n13990 ;
  assign y5268 = ~1'b0 ;
  assign y5269 = ~1'b0 ;
  assign y5270 = n13991 ;
  assign y5271 = n13993 ;
  assign y5272 = ~n13995 ;
  assign y5273 = ~n14000 ;
  assign y5274 = ~n14003 ;
  assign y5275 = ~1'b0 ;
  assign y5276 = ~n14004 ;
  assign y5277 = ~1'b0 ;
  assign y5278 = ~n14006 ;
  assign y5279 = n14008 ;
  assign y5280 = ~1'b0 ;
  assign y5281 = n14009 ;
  assign y5282 = ~1'b0 ;
  assign y5283 = n14013 ;
  assign y5284 = ~1'b0 ;
  assign y5285 = ~n14022 ;
  assign y5286 = ~1'b0 ;
  assign y5287 = ~n14024 ;
  assign y5288 = ~n14025 ;
  assign y5289 = ~n14027 ;
  assign y5290 = n14030 ;
  assign y5291 = ~n14031 ;
  assign y5292 = n14033 ;
  assign y5293 = ~n14035 ;
  assign y5294 = ~1'b0 ;
  assign y5295 = ~1'b0 ;
  assign y5296 = n14036 ;
  assign y5297 = n14038 ;
  assign y5298 = ~1'b0 ;
  assign y5299 = ~1'b0 ;
  assign y5300 = ~1'b0 ;
  assign y5301 = ~1'b0 ;
  assign y5302 = ~n14051 ;
  assign y5303 = n14052 ;
  assign y5304 = ~1'b0 ;
  assign y5305 = n14055 ;
  assign y5306 = n14057 ;
  assign y5307 = ~1'b0 ;
  assign y5308 = ~n14061 ;
  assign y5309 = n14066 ;
  assign y5310 = ~n14075 ;
  assign y5311 = ~n14076 ;
  assign y5312 = ~n14080 ;
  assign y5313 = ~n14081 ;
  assign y5314 = n14084 ;
  assign y5315 = ~n14089 ;
  assign y5316 = n14090 ;
  assign y5317 = n14094 ;
  assign y5318 = ~n14096 ;
  assign y5319 = ~n14098 ;
  assign y5320 = ~n14099 ;
  assign y5321 = ~n14100 ;
  assign y5322 = ~1'b0 ;
  assign y5323 = n2580 ;
  assign y5324 = ~1'b0 ;
  assign y5325 = ~n14103 ;
  assign y5326 = ~n14104 ;
  assign y5327 = ~n14105 ;
  assign y5328 = n14110 ;
  assign y5329 = ~1'b0 ;
  assign y5330 = n14112 ;
  assign y5331 = ~n14116 ;
  assign y5332 = n14117 ;
  assign y5333 = ~n14125 ;
  assign y5334 = n14126 ;
  assign y5335 = ~n14132 ;
  assign y5336 = ~n14133 ;
  assign y5337 = n14138 ;
  assign y5338 = n14139 ;
  assign y5339 = n14140 ;
  assign y5340 = ~n14142 ;
  assign y5341 = ~n14143 ;
  assign y5342 = n14147 ;
  assign y5343 = ~1'b0 ;
  assign y5344 = ~n14151 ;
  assign y5345 = n14152 ;
  assign y5346 = n14153 ;
  assign y5347 = ~n14155 ;
  assign y5348 = ~n14156 ;
  assign y5349 = n14159 ;
  assign y5350 = n14161 ;
  assign y5351 = ~n14162 ;
  assign y5352 = n14165 ;
  assign y5353 = n10155 ;
  assign y5354 = n14171 ;
  assign y5355 = ~n14173 ;
  assign y5356 = n14180 ;
  assign y5357 = ~n14182 ;
  assign y5358 = n14183 ;
  assign y5359 = n14185 ;
  assign y5360 = n14186 ;
  assign y5361 = n14187 ;
  assign y5362 = n14188 ;
  assign y5363 = ~1'b0 ;
  assign y5364 = n318 ;
  assign y5365 = ~1'b0 ;
  assign y5366 = ~1'b0 ;
  assign y5367 = n14191 ;
  assign y5368 = n14192 ;
  assign y5369 = ~1'b0 ;
  assign y5370 = ~1'b0 ;
  assign y5371 = n14193 ;
  assign y5372 = n14194 ;
  assign y5373 = n14199 ;
  assign y5374 = n14206 ;
  assign y5375 = ~1'b0 ;
  assign y5376 = ~n14213 ;
  assign y5377 = ~n14216 ;
  assign y5378 = ~n14217 ;
  assign y5379 = n14219 ;
  assign y5380 = ~n14223 ;
  assign y5381 = ~1'b0 ;
  assign y5382 = ~n14226 ;
  assign y5383 = ~n14228 ;
  assign y5384 = n14236 ;
  assign y5385 = ~n14237 ;
  assign y5386 = ~1'b0 ;
  assign y5387 = ~n14241 ;
  assign y5388 = ~n14243 ;
  assign y5389 = n14253 ;
  assign y5390 = ~1'b0 ;
  assign y5391 = ~n14259 ;
  assign y5392 = ~n14262 ;
  assign y5393 = n14265 ;
  assign y5394 = n14271 ;
  assign y5395 = n14272 ;
  assign y5396 = ~n14274 ;
  assign y5397 = ~n14276 ;
  assign y5398 = ~n14278 ;
  assign y5399 = ~n14283 ;
  assign y5400 = ~n14284 ;
  assign y5401 = ~n14285 ;
  assign y5402 = ~n14292 ;
  assign y5403 = ~1'b0 ;
  assign y5404 = ~n14298 ;
  assign y5405 = n14299 ;
  assign y5406 = ~n14300 ;
  assign y5407 = ~n14303 ;
  assign y5408 = n14310 ;
  assign y5409 = ~n14317 ;
  assign y5410 = ~1'b0 ;
  assign y5411 = n14325 ;
  assign y5412 = n14327 ;
  assign y5413 = ~n14328 ;
  assign y5414 = ~1'b0 ;
  assign y5415 = ~n14331 ;
  assign y5416 = n14333 ;
  assign y5417 = n14335 ;
  assign y5418 = n14337 ;
  assign y5419 = n14339 ;
  assign y5420 = ~n2193 ;
  assign y5421 = ~n14344 ;
  assign y5422 = ~n14345 ;
  assign y5423 = 1'b0 ;
  assign y5424 = ~n14346 ;
  assign y5425 = ~n14348 ;
  assign y5426 = ~n14349 ;
  assign y5427 = ~1'b0 ;
  assign y5428 = ~1'b0 ;
  assign y5429 = n14351 ;
  assign y5430 = ~n14352 ;
  assign y5431 = ~n14354 ;
  assign y5432 = ~n14356 ;
  assign y5433 = ~n14358 ;
  assign y5434 = ~n14359 ;
  assign y5435 = ~n14361 ;
  assign y5436 = ~n14366 ;
  assign y5437 = ~n14369 ;
  assign y5438 = ~n14372 ;
  assign y5439 = n14374 ;
  assign y5440 = ~1'b0 ;
  assign y5441 = ~1'b0 ;
  assign y5442 = ~1'b0 ;
  assign y5443 = n14375 ;
  assign y5444 = n7966 ;
  assign y5445 = n14377 ;
  assign y5446 = ~1'b0 ;
  assign y5447 = ~1'b0 ;
  assign y5448 = n14382 ;
  assign y5449 = ~n14391 ;
  assign y5450 = ~n14395 ;
  assign y5451 = ~1'b0 ;
  assign y5452 = ~n14396 ;
  assign y5453 = n14397 ;
  assign y5454 = ~1'b0 ;
  assign y5455 = n14398 ;
  assign y5456 = ~n14399 ;
  assign y5457 = n14400 ;
  assign y5458 = n14404 ;
  assign y5459 = n14406 ;
  assign y5460 = n14409 ;
  assign y5461 = n14410 ;
  assign y5462 = ~n14412 ;
  assign y5463 = 1'b0 ;
  assign y5464 = n14414 ;
  assign y5465 = ~n14420 ;
  assign y5466 = ~1'b0 ;
  assign y5467 = n14425 ;
  assign y5468 = n14426 ;
  assign y5469 = ~n14431 ;
  assign y5470 = ~1'b0 ;
  assign y5471 = ~n14432 ;
  assign y5472 = ~n14433 ;
  assign y5473 = ~1'b0 ;
  assign y5474 = n14437 ;
  assign y5475 = ~n14441 ;
  assign y5476 = ~n14445 ;
  assign y5477 = n14450 ;
  assign y5478 = ~n14455 ;
  assign y5479 = n14457 ;
  assign y5480 = ~n14463 ;
  assign y5481 = n14467 ;
  assign y5482 = ~1'b0 ;
  assign y5483 = ~1'b0 ;
  assign y5484 = ~n14470 ;
  assign y5485 = ~1'b0 ;
  assign y5486 = ~n14473 ;
  assign y5487 = ~n14477 ;
  assign y5488 = n14481 ;
  assign y5489 = ~n14483 ;
  assign y5490 = ~n14487 ;
  assign y5491 = ~n14488 ;
  assign y5492 = n14489 ;
  assign y5493 = ~n14492 ;
  assign y5494 = n14497 ;
  assign y5495 = ~n14498 ;
  assign y5496 = n14504 ;
  assign y5497 = ~1'b0 ;
  assign y5498 = ~1'b0 ;
  assign y5499 = n14509 ;
  assign y5500 = n14512 ;
  assign y5501 = ~n14516 ;
  assign y5502 = ~1'b0 ;
  assign y5503 = ~n14518 ;
  assign y5504 = ~n14528 ;
  assign y5505 = ~n14529 ;
  assign y5506 = ~n14535 ;
  assign y5507 = ~n14540 ;
  assign y5508 = ~1'b0 ;
  assign y5509 = ~1'b0 ;
  assign y5510 = n14542 ;
  assign y5511 = n14549 ;
  assign y5512 = n14559 ;
  assign y5513 = n14562 ;
  assign y5514 = n14563 ;
  assign y5515 = ~n14564 ;
  assign y5516 = n13052 ;
  assign y5517 = n14566 ;
  assign y5518 = n14569 ;
  assign y5519 = ~n14576 ;
  assign y5520 = ~1'b0 ;
  assign y5521 = ~1'b0 ;
  assign y5522 = ~1'b0 ;
  assign y5523 = ~n14581 ;
  assign y5524 = n14589 ;
  assign y5525 = n14597 ;
  assign y5526 = ~1'b0 ;
  assign y5527 = n14603 ;
  assign y5528 = ~n14606 ;
  assign y5529 = ~n10683 ;
  assign y5530 = n14608 ;
  assign y5531 = ~n14611 ;
  assign y5532 = n14614 ;
  assign y5533 = ~n14619 ;
  assign y5534 = n14623 ;
  assign y5535 = ~n14629 ;
  assign y5536 = ~1'b0 ;
  assign y5537 = ~1'b0 ;
  assign y5538 = ~1'b0 ;
  assign y5539 = n14634 ;
  assign y5540 = n14635 ;
  assign y5541 = n14641 ;
  assign y5542 = n14643 ;
  assign y5543 = ~n14645 ;
  assign y5544 = n14648 ;
  assign y5545 = n14650 ;
  assign y5546 = ~1'b0 ;
  assign y5547 = n14651 ;
  assign y5548 = ~n14652 ;
  assign y5549 = n14654 ;
  assign y5550 = ~1'b0 ;
  assign y5551 = ~n14655 ;
  assign y5552 = ~1'b0 ;
  assign y5553 = ~n14660 ;
  assign y5554 = ~n14662 ;
  assign y5555 = ~1'b0 ;
  assign y5556 = n14663 ;
  assign y5557 = ~1'b0 ;
  assign y5558 = ~n14664 ;
  assign y5559 = ~n14666 ;
  assign y5560 = n6196 ;
  assign y5561 = n14669 ;
  assign y5562 = n14670 ;
  assign y5563 = ~n14673 ;
  assign y5564 = n14674 ;
  assign y5565 = n14677 ;
  assign y5566 = ~1'b0 ;
  assign y5567 = ~n14679 ;
  assign y5568 = n14680 ;
  assign y5569 = n14684 ;
  assign y5570 = ~n14685 ;
  assign y5571 = n14687 ;
  assign y5572 = ~n14688 ;
  assign y5573 = n14690 ;
  assign y5574 = ~n14695 ;
  assign y5575 = n14700 ;
  assign y5576 = ~1'b0 ;
  assign y5577 = n14708 ;
  assign y5578 = n14712 ;
  assign y5579 = ~n14714 ;
  assign y5580 = ~1'b0 ;
  assign y5581 = n14716 ;
  assign y5582 = n14718 ;
  assign y5583 = n14719 ;
  assign y5584 = ~n14721 ;
  assign y5585 = ~1'b0 ;
  assign y5586 = ~1'b0 ;
  assign y5587 = ~n14726 ;
  assign y5588 = ~1'b0 ;
  assign y5589 = ~n14727 ;
  assign y5590 = ~1'b0 ;
  assign y5591 = ~n14729 ;
  assign y5592 = ~n14730 ;
  assign y5593 = ~1'b0 ;
  assign y5594 = ~n14734 ;
  assign y5595 = n14739 ;
  assign y5596 = ~n14743 ;
  assign y5597 = ~n14747 ;
  assign y5598 = n14750 ;
  assign y5599 = ~n14752 ;
  assign y5600 = ~n14756 ;
  assign y5601 = n14761 ;
  assign y5602 = ~1'b0 ;
  assign y5603 = ~n14765 ;
  assign y5604 = ~n14767 ;
  assign y5605 = ~1'b0 ;
  assign y5606 = ~n14772 ;
  assign y5607 = n14774 ;
  assign y5608 = n3403 ;
  assign y5609 = n14776 ;
  assign y5610 = n14785 ;
  assign y5611 = n14790 ;
  assign y5612 = ~n14791 ;
  assign y5613 = n14799 ;
  assign y5614 = n14800 ;
  assign y5615 = n14803 ;
  assign y5616 = ~n14807 ;
  assign y5617 = n14811 ;
  assign y5618 = n14816 ;
  assign y5619 = ~n14817 ;
  assign y5620 = ~1'b0 ;
  assign y5621 = n14821 ;
  assign y5622 = ~n14824 ;
  assign y5623 = ~n14829 ;
  assign y5624 = n14830 ;
  assign y5625 = ~n14832 ;
  assign y5626 = n14834 ;
  assign y5627 = n14837 ;
  assign y5628 = ~n14849 ;
  assign y5629 = n14850 ;
  assign y5630 = ~n14854 ;
  assign y5631 = ~n1123 ;
  assign y5632 = n14857 ;
  assign y5633 = n14859 ;
  assign y5634 = ~n14860 ;
  assign y5635 = ~n14864 ;
  assign y5636 = ~n14868 ;
  assign y5637 = ~n14869 ;
  assign y5638 = n14870 ;
  assign y5639 = ~n14874 ;
  assign y5640 = n14880 ;
  assign y5641 = ~1'b0 ;
  assign y5642 = ~1'b0 ;
  assign y5643 = n14882 ;
  assign y5644 = n14883 ;
  assign y5645 = n14885 ;
  assign y5646 = ~1'b0 ;
  assign y5647 = n14887 ;
  assign y5648 = ~n14889 ;
  assign y5649 = ~n14895 ;
  assign y5650 = n14898 ;
  assign y5651 = ~n14904 ;
  assign y5652 = ~n14906 ;
  assign y5653 = ~n14909 ;
  assign y5654 = ~n14910 ;
  assign y5655 = ~n14912 ;
  assign y5656 = n14913 ;
  assign y5657 = ~n14914 ;
  assign y5658 = ~1'b0 ;
  assign y5659 = n14919 ;
  assign y5660 = n14924 ;
  assign y5661 = ~1'b0 ;
  assign y5662 = ~1'b0 ;
  assign y5663 = n14928 ;
  assign y5664 = n14932 ;
  assign y5665 = ~n14936 ;
  assign y5666 = 1'b0 ;
  assign y5667 = ~n14937 ;
  assign y5668 = n14940 ;
  assign y5669 = n7771 ;
  assign y5670 = n14943 ;
  assign y5671 = ~n14947 ;
  assign y5672 = n14949 ;
  assign y5673 = ~n14951 ;
  assign y5674 = ~n14952 ;
  assign y5675 = ~1'b0 ;
  assign y5676 = ~n14953 ;
  assign y5677 = ~1'b0 ;
  assign y5678 = n14960 ;
  assign y5679 = n14963 ;
  assign y5680 = ~n14964 ;
  assign y5681 = ~n14965 ;
  assign y5682 = ~n14970 ;
  assign y5683 = n14973 ;
  assign y5684 = ~n14975 ;
  assign y5685 = n14980 ;
  assign y5686 = ~1'b0 ;
  assign y5687 = ~1'b0 ;
  assign y5688 = n14983 ;
  assign y5689 = ~n14987 ;
  assign y5690 = ~n14991 ;
  assign y5691 = ~n14992 ;
  assign y5692 = n14993 ;
  assign y5693 = ~n15002 ;
  assign y5694 = n15010 ;
  assign y5695 = ~1'b0 ;
  assign y5696 = ~n15011 ;
  assign y5697 = n15013 ;
  assign y5698 = ~n15014 ;
  assign y5699 = n15015 ;
  assign y5700 = ~n15020 ;
  assign y5701 = n15021 ;
  assign y5702 = ~n15024 ;
  assign y5703 = n15030 ;
  assign y5704 = n15038 ;
  assign y5705 = ~n15042 ;
  assign y5706 = ~n4287 ;
  assign y5707 = ~n15043 ;
  assign y5708 = n15045 ;
  assign y5709 = ~n15046 ;
  assign y5710 = ~n15052 ;
  assign y5711 = n15054 ;
  assign y5712 = n15056 ;
  assign y5713 = n15058 ;
  assign y5714 = ~n15063 ;
  assign y5715 = ~1'b0 ;
  assign y5716 = n15064 ;
  assign y5717 = n15065 ;
  assign y5718 = n15067 ;
  assign y5719 = n15078 ;
  assign y5720 = n15079 ;
  assign y5721 = ~n15080 ;
  assign y5722 = ~n10641 ;
  assign y5723 = ~1'b0 ;
  assign y5724 = ~n15085 ;
  assign y5725 = ~n15091 ;
  assign y5726 = ~1'b0 ;
  assign y5727 = n15099 ;
  assign y5728 = ~n15100 ;
  assign y5729 = ~1'b0 ;
  assign y5730 = ~1'b0 ;
  assign y5731 = n15102 ;
  assign y5732 = ~n15104 ;
  assign y5733 = n15109 ;
  assign y5734 = n15111 ;
  assign y5735 = ~n15112 ;
  assign y5736 = ~n15114 ;
  assign y5737 = ~n15118 ;
  assign y5738 = n15120 ;
  assign y5739 = ~n15126 ;
  assign y5740 = ~1'b0 ;
  assign y5741 = ~n15128 ;
  assign y5742 = ~n15132 ;
  assign y5743 = ~n15139 ;
  assign y5744 = n15145 ;
  assign y5745 = ~n15147 ;
  assign y5746 = ~n15152 ;
  assign y5747 = n15161 ;
  assign y5748 = ~1'b0 ;
  assign y5749 = ~n15166 ;
  assign y5750 = ~n15169 ;
  assign y5751 = ~1'b0 ;
  assign y5752 = ~1'b0 ;
  assign y5753 = ~n15170 ;
  assign y5754 = n15173 ;
  assign y5755 = n15177 ;
  assign y5756 = ~1'b0 ;
  assign y5757 = ~n15178 ;
  assign y5758 = ~n15181 ;
  assign y5759 = ~n15183 ;
  assign y5760 = ~n15184 ;
  assign y5761 = ~n15185 ;
  assign y5762 = ~1'b0 ;
  assign y5763 = n15186 ;
  assign y5764 = ~n15200 ;
  assign y5765 = ~n3862 ;
  assign y5766 = ~n15201 ;
  assign y5767 = ~n15202 ;
  assign y5768 = ~n15206 ;
  assign y5769 = ~1'b0 ;
  assign y5770 = ~n15209 ;
  assign y5771 = 1'b0 ;
  assign y5772 = ~n15211 ;
  assign y5773 = n15214 ;
  assign y5774 = n15215 ;
  assign y5775 = n15218 ;
  assign y5776 = n15220 ;
  assign y5777 = n15227 ;
  assign y5778 = ~n15237 ;
  assign y5779 = n15244 ;
  assign y5780 = ~1'b0 ;
  assign y5781 = ~1'b0 ;
  assign y5782 = n15246 ;
  assign y5783 = ~1'b0 ;
  assign y5784 = ~n15248 ;
  assign y5785 = ~n15249 ;
  assign y5786 = ~1'b0 ;
  assign y5787 = ~1'b0 ;
  assign y5788 = ~n15251 ;
  assign y5789 = ~n15252 ;
  assign y5790 = n15253 ;
  assign y5791 = n15255 ;
  assign y5792 = n15256 ;
  assign y5793 = n15257 ;
  assign y5794 = ~n15258 ;
  assign y5795 = n15259 ;
  assign y5796 = ~n15260 ;
  assign y5797 = ~n15265 ;
  assign y5798 = ~n15268 ;
  assign y5799 = ~n15272 ;
  assign y5800 = n15275 ;
  assign y5801 = ~n15278 ;
  assign y5802 = ~1'b0 ;
  assign y5803 = ~1'b0 ;
  assign y5804 = ~n15280 ;
  assign y5805 = ~n15294 ;
  assign y5806 = ~n15295 ;
  assign y5807 = ~1'b0 ;
  assign y5808 = n15301 ;
  assign y5809 = ~n15304 ;
  assign y5810 = ~1'b0 ;
  assign y5811 = ~1'b0 ;
  assign y5812 = ~1'b0 ;
  assign y5813 = ~1'b0 ;
  assign y5814 = n15305 ;
  assign y5815 = n15307 ;
  assign y5816 = ~n15308 ;
  assign y5817 = ~1'b0 ;
  assign y5818 = ~n15309 ;
  assign y5819 = ~n15315 ;
  assign y5820 = n15316 ;
  assign y5821 = n15317 ;
  assign y5822 = ~1'b0 ;
  assign y5823 = n15325 ;
  assign y5824 = ~1'b0 ;
  assign y5825 = n15330 ;
  assign y5826 = n15331 ;
  assign y5827 = ~1'b0 ;
  assign y5828 = ~n15333 ;
  assign y5829 = n15335 ;
  assign y5830 = ~1'b0 ;
  assign y5831 = n15338 ;
  assign y5832 = n15348 ;
  assign y5833 = ~n15352 ;
  assign y5834 = ~n15354 ;
  assign y5835 = ~n15355 ;
  assign y5836 = n15357 ;
  assign y5837 = n15362 ;
  assign y5838 = n7803 ;
  assign y5839 = ~1'b0 ;
  assign y5840 = 1'b0 ;
  assign y5841 = n4917 ;
  assign y5842 = ~n15366 ;
  assign y5843 = ~1'b0 ;
  assign y5844 = n15367 ;
  assign y5845 = ~1'b0 ;
  assign y5846 = ~n15368 ;
  assign y5847 = ~n15369 ;
  assign y5848 = ~n15370 ;
  assign y5849 = n15371 ;
  assign y5850 = ~n15379 ;
  assign y5851 = n15384 ;
  assign y5852 = ~n15386 ;
  assign y5853 = n15389 ;
  assign y5854 = ~n15393 ;
  assign y5855 = n15394 ;
  assign y5856 = ~n15399 ;
  assign y5857 = ~n15401 ;
  assign y5858 = n1842 ;
  assign y5859 = ~n15404 ;
  assign y5860 = ~n15405 ;
  assign y5861 = n10338 ;
  assign y5862 = n13376 ;
  assign y5863 = ~n15407 ;
  assign y5864 = 1'b0 ;
  assign y5865 = ~1'b0 ;
  assign y5866 = ~n15415 ;
  assign y5867 = n15422 ;
  assign y5868 = ~1'b0 ;
  assign y5869 = ~n15424 ;
  assign y5870 = n15426 ;
  assign y5871 = ~n15428 ;
  assign y5872 = ~1'b0 ;
  assign y5873 = ~n15433 ;
  assign y5874 = ~1'b0 ;
  assign y5875 = ~n15434 ;
  assign y5876 = ~1'b0 ;
  assign y5877 = ~n15437 ;
  assign y5878 = ~1'b0 ;
  assign y5879 = ~n15442 ;
  assign y5880 = ~n15443 ;
  assign y5881 = ~n15446 ;
  assign y5882 = ~1'b0 ;
  assign y5883 = ~1'b0 ;
  assign y5884 = ~n15448 ;
  assign y5885 = ~n15450 ;
  assign y5886 = ~n15454 ;
  assign y5887 = ~n15464 ;
  assign y5888 = n15465 ;
  assign y5889 = n15467 ;
  assign y5890 = n15468 ;
  assign y5891 = n15472 ;
  assign y5892 = ~n15473 ;
  assign y5893 = ~n15475 ;
  assign y5894 = ~1'b0 ;
  assign y5895 = ~n15477 ;
  assign y5896 = n15479 ;
  assign y5897 = ~1'b0 ;
  assign y5898 = n15481 ;
  assign y5899 = ~n15482 ;
  assign y5900 = ~n15484 ;
  assign y5901 = ~n15488 ;
  assign y5902 = n15494 ;
  assign y5903 = ~n15500 ;
  assign y5904 = ~1'b0 ;
  assign y5905 = ~n15507 ;
  assign y5906 = n15508 ;
  assign y5907 = ~n15509 ;
  assign y5908 = n15510 ;
  assign y5909 = n15511 ;
  assign y5910 = ~1'b0 ;
  assign y5911 = ~1'b0 ;
  assign y5912 = ~n15513 ;
  assign y5913 = n15516 ;
  assign y5914 = ~n15520 ;
  assign y5915 = n15521 ;
  assign y5916 = ~1'b0 ;
  assign y5917 = n15526 ;
  assign y5918 = ~n15527 ;
  assign y5919 = ~n15528 ;
  assign y5920 = n15531 ;
  assign y5921 = ~n15532 ;
  assign y5922 = n15539 ;
  assign y5923 = ~n15543 ;
  assign y5924 = ~1'b0 ;
  assign y5925 = ~1'b0 ;
  assign y5926 = n15552 ;
  assign y5927 = ~n15553 ;
  assign y5928 = ~n15554 ;
  assign y5929 = ~n15556 ;
  assign y5930 = ~n15557 ;
  assign y5931 = ~1'b0 ;
  assign y5932 = ~n15559 ;
  assign y5933 = n872 ;
  assign y5934 = ~1'b0 ;
  assign y5935 = n15560 ;
  assign y5936 = ~n15562 ;
  assign y5937 = ~n15568 ;
  assign y5938 = n15570 ;
  assign y5939 = ~n15572 ;
  assign y5940 = n15573 ;
  assign y5941 = ~n15576 ;
  assign y5942 = ~1'b0 ;
  assign y5943 = ~1'b0 ;
  assign y5944 = ~n15577 ;
  assign y5945 = n15578 ;
  assign y5946 = ~n15586 ;
  assign y5947 = ~1'b0 ;
  assign y5948 = ~1'b0 ;
  assign y5949 = ~1'b0 ;
  assign y5950 = ~n231 ;
  assign y5951 = n15589 ;
  assign y5952 = n15590 ;
  assign y5953 = ~n15592 ;
  assign y5954 = ~1'b0 ;
  assign y5955 = n15599 ;
  assign y5956 = n15601 ;
  assign y5957 = ~n15603 ;
  assign y5958 = ~n15604 ;
  assign y5959 = n15608 ;
  assign y5960 = ~1'b0 ;
  assign y5961 = ~1'b0 ;
  assign y5962 = n15616 ;
  assign y5963 = ~n15617 ;
  assign y5964 = ~n15619 ;
  assign y5965 = ~n15623 ;
  assign y5966 = ~n15624 ;
  assign y5967 = n10119 ;
  assign y5968 = n15628 ;
  assign y5969 = ~n15633 ;
  assign y5970 = ~n15634 ;
  assign y5971 = n15638 ;
  assign y5972 = ~1'b0 ;
  assign y5973 = ~1'b0 ;
  assign y5974 = ~1'b0 ;
  assign y5975 = ~1'b0 ;
  assign y5976 = ~n15644 ;
  assign y5977 = ~n15645 ;
  assign y5978 = ~n15646 ;
  assign y5979 = ~1'b0 ;
  assign y5980 = n15649 ;
  assign y5981 = ~1'b0 ;
  assign y5982 = ~n15651 ;
  assign y5983 = n15652 ;
  assign y5984 = n15653 ;
  assign y5985 = n15657 ;
  assign y5986 = n15662 ;
  assign y5987 = n15667 ;
  assign y5988 = n15671 ;
  assign y5989 = ~1'b0 ;
  assign y5990 = n15679 ;
  assign y5991 = ~1'b0 ;
  assign y5992 = n15680 ;
  assign y5993 = n15688 ;
  assign y5994 = ~n15691 ;
  assign y5995 = n15692 ;
  assign y5996 = n15697 ;
  assign y5997 = n15698 ;
  assign y5998 = n13198 ;
  assign y5999 = n15700 ;
  assign y6000 = n15704 ;
  assign y6001 = ~n15709 ;
  assign y6002 = n15713 ;
  assign y6003 = ~1'b0 ;
  assign y6004 = ~1'b0 ;
  assign y6005 = n15715 ;
  assign y6006 = ~1'b0 ;
  assign y6007 = ~1'b0 ;
  assign y6008 = n15716 ;
  assign y6009 = ~n15720 ;
  assign y6010 = ~n15726 ;
  assign y6011 = ~1'b0 ;
  assign y6012 = n15728 ;
  assign y6013 = ~1'b0 ;
  assign y6014 = n15729 ;
  assign y6015 = n15730 ;
  assign y6016 = n15732 ;
  assign y6017 = 1'b0 ;
  assign y6018 = ~n15742 ;
  assign y6019 = n15748 ;
  assign y6020 = ~n15749 ;
  assign y6021 = ~n15751 ;
  assign y6022 = n15756 ;
  assign y6023 = ~n15757 ;
  assign y6024 = ~n14738 ;
  assign y6025 = ~n15760 ;
  assign y6026 = ~n15764 ;
  assign y6027 = ~n15773 ;
  assign y6028 = n15775 ;
  assign y6029 = n15776 ;
  assign y6030 = ~n15777 ;
  assign y6031 = n15778 ;
  assign y6032 = n15779 ;
  assign y6033 = ~1'b0 ;
  assign y6034 = n15782 ;
  assign y6035 = n15790 ;
  assign y6036 = ~n15792 ;
  assign y6037 = ~n15797 ;
  assign y6038 = ~1'b0 ;
  assign y6039 = ~1'b0 ;
  assign y6040 = n15802 ;
  assign y6041 = ~1'b0 ;
  assign y6042 = n15807 ;
  assign y6043 = ~n15808 ;
  assign y6044 = ~n15816 ;
  assign y6045 = n15819 ;
  assign y6046 = n15821 ;
  assign y6047 = n15826 ;
  assign y6048 = ~n15831 ;
  assign y6049 = ~n15832 ;
  assign y6050 = n15838 ;
  assign y6051 = ~n15840 ;
  assign y6052 = n15843 ;
  assign y6053 = ~n15844 ;
  assign y6054 = ~n15847 ;
  assign y6055 = n15849 ;
  assign y6056 = ~n15850 ;
  assign y6057 = ~1'b0 ;
  assign y6058 = ~n15858 ;
  assign y6059 = n15859 ;
  assign y6060 = n15868 ;
  assign y6061 = ~1'b0 ;
  assign y6062 = ~1'b0 ;
  assign y6063 = n15870 ;
  assign y6064 = ~n15872 ;
  assign y6065 = ~n15873 ;
  assign y6066 = ~n15875 ;
  assign y6067 = ~1'b0 ;
  assign y6068 = ~1'b0 ;
  assign y6069 = ~n7892 ;
  assign y6070 = ~n15878 ;
  assign y6071 = n15879 ;
  assign y6072 = ~1'b0 ;
  assign y6073 = ~1'b0 ;
  assign y6074 = ~n5773 ;
  assign y6075 = ~1'b0 ;
  assign y6076 = n15881 ;
  assign y6077 = ~n15884 ;
  assign y6078 = ~1'b0 ;
  assign y6079 = ~1'b0 ;
  assign y6080 = ~n15889 ;
  assign y6081 = n15891 ;
  assign y6082 = ~1'b0 ;
  assign y6083 = n15902 ;
  assign y6084 = ~1'b0 ;
  assign y6085 = ~n15911 ;
  assign y6086 = ~1'b0 ;
  assign y6087 = ~n15912 ;
  assign y6088 = n15913 ;
  assign y6089 = ~n15915 ;
  assign y6090 = n15918 ;
  assign y6091 = n15920 ;
  assign y6092 = ~n15921 ;
  assign y6093 = ~1'b0 ;
  assign y6094 = n15922 ;
  assign y6095 = ~1'b0 ;
  assign y6096 = n15929 ;
  assign y6097 = n15931 ;
  assign y6098 = n15932 ;
  assign y6099 = ~n15937 ;
  assign y6100 = ~n15940 ;
  assign y6101 = ~1'b0 ;
  assign y6102 = n15942 ;
  assign y6103 = ~1'b0 ;
  assign y6104 = ~n15945 ;
  assign y6105 = ~n15947 ;
  assign y6106 = ~1'b0 ;
  assign y6107 = n15948 ;
  assign y6108 = n13545 ;
  assign y6109 = 1'b0 ;
  assign y6110 = ~1'b0 ;
  assign y6111 = ~1'b0 ;
  assign y6112 = n15949 ;
  assign y6113 = ~1'b0 ;
  assign y6114 = ~1'b0 ;
  assign y6115 = n15952 ;
  assign y6116 = n15956 ;
  assign y6117 = ~1'b0 ;
  assign y6118 = 1'b0 ;
  assign y6119 = n15958 ;
  assign y6120 = ~n15964 ;
  assign y6121 = ~n15967 ;
  assign y6122 = n15970 ;
  assign y6123 = n15971 ;
  assign y6124 = n15972 ;
  assign y6125 = n11582 ;
  assign y6126 = 1'b0 ;
  assign y6127 = ~n15974 ;
  assign y6128 = ~n15976 ;
  assign y6129 = n15979 ;
  assign y6130 = n3821 ;
  assign y6131 = n15985 ;
  assign y6132 = ~1'b0 ;
  assign y6133 = n15987 ;
  assign y6134 = ~n15993 ;
  assign y6135 = n15994 ;
  assign y6136 = n15997 ;
  assign y6137 = n15999 ;
  assign y6138 = ~1'b0 ;
  assign y6139 = n16002 ;
  assign y6140 = n16006 ;
  assign y6141 = ~n16007 ;
  assign y6142 = ~n16009 ;
  assign y6143 = n16012 ;
  assign y6144 = n16013 ;
  assign y6145 = ~1'b0 ;
  assign y6146 = ~n16015 ;
  assign y6147 = ~n16019 ;
  assign y6148 = ~n16023 ;
  assign y6149 = ~n16027 ;
  assign y6150 = ~n16034 ;
  assign y6151 = ~n7294 ;
  assign y6152 = ~n16039 ;
  assign y6153 = ~n8689 ;
  assign y6154 = ~n16044 ;
  assign y6155 = ~1'b0 ;
  assign y6156 = n16045 ;
  assign y6157 = ~n16049 ;
  assign y6158 = ~n16050 ;
  assign y6159 = ~n16055 ;
  assign y6160 = n16058 ;
  assign y6161 = n16062 ;
  assign y6162 = ~1'b0 ;
  assign y6163 = n16063 ;
  assign y6164 = ~n16064 ;
  assign y6165 = n16066 ;
  assign y6166 = n16068 ;
  assign y6167 = ~n16072 ;
  assign y6168 = ~n16080 ;
  assign y6169 = n16088 ;
  assign y6170 = x60 ;
  assign y6171 = n16091 ;
  assign y6172 = ~n16095 ;
  assign y6173 = n16098 ;
  assign y6174 = n16102 ;
  assign y6175 = ~n16107 ;
  assign y6176 = n16111 ;
  assign y6177 = ~n16113 ;
  assign y6178 = n16119 ;
  assign y6179 = n10165 ;
  assign y6180 = n16123 ;
  assign y6181 = n16129 ;
  assign y6182 = n16133 ;
  assign y6183 = ~n1995 ;
  assign y6184 = ~n16137 ;
  assign y6185 = n16138 ;
  assign y6186 = ~1'b0 ;
  assign y6187 = n16140 ;
  assign y6188 = ~n16141 ;
  assign y6189 = ~n16142 ;
  assign y6190 = ~n16143 ;
  assign y6191 = ~n16146 ;
  assign y6192 = n16147 ;
  assign y6193 = n11207 ;
  assign y6194 = ~n16148 ;
  assign y6195 = n16150 ;
  assign y6196 = n16155 ;
  assign y6197 = ~1'b0 ;
  assign y6198 = n16157 ;
  assign y6199 = ~n13843 ;
  assign y6200 = ~n16160 ;
  assign y6201 = ~1'b0 ;
  assign y6202 = ~1'b0 ;
  assign y6203 = ~n16162 ;
  assign y6204 = ~1'b0 ;
  assign y6205 = n16163 ;
  assign y6206 = ~n11260 ;
  assign y6207 = n16165 ;
  assign y6208 = n16166 ;
  assign y6209 = ~1'b0 ;
  assign y6210 = n16168 ;
  assign y6211 = ~n16169 ;
  assign y6212 = n16170 ;
  assign y6213 = ~n16177 ;
  assign y6214 = ~1'b0 ;
  assign y6215 = ~n16182 ;
  assign y6216 = ~n16191 ;
  assign y6217 = n16192 ;
  assign y6218 = ~n16198 ;
  assign y6219 = ~1'b0 ;
  assign y6220 = n16199 ;
  assign y6221 = ~1'b0 ;
  assign y6222 = ~n16201 ;
  assign y6223 = ~1'b0 ;
  assign y6224 = n16203 ;
  assign y6225 = 1'b0 ;
  assign y6226 = ~n16213 ;
  assign y6227 = ~1'b0 ;
  assign y6228 = ~n9392 ;
  assign y6229 = ~n16214 ;
  assign y6230 = n16215 ;
  assign y6231 = ~1'b0 ;
  assign y6232 = n16217 ;
  assign y6233 = ~1'b0 ;
  assign y6234 = ~n16223 ;
  assign y6235 = ~n16225 ;
  assign y6236 = ~n16228 ;
  assign y6237 = ~n10464 ;
  assign y6238 = n16234 ;
  assign y6239 = ~n16237 ;
  assign y6240 = ~n16240 ;
  assign y6241 = ~n16245 ;
  assign y6242 = ~n16248 ;
  assign y6243 = n1373 ;
  assign y6244 = n16250 ;
  assign y6245 = ~1'b0 ;
  assign y6246 = ~1'b0 ;
  assign y6247 = ~1'b0 ;
  assign y6248 = ~n16253 ;
  assign y6249 = ~1'b0 ;
  assign y6250 = n16254 ;
  assign y6251 = ~n16255 ;
  assign y6252 = ~n16257 ;
  assign y6253 = ~n16265 ;
  assign y6254 = n16269 ;
  assign y6255 = ~n16271 ;
  assign y6256 = ~1'b0 ;
  assign y6257 = ~n16275 ;
  assign y6258 = ~n16276 ;
  assign y6259 = ~n16281 ;
  assign y6260 = ~n16283 ;
  assign y6261 = n16285 ;
  assign y6262 = ~n16289 ;
  assign y6263 = n16290 ;
  assign y6264 = ~1'b0 ;
  assign y6265 = ~1'b0 ;
  assign y6266 = n16291 ;
  assign y6267 = n16292 ;
  assign y6268 = ~n16293 ;
  assign y6269 = ~1'b0 ;
  assign y6270 = ~n12149 ;
  assign y6271 = ~1'b0 ;
  assign y6272 = ~n16295 ;
  assign y6273 = n16297 ;
  assign y6274 = ~n16300 ;
  assign y6275 = ~n16303 ;
  assign y6276 = ~n16309 ;
  assign y6277 = n16311 ;
  assign y6278 = ~1'b0 ;
  assign y6279 = n16316 ;
  assign y6280 = ~n16320 ;
  assign y6281 = ~n16324 ;
  assign y6282 = ~1'b0 ;
  assign y6283 = ~1'b0 ;
  assign y6284 = ~1'b0 ;
  assign y6285 = ~1'b0 ;
  assign y6286 = n16331 ;
  assign y6287 = n16332 ;
  assign y6288 = ~n16334 ;
  assign y6289 = ~1'b0 ;
  assign y6290 = n16337 ;
  assign y6291 = ~n16338 ;
  assign y6292 = ~n16346 ;
  assign y6293 = n16349 ;
  assign y6294 = ~n16352 ;
  assign y6295 = n16356 ;
  assign y6296 = ~n16364 ;
  assign y6297 = n16371 ;
  assign y6298 = ~n16386 ;
  assign y6299 = n16389 ;
  assign y6300 = 1'b0 ;
  assign y6301 = ~n16390 ;
  assign y6302 = n16391 ;
  assign y6303 = ~n16397 ;
  assign y6304 = n16403 ;
  assign y6305 = ~n16407 ;
  assign y6306 = ~n16414 ;
  assign y6307 = n16416 ;
  assign y6308 = ~1'b0 ;
  assign y6309 = n16421 ;
  assign y6310 = ~1'b0 ;
  assign y6311 = ~n16423 ;
  assign y6312 = n16424 ;
  assign y6313 = n16425 ;
  assign y6314 = ~1'b0 ;
  assign y6315 = ~1'b0 ;
  assign y6316 = ~1'b0 ;
  assign y6317 = ~n16426 ;
  assign y6318 = n16427 ;
  assign y6319 = ~n16429 ;
  assign y6320 = n16430 ;
  assign y6321 = ~1'b0 ;
  assign y6322 = x28 ;
  assign y6323 = 1'b0 ;
  assign y6324 = ~1'b0 ;
  assign y6325 = n16432 ;
  assign y6326 = ~1'b0 ;
  assign y6327 = n16433 ;
  assign y6328 = n16436 ;
  assign y6329 = ~n16437 ;
  assign y6330 = ~1'b0 ;
  assign y6331 = n16439 ;
  assign y6332 = ~n16440 ;
  assign y6333 = ~n16441 ;
  assign y6334 = ~n16442 ;
  assign y6335 = ~1'b0 ;
  assign y6336 = ~n16452 ;
  assign y6337 = ~n16460 ;
  assign y6338 = ~1'b0 ;
  assign y6339 = ~n16463 ;
  assign y6340 = n16467 ;
  assign y6341 = ~n16469 ;
  assign y6342 = n16481 ;
  assign y6343 = n16487 ;
  assign y6344 = n16494 ;
  assign y6345 = n16495 ;
  assign y6346 = n16498 ;
  assign y6347 = n16505 ;
  assign y6348 = n8199 ;
  assign y6349 = n16506 ;
  assign y6350 = ~1'b0 ;
  assign y6351 = ~1'b0 ;
  assign y6352 = n16510 ;
  assign y6353 = n16511 ;
  assign y6354 = ~n16513 ;
  assign y6355 = n16517 ;
  assign y6356 = ~1'b0 ;
  assign y6357 = ~n16522 ;
  assign y6358 = n16526 ;
  assign y6359 = n16533 ;
  assign y6360 = ~n16534 ;
  assign y6361 = ~1'b0 ;
  assign y6362 = ~n16537 ;
  assign y6363 = n16538 ;
  assign y6364 = ~n16540 ;
  assign y6365 = ~1'b0 ;
  assign y6366 = ~n16544 ;
  assign y6367 = n16546 ;
  assign y6368 = n16549 ;
  assign y6369 = ~n16550 ;
  assign y6370 = ~n16551 ;
  assign y6371 = n16552 ;
  assign y6372 = n16557 ;
  assign y6373 = ~n16559 ;
  assign y6374 = ~n16561 ;
  assign y6375 = ~n16567 ;
  assign y6376 = ~n16569 ;
  assign y6377 = ~n16570 ;
  assign y6378 = ~n16571 ;
  assign y6379 = ~n16573 ;
  assign y6380 = n16575 ;
  assign y6381 = ~n220 ;
  assign y6382 = n16582 ;
  assign y6383 = n16585 ;
  assign y6384 = ~1'b0 ;
  assign y6385 = ~1'b0 ;
  assign y6386 = ~1'b0 ;
  assign y6387 = ~n16586 ;
  assign y6388 = 1'b0 ;
  assign y6389 = ~1'b0 ;
  assign y6390 = ~n16588 ;
  assign y6391 = n16590 ;
  assign y6392 = ~n16597 ;
  assign y6393 = ~n16598 ;
  assign y6394 = ~n16601 ;
  assign y6395 = ~n16605 ;
  assign y6396 = ~n16607 ;
  assign y6397 = ~n763 ;
  assign y6398 = ~1'b0 ;
  assign y6399 = ~n16614 ;
  assign y6400 = ~n16615 ;
  assign y6401 = ~n16619 ;
  assign y6402 = n16620 ;
  assign y6403 = ~1'b0 ;
  assign y6404 = ~n16626 ;
  assign y6405 = n16628 ;
  assign y6406 = n16629 ;
  assign y6407 = ~1'b0 ;
  assign y6408 = ~n16630 ;
  assign y6409 = n16631 ;
  assign y6410 = n16636 ;
  assign y6411 = n16639 ;
  assign y6412 = ~n16642 ;
  assign y6413 = n16646 ;
  assign y6414 = ~1'b0 ;
  assign y6415 = ~1'b0 ;
  assign y6416 = n16648 ;
  assign y6417 = ~n16657 ;
  assign y6418 = ~n16659 ;
  assign y6419 = ~n16661 ;
  assign y6420 = ~1'b0 ;
  assign y6421 = ~n16663 ;
  assign y6422 = ~1'b0 ;
  assign y6423 = n16664 ;
  assign y6424 = n16668 ;
  assign y6425 = ~n16669 ;
  assign y6426 = ~n16670 ;
  assign y6427 = ~n16672 ;
  assign y6428 = n16679 ;
  assign y6429 = ~1'b0 ;
  assign y6430 = ~n16681 ;
  assign y6431 = ~n16682 ;
  assign y6432 = n16685 ;
  assign y6433 = n16687 ;
  assign y6434 = ~n16688 ;
  assign y6435 = n16691 ;
  assign y6436 = ~1'b0 ;
  assign y6437 = ~n13789 ;
  assign y6438 = ~n16694 ;
  assign y6439 = n16696 ;
  assign y6440 = n16698 ;
  assign y6441 = ~1'b0 ;
  assign y6442 = ~n16701 ;
  assign y6443 = n16704 ;
  assign y6444 = n16705 ;
  assign y6445 = ~n16706 ;
  assign y6446 = ~n16714 ;
  assign y6447 = n16716 ;
  assign y6448 = n16717 ;
  assign y6449 = ~n16718 ;
  assign y6450 = n16723 ;
  assign y6451 = n16729 ;
  assign y6452 = ~n16731 ;
  assign y6453 = ~1'b0 ;
  assign y6454 = ~n16735 ;
  assign y6455 = ~1'b0 ;
  assign y6456 = n16739 ;
  assign y6457 = n16741 ;
  assign y6458 = ~n16744 ;
  assign y6459 = n16748 ;
  assign y6460 = 1'b0 ;
  assign y6461 = ~n16750 ;
  assign y6462 = n16751 ;
  assign y6463 = ~1'b0 ;
  assign y6464 = ~n16756 ;
  assign y6465 = ~1'b0 ;
  assign y6466 = ~n16758 ;
  assign y6467 = n16759 ;
  assign y6468 = ~n16761 ;
  assign y6469 = n16765 ;
  assign y6470 = ~n16767 ;
  assign y6471 = ~1'b0 ;
  assign y6472 = ~n16768 ;
  assign y6473 = n16769 ;
  assign y6474 = n16770 ;
  assign y6475 = ~n16771 ;
  assign y6476 = ~1'b0 ;
  assign y6477 = ~n16772 ;
  assign y6478 = n16773 ;
  assign y6479 = ~n16777 ;
  assign y6480 = n16778 ;
  assign y6481 = ~1'b0 ;
  assign y6482 = ~n16785 ;
  assign y6483 = ~n16787 ;
  assign y6484 = ~n16788 ;
  assign y6485 = ~n16793 ;
  assign y6486 = ~n16794 ;
  assign y6487 = ~1'b0 ;
  assign y6488 = n16797 ;
  assign y6489 = n16798 ;
  assign y6490 = ~1'b0 ;
  assign y6491 = ~1'b0 ;
  assign y6492 = n16799 ;
  assign y6493 = n16804 ;
  assign y6494 = n16811 ;
  assign y6495 = ~n16812 ;
  assign y6496 = ~1'b0 ;
  assign y6497 = n16816 ;
  assign y6498 = n16818 ;
  assign y6499 = n16819 ;
  assign y6500 = ~1'b0 ;
  assign y6501 = ~1'b0 ;
  assign y6502 = ~1'b0 ;
  assign y6503 = ~n16822 ;
  assign y6504 = ~n16826 ;
  assign y6505 = ~n16827 ;
  assign y6506 = ~n16829 ;
  assign y6507 = n16831 ;
  assign y6508 = n16832 ;
  assign y6509 = n16833 ;
  assign y6510 = n16838 ;
  assign y6511 = ~n16841 ;
  assign y6512 = ~n16843 ;
  assign y6513 = ~n16845 ;
  assign y6514 = ~1'b0 ;
  assign y6515 = ~1'b0 ;
  assign y6516 = ~n1175 ;
  assign y6517 = ~n16850 ;
  assign y6518 = n16853 ;
  assign y6519 = ~1'b0 ;
  assign y6520 = ~1'b0 ;
  assign y6521 = ~n16855 ;
  assign y6522 = n16857 ;
  assign y6523 = n16862 ;
  assign y6524 = n16865 ;
  assign y6525 = n16866 ;
  assign y6526 = ~n16874 ;
  assign y6527 = ~n16875 ;
  assign y6528 = ~1'b0 ;
  assign y6529 = ~n16881 ;
  assign y6530 = n16882 ;
  assign y6531 = ~n16886 ;
  assign y6532 = ~n2597 ;
  assign y6533 = ~n16888 ;
  assign y6534 = ~n16889 ;
  assign y6535 = n16891 ;
  assign y6536 = n16894 ;
  assign y6537 = ~n16897 ;
  assign y6538 = ~1'b0 ;
  assign y6539 = ~1'b0 ;
  assign y6540 = n16899 ;
  assign y6541 = n16902 ;
  assign y6542 = ~n16904 ;
  assign y6543 = ~n16912 ;
  assign y6544 = n16914 ;
  assign y6545 = ~1'b0 ;
  assign y6546 = ~n16916 ;
  assign y6547 = n16920 ;
  assign y6548 = ~n16922 ;
  assign y6549 = ~n16925 ;
  assign y6550 = ~n16927 ;
  assign y6551 = n16931 ;
  assign y6552 = ~n16934 ;
  assign y6553 = ~1'b0 ;
  assign y6554 = ~n16936 ;
  assign y6555 = ~n16938 ;
  assign y6556 = ~n16946 ;
  assign y6557 = n16950 ;
  assign y6558 = ~1'b0 ;
  assign y6559 = ~1'b0 ;
  assign y6560 = n16951 ;
  assign y6561 = ~n16952 ;
  assign y6562 = n16953 ;
  assign y6563 = n16954 ;
  assign y6564 = n16965 ;
  assign y6565 = n16969 ;
  assign y6566 = n16973 ;
  assign y6567 = ~1'b0 ;
  assign y6568 = ~n16978 ;
  assign y6569 = ~n16982 ;
  assign y6570 = ~n16983 ;
  assign y6571 = n3748 ;
  assign y6572 = n16987 ;
  assign y6573 = n16989 ;
  assign y6574 = n16993 ;
  assign y6575 = ~n17000 ;
  assign y6576 = ~1'b0 ;
  assign y6577 = ~1'b0 ;
  assign y6578 = n17001 ;
  assign y6579 = ~n17003 ;
  assign y6580 = ~n17004 ;
  assign y6581 = n17005 ;
  assign y6582 = ~1'b0 ;
  assign y6583 = ~n17013 ;
  assign y6584 = ~n17016 ;
  assign y6585 = n17018 ;
  assign y6586 = n17023 ;
  assign y6587 = ~1'b0 ;
  assign y6588 = n17025 ;
  assign y6589 = ~1'b0 ;
  assign y6590 = n17026 ;
  assign y6591 = ~n17028 ;
  assign y6592 = ~n17029 ;
  assign y6593 = n17030 ;
  assign y6594 = ~1'b0 ;
  assign y6595 = n17032 ;
  assign y6596 = n17036 ;
  assign y6597 = ~1'b0 ;
  assign y6598 = n6749 ;
  assign y6599 = ~n17040 ;
  assign y6600 = ~n17046 ;
  assign y6601 = n17050 ;
  assign y6602 = ~1'b0 ;
  assign y6603 = ~1'b0 ;
  assign y6604 = ~n17051 ;
  assign y6605 = ~1'b0 ;
  assign y6606 = n6806 ;
  assign y6607 = n17053 ;
  assign y6608 = ~n17059 ;
  assign y6609 = n17062 ;
  assign y6610 = ~n17063 ;
  assign y6611 = n17067 ;
  assign y6612 = ~n17068 ;
  assign y6613 = n17071 ;
  assign y6614 = ~n17078 ;
  assign y6615 = n17081 ;
  assign y6616 = ~1'b0 ;
  assign y6617 = ~n17082 ;
  assign y6618 = n17088 ;
  assign y6619 = ~n17096 ;
  assign y6620 = n17098 ;
  assign y6621 = ~n17099 ;
  assign y6622 = ~n4593 ;
  assign y6623 = ~n17103 ;
  assign y6624 = ~n17105 ;
  assign y6625 = n17106 ;
  assign y6626 = n17108 ;
  assign y6627 = ~n17110 ;
  assign y6628 = ~1'b0 ;
  assign y6629 = n17111 ;
  assign y6630 = ~n17122 ;
  assign y6631 = ~n17132 ;
  assign y6632 = ~n17133 ;
  assign y6633 = n17135 ;
  assign y6634 = ~n17138 ;
  assign y6635 = ~n17139 ;
  assign y6636 = 1'b0 ;
  assign y6637 = n17143 ;
  assign y6638 = ~n17146 ;
  assign y6639 = n17151 ;
  assign y6640 = ~n17158 ;
  assign y6641 = ~n17161 ;
  assign y6642 = ~n17162 ;
  assign y6643 = ~n17164 ;
  assign y6644 = ~n17168 ;
  assign y6645 = ~n17169 ;
  assign y6646 = ~n17170 ;
  assign y6647 = ~1'b0 ;
  assign y6648 = ~n17173 ;
  assign y6649 = ~1'b0 ;
  assign y6650 = ~n17174 ;
  assign y6651 = n17178 ;
  assign y6652 = n17194 ;
  assign y6653 = n17201 ;
  assign y6654 = ~n17202 ;
  assign y6655 = n17208 ;
  assign y6656 = n17212 ;
  assign y6657 = ~n17216 ;
  assign y6658 = ~n17217 ;
  assign y6659 = ~1'b0 ;
  assign y6660 = n17218 ;
  assign y6661 = ~n17222 ;
  assign y6662 = 1'b0 ;
  assign y6663 = ~1'b0 ;
  assign y6664 = n17226 ;
  assign y6665 = n17229 ;
  assign y6666 = ~1'b0 ;
  assign y6667 = n17233 ;
  assign y6668 = n17234 ;
  assign y6669 = ~n17239 ;
  assign y6670 = ~n17241 ;
  assign y6671 = ~n17246 ;
  assign y6672 = ~n17253 ;
  assign y6673 = ~n17259 ;
  assign y6674 = ~1'b0 ;
  assign y6675 = n17262 ;
  assign y6676 = ~n17263 ;
  assign y6677 = n17266 ;
  assign y6678 = ~n17267 ;
  assign y6679 = ~n17271 ;
  assign y6680 = ~1'b0 ;
  assign y6681 = ~n17280 ;
  assign y6682 = ~n17285 ;
  assign y6683 = 1'b0 ;
  assign y6684 = ~n17289 ;
  assign y6685 = ~n17295 ;
  assign y6686 = ~1'b0 ;
  assign y6687 = n17296 ;
  assign y6688 = ~n17297 ;
  assign y6689 = ~n17299 ;
  assign y6690 = ~1'b0 ;
  assign y6691 = ~n17301 ;
  assign y6692 = ~n17303 ;
  assign y6693 = ~1'b0 ;
  assign y6694 = ~n17304 ;
  assign y6695 = ~n17323 ;
  assign y6696 = n17326 ;
  assign y6697 = n17337 ;
  assign y6698 = n17345 ;
  assign y6699 = n17347 ;
  assign y6700 = n17351 ;
  assign y6701 = n17352 ;
  assign y6702 = n17376 ;
  assign y6703 = n17377 ;
  assign y6704 = ~1'b0 ;
  assign y6705 = ~n17382 ;
  assign y6706 = ~n17384 ;
  assign y6707 = ~n17388 ;
  assign y6708 = n17392 ;
  assign y6709 = ~1'b0 ;
  assign y6710 = n17393 ;
  assign y6711 = ~1'b0 ;
  assign y6712 = ~n17394 ;
  assign y6713 = ~n17396 ;
  assign y6714 = ~1'b0 ;
  assign y6715 = ~1'b0 ;
  assign y6716 = ~1'b0 ;
  assign y6717 = n17402 ;
  assign y6718 = n17405 ;
  assign y6719 = ~n17411 ;
  assign y6720 = n17416 ;
  assign y6721 = ~n17418 ;
  assign y6722 = n17423 ;
  assign y6723 = n17426 ;
  assign y6724 = ~1'b0 ;
  assign y6725 = ~n17429 ;
  assign y6726 = n17431 ;
  assign y6727 = n17434 ;
  assign y6728 = ~n17439 ;
  assign y6729 = ~n17442 ;
  assign y6730 = ~n17443 ;
  assign y6731 = n17453 ;
  assign y6732 = ~1'b0 ;
  assign y6733 = ~n17455 ;
  assign y6734 = ~n17458 ;
  assign y6735 = n17463 ;
  assign y6736 = ~n17464 ;
  assign y6737 = n17466 ;
  assign y6738 = ~n17471 ;
  assign y6739 = ~1'b0 ;
  assign y6740 = ~1'b0 ;
  assign y6741 = n17475 ;
  assign y6742 = n17477 ;
  assign y6743 = ~n17488 ;
  assign y6744 = n17491 ;
  assign y6745 = ~n17493 ;
  assign y6746 = n17503 ;
  assign y6747 = ~n17508 ;
  assign y6748 = n17511 ;
  assign y6749 = ~1'b0 ;
  assign y6750 = ~1'b0 ;
  assign y6751 = ~n17512 ;
  assign y6752 = ~n17513 ;
  assign y6753 = n17521 ;
  assign y6754 = ~1'b0 ;
  assign y6755 = ~n17525 ;
  assign y6756 = ~1'b0 ;
  assign y6757 = n17526 ;
  assign y6758 = ~n17528 ;
  assign y6759 = ~1'b0 ;
  assign y6760 = n5717 ;
  assign y6761 = ~n17529 ;
  assign y6762 = n17531 ;
  assign y6763 = ~1'b0 ;
  assign y6764 = ~n17535 ;
  assign y6765 = ~1'b0 ;
  assign y6766 = n6530 ;
  assign y6767 = 1'b0 ;
  assign y6768 = n17536 ;
  assign y6769 = ~n17537 ;
  assign y6770 = n17543 ;
  assign y6771 = ~1'b0 ;
  assign y6772 = ~1'b0 ;
  assign y6773 = ~1'b0 ;
  assign y6774 = n17545 ;
  assign y6775 = n17546 ;
  assign y6776 = ~1'b0 ;
  assign y6777 = ~n17548 ;
  assign y6778 = ~n17549 ;
  assign y6779 = n17554 ;
  assign y6780 = ~n17558 ;
  assign y6781 = n17565 ;
  assign y6782 = ~1'b0 ;
  assign y6783 = ~n17567 ;
  assign y6784 = ~1'b0 ;
  assign y6785 = n17570 ;
  assign y6786 = n17572 ;
  assign y6787 = ~n17577 ;
  assign y6788 = ~n17578 ;
  assign y6789 = n17581 ;
  assign y6790 = n17582 ;
  assign y6791 = ~n17584 ;
  assign y6792 = ~n17585 ;
  assign y6793 = n17588 ;
  assign y6794 = ~n17589 ;
  assign y6795 = ~1'b0 ;
  assign y6796 = n17590 ;
  assign y6797 = ~n17595 ;
  assign y6798 = n17597 ;
  assign y6799 = ~n17604 ;
  assign y6800 = n17608 ;
  assign y6801 = ~n17612 ;
  assign y6802 = ~n17620 ;
  assign y6803 = ~1'b0 ;
  assign y6804 = ~n17622 ;
  assign y6805 = ~1'b0 ;
  assign y6806 = n17625 ;
  assign y6807 = ~n17629 ;
  assign y6808 = ~n17630 ;
  assign y6809 = n17634 ;
  assign y6810 = ~1'b0 ;
  assign y6811 = n17635 ;
  assign y6812 = ~n3834 ;
  assign y6813 = n17638 ;
  assign y6814 = n8576 ;
  assign y6815 = ~n17640 ;
  assign y6816 = ~n17644 ;
  assign y6817 = ~n17645 ;
  assign y6818 = ~1'b0 ;
  assign y6819 = n17648 ;
  assign y6820 = n17650 ;
  assign y6821 = ~1'b0 ;
  assign y6822 = ~n17654 ;
  assign y6823 = ~n17657 ;
  assign y6824 = ~n17659 ;
  assign y6825 = ~n17661 ;
  assign y6826 = ~1'b0 ;
  assign y6827 = ~n17662 ;
  assign y6828 = ~n17665 ;
  assign y6829 = ~n11752 ;
  assign y6830 = ~n17669 ;
  assign y6831 = ~1'b0 ;
  assign y6832 = n17671 ;
  assign y6833 = ~1'b0 ;
  assign y6834 = n17672 ;
  assign y6835 = ~1'b0 ;
  assign y6836 = n17673 ;
  assign y6837 = ~n17675 ;
  assign y6838 = n17677 ;
  assign y6839 = ~1'b0 ;
  assign y6840 = ~n17678 ;
  assign y6841 = n17679 ;
  assign y6842 = ~n3763 ;
  assign y6843 = ~1'b0 ;
  assign y6844 = n17682 ;
  assign y6845 = n17683 ;
  assign y6846 = n17687 ;
  assign y6847 = ~n17688 ;
  assign y6848 = n17691 ;
  assign y6849 = ~1'b0 ;
  assign y6850 = ~n17696 ;
  assign y6851 = ~1'b0 ;
  assign y6852 = ~n3263 ;
  assign y6853 = ~n17701 ;
  assign y6854 = n17706 ;
  assign y6855 = n13216 ;
  assign y6856 = ~n17707 ;
  assign y6857 = ~1'b0 ;
  assign y6858 = n17711 ;
  assign y6859 = n17715 ;
  assign y6860 = n17721 ;
  assign y6861 = ~n17723 ;
  assign y6862 = ~n17724 ;
  assign y6863 = n17725 ;
  assign y6864 = ~1'b0 ;
  assign y6865 = ~n17729 ;
  assign y6866 = n17731 ;
  assign y6867 = ~1'b0 ;
  assign y6868 = ~n17732 ;
  assign y6869 = ~n17737 ;
  assign y6870 = ~n17743 ;
  assign y6871 = n17744 ;
  assign y6872 = ~n17748 ;
  assign y6873 = ~n17751 ;
  assign y6874 = n17752 ;
  assign y6875 = ~n17756 ;
  assign y6876 = n17763 ;
  assign y6877 = ~n17765 ;
  assign y6878 = ~n17766 ;
  assign y6879 = ~n17772 ;
  assign y6880 = ~1'b0 ;
  assign y6881 = n17774 ;
  assign y6882 = n17777 ;
  assign y6883 = n17780 ;
  assign y6884 = ~1'b0 ;
  assign y6885 = n17782 ;
  assign y6886 = n17783 ;
  assign y6887 = n17786 ;
  assign y6888 = ~1'b0 ;
  assign y6889 = ~1'b0 ;
  assign y6890 = n17795 ;
  assign y6891 = n17797 ;
  assign y6892 = 1'b0 ;
  assign y6893 = n17800 ;
  assign y6894 = ~n17802 ;
  assign y6895 = ~1'b0 ;
  assign y6896 = n17809 ;
  assign y6897 = ~n17810 ;
  assign y6898 = n17812 ;
  assign y6899 = ~n7663 ;
  assign y6900 = ~1'b0 ;
  assign y6901 = ~n17814 ;
  assign y6902 = ~1'b0 ;
  assign y6903 = n17821 ;
  assign y6904 = n17825 ;
  assign y6905 = ~n17828 ;
  assign y6906 = ~n17831 ;
  assign y6907 = ~n17834 ;
  assign y6908 = ~1'b0 ;
  assign y6909 = ~1'b0 ;
  assign y6910 = ~n17835 ;
  assign y6911 = ~n17839 ;
  assign y6912 = ~1'b0 ;
  assign y6913 = n17840 ;
  assign y6914 = ~n17842 ;
  assign y6915 = ~n17844 ;
  assign y6916 = ~1'b0 ;
  assign y6917 = n17846 ;
  assign y6918 = n17848 ;
  assign y6919 = ~n17849 ;
  assign y6920 = ~n17853 ;
  assign y6921 = n17855 ;
  assign y6922 = n17856 ;
  assign y6923 = n17858 ;
  assign y6924 = ~1'b0 ;
  assign y6925 = ~1'b0 ;
  assign y6926 = n17860 ;
  assign y6927 = ~n17865 ;
  assign y6928 = ~n17867 ;
  assign y6929 = n17868 ;
  assign y6930 = n17874 ;
  assign y6931 = ~n17880 ;
  assign y6932 = ~1'b0 ;
  assign y6933 = n17884 ;
  assign y6934 = ~n17885 ;
  assign y6935 = ~n17889 ;
  assign y6936 = ~n17898 ;
  assign y6937 = n17899 ;
  assign y6938 = ~1'b0 ;
  assign y6939 = ~1'b0 ;
  assign y6940 = ~n17902 ;
  assign y6941 = ~1'b0 ;
  assign y6942 = n17905 ;
  assign y6943 = ~n17906 ;
  assign y6944 = ~n17907 ;
  assign y6945 = n17910 ;
  assign y6946 = n17912 ;
  assign y6947 = ~1'b0 ;
  assign y6948 = ~n17914 ;
  assign y6949 = n17916 ;
  assign y6950 = n17917 ;
  assign y6951 = n17919 ;
  assign y6952 = n17921 ;
  assign y6953 = n17923 ;
  assign y6954 = ~n5393 ;
  assign y6955 = ~1'b0 ;
  assign y6956 = ~1'b0 ;
  assign y6957 = n17924 ;
  assign y6958 = ~n17925 ;
  assign y6959 = n17928 ;
  assign y6960 = ~1'b0 ;
  assign y6961 = n17930 ;
  assign y6962 = ~n17931 ;
  assign y6963 = n17933 ;
  assign y6964 = ~n17937 ;
  assign y6965 = n17948 ;
  assign y6966 = n17950 ;
  assign y6967 = n17951 ;
  assign y6968 = n17956 ;
  assign y6969 = n17962 ;
  assign y6970 = ~n17963 ;
  assign y6971 = n17966 ;
  assign y6972 = n17974 ;
  assign y6973 = n17976 ;
  assign y6974 = n17978 ;
  assign y6975 = ~1'b0 ;
  assign y6976 = ~1'b0 ;
  assign y6977 = ~n17979 ;
  assign y6978 = n17983 ;
  assign y6979 = ~n17989 ;
  assign y6980 = ~1'b0 ;
  assign y6981 = ~n17994 ;
  assign y6982 = n17997 ;
  assign y6983 = n17998 ;
  assign y6984 = ~n18001 ;
  assign y6985 = ~n18007 ;
  assign y6986 = n18009 ;
  assign y6987 = n12783 ;
  assign y6988 = n18023 ;
  assign y6989 = ~n18028 ;
  assign y6990 = ~n18029 ;
  assign y6991 = n18030 ;
  assign y6992 = n18032 ;
  assign y6993 = ~n18034 ;
  assign y6994 = n18039 ;
  assign y6995 = ~n18045 ;
  assign y6996 = n18046 ;
  assign y6997 = ~n18048 ;
  assign y6998 = ~n18056 ;
  assign y6999 = n18059 ;
  assign y7000 = ~n18061 ;
  assign y7001 = ~n18062 ;
  assign y7002 = n18069 ;
  assign y7003 = ~1'b0 ;
  assign y7004 = ~n3345 ;
  assign y7005 = n18070 ;
  assign y7006 = ~1'b0 ;
  assign y7007 = n18071 ;
  assign y7008 = ~n18073 ;
  assign y7009 = ~n18075 ;
  assign y7010 = n18076 ;
  assign y7011 = ~n18081 ;
  assign y7012 = n18083 ;
  assign y7013 = ~n18089 ;
  assign y7014 = n18093 ;
  assign y7015 = n18099 ;
  assign y7016 = ~1'b0 ;
  assign y7017 = ~1'b0 ;
  assign y7018 = ~1'b0 ;
  assign y7019 = ~n18101 ;
  assign y7020 = ~n18103 ;
  assign y7021 = ~1'b0 ;
  assign y7022 = n18104 ;
  assign y7023 = n18105 ;
  assign y7024 = n18106 ;
  assign y7025 = ~1'b0 ;
  assign y7026 = n18109 ;
  assign y7027 = n18114 ;
  assign y7028 = n18116 ;
  assign y7029 = ~n18117 ;
  assign y7030 = ~1'b0 ;
  assign y7031 = ~n18121 ;
  assign y7032 = ~1'b0 ;
  assign y7033 = ~n18123 ;
  assign y7034 = ~n18126 ;
  assign y7035 = n18129 ;
  assign y7036 = ~n18130 ;
  assign y7037 = ~1'b0 ;
  assign y7038 = n18132 ;
  assign y7039 = ~n18133 ;
  assign y7040 = ~1'b0 ;
  assign y7041 = n18136 ;
  assign y7042 = ~n18137 ;
  assign y7043 = ~n18139 ;
  assign y7044 = ~n18140 ;
  assign y7045 = n18142 ;
  assign y7046 = n18143 ;
  assign y7047 = ~n18144 ;
  assign y7048 = n18148 ;
  assign y7049 = n18150 ;
  assign y7050 = ~n18152 ;
  assign y7051 = n18155 ;
  assign y7052 = ~1'b0 ;
  assign y7053 = ~n18158 ;
  assign y7054 = ~n18160 ;
  assign y7055 = n18165 ;
  assign y7056 = n18168 ;
  assign y7057 = ~n18169 ;
  assign y7058 = ~n18171 ;
  assign y7059 = ~1'b0 ;
  assign y7060 = ~n18173 ;
  assign y7061 = ~n18174 ;
  assign y7062 = ~n18178 ;
  assign y7063 = ~n18179 ;
  assign y7064 = ~1'b0 ;
  assign y7065 = ~n18181 ;
  assign y7066 = ~n1595 ;
  assign y7067 = ~n18182 ;
  assign y7068 = n18183 ;
  assign y7069 = ~1'b0 ;
  assign y7070 = ~1'b0 ;
  assign y7071 = n18186 ;
  assign y7072 = ~n18189 ;
  assign y7073 = n18190 ;
  assign y7074 = ~n18191 ;
  assign y7075 = ~n18193 ;
  assign y7076 = n18200 ;
  assign y7077 = ~n18205 ;
  assign y7078 = n18210 ;
  assign y7079 = ~n18223 ;
  assign y7080 = ~n18225 ;
  assign y7081 = ~n18226 ;
  assign y7082 = ~n18232 ;
  assign y7083 = ~n18239 ;
  assign y7084 = ~n18243 ;
  assign y7085 = ~1'b0 ;
  assign y7086 = ~1'b0 ;
  assign y7087 = ~n18248 ;
  assign y7088 = ~n18251 ;
  assign y7089 = ~n18252 ;
  assign y7090 = ~n18254 ;
  assign y7091 = ~1'b0 ;
  assign y7092 = n18255 ;
  assign y7093 = ~n18257 ;
  assign y7094 = n18258 ;
  assign y7095 = n18261 ;
  assign y7096 = n18265 ;
  assign y7097 = ~n18266 ;
  assign y7098 = n18267 ;
  assign y7099 = n18270 ;
  assign y7100 = ~n18272 ;
  assign y7101 = n18275 ;
  assign y7102 = ~1'b0 ;
  assign y7103 = n18276 ;
  assign y7104 = ~n17456 ;
  assign y7105 = ~n18278 ;
  assign y7106 = ~1'b0 ;
  assign y7107 = ~n18279 ;
  assign y7108 = n18281 ;
  assign y7109 = ~n18285 ;
  assign y7110 = n18287 ;
  assign y7111 = ~n18288 ;
  assign y7112 = n18293 ;
  assign y7113 = n18297 ;
  assign y7114 = ~n15089 ;
  assign y7115 = ~1'b0 ;
  assign y7116 = ~n18299 ;
  assign y7117 = ~n18301 ;
  assign y7118 = n18303 ;
  assign y7119 = ~1'b0 ;
  assign y7120 = ~n18306 ;
  assign y7121 = ~n18309 ;
  assign y7122 = n18311 ;
  assign y7123 = ~1'b0 ;
  assign y7124 = n18314 ;
  assign y7125 = ~n18316 ;
  assign y7126 = ~n18318 ;
  assign y7127 = ~n18319 ;
  assign y7128 = ~n18326 ;
  assign y7129 = ~n18327 ;
  assign y7130 = ~n18330 ;
  assign y7131 = n18332 ;
  assign y7132 = n18334 ;
  assign y7133 = n18335 ;
  assign y7134 = n18336 ;
  assign y7135 = n18340 ;
  assign y7136 = n18344 ;
  assign y7137 = n18347 ;
  assign y7138 = n18348 ;
  assign y7139 = ~1'b0 ;
  assign y7140 = ~n18350 ;
  assign y7141 = n18352 ;
  assign y7142 = ~n18355 ;
  assign y7143 = ~n18356 ;
  assign y7144 = ~n18357 ;
  assign y7145 = n18360 ;
  assign y7146 = n18365 ;
  assign y7147 = n18372 ;
  assign y7148 = ~n18373 ;
  assign y7149 = ~n18375 ;
  assign y7150 = ~n18382 ;
  assign y7151 = ~1'b0 ;
  assign y7152 = n18385 ;
  assign y7153 = ~1'b0 ;
  assign y7154 = n18387 ;
  assign y7155 = ~n18388 ;
  assign y7156 = ~1'b0 ;
  assign y7157 = n18392 ;
  assign y7158 = n18393 ;
  assign y7159 = n18394 ;
  assign y7160 = ~n18396 ;
  assign y7161 = n18397 ;
  assign y7162 = ~n18399 ;
  assign y7163 = n18401 ;
  assign y7164 = n18406 ;
  assign y7165 = ~n18407 ;
  assign y7166 = ~n18409 ;
  assign y7167 = ~n4937 ;
  assign y7168 = n18411 ;
  assign y7169 = ~n18413 ;
  assign y7170 = ~n18415 ;
  assign y7171 = ~n18417 ;
  assign y7172 = ~n1936 ;
  assign y7173 = n18418 ;
  assign y7174 = ~1'b0 ;
  assign y7175 = ~1'b0 ;
  assign y7176 = 1'b0 ;
  assign y7177 = n18421 ;
  assign y7178 = n18431 ;
  assign y7179 = n18435 ;
  assign y7180 = n18439 ;
  assign y7181 = ~n18440 ;
  assign y7182 = n18441 ;
  assign y7183 = n18442 ;
  assign y7184 = n18446 ;
  assign y7185 = ~n18447 ;
  assign y7186 = ~n18449 ;
  assign y7187 = n18451 ;
  assign y7188 = ~n18454 ;
  assign y7189 = ~n18456 ;
  assign y7190 = n18459 ;
  assign y7191 = ~n18463 ;
  assign y7192 = ~1'b0 ;
  assign y7193 = ~n18464 ;
  assign y7194 = ~n18467 ;
  assign y7195 = ~n18468 ;
  assign y7196 = ~1'b0 ;
  assign y7197 = ~n18471 ;
  assign y7198 = ~n18476 ;
  assign y7199 = ~n18478 ;
  assign y7200 = ~n18482 ;
  assign y7201 = ~n18483 ;
  assign y7202 = ~n18486 ;
  assign y7203 = ~1'b0 ;
  assign y7204 = n18488 ;
  assign y7205 = ~n18495 ;
  assign y7206 = n18496 ;
  assign y7207 = ~n18497 ;
  assign y7208 = n18498 ;
  assign y7209 = 1'b0 ;
  assign y7210 = ~n18499 ;
  assign y7211 = ~1'b0 ;
  assign y7212 = ~n18501 ;
  assign y7213 = ~n18504 ;
  assign y7214 = n18508 ;
  assign y7215 = n18514 ;
  assign y7216 = ~n18515 ;
  assign y7217 = ~n18516 ;
  assign y7218 = n18517 ;
  assign y7219 = ~1'b0 ;
  assign y7220 = n18522 ;
  assign y7221 = ~n18525 ;
  assign y7222 = ~n18528 ;
  assign y7223 = ~1'b0 ;
  assign y7224 = n18529 ;
  assign y7225 = 1'b0 ;
  assign y7226 = ~1'b0 ;
  assign y7227 = ~1'b0 ;
  assign y7228 = ~n18533 ;
  assign y7229 = ~1'b0 ;
  assign y7230 = ~1'b0 ;
  assign y7231 = ~1'b0 ;
  assign y7232 = n18537 ;
  assign y7233 = n18543 ;
  assign y7234 = n18545 ;
  assign y7235 = ~n18547 ;
  assign y7236 = ~n18550 ;
  assign y7237 = ~1'b0 ;
  assign y7238 = n18553 ;
  assign y7239 = ~n18554 ;
  assign y7240 = n18555 ;
  assign y7241 = n6191 ;
  assign y7242 = n18556 ;
  assign y7243 = ~1'b0 ;
  assign y7244 = n18557 ;
  assign y7245 = ~n18558 ;
  assign y7246 = ~1'b0 ;
  assign y7247 = n18562 ;
  assign y7248 = ~n18564 ;
  assign y7249 = ~n18567 ;
  assign y7250 = ~n18571 ;
  assign y7251 = n18572 ;
  assign y7252 = n18574 ;
  assign y7253 = ~n18577 ;
  assign y7254 = ~n18578 ;
  assign y7255 = n18582 ;
  assign y7256 = ~n18584 ;
  assign y7257 = 1'b0 ;
  assign y7258 = ~1'b0 ;
  assign y7259 = ~n18587 ;
  assign y7260 = ~1'b0 ;
  assign y7261 = ~n18589 ;
  assign y7262 = ~n18590 ;
  assign y7263 = ~n18591 ;
  assign y7264 = ~n18595 ;
  assign y7265 = ~1'b0 ;
  assign y7266 = n18596 ;
  assign y7267 = n18599 ;
  assign y7268 = n18601 ;
  assign y7269 = ~1'b0 ;
  assign y7270 = n18603 ;
  assign y7271 = ~1'b0 ;
  assign y7272 = ~n18606 ;
  assign y7273 = ~n18607 ;
  assign y7274 = ~n18609 ;
  assign y7275 = ~n18610 ;
  assign y7276 = ~n18614 ;
  assign y7277 = n663 ;
  assign y7278 = n18615 ;
  assign y7279 = n18616 ;
  assign y7280 = ~n18617 ;
  assign y7281 = ~n11437 ;
  assign y7282 = n18621 ;
  assign y7283 = ~n18627 ;
  assign y7284 = n18629 ;
  assign y7285 = ~1'b0 ;
  assign y7286 = ~n18630 ;
  assign y7287 = n18631 ;
  assign y7288 = n3070 ;
  assign y7289 = n18632 ;
  assign y7290 = ~n18635 ;
  assign y7291 = ~n18636 ;
  assign y7292 = ~n18638 ;
  assign y7293 = n18640 ;
  assign y7294 = ~1'b0 ;
  assign y7295 = ~n18642 ;
  assign y7296 = ~1'b0 ;
  assign y7297 = n18645 ;
  assign y7298 = n18646 ;
  assign y7299 = ~n18647 ;
  assign y7300 = ~n18652 ;
  assign y7301 = ~n18654 ;
  assign y7302 = ~1'b0 ;
  assign y7303 = ~1'b0 ;
  assign y7304 = n18661 ;
  assign y7305 = ~1'b0 ;
  assign y7306 = ~n18664 ;
  assign y7307 = ~n18665 ;
  assign y7308 = n18666 ;
  assign y7309 = ~n18668 ;
  assign y7310 = ~n18669 ;
  assign y7311 = ~n18671 ;
  assign y7312 = n18672 ;
  assign y7313 = n968 ;
  assign y7314 = n18674 ;
  assign y7315 = ~n18678 ;
  assign y7316 = n5073 ;
  assign y7317 = n18681 ;
  assign y7318 = ~n18682 ;
  assign y7319 = ~n18685 ;
  assign y7320 = n18686 ;
  assign y7321 = ~n18687 ;
  assign y7322 = ~1'b0 ;
  assign y7323 = ~n18690 ;
  assign y7324 = ~1'b0 ;
  assign y7325 = ~1'b0 ;
  assign y7326 = ~n18693 ;
  assign y7327 = n18695 ;
  assign y7328 = ~n18696 ;
  assign y7329 = n18701 ;
  assign y7330 = ~n18706 ;
  assign y7331 = n18708 ;
  assign y7332 = ~n18710 ;
  assign y7333 = ~n18712 ;
  assign y7334 = n18714 ;
  assign y7335 = n18715 ;
  assign y7336 = n18717 ;
  assign y7337 = ~n18721 ;
  assign y7338 = ~n18722 ;
  assign y7339 = n18724 ;
  assign y7340 = 1'b0 ;
  assign y7341 = ~n18727 ;
  assign y7342 = n18736 ;
  assign y7343 = ~n18738 ;
  assign y7344 = n18744 ;
  assign y7345 = ~n18747 ;
  assign y7346 = ~n18749 ;
  assign y7347 = n18750 ;
  assign y7348 = ~1'b0 ;
  assign y7349 = n18754 ;
  assign y7350 = n18757 ;
  assign y7351 = ~n18760 ;
  assign y7352 = n18761 ;
  assign y7353 = ~n18764 ;
  assign y7354 = ~1'b0 ;
  assign y7355 = ~n18765 ;
  assign y7356 = n9704 ;
  assign y7357 = ~n18768 ;
  assign y7358 = n18773 ;
  assign y7359 = ~n18775 ;
  assign y7360 = ~1'b0 ;
  assign y7361 = ~n18778 ;
  assign y7362 = ~n18785 ;
  assign y7363 = ~1'b0 ;
  assign y7364 = ~1'b0 ;
  assign y7365 = ~n18789 ;
  assign y7366 = ~1'b0 ;
  assign y7367 = n18790 ;
  assign y7368 = n18791 ;
  assign y7369 = n18792 ;
  assign y7370 = ~n18793 ;
  assign y7371 = ~n18796 ;
  assign y7372 = ~n18799 ;
  assign y7373 = ~n18800 ;
  assign y7374 = n18801 ;
  assign y7375 = n18803 ;
  assign y7376 = n18804 ;
  assign y7377 = ~n18807 ;
  assign y7378 = ~n18808 ;
  assign y7379 = n18812 ;
  assign y7380 = ~n18813 ;
  assign y7381 = n18815 ;
  assign y7382 = ~n18817 ;
  assign y7383 = n18821 ;
  assign y7384 = ~n18823 ;
  assign y7385 = ~n18825 ;
  assign y7386 = ~n18828 ;
  assign y7387 = ~1'b0 ;
  assign y7388 = n18831 ;
  assign y7389 = ~1'b0 ;
  assign y7390 = ~1'b0 ;
  assign y7391 = ~n18834 ;
  assign y7392 = n18835 ;
  assign y7393 = n18836 ;
  assign y7394 = ~n18839 ;
  assign y7395 = ~1'b0 ;
  assign y7396 = ~n18843 ;
  assign y7397 = ~n18848 ;
  assign y7398 = ~n18849 ;
  assign y7399 = n18851 ;
  assign y7400 = n18852 ;
  assign y7401 = n18853 ;
  assign y7402 = n18855 ;
  assign y7403 = ~n18857 ;
  assign y7404 = ~n18858 ;
  assign y7405 = ~n18859 ;
  assign y7406 = n18863 ;
  assign y7407 = n18867 ;
  assign y7408 = n18870 ;
  assign y7409 = ~1'b0 ;
  assign y7410 = n18873 ;
  assign y7411 = ~n18874 ;
  assign y7412 = n18880 ;
  assign y7413 = ~n18883 ;
  assign y7414 = n18885 ;
  assign y7415 = ~n18888 ;
  assign y7416 = n18895 ;
  assign y7417 = ~n18896 ;
  assign y7418 = ~n18902 ;
  assign y7419 = ~n18904 ;
  assign y7420 = n18907 ;
  assign y7421 = ~n18910 ;
  assign y7422 = n18916 ;
  assign y7423 = ~1'b0 ;
  assign y7424 = ~n18917 ;
  assign y7425 = n18918 ;
  assign y7426 = n18921 ;
  assign y7427 = ~1'b0 ;
  assign y7428 = ~1'b0 ;
  assign y7429 = n18922 ;
  assign y7430 = ~n18923 ;
  assign y7431 = ~n18929 ;
  assign y7432 = n18931 ;
  assign y7433 = ~n18934 ;
  assign y7434 = ~n18936 ;
  assign y7435 = ~n18939 ;
  assign y7436 = n18940 ;
  assign y7437 = n18946 ;
  assign y7438 = n18947 ;
  assign y7439 = n18951 ;
  assign y7440 = n18954 ;
  assign y7441 = ~1'b0 ;
  assign y7442 = ~n18955 ;
  assign y7443 = ~n18957 ;
  assign y7444 = n18959 ;
  assign y7445 = ~n18960 ;
  assign y7446 = ~n18966 ;
  assign y7447 = ~n18970 ;
  assign y7448 = ~1'b0 ;
  assign y7449 = ~1'b0 ;
  assign y7450 = ~n18971 ;
  assign y7451 = n18974 ;
  assign y7452 = n18977 ;
  assign y7453 = 1'b0 ;
  assign y7454 = ~n18979 ;
  assign y7455 = n18980 ;
  assign y7456 = ~n18982 ;
  assign y7457 = ~n18988 ;
  assign y7458 = n18995 ;
  assign y7459 = ~1'b0 ;
  assign y7460 = n18996 ;
  assign y7461 = ~1'b0 ;
  assign y7462 = ~n18998 ;
  assign y7463 = n19002 ;
  assign y7464 = n19003 ;
  assign y7465 = ~1'b0 ;
  assign y7466 = ~n19004 ;
  assign y7467 = ~n19009 ;
  assign y7468 = ~n19011 ;
  assign y7469 = ~n19015 ;
  assign y7470 = ~n19016 ;
  assign y7471 = ~n19019 ;
  assign y7472 = n19020 ;
  assign y7473 = n19023 ;
  assign y7474 = n2383 ;
  assign y7475 = n19026 ;
  assign y7476 = ~n19027 ;
  assign y7477 = n19033 ;
  assign y7478 = ~n19035 ;
  assign y7479 = ~n19036 ;
  assign y7480 = n19038 ;
  assign y7481 = n19041 ;
  assign y7482 = n19042 ;
  assign y7483 = ~n19043 ;
  assign y7484 = ~n19044 ;
  assign y7485 = n19048 ;
  assign y7486 = ~n19050 ;
  assign y7487 = ~n19055 ;
  assign y7488 = n19064 ;
  assign y7489 = ~n19065 ;
  assign y7490 = ~n19066 ;
  assign y7491 = n19069 ;
  assign y7492 = ~n19072 ;
  assign y7493 = ~1'b0 ;
  assign y7494 = n19074 ;
  assign y7495 = n19075 ;
  assign y7496 = ~n19080 ;
  assign y7497 = ~1'b0 ;
  assign y7498 = ~1'b0 ;
  assign y7499 = ~1'b0 ;
  assign y7500 = ~1'b0 ;
  assign y7501 = n19082 ;
  assign y7502 = ~n19087 ;
  assign y7503 = ~n19088 ;
  assign y7504 = n19092 ;
  assign y7505 = ~n19094 ;
  assign y7506 = ~n19096 ;
  assign y7507 = ~1'b0 ;
  assign y7508 = n19098 ;
  assign y7509 = ~n19104 ;
  assign y7510 = ~n19105 ;
  assign y7511 = ~n19109 ;
  assign y7512 = ~n19115 ;
  assign y7513 = ~1'b0 ;
  assign y7514 = n19116 ;
  assign y7515 = ~n19120 ;
  assign y7516 = ~n19121 ;
  assign y7517 = n19122 ;
  assign y7518 = n19123 ;
  assign y7519 = ~n19125 ;
  assign y7520 = ~n19126 ;
  assign y7521 = ~1'b0 ;
  assign y7522 = ~n19130 ;
  assign y7523 = ~n19134 ;
  assign y7524 = n19138 ;
  assign y7525 = n19139 ;
  assign y7526 = ~n19149 ;
  assign y7527 = ~n19155 ;
  assign y7528 = ~n19157 ;
  assign y7529 = ~n19159 ;
  assign y7530 = n5137 ;
  assign y7531 = ~n19160 ;
  assign y7532 = n19165 ;
  assign y7533 = ~1'b0 ;
  assign y7534 = ~n19166 ;
  assign y7535 = ~1'b0 ;
  assign y7536 = n19168 ;
  assign y7537 = ~n19170 ;
  assign y7538 = ~n19175 ;
  assign y7539 = ~n19178 ;
  assign y7540 = n19179 ;
  assign y7541 = ~n19182 ;
  assign y7542 = ~n19183 ;
  assign y7543 = ~1'b0 ;
  assign y7544 = n19186 ;
  assign y7545 = ~n19189 ;
  assign y7546 = n19191 ;
  assign y7547 = ~1'b0 ;
  assign y7548 = n19195 ;
  assign y7549 = n19199 ;
  assign y7550 = n19206 ;
  assign y7551 = ~n19208 ;
  assign y7552 = n19210 ;
  assign y7553 = ~1'b0 ;
  assign y7554 = ~n19213 ;
  assign y7555 = n19214 ;
  assign y7556 = ~n19216 ;
  assign y7557 = n19217 ;
  assign y7558 = ~1'b0 ;
  assign y7559 = n19218 ;
  assign y7560 = n19220 ;
  assign y7561 = ~n19223 ;
  assign y7562 = ~n19225 ;
  assign y7563 = ~n19229 ;
  assign y7564 = n19230 ;
  assign y7565 = n19233 ;
  assign y7566 = ~n19236 ;
  assign y7567 = ~1'b0 ;
  assign y7568 = ~1'b0 ;
  assign y7569 = ~1'b0 ;
  assign y7570 = 1'b0 ;
  assign y7571 = ~n19237 ;
  assign y7572 = n19239 ;
  assign y7573 = ~1'b0 ;
  assign y7574 = n19241 ;
  assign y7575 = n19245 ;
  assign y7576 = n19249 ;
  assign y7577 = n19250 ;
  assign y7578 = ~n19252 ;
  assign y7579 = n19255 ;
  assign y7580 = n19261 ;
  assign y7581 = n19264 ;
  assign y7582 = n19267 ;
  assign y7583 = n19269 ;
  assign y7584 = ~1'b0 ;
  assign y7585 = ~1'b0 ;
  assign y7586 = ~n19270 ;
  assign y7587 = n19272 ;
  assign y7588 = ~n19273 ;
  assign y7589 = ~n19274 ;
  assign y7590 = ~n19276 ;
  assign y7591 = ~n19277 ;
  assign y7592 = ~n19279 ;
  assign y7593 = 1'b0 ;
  assign y7594 = n19281 ;
  assign y7595 = ~n19282 ;
  assign y7596 = n19283 ;
  assign y7597 = ~1'b0 ;
  assign y7598 = n19285 ;
  assign y7599 = ~1'b0 ;
  assign y7600 = ~1'b0 ;
  assign y7601 = n19288 ;
  assign y7602 = ~n19290 ;
  assign y7603 = ~n19292 ;
  assign y7604 = ~1'b0 ;
  assign y7605 = ~n19295 ;
  assign y7606 = n19297 ;
  assign y7607 = ~1'b0 ;
  assign y7608 = n19307 ;
  assign y7609 = ~n19310 ;
  assign y7610 = n19316 ;
  assign y7611 = ~1'b0 ;
  assign y7612 = 1'b0 ;
  assign y7613 = ~1'b0 ;
  assign y7614 = n19323 ;
  assign y7615 = n19325 ;
  assign y7616 = ~n19327 ;
  assign y7617 = ~n19332 ;
  assign y7618 = ~1'b0 ;
  assign y7619 = ~n19334 ;
  assign y7620 = ~n19338 ;
  assign y7621 = ~n19340 ;
  assign y7622 = ~n19341 ;
  assign y7623 = n19347 ;
  assign y7624 = n19350 ;
  assign y7625 = n19351 ;
  assign y7626 = ~1'b0 ;
  assign y7627 = ~n19352 ;
  assign y7628 = ~n19355 ;
  assign y7629 = ~1'b0 ;
  assign y7630 = ~n19357 ;
  assign y7631 = n19358 ;
  assign y7632 = n19359 ;
  assign y7633 = ~n19361 ;
  assign y7634 = 1'b0 ;
  assign y7635 = ~1'b0 ;
  assign y7636 = ~n19363 ;
  assign y7637 = n19365 ;
  assign y7638 = ~1'b0 ;
  assign y7639 = n9066 ;
  assign y7640 = n19367 ;
  assign y7641 = n19374 ;
  assign y7642 = ~1'b0 ;
  assign y7643 = ~1'b0 ;
  assign y7644 = ~1'b0 ;
  assign y7645 = n19378 ;
  assign y7646 = n19383 ;
  assign y7647 = ~n19384 ;
  assign y7648 = ~n19386 ;
  assign y7649 = n19393 ;
  assign y7650 = ~n19396 ;
  assign y7651 = ~n5170 ;
  assign y7652 = n19423 ;
  assign y7653 = ~1'b0 ;
  assign y7654 = n19424 ;
  assign y7655 = ~n19426 ;
  assign y7656 = ~n19435 ;
  assign y7657 = ~1'b0 ;
  assign y7658 = n19438 ;
  assign y7659 = ~n19440 ;
  assign y7660 = ~n19442 ;
  assign y7661 = ~n19443 ;
  assign y7662 = ~1'b0 ;
  assign y7663 = n19444 ;
  assign y7664 = ~n19455 ;
  assign y7665 = n19462 ;
  assign y7666 = ~n19463 ;
  assign y7667 = n19464 ;
  assign y7668 = ~n19470 ;
  assign y7669 = n19472 ;
  assign y7670 = ~n19481 ;
  assign y7671 = n19484 ;
  assign y7672 = n19485 ;
  assign y7673 = ~1'b0 ;
  assign y7674 = n19486 ;
  assign y7675 = ~1'b0 ;
  assign y7676 = ~1'b0 ;
  assign y7677 = ~1'b0 ;
  assign y7678 = ~n19487 ;
  assign y7679 = ~1'b0 ;
  assign y7680 = n19495 ;
  assign y7681 = ~1'b0 ;
  assign y7682 = ~n19497 ;
  assign y7683 = ~n19501 ;
  assign y7684 = n19503 ;
  assign y7685 = ~1'b0 ;
  assign y7686 = ~n19504 ;
  assign y7687 = n19505 ;
  assign y7688 = n19512 ;
  assign y7689 = n19517 ;
  assign y7690 = ~1'b0 ;
  assign y7691 = ~n19518 ;
  assign y7692 = ~n19519 ;
  assign y7693 = ~1'b0 ;
  assign y7694 = ~n19521 ;
  assign y7695 = n19523 ;
  assign y7696 = ~n19526 ;
  assign y7697 = n19527 ;
  assign y7698 = n19530 ;
  assign y7699 = ~1'b0 ;
  assign y7700 = n19533 ;
  assign y7701 = ~n19538 ;
  assign y7702 = n19542 ;
  assign y7703 = ~n19548 ;
  assign y7704 = ~1'b0 ;
  assign y7705 = n9618 ;
  assign y7706 = ~1'b0 ;
  assign y7707 = n19549 ;
  assign y7708 = ~1'b0 ;
  assign y7709 = ~1'b0 ;
  assign y7710 = ~n19551 ;
  assign y7711 = n19556 ;
  assign y7712 = ~n19557 ;
  assign y7713 = n19559 ;
  assign y7714 = ~n19562 ;
  assign y7715 = ~n19568 ;
  assign y7716 = n19570 ;
  assign y7717 = ~n19574 ;
  assign y7718 = 1'b0 ;
  assign y7719 = ~n19578 ;
  assign y7720 = ~n19579 ;
  assign y7721 = ~n19580 ;
  assign y7722 = ~n19581 ;
  assign y7723 = ~n19583 ;
  assign y7724 = n19586 ;
  assign y7725 = ~n19589 ;
  assign y7726 = ~1'b0 ;
  assign y7727 = ~n19590 ;
  assign y7728 = ~n19597 ;
  assign y7729 = n19600 ;
  assign y7730 = n19604 ;
  assign y7731 = ~n19606 ;
  assign y7732 = n19610 ;
  assign y7733 = n19613 ;
  assign y7734 = n19616 ;
  assign y7735 = ~n19621 ;
  assign y7736 = ~n19628 ;
  assign y7737 = ~n19629 ;
  assign y7738 = ~n19630 ;
  assign y7739 = ~1'b0 ;
  assign y7740 = n19632 ;
  assign y7741 = ~n19638 ;
  assign y7742 = ~n19639 ;
  assign y7743 = n19640 ;
  assign y7744 = ~1'b0 ;
  assign y7745 = ~n19643 ;
  assign y7746 = ~1'b0 ;
  assign y7747 = ~n19649 ;
  assign y7748 = n19651 ;
  assign y7749 = ~n19657 ;
  assign y7750 = ~1'b0 ;
  assign y7751 = ~n19658 ;
  assign y7752 = n19659 ;
  assign y7753 = ~1'b0 ;
  assign y7754 = ~n19661 ;
  assign y7755 = ~1'b0 ;
  assign y7756 = ~n19666 ;
  assign y7757 = ~1'b0 ;
  assign y7758 = ~n19672 ;
  assign y7759 = n19674 ;
  assign y7760 = n19676 ;
  assign y7761 = n19677 ;
  assign y7762 = ~n19681 ;
  assign y7763 = n19684 ;
  assign y7764 = ~1'b0 ;
  assign y7765 = ~n19688 ;
  assign y7766 = n19690 ;
  assign y7767 = ~1'b0 ;
  assign y7768 = n19692 ;
  assign y7769 = n6675 ;
  assign y7770 = n19700 ;
  assign y7771 = ~n19701 ;
  assign y7772 = ~n19705 ;
  assign y7773 = ~1'b0 ;
  assign y7774 = ~n19707 ;
  assign y7775 = ~1'b0 ;
  assign y7776 = ~1'b0 ;
  assign y7777 = ~n19710 ;
  assign y7778 = ~n19712 ;
  assign y7779 = n19713 ;
  assign y7780 = ~n19714 ;
  assign y7781 = ~n5123 ;
  assign y7782 = ~n19718 ;
  assign y7783 = ~1'b0 ;
  assign y7784 = ~1'b0 ;
  assign y7785 = ~1'b0 ;
  assign y7786 = ~1'b0 ;
  assign y7787 = ~n6370 ;
  assign y7788 = n19722 ;
  assign y7789 = n19725 ;
  assign y7790 = ~n13716 ;
  assign y7791 = ~1'b0 ;
  assign y7792 = n19728 ;
  assign y7793 = ~n9791 ;
  assign y7794 = ~n14824 ;
  assign y7795 = ~n19729 ;
  assign y7796 = ~n19730 ;
  assign y7797 = ~1'b0 ;
  assign y7798 = ~1'b0 ;
  assign y7799 = ~n19732 ;
  assign y7800 = ~1'b0 ;
  assign y7801 = ~n19733 ;
  assign y7802 = ~1'b0 ;
  assign y7803 = ~n19736 ;
  assign y7804 = ~n19737 ;
  assign y7805 = ~n19741 ;
  assign y7806 = n19743 ;
  assign y7807 = ~n19744 ;
  assign y7808 = n19746 ;
  assign y7809 = ~n19748 ;
  assign y7810 = n19750 ;
  assign y7811 = ~n19751 ;
  assign y7812 = ~1'b0 ;
  assign y7813 = n19753 ;
  assign y7814 = ~1'b0 ;
  assign y7815 = ~n6421 ;
  assign y7816 = ~1'b0 ;
  assign y7817 = n19758 ;
  assign y7818 = n19764 ;
  assign y7819 = ~n19768 ;
  assign y7820 = ~n19769 ;
  assign y7821 = ~1'b0 ;
  assign y7822 = ~1'b0 ;
  assign y7823 = ~n19772 ;
  assign y7824 = n19777 ;
  assign y7825 = ~1'b0 ;
  assign y7826 = ~1'b0 ;
  assign y7827 = n19780 ;
  assign y7828 = ~n19784 ;
  assign y7829 = ~n19785 ;
  assign y7830 = ~1'b0 ;
  assign y7831 = ~1'b0 ;
  assign y7832 = ~1'b0 ;
  assign y7833 = ~n19788 ;
  assign y7834 = ~1'b0 ;
  assign y7835 = n19791 ;
  assign y7836 = n19793 ;
  assign y7837 = ~n19797 ;
  assign y7838 = n19799 ;
  assign y7839 = ~n19803 ;
  assign y7840 = ~1'b0 ;
  assign y7841 = ~1'b0 ;
  assign y7842 = n19804 ;
  assign y7843 = ~1'b0 ;
  assign y7844 = n19808 ;
  assign y7845 = ~n19362 ;
  assign y7846 = ~1'b0 ;
  assign y7847 = ~1'b0 ;
  assign y7848 = n19809 ;
  assign y7849 = n19811 ;
  assign y7850 = n19817 ;
  assign y7851 = ~1'b0 ;
  assign y7852 = ~n19818 ;
  assign y7853 = n19822 ;
  assign y7854 = n19828 ;
  assign y7855 = ~n19829 ;
  assign y7856 = n19832 ;
  assign y7857 = ~n8286 ;
  assign y7858 = ~n19836 ;
  assign y7859 = n16355 ;
  assign y7860 = ~n19840 ;
  assign y7861 = ~n19841 ;
  assign y7862 = n19845 ;
  assign y7863 = ~n19848 ;
  assign y7864 = ~1'b0 ;
  assign y7865 = ~1'b0 ;
  assign y7866 = ~1'b0 ;
  assign y7867 = ~1'b0 ;
  assign y7868 = ~n19856 ;
  assign y7869 = n19857 ;
  assign y7870 = n19859 ;
  assign y7871 = 1'b0 ;
  assign y7872 = ~1'b0 ;
  assign y7873 = ~1'b0 ;
  assign y7874 = n19862 ;
  assign y7875 = ~n19865 ;
  assign y7876 = ~n19869 ;
  assign y7877 = ~n19871 ;
  assign y7878 = n11811 ;
  assign y7879 = ~n19872 ;
  assign y7880 = n19873 ;
  assign y7881 = n19877 ;
  assign y7882 = ~n19879 ;
  assign y7883 = n19884 ;
  assign y7884 = ~n19890 ;
  assign y7885 = n19893 ;
  assign y7886 = n19894 ;
  assign y7887 = ~1'b0 ;
  assign y7888 = n19895 ;
  assign y7889 = n19897 ;
  assign y7890 = ~n19898 ;
  assign y7891 = ~n19899 ;
  assign y7892 = ~n19901 ;
  assign y7893 = ~n19902 ;
  assign y7894 = n19910 ;
  assign y7895 = ~n19913 ;
  assign y7896 = n19916 ;
  assign y7897 = ~1'b0 ;
  assign y7898 = ~1'b0 ;
  assign y7899 = ~1'b0 ;
  assign y7900 = ~n19919 ;
  assign y7901 = ~n10372 ;
  assign y7902 = n19922 ;
  assign y7903 = ~n19924 ;
  assign y7904 = n19928 ;
  assign y7905 = ~1'b0 ;
  assign y7906 = n19936 ;
  assign y7907 = ~n19940 ;
  assign y7908 = n19941 ;
  assign y7909 = ~n19945 ;
  assign y7910 = n19948 ;
  assign y7911 = ~n19950 ;
  assign y7912 = ~n19955 ;
  assign y7913 = ~n19956 ;
  assign y7914 = n19957 ;
  assign y7915 = ~1'b0 ;
  assign y7916 = n19960 ;
  assign y7917 = n19962 ;
  assign y7918 = ~n19964 ;
  assign y7919 = n19965 ;
  assign y7920 = n19968 ;
  assign y7921 = n19972 ;
  assign y7922 = n19975 ;
  assign y7923 = n19977 ;
  assign y7924 = n19983 ;
  assign y7925 = ~1'b0 ;
  assign y7926 = n19984 ;
  assign y7927 = n19986 ;
  assign y7928 = n19988 ;
  assign y7929 = ~n19990 ;
  assign y7930 = ~1'b0 ;
  assign y7931 = ~n20006 ;
  assign y7932 = n20008 ;
  assign y7933 = n20012 ;
  assign y7934 = n20013 ;
  assign y7935 = ~n20015 ;
  assign y7936 = ~1'b0 ;
  assign y7937 = ~n20018 ;
  assign y7938 = n20019 ;
  assign y7939 = ~n20020 ;
  assign y7940 = ~1'b0 ;
  assign y7941 = n20025 ;
  assign y7942 = n20026 ;
  assign y7943 = ~n20028 ;
  assign y7944 = 1'b0 ;
  assign y7945 = n20030 ;
  assign y7946 = ~1'b0 ;
  assign y7947 = n20033 ;
  assign y7948 = n20036 ;
  assign y7949 = ~n20040 ;
  assign y7950 = ~1'b0 ;
  assign y7951 = n20041 ;
  assign y7952 = ~1'b0 ;
  assign y7953 = ~n20042 ;
  assign y7954 = ~1'b0 ;
  assign y7955 = n20046 ;
  assign y7956 = ~n20049 ;
  assign y7957 = n20050 ;
  assign y7958 = ~n20053 ;
  assign y7959 = ~n20056 ;
  assign y7960 = ~1'b0 ;
  assign y7961 = n20058 ;
  assign y7962 = n20060 ;
  assign y7963 = ~n20061 ;
  assign y7964 = ~n20063 ;
  assign y7965 = ~n9458 ;
  assign y7966 = n20065 ;
  assign y7967 = ~n20066 ;
  assign y7968 = n20068 ;
  assign y7969 = ~n20069 ;
  assign y7970 = ~n20071 ;
  assign y7971 = ~1'b0 ;
  assign y7972 = ~n20073 ;
  assign y7973 = ~n20074 ;
  assign y7974 = ~n20075 ;
  assign y7975 = ~n20077 ;
  assign y7976 = ~n20078 ;
  assign y7977 = ~n20085 ;
  assign y7978 = n20087 ;
  assign y7979 = ~1'b0 ;
  assign y7980 = n20089 ;
  assign y7981 = ~1'b0 ;
  assign y7982 = n20090 ;
  assign y7983 = ~n20092 ;
  assign y7984 = n20101 ;
  assign y7985 = ~n20107 ;
  assign y7986 = ~n11596 ;
  assign y7987 = ~1'b0 ;
  assign y7988 = n20110 ;
  assign y7989 = ~n20115 ;
  assign y7990 = n20120 ;
  assign y7991 = ~1'b0 ;
  assign y7992 = n20121 ;
  assign y7993 = n20122 ;
  assign y7994 = n20125 ;
  assign y7995 = n20126 ;
  assign y7996 = n20127 ;
  assign y7997 = ~n20129 ;
  assign y7998 = n20131 ;
  assign y7999 = ~n545 ;
  assign y8000 = ~n20132 ;
  assign y8001 = n20133 ;
  assign y8002 = ~n20134 ;
  assign y8003 = ~n20142 ;
  assign y8004 = ~1'b0 ;
  assign y8005 = ~1'b0 ;
  assign y8006 = ~n20143 ;
  assign y8007 = ~n20144 ;
  assign y8008 = ~1'b0 ;
  assign y8009 = n20145 ;
  assign y8010 = ~1'b0 ;
  assign y8011 = ~n20147 ;
  assign y8012 = n20149 ;
  assign y8013 = ~n20150 ;
  assign y8014 = ~n20153 ;
  assign y8015 = n20154 ;
  assign y8016 = n20156 ;
  assign y8017 = ~1'b0 ;
  assign y8018 = n20157 ;
  assign y8019 = ~n20159 ;
  assign y8020 = ~n20160 ;
  assign y8021 = ~n20163 ;
  assign y8022 = n20165 ;
  assign y8023 = ~1'b0 ;
  assign y8024 = n20166 ;
  assign y8025 = n20171 ;
  assign y8026 = ~1'b0 ;
  assign y8027 = ~1'b0 ;
  assign y8028 = ~n20174 ;
  assign y8029 = n20179 ;
  assign y8030 = n20186 ;
  assign y8031 = n20188 ;
  assign y8032 = n20194 ;
  assign y8033 = ~n20199 ;
  assign y8034 = ~n20203 ;
  assign y8035 = ~n20207 ;
  assign y8036 = n20212 ;
  assign y8037 = ~n20213 ;
  assign y8038 = n20215 ;
  assign y8039 = ~n20220 ;
  assign y8040 = ~n20222 ;
  assign y8041 = n20225 ;
  assign y8042 = n20227 ;
  assign y8043 = n20234 ;
  assign y8044 = ~n20238 ;
  assign y8045 = ~1'b0 ;
  assign y8046 = ~1'b0 ;
  assign y8047 = ~n20242 ;
  assign y8048 = ~1'b0 ;
  assign y8049 = ~n20244 ;
  assign y8050 = ~n20245 ;
  assign y8051 = n20248 ;
  assign y8052 = ~n5513 ;
  assign y8053 = ~1'b0 ;
  assign y8054 = ~n20250 ;
  assign y8055 = ~n20254 ;
  assign y8056 = ~n18598 ;
  assign y8057 = n20257 ;
  assign y8058 = ~n20261 ;
  assign y8059 = ~n20263 ;
  assign y8060 = ~1'b0 ;
  assign y8061 = ~n20265 ;
  assign y8062 = ~1'b0 ;
  assign y8063 = ~n791 ;
  assign y8064 = n20266 ;
  assign y8065 = n20269 ;
  assign y8066 = n20273 ;
  assign y8067 = ~n20277 ;
  assign y8068 = ~n20281 ;
  assign y8069 = ~n20283 ;
  assign y8070 = n20286 ;
  assign y8071 = n20287 ;
  assign y8072 = ~n20289 ;
  assign y8073 = ~n20292 ;
  assign y8074 = ~n20295 ;
  assign y8075 = ~1'b0 ;
  assign y8076 = ~n20298 ;
  assign y8077 = n20304 ;
  assign y8078 = ~n20309 ;
  assign y8079 = ~1'b0 ;
  assign y8080 = ~1'b0 ;
  assign y8081 = n20312 ;
  assign y8082 = n20315 ;
  assign y8083 = ~n11103 ;
  assign y8084 = ~n20316 ;
  assign y8085 = ~n20317 ;
  assign y8086 = n20321 ;
  assign y8087 = n20322 ;
  assign y8088 = ~1'b0 ;
  assign y8089 = 1'b0 ;
  assign y8090 = ~n20324 ;
  assign y8091 = n2520 ;
  assign y8092 = n20326 ;
  assign y8093 = n20327 ;
  assign y8094 = ~n20328 ;
  assign y8095 = ~1'b0 ;
  assign y8096 = ~1'b0 ;
  assign y8097 = n20332 ;
  assign y8098 = n20337 ;
  assign y8099 = ~n20342 ;
  assign y8100 = ~1'b0 ;
  assign y8101 = n20344 ;
  assign y8102 = ~n20347 ;
  assign y8103 = ~1'b0 ;
  assign y8104 = n20348 ;
  assign y8105 = n20349 ;
  assign y8106 = ~1'b0 ;
  assign y8107 = ~n20354 ;
  assign y8108 = n20355 ;
  assign y8109 = ~n20357 ;
  assign y8110 = n20358 ;
  assign y8111 = n20369 ;
  assign y8112 = ~n20370 ;
  assign y8113 = n20374 ;
  assign y8114 = ~n20377 ;
  assign y8115 = ~n20378 ;
  assign y8116 = n20379 ;
  assign y8117 = n20384 ;
  assign y8118 = ~n20387 ;
  assign y8119 = ~1'b0 ;
  assign y8120 = ~n20390 ;
  assign y8121 = n20391 ;
  assign y8122 = ~n20394 ;
  assign y8123 = ~n20395 ;
  assign y8124 = n20400 ;
  assign y8125 = ~n20401 ;
  assign y8126 = ~n20403 ;
  assign y8127 = n20406 ;
  assign y8128 = ~n20407 ;
  assign y8129 = n20408 ;
  assign y8130 = ~n20411 ;
  assign y8131 = ~n20414 ;
  assign y8132 = n20418 ;
  assign y8133 = ~n20422 ;
  assign y8134 = ~1'b0 ;
  assign y8135 = ~1'b0 ;
  assign y8136 = ~n20426 ;
  assign y8137 = ~1'b0 ;
  assign y8138 = ~n20428 ;
  assign y8139 = n20429 ;
  assign y8140 = ~n20430 ;
  assign y8141 = ~1'b0 ;
  assign y8142 = ~n20433 ;
  assign y8143 = n20436 ;
  assign y8144 = n20437 ;
  assign y8145 = ~n20438 ;
  assign y8146 = ~1'b0 ;
  assign y8147 = ~1'b0 ;
  assign y8148 = n20442 ;
  assign y8149 = ~1'b0 ;
  assign y8150 = ~1'b0 ;
  assign y8151 = ~n20447 ;
  assign y8152 = n20456 ;
  assign y8153 = ~n20459 ;
  assign y8154 = ~n20461 ;
  assign y8155 = ~n20464 ;
  assign y8156 = ~1'b0 ;
  assign y8157 = ~n20466 ;
  assign y8158 = n20475 ;
  assign y8159 = n20477 ;
  assign y8160 = ~n20478 ;
  assign y8161 = n20479 ;
  assign y8162 = ~1'b0 ;
  assign y8163 = ~n20488 ;
  assign y8164 = ~n20491 ;
  assign y8165 = n20493 ;
  assign y8166 = ~1'b0 ;
  assign y8167 = ~1'b0 ;
  assign y8168 = ~1'b0 ;
  assign y8169 = n20494 ;
  assign y8170 = ~n20496 ;
  assign y8171 = ~1'b0 ;
  assign y8172 = ~n20499 ;
  assign y8173 = n20504 ;
  assign y8174 = ~n20505 ;
  assign y8175 = ~n20507 ;
  assign y8176 = n20517 ;
  assign y8177 = ~1'b0 ;
  assign y8178 = ~1'b0 ;
  assign y8179 = ~1'b0 ;
  assign y8180 = n20519 ;
  assign y8181 = ~n20521 ;
  assign y8182 = ~n20524 ;
  assign y8183 = ~n20528 ;
  assign y8184 = ~n20529 ;
  assign y8185 = n20531 ;
  assign y8186 = ~n20538 ;
  assign y8187 = ~n20543 ;
  assign y8188 = ~n20547 ;
  assign y8189 = n20550 ;
  assign y8190 = ~1'b0 ;
  assign y8191 = ~1'b0 ;
  assign y8192 = ~1'b0 ;
  assign y8193 = ~n20554 ;
  assign y8194 = ~n20557 ;
  assign y8195 = ~1'b0 ;
  assign y8196 = ~n20559 ;
  assign y8197 = ~n20561 ;
  assign y8198 = ~n20562 ;
  assign y8199 = n20566 ;
  assign y8200 = ~1'b0 ;
  assign y8201 = n20574 ;
  assign y8202 = ~n20579 ;
  assign y8203 = n20580 ;
  assign y8204 = ~n20584 ;
  assign y8205 = ~n20586 ;
  assign y8206 = ~n20589 ;
  assign y8207 = ~n20590 ;
  assign y8208 = n20591 ;
  assign y8209 = n20597 ;
  assign y8210 = ~n20600 ;
  assign y8211 = n20601 ;
  assign y8212 = ~1'b0 ;
  assign y8213 = ~n20605 ;
  assign y8214 = n20607 ;
  assign y8215 = n20615 ;
  assign y8216 = ~1'b0 ;
  assign y8217 = n20617 ;
  assign y8218 = ~n20619 ;
  assign y8219 = n20621 ;
  assign y8220 = ~n20622 ;
  assign y8221 = n20624 ;
  assign y8222 = n20626 ;
  assign y8223 = n6744 ;
  assign y8224 = n20627 ;
  assign y8225 = n20629 ;
  assign y8226 = n20630 ;
  assign y8227 = 1'b0 ;
  assign y8228 = n20632 ;
  assign y8229 = n20634 ;
  assign y8230 = n20635 ;
  assign y8231 = ~n20637 ;
  assign y8232 = ~n20638 ;
  assign y8233 = n20642 ;
  assign y8234 = 1'b0 ;
  assign y8235 = ~1'b0 ;
  assign y8236 = ~n20648 ;
  assign y8237 = ~n20652 ;
  assign y8238 = n20654 ;
  assign y8239 = ~n20657 ;
  assign y8240 = ~1'b0 ;
  assign y8241 = ~n20658 ;
  assign y8242 = ~n20659 ;
  assign y8243 = n20660 ;
  assign y8244 = ~n20666 ;
  assign y8245 = ~1'b0 ;
  assign y8246 = n20673 ;
  assign y8247 = ~n20678 ;
  assign y8248 = ~1'b0 ;
  assign y8249 = 1'b0 ;
  assign y8250 = n20679 ;
  assign y8251 = n20684 ;
  assign y8252 = n20685 ;
  assign y8253 = ~n20686 ;
  assign y8254 = n20687 ;
  assign y8255 = n20689 ;
  assign y8256 = ~1'b0 ;
  assign y8257 = ~n20695 ;
  assign y8258 = ~n20697 ;
  assign y8259 = n15673 ;
  assign y8260 = n20701 ;
  assign y8261 = ~n20705 ;
  assign y8262 = ~n20707 ;
  assign y8263 = ~n20708 ;
  assign y8264 = n20709 ;
  assign y8265 = ~n20713 ;
  assign y8266 = ~1'b0 ;
  assign y8267 = ~n20715 ;
  assign y8268 = n20716 ;
  assign y8269 = ~1'b0 ;
  assign y8270 = n20725 ;
  assign y8271 = ~n20726 ;
  assign y8272 = n20728 ;
  assign y8273 = ~n20730 ;
  assign y8274 = n20734 ;
  assign y8275 = ~n20736 ;
  assign y8276 = n20741 ;
  assign y8277 = ~n20743 ;
  assign y8278 = n20744 ;
  assign y8279 = n20747 ;
  assign y8280 = ~n20748 ;
  assign y8281 = ~1'b0 ;
  assign y8282 = ~n20751 ;
  assign y8283 = ~1'b0 ;
  assign y8284 = n20755 ;
  assign y8285 = ~1'b0 ;
  assign y8286 = ~1'b0 ;
  assign y8287 = n20756 ;
  assign y8288 = n20763 ;
  assign y8289 = ~1'b0 ;
  assign y8290 = ~1'b0 ;
  assign y8291 = ~n20765 ;
  assign y8292 = ~1'b0 ;
  assign y8293 = ~n20770 ;
  assign y8294 = n20771 ;
  assign y8295 = n20776 ;
  assign y8296 = ~1'b0 ;
  assign y8297 = ~n20779 ;
  assign y8298 = ~1'b0 ;
  assign y8299 = ~n20780 ;
  assign y8300 = ~n20783 ;
  assign y8301 = n20784 ;
  assign y8302 = ~n20786 ;
  assign y8303 = ~n20790 ;
  assign y8304 = ~n20792 ;
  assign y8305 = n20794 ;
  assign y8306 = ~1'b0 ;
  assign y8307 = ~n4510 ;
  assign y8308 = ~1'b0 ;
  assign y8309 = ~n20797 ;
  assign y8310 = ~n20800 ;
  assign y8311 = ~1'b0 ;
  assign y8312 = n20802 ;
  assign y8313 = n20804 ;
  assign y8314 = n20806 ;
  assign y8315 = ~n20808 ;
  assign y8316 = ~n20811 ;
  assign y8317 = n20812 ;
  assign y8318 = ~n20817 ;
  assign y8319 = n20822 ;
  assign y8320 = n20825 ;
  assign y8321 = n20829 ;
  assign y8322 = ~1'b0 ;
  assign y8323 = ~1'b0 ;
  assign y8324 = ~n20830 ;
  assign y8325 = 1'b0 ;
  assign y8326 = ~n20832 ;
  assign y8327 = ~1'b0 ;
  assign y8328 = ~n20835 ;
  assign y8329 = n20841 ;
  assign y8330 = n20845 ;
  assign y8331 = n20848 ;
  assign y8332 = n20853 ;
  assign y8333 = n20855 ;
  assign y8334 = ~n20857 ;
  assign y8335 = n20859 ;
  assign y8336 = ~n20864 ;
  assign y8337 = ~1'b0 ;
  assign y8338 = ~1'b0 ;
  assign y8339 = ~n20870 ;
  assign y8340 = n20872 ;
  assign y8341 = n20875 ;
  assign y8342 = ~n20876 ;
  assign y8343 = ~1'b0 ;
  assign y8344 = n20880 ;
  assign y8345 = n20882 ;
  assign y8346 = ~1'b0 ;
  assign y8347 = n20888 ;
  assign y8348 = ~n20892 ;
  assign y8349 = n20893 ;
  assign y8350 = ~1'b0 ;
  assign y8351 = ~n20895 ;
  assign y8352 = ~n20897 ;
  assign y8353 = ~n20898 ;
  assign y8354 = n20900 ;
  assign y8355 = ~n20901 ;
  assign y8356 = n20902 ;
  assign y8357 = ~n20903 ;
  assign y8358 = ~n10186 ;
  assign y8359 = ~n20905 ;
  assign y8360 = ~n20906 ;
  assign y8361 = ~1'b0 ;
  assign y8362 = n20908 ;
  assign y8363 = ~n20910 ;
  assign y8364 = n20916 ;
  assign y8365 = ~n20917 ;
  assign y8366 = ~1'b0 ;
  assign y8367 = n20921 ;
  assign y8368 = n20922 ;
  assign y8369 = ~n20924 ;
  assign y8370 = ~n20925 ;
  assign y8371 = n20927 ;
  assign y8372 = ~n20928 ;
  assign y8373 = ~n20929 ;
  assign y8374 = n20931 ;
  assign y8375 = ~1'b0 ;
  assign y8376 = ~n4628 ;
  assign y8377 = ~1'b0 ;
  assign y8378 = n20932 ;
  assign y8379 = n5135 ;
  assign y8380 = ~n20933 ;
  assign y8381 = n20935 ;
  assign y8382 = n20941 ;
  assign y8383 = ~1'b0 ;
  assign y8384 = ~1'b0 ;
  assign y8385 = n20945 ;
  assign y8386 = n20947 ;
  assign y8387 = n20951 ;
  assign y8388 = ~1'b0 ;
  assign y8389 = n20952 ;
  assign y8390 = n20959 ;
  assign y8391 = n20960 ;
  assign y8392 = n20963 ;
  assign y8393 = n20964 ;
  assign y8394 = ~n20967 ;
  assign y8395 = n20972 ;
  assign y8396 = ~n20974 ;
  assign y8397 = ~n20975 ;
  assign y8398 = ~n20978 ;
  assign y8399 = ~1'b0 ;
  assign y8400 = ~1'b0 ;
  assign y8401 = ~n20983 ;
  assign y8402 = n20984 ;
  assign y8403 = n20988 ;
  assign y8404 = ~1'b0 ;
  assign y8405 = n20993 ;
  assign y8406 = ~n20996 ;
  assign y8407 = n20998 ;
  assign y8408 = ~n3274 ;
  assign y8409 = ~n21001 ;
  assign y8410 = ~n21004 ;
  assign y8411 = ~n21008 ;
  assign y8412 = n21015 ;
  assign y8413 = n21018 ;
  assign y8414 = ~n21030 ;
  assign y8415 = n21031 ;
  assign y8416 = n21033 ;
  assign y8417 = n21036 ;
  assign y8418 = ~n21038 ;
  assign y8419 = ~1'b0 ;
  assign y8420 = ~1'b0 ;
  assign y8421 = ~1'b0 ;
  assign y8422 = n21040 ;
  assign y8423 = n21043 ;
  assign y8424 = n21044 ;
  assign y8425 = n21046 ;
  assign y8426 = n21049 ;
  assign y8427 = n21051 ;
  assign y8428 = ~n21059 ;
  assign y8429 = ~n21062 ;
  assign y8430 = ~n21066 ;
  assign y8431 = n21071 ;
  assign y8432 = ~n21072 ;
  assign y8433 = n21073 ;
  assign y8434 = ~1'b0 ;
  assign y8435 = ~n21075 ;
  assign y8436 = ~n21078 ;
  assign y8437 = ~n21082 ;
  assign y8438 = n21084 ;
  assign y8439 = n7428 ;
  assign y8440 = 1'b0 ;
  assign y8441 = n21087 ;
  assign y8442 = ~1'b0 ;
  assign y8443 = n21090 ;
  assign y8444 = n21093 ;
  assign y8445 = ~n16482 ;
  assign y8446 = ~n21098 ;
  assign y8447 = ~n21103 ;
  assign y8448 = ~1'b0 ;
  assign y8449 = n21104 ;
  assign y8450 = ~n6583 ;
  assign y8451 = n21107 ;
  assign y8452 = ~n21108 ;
  assign y8453 = n21110 ;
  assign y8454 = ~1'b0 ;
  assign y8455 = n21117 ;
  assign y8456 = ~1'b0 ;
  assign y8457 = n21118 ;
  assign y8458 = n21120 ;
  assign y8459 = n21121 ;
  assign y8460 = n21122 ;
  assign y8461 = ~1'b0 ;
  assign y8462 = ~1'b0 ;
  assign y8463 = n21125 ;
  assign y8464 = ~n21129 ;
  assign y8465 = ~n21132 ;
  assign y8466 = n21133 ;
  assign y8467 = ~1'b0 ;
  assign y8468 = n21135 ;
  assign y8469 = n21136 ;
  assign y8470 = n21138 ;
  assign y8471 = n21140 ;
  assign y8472 = ~n21143 ;
  assign y8473 = ~n21144 ;
  assign y8474 = ~1'b0 ;
  assign y8475 = n21145 ;
  assign y8476 = n21146 ;
  assign y8477 = n21147 ;
  assign y8478 = n21149 ;
  assign y8479 = ~n21150 ;
  assign y8480 = ~n21151 ;
  assign y8481 = ~1'b0 ;
  assign y8482 = 1'b0 ;
  assign y8483 = n21152 ;
  assign y8484 = ~n21154 ;
  assign y8485 = ~n21157 ;
  assign y8486 = ~n21158 ;
  assign y8487 = ~n21159 ;
  assign y8488 = n21161 ;
  assign y8489 = ~n21162 ;
  assign y8490 = ~n21164 ;
  assign y8491 = ~n21167 ;
  assign y8492 = ~n21168 ;
  assign y8493 = ~n21169 ;
  assign y8494 = ~n21171 ;
  assign y8495 = n21172 ;
  assign y8496 = n21174 ;
  assign y8497 = n21175 ;
  assign y8498 = ~1'b0 ;
  assign y8499 = ~n21177 ;
  assign y8500 = ~1'b0 ;
  assign y8501 = ~n21179 ;
  assign y8502 = ~n21180 ;
  assign y8503 = n21186 ;
  assign y8504 = n21190 ;
  assign y8505 = ~1'b0 ;
  assign y8506 = ~n21193 ;
  assign y8507 = ~n21200 ;
  assign y8508 = ~1'b0 ;
  assign y8509 = ~1'b0 ;
  assign y8510 = n21202 ;
  assign y8511 = ~n21204 ;
  assign y8512 = ~n21207 ;
  assign y8513 = n21208 ;
  assign y8514 = ~1'b0 ;
  assign y8515 = n21209 ;
  assign y8516 = n21212 ;
  assign y8517 = ~1'b0 ;
  assign y8518 = ~n21213 ;
  assign y8519 = ~n21217 ;
  assign y8520 = n15478 ;
  assign y8521 = ~1'b0 ;
  assign y8522 = ~1'b0 ;
  assign y8523 = ~n21220 ;
  assign y8524 = ~n21222 ;
  assign y8525 = ~n21223 ;
  assign y8526 = n21225 ;
  assign y8527 = ~n21226 ;
  assign y8528 = n21228 ;
  assign y8529 = ~n13203 ;
  assign y8530 = ~n21229 ;
  assign y8531 = ~n21230 ;
  assign y8532 = ~n21231 ;
  assign y8533 = n21235 ;
  assign y8534 = n21240 ;
  assign y8535 = ~1'b0 ;
  assign y8536 = ~1'b0 ;
  assign y8537 = n21242 ;
  assign y8538 = ~n21243 ;
  assign y8539 = ~n21248 ;
  assign y8540 = ~n21251 ;
  assign y8541 = ~n17730 ;
  assign y8542 = n13334 ;
  assign y8543 = 1'b0 ;
  assign y8544 = ~n21255 ;
  assign y8545 = ~n21260 ;
  assign y8546 = ~n21262 ;
  assign y8547 = ~n21266 ;
  assign y8548 = ~n21269 ;
  assign y8549 = ~n21274 ;
  assign y8550 = n21277 ;
  assign y8551 = ~1'b0 ;
  assign y8552 = ~n21279 ;
  assign y8553 = ~n21282 ;
  assign y8554 = n21285 ;
  assign y8555 = ~n21290 ;
  assign y8556 = n21294 ;
  assign y8557 = n21300 ;
  assign y8558 = ~n21306 ;
  assign y8559 = ~1'b0 ;
  assign y8560 = ~n21314 ;
  assign y8561 = n21316 ;
  assign y8562 = n21319 ;
  assign y8563 = ~1'b0 ;
  assign y8564 = ~1'b0 ;
  assign y8565 = n21324 ;
  assign y8566 = n21326 ;
  assign y8567 = n21329 ;
  assign y8568 = ~1'b0 ;
  assign y8569 = ~1'b0 ;
  assign y8570 = n21330 ;
  assign y8571 = n21334 ;
  assign y8572 = ~n21335 ;
  assign y8573 = ~n21336 ;
  assign y8574 = n21338 ;
  assign y8575 = n21340 ;
  assign y8576 = ~n21342 ;
  assign y8577 = ~1'b0 ;
  assign y8578 = ~n21344 ;
  assign y8579 = ~1'b0 ;
  assign y8580 = n21346 ;
  assign y8581 = n21349 ;
  assign y8582 = ~n21351 ;
  assign y8583 = n21353 ;
  assign y8584 = ~n21356 ;
  assign y8585 = ~n4310 ;
  assign y8586 = ~n21359 ;
  assign y8587 = ~1'b0 ;
  assign y8588 = ~n21360 ;
  assign y8589 = ~n21362 ;
  assign y8590 = n21363 ;
  assign y8591 = n21364 ;
  assign y8592 = ~n21365 ;
  assign y8593 = n21366 ;
  assign y8594 = n21371 ;
  assign y8595 = ~1'b0 ;
  assign y8596 = ~1'b0 ;
  assign y8597 = n21372 ;
  assign y8598 = ~n21380 ;
  assign y8599 = n21381 ;
  assign y8600 = n21384 ;
  assign y8601 = n21389 ;
  assign y8602 = ~1'b0 ;
  assign y8603 = ~1'b0 ;
  assign y8604 = ~n21390 ;
  assign y8605 = n21391 ;
  assign y8606 = n21393 ;
  assign y8607 = ~n21396 ;
  assign y8608 = ~n19828 ;
  assign y8609 = n21397 ;
  assign y8610 = ~x39 ;
  assign y8611 = ~n21398 ;
  assign y8612 = ~n21399 ;
  assign y8613 = n21401 ;
  assign y8614 = n21404 ;
  assign y8615 = n21409 ;
  assign y8616 = ~1'b0 ;
  assign y8617 = ~n21410 ;
  assign y8618 = n21411 ;
  assign y8619 = n9940 ;
  assign y8620 = ~1'b0 ;
  assign y8621 = ~n21414 ;
  assign y8622 = n21416 ;
  assign y8623 = ~1'b0 ;
  assign y8624 = ~n21417 ;
  assign y8625 = ~n21418 ;
  assign y8626 = n21425 ;
  assign y8627 = n21427 ;
  assign y8628 = n21429 ;
  assign y8629 = n21431 ;
  assign y8630 = n21434 ;
  assign y8631 = ~1'b0 ;
  assign y8632 = n21435 ;
  assign y8633 = ~1'b0 ;
  assign y8634 = n21438 ;
  assign y8635 = n21440 ;
  assign y8636 = 1'b0 ;
  assign y8637 = ~n21442 ;
  assign y8638 = ~n21450 ;
  assign y8639 = ~n21451 ;
  assign y8640 = n21453 ;
  assign y8641 = ~1'b0 ;
  assign y8642 = n21457 ;
  assign y8643 = ~n21461 ;
  assign y8644 = ~n21466 ;
  assign y8645 = ~n21474 ;
  assign y8646 = ~1'b0 ;
  assign y8647 = ~n21478 ;
  assign y8648 = n21481 ;
  assign y8649 = n21482 ;
  assign y8650 = n21488 ;
  assign y8651 = ~n21489 ;
  assign y8652 = ~n21493 ;
  assign y8653 = n21494 ;
  assign y8654 = ~n21495 ;
  assign y8655 = ~1'b0 ;
  assign y8656 = ~n21497 ;
  assign y8657 = ~n21502 ;
  assign y8658 = n21504 ;
  assign y8659 = ~n21510 ;
  assign y8660 = ~n21515 ;
  assign y8661 = ~n21518 ;
  assign y8662 = n21520 ;
  assign y8663 = ~1'b0 ;
  assign y8664 = ~n21521 ;
  assign y8665 = ~n21522 ;
  assign y8666 = n21523 ;
  assign y8667 = ~n21524 ;
  assign y8668 = ~n21530 ;
  assign y8669 = n21535 ;
  assign y8670 = ~n21540 ;
  assign y8671 = n21544 ;
  assign y8672 = n21546 ;
  assign y8673 = n21547 ;
  assign y8674 = n21549 ;
  assign y8675 = n21553 ;
  assign y8676 = ~1'b0 ;
  assign y8677 = ~1'b0 ;
  assign y8678 = ~n18296 ;
  assign y8679 = ~n21556 ;
  assign y8680 = ~n21562 ;
  assign y8681 = ~n21569 ;
  assign y8682 = ~n21570 ;
  assign y8683 = ~n21573 ;
  assign y8684 = n21577 ;
  assign y8685 = ~n21579 ;
  assign y8686 = n21582 ;
  assign y8687 = n21583 ;
  assign y8688 = ~n21585 ;
  assign y8689 = n21586 ;
  assign y8690 = 1'b0 ;
  assign y8691 = ~1'b0 ;
  assign y8692 = ~1'b0 ;
  assign y8693 = ~1'b0 ;
  assign y8694 = ~1'b0 ;
  assign y8695 = n4014 ;
  assign y8696 = ~n21587 ;
  assign y8697 = ~n21589 ;
  assign y8698 = n21590 ;
  assign y8699 = ~1'b0 ;
  assign y8700 = ~n12201 ;
  assign y8701 = ~n21595 ;
  assign y8702 = ~n21597 ;
  assign y8703 = ~1'b0 ;
  assign y8704 = ~1'b0 ;
  assign y8705 = ~n21599 ;
  assign y8706 = ~1'b0 ;
  assign y8707 = n21600 ;
  assign y8708 = ~n21603 ;
  assign y8709 = ~n11147 ;
  assign y8710 = ~n21605 ;
  assign y8711 = ~n21606 ;
  assign y8712 = n21608 ;
  assign y8713 = ~1'b0 ;
  assign y8714 = ~n21611 ;
  assign y8715 = n21614 ;
  assign y8716 = ~n21618 ;
  assign y8717 = ~n21621 ;
  assign y8718 = n21622 ;
  assign y8719 = n21624 ;
  assign y8720 = n21629 ;
  assign y8721 = ~n21630 ;
  assign y8722 = n21632 ;
  assign y8723 = ~1'b0 ;
  assign y8724 = ~n21635 ;
  assign y8725 = ~n21637 ;
  assign y8726 = ~n21640 ;
  assign y8727 = ~n21642 ;
  assign y8728 = n21643 ;
  assign y8729 = ~n21644 ;
  assign y8730 = ~n21648 ;
  assign y8731 = ~1'b0 ;
  assign y8732 = ~1'b0 ;
  assign y8733 = ~1'b0 ;
  assign y8734 = ~1'b0 ;
  assign y8735 = ~n21656 ;
  assign y8736 = n21659 ;
  assign y8737 = ~n21661 ;
  assign y8738 = n21664 ;
  assign y8739 = ~1'b0 ;
  assign y8740 = n21665 ;
  assign y8741 = ~n21670 ;
  assign y8742 = ~1'b0 ;
  assign y8743 = n21673 ;
  assign y8744 = n21676 ;
  assign y8745 = n21679 ;
  assign y8746 = ~n21680 ;
  assign y8747 = n21682 ;
  assign y8748 = n21688 ;
  assign y8749 = n21690 ;
  assign y8750 = ~n21691 ;
  assign y8751 = n21695 ;
  assign y8752 = ~1'b0 ;
  assign y8753 = n21703 ;
  assign y8754 = n21706 ;
  assign y8755 = n10260 ;
  assign y8756 = n21711 ;
  assign y8757 = ~n6320 ;
  assign y8758 = ~1'b0 ;
  assign y8759 = ~n21719 ;
  assign y8760 = n21723 ;
  assign y8761 = n21725 ;
  assign y8762 = ~n21727 ;
  assign y8763 = n21728 ;
  assign y8764 = ~n21732 ;
  assign y8765 = n21734 ;
  assign y8766 = n21736 ;
  assign y8767 = ~n21740 ;
  assign y8768 = ~n21744 ;
  assign y8769 = ~n21747 ;
  assign y8770 = ~n21748 ;
  assign y8771 = n21753 ;
  assign y8772 = ~n21756 ;
  assign y8773 = ~n21758 ;
  assign y8774 = 1'b0 ;
  assign y8775 = ~1'b0 ;
  assign y8776 = n21760 ;
  assign y8777 = ~n21762 ;
  assign y8778 = ~n3988 ;
  assign y8779 = ~1'b0 ;
  assign y8780 = ~1'b0 ;
  assign y8781 = ~n21771 ;
  assign y8782 = ~n21773 ;
  assign y8783 = n21781 ;
  assign y8784 = ~n21789 ;
  assign y8785 = ~n21790 ;
  assign y8786 = ~1'b0 ;
  assign y8787 = ~1'b0 ;
  assign y8788 = ~1'b0 ;
  assign y8789 = n20157 ;
  assign y8790 = ~n21795 ;
  assign y8791 = n21799 ;
  assign y8792 = n21800 ;
  assign y8793 = n21801 ;
  assign y8794 = ~n21804 ;
  assign y8795 = ~n21808 ;
  assign y8796 = ~1'b0 ;
  assign y8797 = ~1'b0 ;
  assign y8798 = n2933 ;
  assign y8799 = ~n21811 ;
  assign y8800 = ~n21817 ;
  assign y8801 = ~n21819 ;
  assign y8802 = n21820 ;
  assign y8803 = n21823 ;
  assign y8804 = ~1'b0 ;
  assign y8805 = ~1'b0 ;
  assign y8806 = ~1'b0 ;
  assign y8807 = ~n21825 ;
  assign y8808 = ~1'b0 ;
  assign y8809 = n21830 ;
  assign y8810 = n21833 ;
  assign y8811 = n21840 ;
  assign y8812 = n21844 ;
  assign y8813 = ~n21845 ;
  assign y8814 = ~n21846 ;
  assign y8815 = n21847 ;
  assign y8816 = ~n21849 ;
  assign y8817 = ~n21852 ;
  assign y8818 = ~n21853 ;
  assign y8819 = ~n21854 ;
  assign y8820 = n21857 ;
  assign y8821 = ~1'b0 ;
  assign y8822 = ~1'b0 ;
  assign y8823 = ~1'b0 ;
  assign y8824 = ~n21861 ;
  assign y8825 = ~1'b0 ;
  assign y8826 = n21862 ;
  assign y8827 = n21865 ;
  assign y8828 = n21867 ;
  assign y8829 = ~n21868 ;
  assign y8830 = ~n21870 ;
  assign y8831 = ~1'b0 ;
  assign y8832 = ~n21871 ;
  assign y8833 = n21872 ;
  assign y8834 = ~n21877 ;
  assign y8835 = n21879 ;
  assign y8836 = ~n21883 ;
  assign y8837 = ~n21887 ;
  assign y8838 = ~n21891 ;
  assign y8839 = n21892 ;
  assign y8840 = n21896 ;
  assign y8841 = ~n21897 ;
  assign y8842 = ~n21904 ;
  assign y8843 = n21908 ;
  assign y8844 = n21912 ;
  assign y8845 = ~1'b0 ;
  assign y8846 = ~1'b0 ;
  assign y8847 = ~1'b0 ;
  assign y8848 = n21914 ;
  assign y8849 = n21917 ;
  assign y8850 = n21923 ;
  assign y8851 = ~n21927 ;
  assign y8852 = ~n21929 ;
  assign y8853 = ~n11536 ;
  assign y8854 = ~n21931 ;
  assign y8855 = ~n21933 ;
  assign y8856 = ~1'b0 ;
  assign y8857 = ~n21936 ;
  assign y8858 = ~n21938 ;
  assign y8859 = ~n21940 ;
  assign y8860 = ~n21942 ;
  assign y8861 = ~n21947 ;
  assign y8862 = ~n11402 ;
  assign y8863 = n21949 ;
  assign y8864 = ~n21951 ;
  assign y8865 = ~n21953 ;
  assign y8866 = n9544 ;
  assign y8867 = ~1'b0 ;
  assign y8868 = n21955 ;
  assign y8869 = 1'b0 ;
  assign y8870 = n21960 ;
  assign y8871 = ~n21962 ;
  assign y8872 = ~n21963 ;
  assign y8873 = ~n21969 ;
  assign y8874 = ~n21970 ;
  assign y8875 = ~1'b0 ;
  assign y8876 = ~n21972 ;
  assign y8877 = ~n21974 ;
  assign y8878 = n21975 ;
  assign y8879 = ~n21978 ;
  assign y8880 = ~n21983 ;
  assign y8881 = ~n21984 ;
  assign y8882 = ~n21985 ;
  assign y8883 = n21991 ;
  assign y8884 = ~1'b0 ;
  assign y8885 = ~1'b0 ;
  assign y8886 = n15149 ;
  assign y8887 = ~n21992 ;
  assign y8888 = ~n7311 ;
  assign y8889 = n21994 ;
  assign y8890 = ~1'b0 ;
  assign y8891 = n21995 ;
  assign y8892 = ~n21996 ;
  assign y8893 = n21999 ;
  assign y8894 = n22000 ;
  assign y8895 = n22001 ;
  assign y8896 = ~1'b0 ;
  assign y8897 = ~n22002 ;
  assign y8898 = ~1'b0 ;
  assign y8899 = ~n22003 ;
  assign y8900 = n22004 ;
  assign y8901 = n22006 ;
  assign y8902 = ~n22007 ;
  assign y8903 = n22009 ;
  assign y8904 = ~n22011 ;
  assign y8905 = n22016 ;
  assign y8906 = n22017 ;
  assign y8907 = n22021 ;
  assign y8908 = n22022 ;
  assign y8909 = ~n22029 ;
  assign y8910 = ~1'b0 ;
  assign y8911 = ~1'b0 ;
  assign y8912 = n22034 ;
  assign y8913 = n22036 ;
  assign y8914 = ~n22041 ;
  assign y8915 = ~n22043 ;
  assign y8916 = ~1'b0 ;
  assign y8917 = ~n22044 ;
  assign y8918 = n22045 ;
  assign y8919 = ~n22047 ;
  assign y8920 = ~n22052 ;
  assign y8921 = ~n22053 ;
  assign y8922 = ~n22055 ;
  assign y8923 = n22059 ;
  assign y8924 = ~1'b0 ;
  assign y8925 = ~n22062 ;
  assign y8926 = n22064 ;
  assign y8927 = n22066 ;
  assign y8928 = ~1'b0 ;
  assign y8929 = n22067 ;
  assign y8930 = ~n22069 ;
  assign y8931 = ~1'b0 ;
  assign y8932 = n22073 ;
  assign y8933 = n22074 ;
  assign y8934 = ~n22076 ;
  assign y8935 = n22077 ;
  assign y8936 = ~n22078 ;
  assign y8937 = ~n22080 ;
  assign y8938 = ~n22082 ;
  assign y8939 = ~n22086 ;
  assign y8940 = ~n22088 ;
  assign y8941 = ~1'b0 ;
  assign y8942 = n22090 ;
  assign y8943 = ~n22091 ;
  assign y8944 = ~n22092 ;
  assign y8945 = ~n22094 ;
  assign y8946 = n22095 ;
  assign y8947 = n22096 ;
  assign y8948 = ~1'b0 ;
  assign y8949 = ~n4887 ;
  assign y8950 = ~n22097 ;
  assign y8951 = n22098 ;
  assign y8952 = n22100 ;
  assign y8953 = ~n22103 ;
  assign y8954 = ~n4593 ;
  assign y8955 = ~n22104 ;
  assign y8956 = ~1'b0 ;
  assign y8957 = ~n22107 ;
  assign y8958 = n22109 ;
  assign y8959 = n22111 ;
  assign y8960 = n22112 ;
  assign y8961 = n22115 ;
  assign y8962 = ~n22116 ;
  assign y8963 = ~n22117 ;
  assign y8964 = n22119 ;
  assign y8965 = ~n22121 ;
  assign y8966 = ~1'b0 ;
  assign y8967 = ~1'b0 ;
  assign y8968 = n22123 ;
  assign y8969 = n22125 ;
  assign y8970 = n22127 ;
  assign y8971 = n22128 ;
  assign y8972 = n22129 ;
  assign y8973 = n19405 ;
  assign y8974 = ~n22133 ;
  assign y8975 = n22134 ;
  assign y8976 = n22137 ;
  assign y8977 = ~1'b0 ;
  assign y8978 = ~n22139 ;
  assign y8979 = ~n22140 ;
  assign y8980 = n22141 ;
  assign y8981 = n22142 ;
  assign y8982 = n22146 ;
  assign y8983 = n22151 ;
  assign y8984 = n14665 ;
  assign y8985 = n22152 ;
  assign y8986 = ~n22153 ;
  assign y8987 = n22155 ;
  assign y8988 = ~n22165 ;
  assign y8989 = n22170 ;
  assign y8990 = ~n438 ;
  assign y8991 = ~n22174 ;
  assign y8992 = 1'b0 ;
  assign y8993 = ~n22175 ;
  assign y8994 = ~1'b0 ;
  assign y8995 = n22177 ;
  assign y8996 = ~1'b0 ;
  assign y8997 = ~1'b0 ;
  assign y8998 = ~n22180 ;
  assign y8999 = ~n22182 ;
  assign y9000 = n22185 ;
  assign y9001 = ~n22187 ;
  assign y9002 = ~n22191 ;
  assign y9003 = n22192 ;
  assign y9004 = ~n22193 ;
  assign y9005 = ~n22194 ;
  assign y9006 = ~n22196 ;
  assign y9007 = ~n22198 ;
  assign y9008 = n22200 ;
  assign y9009 = ~n22202 ;
  assign y9010 = ~1'b0 ;
  assign y9011 = ~n22203 ;
  assign y9012 = ~n22205 ;
  assign y9013 = ~n22206 ;
  assign y9014 = n22215 ;
  assign y9015 = ~n22216 ;
  assign y9016 = ~n22218 ;
  assign y9017 = ~1'b0 ;
  assign y9018 = ~n22224 ;
  assign y9019 = n22227 ;
  assign y9020 = n22230 ;
  assign y9021 = ~n22233 ;
  assign y9022 = n22238 ;
  assign y9023 = n22240 ;
  assign y9024 = ~1'b0 ;
  assign y9025 = n22248 ;
  assign y9026 = n22249 ;
  assign y9027 = n22255 ;
  assign y9028 = ~1'b0 ;
  assign y9029 = ~n22256 ;
  assign y9030 = ~n22262 ;
  assign y9031 = ~n22263 ;
  assign y9032 = ~1'b0 ;
  assign y9033 = n22264 ;
  assign y9034 = ~n22265 ;
  assign y9035 = ~1'b0 ;
  assign y9036 = ~n22266 ;
  assign y9037 = ~n22267 ;
  assign y9038 = ~n22269 ;
  assign y9039 = n22272 ;
  assign y9040 = ~1'b0 ;
  assign y9041 = ~n22277 ;
  assign y9042 = ~n22278 ;
  assign y9043 = n22280 ;
  assign y9044 = ~n22281 ;
  assign y9045 = ~n22290 ;
  assign y9046 = n20655 ;
  assign y9047 = n22295 ;
  assign y9048 = ~1'b0 ;
  assign y9049 = ~n22297 ;
  assign y9050 = ~1'b0 ;
  assign y9051 = ~n22300 ;
  assign y9052 = n22302 ;
  assign y9053 = n22304 ;
  assign y9054 = ~n22308 ;
  assign y9055 = ~n17727 ;
  assign y9056 = ~n22311 ;
  assign y9057 = ~n22316 ;
  assign y9058 = ~1'b0 ;
  assign y9059 = ~1'b0 ;
  assign y9060 = n22325 ;
  assign y9061 = ~1'b0 ;
  assign y9062 = ~1'b0 ;
  assign y9063 = ~n22328 ;
  assign y9064 = n22331 ;
  assign y9065 = n22334 ;
  assign y9066 = ~n22335 ;
  assign y9067 = n22343 ;
  assign y9068 = ~n22345 ;
  assign y9069 = ~1'b0 ;
  assign y9070 = n22356 ;
  assign y9071 = ~n22358 ;
  assign y9072 = ~n22360 ;
  assign y9073 = n22362 ;
  assign y9074 = ~1'b0 ;
  assign y9075 = ~1'b0 ;
  assign y9076 = ~1'b0 ;
  assign y9077 = n22366 ;
  assign y9078 = ~n5745 ;
  assign y9079 = ~n22369 ;
  assign y9080 = n22371 ;
  assign y9081 = 1'b0 ;
  assign y9082 = ~n22372 ;
  assign y9083 = ~1'b0 ;
  assign y9084 = n22373 ;
  assign y9085 = n22376 ;
  assign y9086 = ~1'b0 ;
  assign y9087 = ~n22378 ;
  assign y9088 = ~n22379 ;
  assign y9089 = n16900 ;
  assign y9090 = ~n22380 ;
  assign y9091 = ~n22389 ;
  assign y9092 = ~1'b0 ;
  assign y9093 = n22391 ;
  assign y9094 = ~1'b0 ;
  assign y9095 = n22395 ;
  assign y9096 = n302 ;
  assign y9097 = n22396 ;
  assign y9098 = ~n22399 ;
  assign y9099 = ~n10335 ;
  assign y9100 = n22404 ;
  assign y9101 = ~n22405 ;
  assign y9102 = ~n22407 ;
  assign y9103 = ~1'b0 ;
  assign y9104 = n22409 ;
  assign y9105 = n22413 ;
  assign y9106 = ~1'b0 ;
  assign y9107 = n22415 ;
  assign y9108 = ~1'b0 ;
  assign y9109 = ~n22421 ;
  assign y9110 = ~1'b0 ;
  assign y9111 = ~n22423 ;
  assign y9112 = n22424 ;
  assign y9113 = ~n22428 ;
  assign y9114 = ~n22431 ;
  assign y9115 = ~n22432 ;
  assign y9116 = n22436 ;
  assign y9117 = n1175 ;
  assign y9118 = n22438 ;
  assign y9119 = n22439 ;
  assign y9120 = ~1'b0 ;
  assign y9121 = ~n22443 ;
  assign y9122 = ~n22448 ;
  assign y9123 = ~n22449 ;
  assign y9124 = n22452 ;
  assign y9125 = ~n22453 ;
  assign y9126 = n8794 ;
  assign y9127 = ~n22455 ;
  assign y9128 = ~n22456 ;
  assign y9129 = n22457 ;
  assign y9130 = n22460 ;
  assign y9131 = n22463 ;
  assign y9132 = ~n22464 ;
  assign y9133 = ~n22466 ;
  assign y9134 = ~n22468 ;
  assign y9135 = n22472 ;
  assign y9136 = n22475 ;
  assign y9137 = ~n22477 ;
  assign y9138 = ~n22479 ;
  assign y9139 = n22485 ;
  assign y9140 = ~1'b0 ;
  assign y9141 = n22492 ;
  assign y9142 = n22493 ;
  assign y9143 = ~n22494 ;
  assign y9144 = n22495 ;
  assign y9145 = n22496 ;
  assign y9146 = ~1'b0 ;
  assign y9147 = ~n22502 ;
  assign y9148 = n22506 ;
  assign y9149 = ~1'b0 ;
  assign y9150 = ~1'b0 ;
  assign y9151 = n22508 ;
  assign y9152 = ~1'b0 ;
  assign y9153 = ~n22509 ;
  assign y9154 = ~n22515 ;
  assign y9155 = ~1'b0 ;
  assign y9156 = ~n22517 ;
  assign y9157 = ~n22519 ;
  assign y9158 = ~1'b0 ;
  assign y9159 = ~1'b0 ;
  assign y9160 = n22522 ;
  assign y9161 = ~n22525 ;
  assign y9162 = ~n22526 ;
  assign y9163 = ~n22529 ;
  assign y9164 = ~1'b0 ;
  assign y9165 = n22535 ;
  assign y9166 = ~n22536 ;
  assign y9167 = ~n22538 ;
  assign y9168 = n22541 ;
  assign y9169 = n22542 ;
  assign y9170 = n22545 ;
  assign y9171 = ~1'b0 ;
  assign y9172 = n22547 ;
  assign y9173 = n17803 ;
  assign y9174 = n22550 ;
  assign y9175 = ~n22551 ;
  assign y9176 = n22555 ;
  assign y9177 = ~n22556 ;
  assign y9178 = ~n22557 ;
  assign y9179 = n22562 ;
  assign y9180 = n22567 ;
  assign y9181 = ~1'b0 ;
  assign y9182 = ~n22569 ;
  assign y9183 = n22570 ;
  assign y9184 = n22572 ;
  assign y9185 = ~n22574 ;
  assign y9186 = n22575 ;
  assign y9187 = ~n22580 ;
  assign y9188 = n22582 ;
  assign y9189 = n22588 ;
  assign y9190 = ~1'b0 ;
  assign y9191 = ~1'b0 ;
  assign y9192 = ~n22591 ;
  assign y9193 = n22592 ;
  assign y9194 = ~n22598 ;
  assign y9195 = ~n22601 ;
  assign y9196 = n22602 ;
  assign y9197 = ~n22603 ;
  assign y9198 = n22606 ;
  assign y9199 = n22607 ;
  assign y9200 = n22608 ;
  assign y9201 = n22610 ;
  assign y9202 = ~n22613 ;
  assign y9203 = ~1'b0 ;
  assign y9204 = ~1'b0 ;
  assign y9205 = ~n22614 ;
  assign y9206 = ~n22615 ;
  assign y9207 = ~1'b0 ;
  assign y9208 = ~n22618 ;
  assign y9209 = ~1'b0 ;
  assign y9210 = ~n22622 ;
  assign y9211 = n22623 ;
  assign y9212 = ~n22625 ;
  assign y9213 = ~n22628 ;
  assign y9214 = ~n22633 ;
  assign y9215 = n22635 ;
  assign y9216 = ~1'b0 ;
  assign y9217 = n22637 ;
  assign y9218 = ~n22639 ;
  assign y9219 = n22640 ;
  assign y9220 = ~n22645 ;
  assign y9221 = ~n22646 ;
  assign y9222 = ~1'b0 ;
  assign y9223 = n22650 ;
  assign y9224 = ~n22652 ;
  assign y9225 = n22655 ;
  assign y9226 = ~1'b0 ;
  assign y9227 = ~1'b0 ;
  assign y9228 = ~n22662 ;
  assign y9229 = ~n22663 ;
  assign y9230 = ~n22664 ;
  assign y9231 = ~1'b0 ;
  assign y9232 = ~n22666 ;
  assign y9233 = ~1'b0 ;
  assign y9234 = n22670 ;
  assign y9235 = ~1'b0 ;
  assign y9236 = n22673 ;
  assign y9237 = ~n11892 ;
  assign y9238 = n22674 ;
  assign y9239 = ~1'b0 ;
  assign y9240 = ~n22676 ;
  assign y9241 = ~1'b0 ;
  assign y9242 = ~1'b0 ;
  assign y9243 = n22678 ;
  assign y9244 = n22680 ;
  assign y9245 = n22683 ;
  assign y9246 = ~n22687 ;
  assign y9247 = n22694 ;
  assign y9248 = ~n22695 ;
  assign y9249 = ~n22696 ;
  assign y9250 = n22699 ;
  assign y9251 = ~n22700 ;
  assign y9252 = ~n22702 ;
  assign y9253 = ~n22703 ;
  assign y9254 = ~n22706 ;
  assign y9255 = ~n22707 ;
  assign y9256 = ~n22712 ;
  assign y9257 = n22713 ;
  assign y9258 = ~n22717 ;
  assign y9259 = ~1'b0 ;
  assign y9260 = ~1'b0 ;
  assign y9261 = ~n22719 ;
  assign y9262 = ~n1918 ;
  assign y9263 = n19331 ;
  assign y9264 = ~n22720 ;
  assign y9265 = ~1'b0 ;
  assign y9266 = ~n22722 ;
  assign y9267 = ~1'b0 ;
  assign y9268 = n22723 ;
  assign y9269 = ~n22724 ;
  assign y9270 = 1'b0 ;
  assign y9271 = n22726 ;
  assign y9272 = n22728 ;
  assign y9273 = n22735 ;
  assign y9274 = n22737 ;
  assign y9275 = ~n22739 ;
  assign y9276 = n22745 ;
  assign y9277 = ~1'b0 ;
  assign y9278 = ~n22749 ;
  assign y9279 = n22752 ;
  assign y9280 = n22753 ;
  assign y9281 = ~n22757 ;
  assign y9282 = ~n12504 ;
  assign y9283 = n22761 ;
  assign y9284 = ~n22765 ;
  assign y9285 = n22768 ;
  assign y9286 = n22770 ;
  assign y9287 = n22772 ;
  assign y9288 = ~n22778 ;
  assign y9289 = ~n22779 ;
  assign y9290 = ~n22781 ;
  assign y9291 = ~1'b0 ;
  assign y9292 = n22786 ;
  assign y9293 = ~1'b0 ;
  assign y9294 = ~n10736 ;
  assign y9295 = ~n22787 ;
  assign y9296 = ~n22791 ;
  assign y9297 = n22792 ;
  assign y9298 = ~n22794 ;
  assign y9299 = ~1'b0 ;
  assign y9300 = ~n22795 ;
  assign y9301 = n22798 ;
  assign y9302 = ~1'b0 ;
  assign y9303 = ~1'b0 ;
  assign y9304 = n22800 ;
  assign y9305 = n22801 ;
  assign y9306 = n22802 ;
  assign y9307 = ~n22805 ;
  assign y9308 = ~n22808 ;
  assign y9309 = n22816 ;
  assign y9310 = ~n22817 ;
  assign y9311 = ~n22819 ;
  assign y9312 = ~1'b0 ;
  assign y9313 = ~n22821 ;
  assign y9314 = n22824 ;
  assign y9315 = ~1'b0 ;
  assign y9316 = n13401 ;
  assign y9317 = n22825 ;
  assign y9318 = 1'b0 ;
  assign y9319 = ~1'b0 ;
  assign y9320 = n22829 ;
  assign y9321 = n22834 ;
  assign y9322 = n22835 ;
  assign y9323 = n22836 ;
  assign y9324 = ~1'b0 ;
  assign y9325 = ~n22840 ;
  assign y9326 = n22843 ;
  assign y9327 = ~n22846 ;
  assign y9328 = ~n19013 ;
  assign y9329 = ~n22847 ;
  assign y9330 = ~n22849 ;
  assign y9331 = ~n22851 ;
  assign y9332 = ~n22853 ;
  assign y9333 = n22855 ;
  assign y9334 = ~n22856 ;
  assign y9335 = ~n22862 ;
  assign y9336 = ~n22864 ;
  assign y9337 = n22865 ;
  assign y9338 = ~1'b0 ;
  assign y9339 = ~n22871 ;
  assign y9340 = n22873 ;
  assign y9341 = n22876 ;
  assign y9342 = ~n22877 ;
  assign y9343 = n22881 ;
  assign y9344 = n22887 ;
  assign y9345 = ~n22889 ;
  assign y9346 = ~n22892 ;
  assign y9347 = ~1'b0 ;
  assign y9348 = n22894 ;
  assign y9349 = n22896 ;
  assign y9350 = ~n22897 ;
  assign y9351 = ~n22898 ;
  assign y9352 = ~n22900 ;
  assign y9353 = ~1'b0 ;
  assign y9354 = n22904 ;
  assign y9355 = ~n22907 ;
  assign y9356 = 1'b0 ;
  assign y9357 = n22908 ;
  assign y9358 = ~n22909 ;
  assign y9359 = 1'b0 ;
  assign y9360 = n22910 ;
  assign y9361 = n22911 ;
  assign y9362 = ~1'b0 ;
  assign y9363 = ~1'b0 ;
  assign y9364 = ~1'b0 ;
  assign y9365 = ~1'b0 ;
  assign y9366 = n22917 ;
  assign y9367 = ~n22928 ;
  assign y9368 = ~n22931 ;
  assign y9369 = n22934 ;
  assign y9370 = ~1'b0 ;
  assign y9371 = n3141 ;
  assign y9372 = ~n22937 ;
  assign y9373 = n22939 ;
  assign y9374 = n22940 ;
  assign y9375 = n22942 ;
  assign y9376 = n22943 ;
  assign y9377 = ~n22944 ;
  assign y9378 = ~n22948 ;
  assign y9379 = n22949 ;
  assign y9380 = ~n22951 ;
  assign y9381 = n22959 ;
  assign y9382 = n22960 ;
  assign y9383 = ~1'b0 ;
  assign y9384 = ~n22966 ;
  assign y9385 = ~n22967 ;
  assign y9386 = ~n22972 ;
  assign y9387 = ~n22973 ;
  assign y9388 = ~1'b0 ;
  assign y9389 = ~1'b0 ;
  assign y9390 = n22974 ;
  assign y9391 = ~1'b0 ;
  assign y9392 = n22979 ;
  assign y9393 = n22984 ;
  assign y9394 = n12520 ;
  assign y9395 = n22531 ;
  assign y9396 = n22988 ;
  assign y9397 = ~n22989 ;
  assign y9398 = n8334 ;
  assign y9399 = ~1'b0 ;
  assign y9400 = n22990 ;
  assign y9401 = n22992 ;
  assign y9402 = ~1'b0 ;
  assign y9403 = ~n22993 ;
  assign y9404 = ~n22994 ;
  assign y9405 = ~n22995 ;
  assign y9406 = n22996 ;
  assign y9407 = ~n22998 ;
  assign y9408 = ~1'b0 ;
  assign y9409 = n22999 ;
  assign y9410 = ~n23001 ;
  assign y9411 = ~n23007 ;
  assign y9412 = n23008 ;
  assign y9413 = 1'b0 ;
  assign y9414 = ~n23011 ;
  assign y9415 = n23012 ;
  assign y9416 = ~n23013 ;
  assign y9417 = ~1'b0 ;
  assign y9418 = n23017 ;
  assign y9419 = ~n23018 ;
  assign y9420 = n23024 ;
  assign y9421 = ~n23026 ;
  assign y9422 = ~1'b0 ;
  assign y9423 = ~n23028 ;
  assign y9424 = n23029 ;
  assign y9425 = n23030 ;
  assign y9426 = n23035 ;
  assign y9427 = n23038 ;
  assign y9428 = ~n23040 ;
  assign y9429 = ~1'b0 ;
  assign y9430 = n23043 ;
  assign y9431 = ~n23047 ;
  assign y9432 = ~1'b0 ;
  assign y9433 = n23049 ;
  assign y9434 = n23051 ;
  assign y9435 = ~n23052 ;
  assign y9436 = ~n23053 ;
  assign y9437 = n23056 ;
  assign y9438 = n23059 ;
  assign y9439 = ~1'b0 ;
  assign y9440 = n23061 ;
  assign y9441 = ~n23065 ;
  assign y9442 = n23066 ;
  assign y9443 = ~1'b0 ;
  assign y9444 = n23067 ;
  assign y9445 = ~n23068 ;
  assign y9446 = n23073 ;
  assign y9447 = ~n23075 ;
  assign y9448 = n23078 ;
  assign y9449 = ~n23080 ;
  assign y9450 = ~1'b0 ;
  assign y9451 = ~1'b0 ;
  assign y9452 = ~1'b0 ;
  assign y9453 = ~n23086 ;
  assign y9454 = n23087 ;
  assign y9455 = n23090 ;
  assign y9456 = ~n23092 ;
  assign y9457 = ~n23095 ;
  assign y9458 = ~n23099 ;
  assign y9459 = ~n23100 ;
  assign y9460 = n23103 ;
  assign y9461 = 1'b0 ;
  assign y9462 = ~1'b0 ;
  assign y9463 = ~n23107 ;
  assign y9464 = ~n23111 ;
  assign y9465 = n23114 ;
  assign y9466 = n23116 ;
  assign y9467 = n23119 ;
  assign y9468 = n23123 ;
  assign y9469 = ~1'b0 ;
  assign y9470 = n23124 ;
  assign y9471 = ~1'b0 ;
  assign y9472 = ~1'b0 ;
  assign y9473 = n23127 ;
  assign y9474 = n23129 ;
  assign y9475 = n23130 ;
  assign y9476 = ~n23131 ;
  assign y9477 = n23133 ;
  assign y9478 = ~n23134 ;
  assign y9479 = n23136 ;
  assign y9480 = ~1'b0 ;
  assign y9481 = ~n23137 ;
  assign y9482 = ~1'b0 ;
  assign y9483 = n23140 ;
  assign y9484 = n23146 ;
  assign y9485 = n23150 ;
  assign y9486 = ~1'b0 ;
  assign y9487 = n23153 ;
  assign y9488 = ~n23154 ;
  assign y9489 = n23156 ;
  assign y9490 = n23160 ;
  assign y9491 = ~n23161 ;
  assign y9492 = n3883 ;
  assign y9493 = ~n23163 ;
  assign y9494 = n23165 ;
  assign y9495 = ~n23167 ;
  assign y9496 = ~n23170 ;
  assign y9497 = ~n23173 ;
  assign y9498 = n23175 ;
  assign y9499 = n23180 ;
  assign y9500 = ~n23181 ;
  assign y9501 = n23183 ;
  assign y9502 = n23184 ;
  assign y9503 = ~1'b0 ;
  assign y9504 = ~n23187 ;
  assign y9505 = n23191 ;
  assign y9506 = n1518 ;
  assign y9507 = ~1'b0 ;
  assign y9508 = ~n23192 ;
  assign y9509 = ~n23194 ;
  assign y9510 = ~1'b0 ;
  assign y9511 = n23196 ;
  assign y9512 = ~n23198 ;
  assign y9513 = ~1'b0 ;
  assign y9514 = ~n23202 ;
  assign y9515 = ~n23203 ;
  assign y9516 = ~1'b0 ;
  assign y9517 = n23209 ;
  assign y9518 = ~1'b0 ;
  assign y9519 = ~n23212 ;
  assign y9520 = n23217 ;
  assign y9521 = ~n23219 ;
  assign y9522 = n23220 ;
  assign y9523 = ~n23225 ;
  assign y9524 = n23227 ;
  assign y9525 = ~1'b0 ;
  assign y9526 = ~n23229 ;
  assign y9527 = ~1'b0 ;
  assign y9528 = n23231 ;
  assign y9529 = n23233 ;
  assign y9530 = n23237 ;
  assign y9531 = ~n23238 ;
  assign y9532 = n23240 ;
  assign y9533 = ~n23245 ;
  assign y9534 = ~n23246 ;
  assign y9535 = ~n23250 ;
  assign y9536 = n23251 ;
  assign y9537 = ~n23254 ;
  assign y9538 = ~n23256 ;
  assign y9539 = ~1'b0 ;
  assign y9540 = ~1'b0 ;
  assign y9541 = n23259 ;
  assign y9542 = ~n23260 ;
  assign y9543 = ~n23261 ;
  assign y9544 = ~1'b0 ;
  assign y9545 = n23267 ;
  assign y9546 = ~n17342 ;
  assign y9547 = ~n23268 ;
  assign y9548 = ~n23269 ;
  assign y9549 = n23271 ;
  assign y9550 = ~n23274 ;
  assign y9551 = n23277 ;
  assign y9552 = ~1'b0 ;
  assign y9553 = n23280 ;
  assign y9554 = ~n23281 ;
  assign y9555 = ~n23283 ;
  assign y9556 = ~n23285 ;
  assign y9557 = ~1'b0 ;
  assign y9558 = n23287 ;
  assign y9559 = n23289 ;
  assign y9560 = ~n23291 ;
  assign y9561 = n23294 ;
  assign y9562 = ~n4455 ;
  assign y9563 = ~n23295 ;
  assign y9564 = ~n23297 ;
  assign y9565 = n23298 ;
  assign y9566 = ~n23299 ;
  assign y9567 = ~n23300 ;
  assign y9568 = ~n23309 ;
  assign y9569 = n23312 ;
  assign y9570 = ~1'b0 ;
  assign y9571 = n23313 ;
  assign y9572 = ~n23315 ;
  assign y9573 = ~1'b0 ;
  assign y9574 = ~n23316 ;
  assign y9575 = ~n23317 ;
  assign y9576 = 1'b0 ;
  assign y9577 = n2728 ;
  assign y9578 = n23321 ;
  assign y9579 = ~1'b0 ;
  assign y9580 = ~1'b0 ;
  assign y9581 = ~1'b0 ;
  assign y9582 = ~1'b0 ;
  assign y9583 = ~1'b0 ;
  assign y9584 = n23324 ;
  assign y9585 = n23328 ;
  assign y9586 = ~n23329 ;
  assign y9587 = ~n23330 ;
  assign y9588 = n23332 ;
  assign y9589 = n23334 ;
  assign y9590 = ~1'b0 ;
  assign y9591 = n23335 ;
  assign y9592 = ~1'b0 ;
  assign y9593 = ~n23337 ;
  assign y9594 = n23341 ;
  assign y9595 = n23347 ;
  assign y9596 = ~n23348 ;
  assign y9597 = n23351 ;
  assign y9598 = ~n23352 ;
  assign y9599 = ~n20716 ;
  assign y9600 = n2388 ;
  assign y9601 = n23359 ;
  assign y9602 = ~n23360 ;
  assign y9603 = n8231 ;
  assign y9604 = ~n23364 ;
  assign y9605 = n23367 ;
  assign y9606 = ~n23368 ;
  assign y9607 = n23373 ;
  assign y9608 = ~1'b0 ;
  assign y9609 = ~1'b0 ;
  assign y9610 = n23374 ;
  assign y9611 = ~n23376 ;
  assign y9612 = ~n23378 ;
  assign y9613 = n23379 ;
  assign y9614 = n23387 ;
  assign y9615 = ~n23388 ;
  assign y9616 = n23389 ;
  assign y9617 = ~n23390 ;
  assign y9618 = ~1'b0 ;
  assign y9619 = ~n23392 ;
  assign y9620 = n23396 ;
  assign y9621 = n23397 ;
  assign y9622 = ~n23400 ;
  assign y9623 = ~1'b0 ;
  assign y9624 = n23401 ;
  assign y9625 = n23404 ;
  assign y9626 = n23405 ;
  assign y9627 = n23407 ;
  assign y9628 = ~1'b0 ;
  assign y9629 = ~n23409 ;
  assign y9630 = n23411 ;
  assign y9631 = ~n23412 ;
  assign y9632 = ~n23415 ;
  assign y9633 = n23416 ;
  assign y9634 = n23420 ;
  assign y9635 = n23424 ;
  assign y9636 = ~n23425 ;
  assign y9637 = ~1'b0 ;
  assign y9638 = ~1'b0 ;
  assign y9639 = n23427 ;
  assign y9640 = ~1'b0 ;
  assign y9641 = n22351 ;
  assign y9642 = ~n23434 ;
  assign y9643 = n23437 ;
  assign y9644 = n23438 ;
  assign y9645 = n23441 ;
  assign y9646 = ~n23444 ;
  assign y9647 = n23445 ;
  assign y9648 = ~n23447 ;
  assign y9649 = ~n23453 ;
  assign y9650 = ~1'b0 ;
  assign y9651 = ~n23458 ;
  assign y9652 = n23459 ;
  assign y9653 = ~n23461 ;
  assign y9654 = ~n23462 ;
  assign y9655 = ~n23464 ;
  assign y9656 = ~n23465 ;
  assign y9657 = ~1'b0 ;
  assign y9658 = ~n23471 ;
  assign y9659 = ~n23473 ;
  assign y9660 = ~1'b0 ;
  assign y9661 = ~1'b0 ;
  assign y9662 = ~1'b0 ;
  assign y9663 = n23475 ;
  assign y9664 = ~n23477 ;
  assign y9665 = n6205 ;
  assign y9666 = ~n1192 ;
  assign y9667 = ~n23479 ;
  assign y9668 = ~n23485 ;
  assign y9669 = n23494 ;
  assign y9670 = ~1'b0 ;
  assign y9671 = ~n23495 ;
  assign y9672 = ~1'b0 ;
  assign y9673 = n23497 ;
  assign y9674 = ~n23501 ;
  assign y9675 = n23506 ;
  assign y9676 = n23508 ;
  assign y9677 = ~n23514 ;
  assign y9678 = n23517 ;
  assign y9679 = ~n23521 ;
  assign y9680 = ~1'b0 ;
  assign y9681 = ~n23522 ;
  assign y9682 = ~n23525 ;
  assign y9683 = ~n23526 ;
  assign y9684 = n23527 ;
  assign y9685 = n23530 ;
  assign y9686 = ~n23531 ;
  assign y9687 = ~1'b0 ;
  assign y9688 = n23533 ;
  assign y9689 = n23537 ;
  assign y9690 = n23539 ;
  assign y9691 = n23541 ;
  assign y9692 = ~n23543 ;
  assign y9693 = ~n23546 ;
  assign y9694 = ~1'b0 ;
  assign y9695 = ~1'b0 ;
  assign y9696 = ~n23549 ;
  assign y9697 = n23550 ;
  assign y9698 = n23552 ;
  assign y9699 = ~n23554 ;
  assign y9700 = ~n23557 ;
  assign y9701 = ~n23558 ;
  assign y9702 = ~n23560 ;
  assign y9703 = ~n23563 ;
  assign y9704 = n23564 ;
  assign y9705 = n23566 ;
  assign y9706 = ~n23568 ;
  assign y9707 = n8491 ;
  assign y9708 = n23573 ;
  assign y9709 = ~n23574 ;
  assign y9710 = n23577 ;
  assign y9711 = n23578 ;
  assign y9712 = ~n23579 ;
  assign y9713 = ~1'b0 ;
  assign y9714 = n23581 ;
  assign y9715 = n23582 ;
  assign y9716 = ~n23584 ;
  assign y9717 = n23588 ;
  assign y9718 = n23589 ;
  assign y9719 = n23590 ;
  assign y9720 = ~n23594 ;
  assign y9721 = ~1'b0 ;
  assign y9722 = ~n23595 ;
  assign y9723 = n23599 ;
  assign y9724 = n23601 ;
  assign y9725 = n23603 ;
  assign y9726 = n23612 ;
  assign y9727 = ~n23613 ;
  assign y9728 = ~n23616 ;
  assign y9729 = ~1'b0 ;
  assign y9730 = ~1'b0 ;
  assign y9731 = ~1'b0 ;
  assign y9732 = ~n23618 ;
  assign y9733 = ~n23619 ;
  assign y9734 = ~n23626 ;
  assign y9735 = ~n23627 ;
  assign y9736 = n23630 ;
  assign y9737 = ~1'b0 ;
  assign y9738 = ~n23631 ;
  assign y9739 = ~1'b0 ;
  assign y9740 = n23632 ;
  assign y9741 = ~n23634 ;
  assign y9742 = ~n23638 ;
  assign y9743 = ~n23640 ;
  assign y9744 = n9292 ;
  assign y9745 = ~1'b0 ;
  assign y9746 = n23643 ;
  assign y9747 = ~1'b0 ;
  assign y9748 = ~n23644 ;
  assign y9749 = ~n23646 ;
  assign y9750 = ~n23649 ;
  assign y9751 = n23650 ;
  assign y9752 = ~1'b0 ;
  assign y9753 = ~1'b0 ;
  assign y9754 = n23652 ;
  assign y9755 = ~n23655 ;
  assign y9756 = n23664 ;
  assign y9757 = n23667 ;
  assign y9758 = n23673 ;
  assign y9759 = ~n23674 ;
  assign y9760 = 1'b0 ;
  assign y9761 = ~1'b0 ;
  assign y9762 = ~1'b0 ;
  assign y9763 = ~1'b0 ;
  assign y9764 = n23681 ;
  assign y9765 = 1'b0 ;
  assign y9766 = n23683 ;
  assign y9767 = n23686 ;
  assign y9768 = n23689 ;
  assign y9769 = ~n23690 ;
  assign y9770 = ~1'b0 ;
  assign y9771 = ~n23694 ;
  assign y9772 = ~n23697 ;
  assign y9773 = n23699 ;
  assign y9774 = ~n23700 ;
  assign y9775 = n23702 ;
  assign y9776 = ~n16056 ;
  assign y9777 = ~n23708 ;
  assign y9778 = n23712 ;
  assign y9779 = ~n23715 ;
  assign y9780 = n23717 ;
  assign y9781 = ~1'b0 ;
  assign y9782 = ~1'b0 ;
  assign y9783 = n23718 ;
  assign y9784 = ~n23722 ;
  assign y9785 = n23729 ;
  assign y9786 = n23730 ;
  assign y9787 = n23732 ;
  assign y9788 = ~n7010 ;
  assign y9789 = ~1'b0 ;
  assign y9790 = ~1'b0 ;
  assign y9791 = n23739 ;
  assign y9792 = n9343 ;
  assign y9793 = n23740 ;
  assign y9794 = n23741 ;
  assign y9795 = ~n23742 ;
  assign y9796 = ~1'b0 ;
  assign y9797 = n14393 ;
  assign y9798 = ~1'b0 ;
  assign y9799 = ~1'b0 ;
  assign y9800 = ~n17856 ;
  assign y9801 = ~1'b0 ;
  assign y9802 = n23748 ;
  assign y9803 = n23751 ;
  assign y9804 = ~n23753 ;
  assign y9805 = ~n23755 ;
  assign y9806 = ~1'b0 ;
  assign y9807 = ~n23756 ;
  assign y9808 = ~1'b0 ;
  assign y9809 = ~n23758 ;
  assign y9810 = ~1'b0 ;
  assign y9811 = ~n23759 ;
  assign y9812 = n23770 ;
  assign y9813 = n23771 ;
  assign y9814 = ~n23709 ;
  assign y9815 = ~n23773 ;
  assign y9816 = n23775 ;
  assign y9817 = ~1'b0 ;
  assign y9818 = ~n23778 ;
  assign y9819 = n23782 ;
  assign y9820 = ~1'b0 ;
  assign y9821 = n23783 ;
  assign y9822 = n23784 ;
  assign y9823 = ~1'b0 ;
  assign y9824 = ~n23788 ;
  assign y9825 = ~n23790 ;
  assign y9826 = ~n23792 ;
  assign y9827 = ~n23795 ;
  assign y9828 = ~1'b0 ;
  assign y9829 = ~n7162 ;
  assign y9830 = ~n23796 ;
  assign y9831 = ~1'b0 ;
  assign y9832 = n23798 ;
  assign y9833 = ~1'b0 ;
  assign y9834 = ~n23803 ;
  assign y9835 = ~n23807 ;
  assign y9836 = ~n23809 ;
  assign y9837 = ~n23813 ;
  assign y9838 = ~1'b0 ;
  assign y9839 = n23816 ;
  assign y9840 = ~n23818 ;
  assign y9841 = ~n23820 ;
  assign y9842 = ~n23821 ;
  assign y9843 = ~1'b0 ;
  assign y9844 = n23822 ;
  assign y9845 = n23826 ;
  assign y9846 = n23827 ;
  assign y9847 = ~n23834 ;
  assign y9848 = ~n23838 ;
  assign y9849 = n23843 ;
  assign y9850 = ~n23845 ;
  assign y9851 = n23847 ;
  assign y9852 = ~1'b0 ;
  assign y9853 = ~1'b0 ;
  assign y9854 = ~n23852 ;
  assign y9855 = ~1'b0 ;
  assign y9856 = ~n23853 ;
  assign y9857 = ~1'b0 ;
  assign y9858 = n23855 ;
  assign y9859 = ~1'b0 ;
  assign y9860 = ~1'b0 ;
  assign y9861 = ~n23856 ;
  assign y9862 = ~1'b0 ;
  assign y9863 = n1653 ;
  assign y9864 = n23858 ;
  assign y9865 = ~n23862 ;
  assign y9866 = ~n23865 ;
  assign y9867 = n2171 ;
  assign y9868 = ~n23867 ;
  assign y9869 = ~1'b0 ;
  assign y9870 = n23868 ;
  assign y9871 = ~n23871 ;
  assign y9872 = ~n23874 ;
  assign y9873 = ~n23876 ;
  assign y9874 = n23880 ;
  assign y9875 = n23882 ;
  assign y9876 = 1'b0 ;
  assign y9877 = n23884 ;
  assign y9878 = ~n23886 ;
  assign y9879 = n23888 ;
  assign y9880 = ~n23889 ;
  assign y9881 = n23891 ;
  assign y9882 = n23892 ;
  assign y9883 = n23896 ;
  assign y9884 = n23897 ;
  assign y9885 = n23900 ;
  assign y9886 = ~1'b0 ;
  assign y9887 = n15756 ;
  assign y9888 = ~n23907 ;
  assign y9889 = n23908 ;
  assign y9890 = n23909 ;
  assign y9891 = ~n23913 ;
  assign y9892 = ~n23914 ;
  assign y9893 = n23916 ;
  assign y9894 = ~1'b0 ;
  assign y9895 = ~1'b0 ;
  assign y9896 = ~1'b0 ;
  assign y9897 = ~n23921 ;
  assign y9898 = ~1'b0 ;
  assign y9899 = ~n23923 ;
  assign y9900 = ~n21126 ;
  assign y9901 = ~n23924 ;
  assign y9902 = n23925 ;
  assign y9903 = ~n23926 ;
  assign y9904 = n23929 ;
  assign y9905 = ~n4890 ;
  assign y9906 = ~n23931 ;
  assign y9907 = ~n23932 ;
  assign y9908 = ~1'b0 ;
  assign y9909 = n23933 ;
  assign y9910 = n23934 ;
  assign y9911 = n23935 ;
  assign y9912 = n23939 ;
  assign y9913 = n23941 ;
  assign y9914 = n23943 ;
  assign y9915 = n23944 ;
  assign y9916 = ~n23947 ;
  assign y9917 = ~1'b0 ;
  assign y9918 = ~n23948 ;
  assign y9919 = ~n23949 ;
  assign y9920 = n23950 ;
  assign y9921 = ~n23951 ;
  assign y9922 = ~n23954 ;
  assign y9923 = n23956 ;
  assign y9924 = ~n23957 ;
  assign y9925 = ~n23963 ;
  assign y9926 = ~n23971 ;
  assign y9927 = ~n23973 ;
  assign y9928 = n23974 ;
  assign y9929 = ~n23978 ;
  assign y9930 = n23982 ;
  assign y9931 = ~1'b0 ;
  assign y9932 = ~1'b0 ;
  assign y9933 = n23988 ;
  assign y9934 = ~n23994 ;
  assign y9935 = ~n24000 ;
  assign y9936 = n24001 ;
  assign y9937 = ~n24002 ;
  assign y9938 = ~n24004 ;
  assign y9939 = ~n24006 ;
  assign y9940 = n24008 ;
  assign y9941 = n2371 ;
  assign y9942 = ~1'b0 ;
  assign y9943 = ~n24009 ;
  assign y9944 = ~1'b0 ;
  assign y9945 = ~n24012 ;
  assign y9946 = n24014 ;
  assign y9947 = n24020 ;
  assign y9948 = ~n24021 ;
  assign y9949 = ~n24024 ;
  assign y9950 = n24028 ;
  assign y9951 = n24030 ;
  assign y9952 = ~n24032 ;
  assign y9953 = ~n24033 ;
  assign y9954 = ~n24038 ;
  assign y9955 = ~n24042 ;
  assign y9956 = n24045 ;
  assign y9957 = ~n24047 ;
  assign y9958 = ~n24048 ;
  assign y9959 = ~n24051 ;
  assign y9960 = n24052 ;
  assign y9961 = ~n24053 ;
  assign y9962 = ~n24059 ;
  assign y9963 = ~1'b0 ;
  assign y9964 = ~n24062 ;
  assign y9965 = ~n24063 ;
  assign y9966 = n24065 ;
  assign y9967 = ~n24069 ;
  assign y9968 = ~n24070 ;
  assign y9969 = 1'b0 ;
  assign y9970 = ~n24072 ;
  assign y9971 = ~n24073 ;
  assign y9972 = n24078 ;
  assign y9973 = ~1'b0 ;
  assign y9974 = n24083 ;
  assign y9975 = n24085 ;
  assign y9976 = n24087 ;
  assign y9977 = ~n24090 ;
  assign y9978 = n2753 ;
  assign y9979 = ~n24093 ;
  assign y9980 = n24103 ;
  assign y9981 = ~n24105 ;
  assign y9982 = n24111 ;
  assign y9983 = ~1'b0 ;
  assign y9984 = ~1'b0 ;
  assign y9985 = ~1'b0 ;
  assign y9986 = ~n24113 ;
  assign y9987 = n24116 ;
  assign y9988 = ~n24118 ;
  assign y9989 = ~n24120 ;
  assign y9990 = ~n24122 ;
  assign y9991 = ~1'b0 ;
  assign y9992 = ~n24124 ;
  assign y9993 = ~1'b0 ;
  assign y9994 = n24126 ;
  assign y9995 = ~n24130 ;
  assign y9996 = ~1'b0 ;
  assign y9997 = n22488 ;
  assign y9998 = n24131 ;
  assign y9999 = ~n24132 ;
  assign y10000 = n24134 ;
  assign y10001 = ~1'b0 ;
  assign y10002 = ~n24135 ;
  assign y10003 = n24139 ;
  assign y10004 = ~1'b0 ;
  assign y10005 = n10464 ;
  assign y10006 = n24142 ;
  assign y10007 = n24144 ;
  assign y10008 = n24148 ;
  assign y10009 = n24154 ;
  assign y10010 = ~n24156 ;
  assign y10011 = n24157 ;
  assign y10012 = ~n24158 ;
  assign y10013 = ~n24160 ;
  assign y10014 = ~n24165 ;
  assign y10015 = n24166 ;
  assign y10016 = ~n24169 ;
  assign y10017 = ~n24171 ;
  assign y10018 = ~n24172 ;
  assign y10019 = ~n24173 ;
  assign y10020 = ~n4224 ;
  assign y10021 = n24174 ;
  assign y10022 = ~n24177 ;
  assign y10023 = ~n24178 ;
  assign y10024 = ~n24179 ;
  assign y10025 = ~1'b0 ;
  assign y10026 = ~n24184 ;
  assign y10027 = ~n24187 ;
  assign y10028 = ~n24188 ;
  assign y10029 = ~n24191 ;
  assign y10030 = n24192 ;
  assign y10031 = ~n24194 ;
  assign y10032 = ~1'b0 ;
  assign y10033 = ~n24196 ;
  assign y10034 = ~n24203 ;
  assign y10035 = ~n24205 ;
  assign y10036 = n24208 ;
  assign y10037 = ~n24211 ;
  assign y10038 = ~1'b0 ;
  assign y10039 = ~n24213 ;
  assign y10040 = ~n24214 ;
  assign y10041 = ~1'b0 ;
  assign y10042 = ~n24216 ;
  assign y10043 = ~n24217 ;
  assign y10044 = ~n15033 ;
  assign y10045 = ~n24218 ;
  assign y10046 = ~n24222 ;
  assign y10047 = ~1'b0 ;
  assign y10048 = ~1'b0 ;
  assign y10049 = ~n24227 ;
  assign y10050 = n24228 ;
  assign y10051 = n24233 ;
  assign y10052 = n24235 ;
  assign y10053 = ~n24238 ;
  assign y10054 = n24240 ;
  assign y10055 = ~n1104 ;
  assign y10056 = ~1'b0 ;
  assign y10057 = n17209 ;
  assign y10058 = ~n24241 ;
  assign y10059 = ~n24243 ;
  assign y10060 = ~1'b0 ;
  assign y10061 = n24246 ;
  assign y10062 = n24247 ;
  assign y10063 = ~n24250 ;
  assign y10064 = ~n24251 ;
  assign y10065 = ~n24257 ;
  assign y10066 = ~1'b0 ;
  assign y10067 = ~1'b0 ;
  assign y10068 = ~1'b0 ;
  assign y10069 = ~n24259 ;
  assign y10070 = n24261 ;
  assign y10071 = n4085 ;
  assign y10072 = ~n24262 ;
  assign y10073 = ~n13772 ;
  assign y10074 = ~1'b0 ;
  assign y10075 = ~1'b0 ;
  assign y10076 = ~1'b0 ;
  assign y10077 = ~1'b0 ;
  assign y10078 = ~1'b0 ;
  assign y10079 = ~n24265 ;
  assign y10080 = n24267 ;
  assign y10081 = ~n24270 ;
  assign y10082 = n24272 ;
  assign y10083 = n24274 ;
  assign y10084 = ~n24275 ;
  assign y10085 = ~1'b0 ;
  assign y10086 = ~n24276 ;
  assign y10087 = ~1'b0 ;
  assign y10088 = ~n24279 ;
  assign y10089 = n24281 ;
  assign y10090 = n24284 ;
  assign y10091 = ~n24285 ;
  assign y10092 = ~n24290 ;
  assign y10093 = n24293 ;
  assign y10094 = n24298 ;
  assign y10095 = ~1'b0 ;
  assign y10096 = ~1'b0 ;
  assign y10097 = ~n24302 ;
  assign y10098 = ~n24303 ;
  assign y10099 = ~n24304 ;
  assign y10100 = ~n24308 ;
  assign y10101 = n24313 ;
  assign y10102 = ~n24316 ;
  assign y10103 = n24318 ;
  assign y10104 = n24320 ;
  assign y10105 = n24324 ;
  assign y10106 = ~n24325 ;
  assign y10107 = n24327 ;
  assign y10108 = ~n24331 ;
  assign y10109 = ~n24332 ;
  assign y10110 = n24333 ;
  assign y10111 = ~1'b0 ;
  assign y10112 = n24337 ;
  assign y10113 = ~n24339 ;
  assign y10114 = n24341 ;
  assign y10115 = n24342 ;
  assign y10116 = ~n24344 ;
  assign y10117 = n24345 ;
  assign y10118 = n24346 ;
  assign y10119 = n24355 ;
  assign y10120 = ~n24357 ;
  assign y10121 = ~n12231 ;
  assign y10122 = ~1'b0 ;
  assign y10123 = ~1'b0 ;
  assign y10124 = n24359 ;
  assign y10125 = n24361 ;
  assign y10126 = ~n24366 ;
  assign y10127 = n24370 ;
  assign y10128 = n24371 ;
  assign y10129 = ~n24373 ;
  assign y10130 = n24377 ;
  assign y10131 = ~1'b0 ;
  assign y10132 = 1'b0 ;
  assign y10133 = n24378 ;
  assign y10134 = n24379 ;
  assign y10135 = ~n24383 ;
  assign y10136 = ~1'b0 ;
  assign y10137 = ~n24387 ;
  assign y10138 = ~n24390 ;
  assign y10139 = ~n24393 ;
  assign y10140 = ~n24396 ;
  assign y10141 = ~1'b0 ;
  assign y10142 = ~n24399 ;
  assign y10143 = n24401 ;
  assign y10144 = n24404 ;
  assign y10145 = n24405 ;
  assign y10146 = ~n24410 ;
  assign y10147 = ~1'b0 ;
  assign y10148 = ~n24414 ;
  assign y10149 = ~n24419 ;
  assign y10150 = ~1'b0 ;
  assign y10151 = ~n24422 ;
  assign y10152 = n24423 ;
  assign y10153 = ~1'b0 ;
  assign y10154 = ~n24424 ;
  assign y10155 = n24426 ;
  assign y10156 = ~1'b0 ;
  assign y10157 = ~1'b0 ;
  assign y10158 = n24429 ;
  assign y10159 = ~1'b0 ;
  assign y10160 = n24430 ;
  assign y10161 = n24433 ;
  assign y10162 = ~n24434 ;
  assign y10163 = ~1'b0 ;
  assign y10164 = ~1'b0 ;
  assign y10165 = n24436 ;
  assign y10166 = ~n24438 ;
  assign y10167 = n24441 ;
  assign y10168 = ~n24444 ;
  assign y10169 = n24445 ;
  assign y10170 = ~n24446 ;
  assign y10171 = ~n11927 ;
  assign y10172 = n24448 ;
  assign y10173 = ~n9538 ;
  assign y10174 = ~n24453 ;
  assign y10175 = ~n24457 ;
  assign y10176 = ~1'b0 ;
  assign y10177 = ~n24460 ;
  assign y10178 = n24467 ;
  assign y10179 = n24469 ;
  assign y10180 = n24470 ;
  assign y10181 = n9314 ;
  assign y10182 = ~n24472 ;
  assign y10183 = n2853 ;
  assign y10184 = n24474 ;
  assign y10185 = n24476 ;
  assign y10186 = ~n24487 ;
  assign y10187 = ~n24492 ;
  assign y10188 = ~n24495 ;
  assign y10189 = ~n24500 ;
  assign y10190 = ~1'b0 ;
  assign y10191 = n24502 ;
  assign y10192 = ~n24506 ;
  assign y10193 = ~n24510 ;
  assign y10194 = n9068 ;
  assign y10195 = ~1'b0 ;
  assign y10196 = ~n24512 ;
  assign y10197 = n15377 ;
  assign y10198 = ~n24514 ;
  assign y10199 = ~1'b0 ;
  assign y10200 = n24515 ;
  assign y10201 = ~1'b0 ;
  assign y10202 = ~1'b0 ;
  assign y10203 = ~n10791 ;
  assign y10204 = ~n11725 ;
  assign y10205 = n24516 ;
  assign y10206 = n24517 ;
  assign y10207 = n24518 ;
  assign y10208 = n24521 ;
  assign y10209 = ~n24522 ;
  assign y10210 = ~1'b0 ;
  assign y10211 = ~n24527 ;
  assign y10212 = ~1'b0 ;
  assign y10213 = ~1'b0 ;
  assign y10214 = n24531 ;
  assign y10215 = ~n24533 ;
  assign y10216 = ~n24535 ;
  assign y10217 = ~n24540 ;
  assign y10218 = ~n24541 ;
  assign y10219 = n24543 ;
  assign y10220 = ~1'b0 ;
  assign y10221 = n24546 ;
  assign y10222 = ~n24553 ;
  assign y10223 = ~n24556 ;
  assign y10224 = n24557 ;
  assign y10225 = ~n24558 ;
  assign y10226 = ~n24559 ;
  assign y10227 = ~n24564 ;
  assign y10228 = ~1'b0 ;
  assign y10229 = n24568 ;
  assign y10230 = ~n24569 ;
  assign y10231 = n24570 ;
  assign y10232 = ~n24571 ;
  assign y10233 = n24575 ;
  assign y10234 = ~n24577 ;
  assign y10235 = ~1'b0 ;
  assign y10236 = n24579 ;
  assign y10237 = n24581 ;
  assign y10238 = n24583 ;
  assign y10239 = ~n24586 ;
  assign y10240 = ~n24591 ;
  assign y10241 = n24597 ;
  assign y10242 = ~n24600 ;
  assign y10243 = ~1'b0 ;
  assign y10244 = ~n24602 ;
  assign y10245 = ~n24604 ;
  assign y10246 = n16346 ;
  assign y10247 = ~n24605 ;
  assign y10248 = n24607 ;
  assign y10249 = ~n24609 ;
  assign y10250 = ~n9788 ;
  assign y10251 = ~n11682 ;
  assign y10252 = ~n24615 ;
  assign y10253 = n24619 ;
  assign y10254 = ~n24621 ;
  assign y10255 = n24630 ;
  assign y10256 = ~1'b0 ;
  assign y10257 = n24632 ;
  assign y10258 = ~1'b0 ;
  assign y10259 = n24635 ;
  assign y10260 = ~n24640 ;
  assign y10261 = ~n24641 ;
  assign y10262 = ~n24643 ;
  assign y10263 = ~1'b0 ;
  assign y10264 = n24649 ;
  assign y10265 = ~n24652 ;
  assign y10266 = ~n24654 ;
  assign y10267 = ~n24656 ;
  assign y10268 = ~n24657 ;
  assign y10269 = n24659 ;
  assign y10270 = ~n24660 ;
  assign y10271 = ~n24661 ;
  assign y10272 = ~1'b0 ;
  assign y10273 = ~n24666 ;
  assign y10274 = n24667 ;
  assign y10275 = n24672 ;
  assign y10276 = n24673 ;
  assign y10277 = ~n24674 ;
  assign y10278 = ~n24676 ;
  assign y10279 = n24677 ;
  assign y10280 = ~1'b0 ;
  assign y10281 = ~n24678 ;
  assign y10282 = n11374 ;
  assign y10283 = ~n24679 ;
  assign y10284 = n24684 ;
  assign y10285 = n24686 ;
  assign y10286 = n24689 ;
  assign y10287 = n11863 ;
  assign y10288 = n24693 ;
  assign y10289 = n24694 ;
  assign y10290 = 1'b0 ;
  assign y10291 = ~1'b0 ;
  assign y10292 = ~1'b0 ;
  assign y10293 = ~n24696 ;
  assign y10294 = ~1'b0 ;
  assign y10295 = ~1'b0 ;
  assign y10296 = n24699 ;
  assign y10297 = n24700 ;
  assign y10298 = ~1'b0 ;
  assign y10299 = n24702 ;
  assign y10300 = ~n24705 ;
  assign y10301 = ~1'b0 ;
  assign y10302 = n24707 ;
  assign y10303 = ~1'b0 ;
  assign y10304 = ~n24712 ;
  assign y10305 = n1430 ;
  assign y10306 = ~n24714 ;
  assign y10307 = n8004 ;
  assign y10308 = ~1'b0 ;
  assign y10309 = n24715 ;
  assign y10310 = ~1'b0 ;
  assign y10311 = n24720 ;
  assign y10312 = ~1'b0 ;
  assign y10313 = n24721 ;
  assign y10314 = ~1'b0 ;
  assign y10315 = n24722 ;
  assign y10316 = n24727 ;
  assign y10317 = n24729 ;
  assign y10318 = ~1'b0 ;
  assign y10319 = ~n24731 ;
  assign y10320 = ~1'b0 ;
  assign y10321 = n24735 ;
  assign y10322 = ~n24740 ;
  assign y10323 = ~n24741 ;
  assign y10324 = n24744 ;
  assign y10325 = ~1'b0 ;
  assign y10326 = n24747 ;
  assign y10327 = ~1'b0 ;
  assign y10328 = n24748 ;
  assign y10329 = n24749 ;
  assign y10330 = n24751 ;
  assign y10331 = n24754 ;
  assign y10332 = n24755 ;
  assign y10333 = n1123 ;
  assign y10334 = n24756 ;
  assign y10335 = ~1'b0 ;
  assign y10336 = ~n24758 ;
  assign y10337 = ~n24761 ;
  assign y10338 = n24763 ;
  assign y10339 = n24765 ;
  assign y10340 = ~n24766 ;
  assign y10341 = n24768 ;
  assign y10342 = n24771 ;
  assign y10343 = ~n24775 ;
  assign y10344 = n24777 ;
  assign y10345 = ~1'b0 ;
  assign y10346 = n24779 ;
  assign y10347 = n24787 ;
  assign y10348 = n24790 ;
  assign y10349 = ~n24794 ;
  assign y10350 = n24796 ;
  assign y10351 = n24797 ;
  assign y10352 = ~n24799 ;
  assign y10353 = n24802 ;
  assign y10354 = ~1'b0 ;
  assign y10355 = ~1'b0 ;
  assign y10356 = ~n24808 ;
  assign y10357 = ~n24810 ;
  assign y10358 = n24812 ;
  assign y10359 = ~n24813 ;
  assign y10360 = ~n24819 ;
  assign y10361 = ~n24820 ;
  assign y10362 = n24823 ;
  assign y10363 = ~n24825 ;
  assign y10364 = ~1'b0 ;
  assign y10365 = ~n24827 ;
  assign y10366 = ~n24828 ;
  assign y10367 = ~1'b0 ;
  assign y10368 = n24831 ;
  assign y10369 = ~1'b0 ;
  assign y10370 = ~n24832 ;
  assign y10371 = ~1'b0 ;
  assign y10372 = n24834 ;
  assign y10373 = ~n24835 ;
  assign y10374 = ~1'b0 ;
  assign y10375 = ~n24837 ;
  assign y10376 = ~n24839 ;
  assign y10377 = n24841 ;
  assign y10378 = ~n24847 ;
  assign y10379 = ~n24848 ;
  assign y10380 = ~n24849 ;
  assign y10381 = ~n24852 ;
  assign y10382 = ~1'b0 ;
  assign y10383 = n24856 ;
  assign y10384 = ~1'b0 ;
  assign y10385 = ~1'b0 ;
  assign y10386 = n24857 ;
  assign y10387 = ~n24862 ;
  assign y10388 = n24865 ;
  assign y10389 = ~1'b0 ;
  assign y10390 = ~1'b0 ;
  assign y10391 = n24866 ;
  assign y10392 = ~n24868 ;
  assign y10393 = n24869 ;
  assign y10394 = ~1'b0 ;
  assign y10395 = n5933 ;
  assign y10396 = ~n24870 ;
  assign y10397 = ~n24871 ;
  assign y10398 = n24873 ;
  assign y10399 = n24875 ;
  assign y10400 = ~n24880 ;
  assign y10401 = n24887 ;
  assign y10402 = 1'b0 ;
  assign y10403 = ~n24892 ;
  assign y10404 = n24897 ;
  assign y10405 = ~n22970 ;
  assign y10406 = n24898 ;
  assign y10407 = n4737 ;
  assign y10408 = n24899 ;
  assign y10409 = n24900 ;
  assign y10410 = ~n24902 ;
  assign y10411 = ~1'b0 ;
  assign y10412 = ~n24905 ;
  assign y10413 = ~n1160 ;
  assign y10414 = n24907 ;
  assign y10415 = ~1'b0 ;
  assign y10416 = ~1'b0 ;
  assign y10417 = ~1'b0 ;
  assign y10418 = ~1'b0 ;
  assign y10419 = n24910 ;
  assign y10420 = n24912 ;
  assign y10421 = n24913 ;
  assign y10422 = n24916 ;
  assign y10423 = ~n24919 ;
  assign y10424 = ~n643 ;
  assign y10425 = n24920 ;
  assign y10426 = n24922 ;
  assign y10427 = ~n24924 ;
  assign y10428 = n24926 ;
  assign y10429 = n24936 ;
  assign y10430 = n24938 ;
  assign y10431 = n8562 ;
  assign y10432 = ~n24940 ;
  assign y10433 = n24941 ;
  assign y10434 = ~n24946 ;
  assign y10435 = ~1'b0 ;
  assign y10436 = ~1'b0 ;
  assign y10437 = ~n24950 ;
  assign y10438 = ~n24953 ;
  assign y10439 = n24954 ;
  assign y10440 = ~1'b0 ;
  assign y10441 = ~n24956 ;
  assign y10442 = n24957 ;
  assign y10443 = ~n24962 ;
  assign y10444 = n24963 ;
  assign y10445 = 1'b0 ;
  assign y10446 = n24965 ;
  assign y10447 = 1'b0 ;
  assign y10448 = ~n24966 ;
  assign y10449 = ~1'b0 ;
  assign y10450 = n24969 ;
  assign y10451 = ~n24970 ;
  assign y10452 = ~n24973 ;
  assign y10453 = ~n24974 ;
  assign y10454 = ~n24976 ;
  assign y10455 = ~n24978 ;
  assign y10456 = n24979 ;
  assign y10457 = ~1'b0 ;
  assign y10458 = ~n24984 ;
  assign y10459 = n24987 ;
  assign y10460 = ~n24989 ;
  assign y10461 = ~1'b0 ;
  assign y10462 = ~1'b0 ;
  assign y10463 = ~n24996 ;
  assign y10464 = n25002 ;
  assign y10465 = 1'b0 ;
  assign y10466 = n25003 ;
  assign y10467 = n25004 ;
  assign y10468 = n25016 ;
  assign y10469 = n25017 ;
  assign y10470 = n25019 ;
  assign y10471 = n25022 ;
  assign y10472 = ~1'b0 ;
  assign y10473 = ~n25027 ;
  assign y10474 = n25030 ;
  assign y10475 = ~1'b0 ;
  assign y10476 = n25033 ;
  assign y10477 = ~n6053 ;
  assign y10478 = n25036 ;
  assign y10479 = ~n25043 ;
  assign y10480 = ~1'b0 ;
  assign y10481 = ~1'b0 ;
  assign y10482 = ~n25048 ;
  assign y10483 = ~n25050 ;
  assign y10484 = ~n25051 ;
  assign y10485 = ~1'b0 ;
  assign y10486 = n25058 ;
  assign y10487 = ~n25061 ;
  assign y10488 = n25063 ;
  assign y10489 = ~n25066 ;
  assign y10490 = ~n25068 ;
  assign y10491 = ~n25069 ;
  assign y10492 = ~n25071 ;
  assign y10493 = ~n25072 ;
  assign y10494 = ~n25073 ;
  assign y10495 = n25075 ;
  assign y10496 = n25078 ;
  assign y10497 = n25081 ;
  assign y10498 = n25085 ;
  assign y10499 = n25089 ;
  assign y10500 = ~n25091 ;
  assign y10501 = 1'b0 ;
  assign y10502 = n25093 ;
  assign y10503 = ~n25096 ;
  assign y10504 = ~n25100 ;
  assign y10505 = ~n25101 ;
  assign y10506 = n25103 ;
  assign y10507 = n25109 ;
  assign y10508 = n25111 ;
  assign y10509 = n25113 ;
  assign y10510 = ~n25115 ;
  assign y10511 = ~n25117 ;
  assign y10512 = ~n25118 ;
  assign y10513 = ~1'b0 ;
  assign y10514 = n25119 ;
  assign y10515 = ~n9752 ;
  assign y10516 = ~n25121 ;
  assign y10517 = ~n25122 ;
  assign y10518 = ~n25124 ;
  assign y10519 = ~n25126 ;
  assign y10520 = n19075 ;
  assign y10521 = ~n25128 ;
  assign y10522 = ~n3046 ;
  assign y10523 = ~1'b0 ;
  assign y10524 = n25129 ;
  assign y10525 = ~n25133 ;
  assign y10526 = n25134 ;
  assign y10527 = ~n25137 ;
  assign y10528 = ~1'b0 ;
  assign y10529 = ~1'b0 ;
  assign y10530 = ~1'b0 ;
  assign y10531 = ~n25139 ;
  assign y10532 = ~n25150 ;
  assign y10533 = ~n25152 ;
  assign y10534 = ~n25153 ;
  assign y10535 = ~n25156 ;
  assign y10536 = n25158 ;
  assign y10537 = ~1'b0 ;
  assign y10538 = n25160 ;
  assign y10539 = ~1'b0 ;
  assign y10540 = ~1'b0 ;
  assign y10541 = ~n25162 ;
  assign y10542 = ~1'b0 ;
  assign y10543 = n25163 ;
  assign y10544 = ~n4235 ;
  assign y10545 = n25167 ;
  assign y10546 = ~n25169 ;
  assign y10547 = ~n25170 ;
  assign y10548 = ~n25171 ;
  assign y10549 = n25173 ;
  assign y10550 = ~1'b0 ;
  assign y10551 = n25174 ;
  assign y10552 = n25175 ;
  assign y10553 = ~n25176 ;
  assign y10554 = ~n25177 ;
  assign y10555 = n25180 ;
  assign y10556 = n25181 ;
  assign y10557 = ~n25183 ;
  assign y10558 = n17292 ;
  assign y10559 = ~1'b0 ;
  assign y10560 = n25184 ;
  assign y10561 = ~n25186 ;
  assign y10562 = ~n25187 ;
  assign y10563 = n11177 ;
  assign y10564 = n25190 ;
  assign y10565 = n25191 ;
  assign y10566 = n25193 ;
  assign y10567 = ~1'b0 ;
  assign y10568 = n25197 ;
  assign y10569 = ~1'b0 ;
  assign y10570 = ~n25199 ;
  assign y10571 = n8086 ;
  assign y10572 = ~n25200 ;
  assign y10573 = n16466 ;
  assign y10574 = ~n25202 ;
  assign y10575 = n20936 ;
  assign y10576 = ~n25204 ;
  assign y10577 = ~n25206 ;
  assign y10578 = ~1'b0 ;
  assign y10579 = ~1'b0 ;
  assign y10580 = ~n25209 ;
  assign y10581 = n25212 ;
  assign y10582 = ~n25213 ;
  assign y10583 = ~n25214 ;
  assign y10584 = ~1'b0 ;
  assign y10585 = ~n25216 ;
  assign y10586 = n25217 ;
  assign y10587 = ~n25221 ;
  assign y10588 = ~1'b0 ;
  assign y10589 = ~n25223 ;
  assign y10590 = ~n25224 ;
  assign y10591 = ~n25226 ;
  assign y10592 = n25229 ;
  assign y10593 = ~n25230 ;
  assign y10594 = ~1'b0 ;
  assign y10595 = n25232 ;
  assign y10596 = 1'b0 ;
  assign y10597 = ~1'b0 ;
  assign y10598 = ~1'b0 ;
  assign y10599 = ~n25234 ;
  assign y10600 = ~1'b0 ;
  assign y10601 = ~1'b0 ;
  assign y10602 = n25235 ;
  assign y10603 = ~n25236 ;
  assign y10604 = ~1'b0 ;
  assign y10605 = n25238 ;
  assign y10606 = n25239 ;
  assign y10607 = n25242 ;
  assign y10608 = ~n25244 ;
  assign y10609 = ~n25246 ;
  assign y10610 = n25251 ;
  assign y10611 = ~n25253 ;
  assign y10612 = n25255 ;
  assign y10613 = ~1'b0 ;
  assign y10614 = ~1'b0 ;
  assign y10615 = ~x78 ;
  assign y10616 = n25257 ;
  assign y10617 = ~n25261 ;
  assign y10618 = ~n25263 ;
  assign y10619 = ~n25264 ;
  assign y10620 = ~n25267 ;
  assign y10621 = n25268 ;
  assign y10622 = n25269 ;
  assign y10623 = ~n25270 ;
  assign y10624 = n25272 ;
  assign y10625 = n25274 ;
  assign y10626 = n25278 ;
  assign y10627 = n1678 ;
  assign y10628 = n25279 ;
  assign y10629 = ~n25283 ;
  assign y10630 = ~n25285 ;
  assign y10631 = ~n25290 ;
  assign y10632 = ~1'b0 ;
  assign y10633 = n25291 ;
  assign y10634 = ~n25292 ;
  assign y10635 = n25294 ;
  assign y10636 = n25295 ;
  assign y10637 = ~n25296 ;
  assign y10638 = n25301 ;
  assign y10639 = n25303 ;
  assign y10640 = ~1'b0 ;
  assign y10641 = ~1'b0 ;
  assign y10642 = ~1'b0 ;
  assign y10643 = ~n25310 ;
  assign y10644 = ~n25314 ;
  assign y10645 = ~n25316 ;
  assign y10646 = n25317 ;
  assign y10647 = n25318 ;
  assign y10648 = ~n25325 ;
  assign y10649 = ~n25326 ;
  assign y10650 = n25334 ;
  assign y10651 = ~n25335 ;
  assign y10652 = 1'b0 ;
  assign y10653 = n25336 ;
  assign y10654 = ~1'b0 ;
  assign y10655 = n25337 ;
  assign y10656 = ~1'b0 ;
  assign y10657 = n25338 ;
  assign y10658 = ~n25339 ;
  assign y10659 = n25340 ;
  assign y10660 = ~1'b0 ;
  assign y10661 = n25343 ;
  assign y10662 = n25345 ;
  assign y10663 = n25346 ;
  assign y10664 = ~1'b0 ;
  assign y10665 = ~n25355 ;
  assign y10666 = ~n25358 ;
  assign y10667 = n25359 ;
  assign y10668 = n25364 ;
  assign y10669 = n25367 ;
  assign y10670 = ~n25371 ;
  assign y10671 = ~n25375 ;
  assign y10672 = ~1'b0 ;
  assign y10673 = n25377 ;
  assign y10674 = n25378 ;
  assign y10675 = n25383 ;
  assign y10676 = n637 ;
  assign y10677 = ~n25384 ;
  assign y10678 = ~n23570 ;
  assign y10679 = n25386 ;
  assign y10680 = ~1'b0 ;
  assign y10681 = ~n25388 ;
  assign y10682 = ~1'b0 ;
  assign y10683 = ~1'b0 ;
  assign y10684 = n17066 ;
  assign y10685 = ~n25389 ;
  assign y10686 = n25390 ;
  assign y10687 = ~n25391 ;
  assign y10688 = n25394 ;
  assign y10689 = n25396 ;
  assign y10690 = ~n25398 ;
  assign y10691 = n17484 ;
  assign y10692 = ~n25399 ;
  assign y10693 = ~n25401 ;
  assign y10694 = n25402 ;
  assign y10695 = ~n25405 ;
  assign y10696 = ~n25406 ;
  assign y10697 = n25407 ;
  assign y10698 = ~n25410 ;
  assign y10699 = ~n25413 ;
  assign y10700 = n25417 ;
  assign y10701 = ~1'b0 ;
  assign y10702 = ~1'b0 ;
  assign y10703 = n25423 ;
  assign y10704 = ~n25425 ;
  assign y10705 = n25430 ;
  assign y10706 = ~n25431 ;
  assign y10707 = ~1'b0 ;
  assign y10708 = n25432 ;
  assign y10709 = ~1'b0 ;
  assign y10710 = n25435 ;
  assign y10711 = ~1'b0 ;
  assign y10712 = ~n25436 ;
  assign y10713 = n25439 ;
  assign y10714 = n25443 ;
  assign y10715 = ~n850 ;
  assign y10716 = ~n25445 ;
  assign y10717 = ~1'b0 ;
  assign y10718 = ~1'b0 ;
  assign y10719 = ~1'b0 ;
  assign y10720 = ~n25449 ;
  assign y10721 = ~n18160 ;
  assign y10722 = n25450 ;
  assign y10723 = ~n25451 ;
  assign y10724 = ~n25453 ;
  assign y10725 = n25459 ;
  assign y10726 = ~n25460 ;
  assign y10727 = ~n25461 ;
  assign y10728 = ~1'b0 ;
  assign y10729 = ~n25463 ;
  assign y10730 = n25465 ;
  assign y10731 = ~n25467 ;
  assign y10732 = ~n25468 ;
  assign y10733 = n25470 ;
  assign y10734 = n25473 ;
  assign y10735 = ~n25477 ;
  assign y10736 = ~1'b0 ;
  assign y10737 = ~1'b0 ;
  assign y10738 = ~n25481 ;
  assign y10739 = n25482 ;
  assign y10740 = ~n25484 ;
  assign y10741 = ~x98 ;
  assign y10742 = ~n25486 ;
  assign y10743 = ~1'b0 ;
  assign y10744 = ~n25488 ;
  assign y10745 = n25490 ;
  assign y10746 = n25492 ;
  assign y10747 = n25494 ;
  assign y10748 = ~1'b0 ;
  assign y10749 = ~n25498 ;
  assign y10750 = n25503 ;
  assign y10751 = ~n25506 ;
  assign y10752 = ~1'b0 ;
  assign y10753 = n14317 ;
  assign y10754 = n25509 ;
  assign y10755 = n25510 ;
  assign y10756 = ~n25512 ;
  assign y10757 = ~n25515 ;
  assign y10758 = ~1'b0 ;
  assign y10759 = n4839 ;
  assign y10760 = ~n25516 ;
  assign y10761 = ~1'b0 ;
  assign y10762 = ~n25517 ;
  assign y10763 = n25518 ;
  assign y10764 = ~n25519 ;
  assign y10765 = n25524 ;
  assign y10766 = ~1'b0 ;
  assign y10767 = ~1'b0 ;
  assign y10768 = ~n25525 ;
  assign y10769 = ~n25527 ;
  assign y10770 = ~n25530 ;
  assign y10771 = ~n25531 ;
  assign y10772 = ~n25533 ;
  assign y10773 = n25534 ;
  assign y10774 = ~1'b0 ;
  assign y10775 = ~n25536 ;
  assign y10776 = ~1'b0 ;
  assign y10777 = ~1'b0 ;
  assign y10778 = ~n25537 ;
  assign y10779 = n25547 ;
  assign y10780 = n25552 ;
  assign y10781 = ~n25559 ;
  assign y10782 = n25563 ;
  assign y10783 = ~n25565 ;
  assign y10784 = ~n25568 ;
  assign y10785 = ~1'b0 ;
  assign y10786 = ~1'b0 ;
  assign y10787 = ~n25572 ;
  assign y10788 = ~n25574 ;
  assign y10789 = ~n25577 ;
  assign y10790 = ~n25580 ;
  assign y10791 = ~n661 ;
  assign y10792 = ~1'b0 ;
  assign y10793 = ~n25584 ;
  assign y10794 = ~n25585 ;
  assign y10795 = n25586 ;
  assign y10796 = ~1'b0 ;
  assign y10797 = ~n25589 ;
  assign y10798 = ~n25592 ;
  assign y10799 = ~n25593 ;
  assign y10800 = ~n25596 ;
  assign y10801 = ~n25598 ;
  assign y10802 = n25599 ;
  assign y10803 = ~n25601 ;
  assign y10804 = ~n25604 ;
  assign y10805 = n25605 ;
  assign y10806 = n25607 ;
  assign y10807 = n25608 ;
  assign y10808 = ~1'b0 ;
  assign y10809 = ~n25609 ;
  assign y10810 = ~n25610 ;
  assign y10811 = n25613 ;
  assign y10812 = ~n5155 ;
  assign y10813 = ~1'b0 ;
  assign y10814 = ~1'b0 ;
  assign y10815 = ~n25618 ;
  assign y10816 = n25621 ;
  assign y10817 = ~1'b0 ;
  assign y10818 = n25623 ;
  assign y10819 = ~n25625 ;
  assign y10820 = ~n25626 ;
  assign y10821 = ~n25631 ;
  assign y10822 = ~1'b0 ;
  assign y10823 = ~1'b0 ;
  assign y10824 = ~1'b0 ;
  assign y10825 = n25633 ;
  assign y10826 = ~1'b0 ;
  assign y10827 = ~n25637 ;
  assign y10828 = ~1'b0 ;
  assign y10829 = n25638 ;
  assign y10830 = ~n25641 ;
  assign y10831 = ~n25642 ;
  assign y10832 = ~n25646 ;
  assign y10833 = ~1'b0 ;
  assign y10834 = 1'b0 ;
  assign y10835 = ~n25649 ;
  assign y10836 = n25653 ;
  assign y10837 = ~1'b0 ;
  assign y10838 = ~1'b0 ;
  assign y10839 = ~n25655 ;
  assign y10840 = n25658 ;
  assign y10841 = n25661 ;
  assign y10842 = ~1'b0 ;
  assign y10843 = n25662 ;
  assign y10844 = n25664 ;
  assign y10845 = ~n25665 ;
  assign y10846 = ~n25666 ;
  assign y10847 = ~1'b0 ;
  assign y10848 = ~1'b0 ;
  assign y10849 = n25667 ;
  assign y10850 = n25668 ;
  assign y10851 = n25669 ;
  assign y10852 = ~n25672 ;
  assign y10853 = n25673 ;
  assign y10854 = ~n16445 ;
  assign y10855 = ~1'b0 ;
  assign y10856 = n25674 ;
  assign y10857 = n25676 ;
  assign y10858 = ~n25678 ;
  assign y10859 = ~n25679 ;
  assign y10860 = ~n25680 ;
  assign y10861 = ~n25688 ;
  assign y10862 = ~n25689 ;
  assign y10863 = n25690 ;
  assign y10864 = ~1'b0 ;
  assign y10865 = n25694 ;
  assign y10866 = n25700 ;
  assign y10867 = ~n25702 ;
  assign y10868 = n25705 ;
  assign y10869 = n25707 ;
  assign y10870 = n25710 ;
  assign y10871 = n25712 ;
  assign y10872 = ~n25714 ;
  assign y10873 = ~1'b0 ;
  assign y10874 = ~1'b0 ;
  assign y10875 = ~n25715 ;
  assign y10876 = n25720 ;
  assign y10877 = n25723 ;
  assign y10878 = ~n12138 ;
  assign y10879 = ~1'b0 ;
  assign y10880 = n25724 ;
  assign y10881 = n25725 ;
  assign y10882 = ~n25726 ;
  assign y10883 = ~n25727 ;
  assign y10884 = ~n25729 ;
  assign y10885 = ~n25731 ;
  assign y10886 = n25733 ;
  assign y10887 = ~1'b0 ;
  assign y10888 = n25734 ;
  assign y10889 = n25742 ;
  assign y10890 = ~n6286 ;
  assign y10891 = ~n25743 ;
  assign y10892 = ~1'b0 ;
  assign y10893 = ~n25745 ;
  assign y10894 = ~n25749 ;
  assign y10895 = n25750 ;
  assign y10896 = ~n25757 ;
  assign y10897 = n25762 ;
  assign y10898 = n25764 ;
  assign y10899 = ~n25767 ;
  assign y10900 = n25768 ;
  assign y10901 = ~1'b0 ;
  assign y10902 = ~1'b0 ;
  assign y10903 = ~1'b0 ;
  assign y10904 = n25769 ;
  assign y10905 = n25770 ;
  assign y10906 = ~n25772 ;
  assign y10907 = ~n25774 ;
  assign y10908 = n25775 ;
  assign y10909 = n25777 ;
  assign y10910 = ~n25779 ;
  assign y10911 = ~1'b0 ;
  assign y10912 = ~n25782 ;
  assign y10913 = n25783 ;
  assign y10914 = ~1'b0 ;
  assign y10915 = ~n25785 ;
  assign y10916 = ~n25787 ;
  assign y10917 = n25789 ;
  assign y10918 = n25791 ;
  assign y10919 = n25793 ;
  assign y10920 = ~1'b0 ;
  assign y10921 = ~1'b0 ;
  assign y10922 = ~1'b0 ;
  assign y10923 = ~n25794 ;
  assign y10924 = n25795 ;
  assign y10925 = ~n25797 ;
  assign y10926 = ~n25801 ;
  assign y10927 = n25802 ;
  assign y10928 = n25803 ;
  assign y10929 = ~1'b0 ;
  assign y10930 = ~1'b0 ;
  assign y10931 = n25805 ;
  assign y10932 = ~1'b0 ;
  assign y10933 = ~n25807 ;
  assign y10934 = n25809 ;
  assign y10935 = ~n25810 ;
  assign y10936 = ~n25811 ;
  assign y10937 = ~n25815 ;
  assign y10938 = ~n25816 ;
  assign y10939 = ~1'b0 ;
  assign y10940 = n25817 ;
  assign y10941 = ~n25819 ;
  assign y10942 = ~n25826 ;
  assign y10943 = ~1'b0 ;
  assign y10944 = n25830 ;
  assign y10945 = ~n25831 ;
  assign y10946 = n25833 ;
  assign y10947 = ~n25834 ;
  assign y10948 = ~n25839 ;
  assign y10949 = ~n25840 ;
  assign y10950 = ~n25841 ;
  assign y10951 = ~n25843 ;
  assign y10952 = ~n25846 ;
  assign y10953 = n25847 ;
  assign y10954 = ~n25850 ;
  assign y10955 = ~1'b0 ;
  assign y10956 = ~n25852 ;
  assign y10957 = n25856 ;
  assign y10958 = n25857 ;
  assign y10959 = n25860 ;
  assign y10960 = ~1'b0 ;
  assign y10961 = ~1'b0 ;
  assign y10962 = ~1'b0 ;
  assign y10963 = ~n19053 ;
  assign y10964 = ~1'b0 ;
  assign y10965 = n25865 ;
  assign y10966 = ~1'b0 ;
  assign y10967 = n25868 ;
  assign y10968 = ~n25872 ;
  assign y10969 = n25874 ;
  assign y10970 = ~1'b0 ;
  assign y10971 = n25876 ;
  assign y10972 = n25881 ;
  assign y10973 = ~n25885 ;
  assign y10974 = n25887 ;
  assign y10975 = ~n25891 ;
  assign y10976 = n25894 ;
  assign y10977 = ~n25896 ;
  assign y10978 = n25897 ;
  assign y10979 = ~n25900 ;
  assign y10980 = ~n25903 ;
  assign y10981 = ~1'b0 ;
  assign y10982 = ~n25904 ;
  assign y10983 = n25906 ;
  assign y10984 = n25908 ;
  assign y10985 = n25912 ;
  assign y10986 = ~n25913 ;
  assign y10987 = ~n25920 ;
  assign y10988 = n25922 ;
  assign y10989 = ~1'b0 ;
  assign y10990 = n25927 ;
  assign y10991 = n25928 ;
  assign y10992 = ~n25930 ;
  assign y10993 = n25931 ;
  assign y10994 = n25932 ;
  assign y10995 = ~n25933 ;
  assign y10996 = ~n25934 ;
  assign y10997 = n25940 ;
  assign y10998 = ~n25942 ;
  assign y10999 = n25944 ;
  assign y11000 = ~n1960 ;
  assign y11001 = ~1'b0 ;
  assign y11002 = n25946 ;
  assign y11003 = ~1'b0 ;
  assign y11004 = n9764 ;
  assign y11005 = ~n25960 ;
  assign y11006 = ~n25963 ;
  assign y11007 = n25964 ;
  assign y11008 = ~n25966 ;
  assign y11009 = n25969 ;
  assign y11010 = n25972 ;
  assign y11011 = 1'b0 ;
  assign y11012 = n25973 ;
  assign y11013 = ~1'b0 ;
  assign y11014 = ~n25978 ;
  assign y11015 = n25981 ;
  assign y11016 = n25982 ;
  assign y11017 = n25986 ;
  assign y11018 = n25990 ;
  assign y11019 = n25991 ;
  assign y11020 = n25993 ;
  assign y11021 = ~n25996 ;
  assign y11022 = n1118 ;
  assign y11023 = ~n25997 ;
  assign y11024 = ~n26000 ;
  assign y11025 = ~n26003 ;
  assign y11026 = ~n26006 ;
  assign y11027 = n26011 ;
  assign y11028 = n26014 ;
  assign y11029 = ~n26016 ;
  assign y11030 = ~n26018 ;
  assign y11031 = ~n26020 ;
  assign y11032 = ~n26022 ;
  assign y11033 = n7301 ;
  assign y11034 = ~1'b0 ;
  assign y11035 = n26024 ;
  assign y11036 = n26029 ;
  assign y11037 = n26033 ;
  assign y11038 = n26036 ;
  assign y11039 = n26038 ;
  assign y11040 = n26039 ;
  assign y11041 = n26040 ;
  assign y11042 = n26043 ;
  assign y11043 = ~n26044 ;
  assign y11044 = n26045 ;
  assign y11045 = n26047 ;
  assign y11046 = ~n26054 ;
  assign y11047 = n26055 ;
  assign y11048 = n26057 ;
  assign y11049 = n26061 ;
  assign y11050 = n26063 ;
  assign y11051 = ~n26065 ;
  assign y11052 = ~n26069 ;
  assign y11053 = ~n26070 ;
  assign y11054 = n26079 ;
  assign y11055 = n26081 ;
  assign y11056 = ~n26085 ;
  assign y11057 = ~n26089 ;
  assign y11058 = ~n26090 ;
  assign y11059 = 1'b0 ;
  assign y11060 = n26092 ;
  assign y11061 = ~1'b0 ;
  assign y11062 = ~n26094 ;
  assign y11063 = ~n26099 ;
  assign y11064 = ~n6079 ;
  assign y11065 = ~n26102 ;
  assign y11066 = ~1'b0 ;
  assign y11067 = ~1'b0 ;
  assign y11068 = 1'b0 ;
  assign y11069 = n26106 ;
  assign y11070 = ~n26108 ;
  assign y11071 = ~n26111 ;
  assign y11072 = ~1'b0 ;
  assign y11073 = n26114 ;
  assign y11074 = ~n26119 ;
  assign y11075 = ~n26121 ;
  assign y11076 = ~n26122 ;
  assign y11077 = ~1'b0 ;
  assign y11078 = n26123 ;
  assign y11079 = ~1'b0 ;
  assign y11080 = ~n26124 ;
  assign y11081 = n26127 ;
  assign y11082 = n26132 ;
  assign y11083 = n26133 ;
  assign y11084 = n3640 ;
  assign y11085 = n26135 ;
  assign y11086 = n25635 ;
  assign y11087 = n26136 ;
  assign y11088 = ~n26137 ;
  assign y11089 = n26142 ;
  assign y11090 = ~1'b0 ;
  assign y11091 = ~n1695 ;
  assign y11092 = ~n25225 ;
  assign y11093 = ~n26145 ;
  assign y11094 = ~n9767 ;
  assign y11095 = n26147 ;
  assign y11096 = ~n26149 ;
  assign y11097 = ~1'b0 ;
  assign y11098 = n11430 ;
  assign y11099 = ~1'b0 ;
  assign y11100 = ~n26151 ;
  assign y11101 = ~1'b0 ;
  assign y11102 = ~n26153 ;
  assign y11103 = n26155 ;
  assign y11104 = n26157 ;
  assign y11105 = n26161 ;
  assign y11106 = ~n26165 ;
  assign y11107 = n1288 ;
  assign y11108 = ~n26173 ;
  assign y11109 = n26176 ;
  assign y11110 = ~1'b0 ;
  assign y11111 = n26179 ;
  assign y11112 = ~n26181 ;
  assign y11113 = ~n17171 ;
  assign y11114 = n26183 ;
  assign y11115 = n26186 ;
  assign y11116 = n26195 ;
  assign y11117 = ~n26196 ;
  assign y11118 = ~n6664 ;
  assign y11119 = ~1'b0 ;
  assign y11120 = ~1'b0 ;
  assign y11121 = n26198 ;
  assign y11122 = ~1'b0 ;
  assign y11123 = ~n26201 ;
  assign y11124 = n26203 ;
  assign y11125 = ~n26206 ;
  assign y11126 = ~n26209 ;
  assign y11127 = ~n26211 ;
  assign y11128 = ~1'b0 ;
  assign y11129 = ~1'b0 ;
  assign y11130 = ~1'b0 ;
  assign y11131 = n26214 ;
  assign y11132 = n26216 ;
  assign y11133 = ~1'b0 ;
  assign y11134 = n26219 ;
  assign y11135 = ~n26222 ;
  assign y11136 = ~1'b0 ;
  assign y11137 = ~1'b0 ;
  assign y11138 = ~1'b0 ;
  assign y11139 = ~n26225 ;
  assign y11140 = ~1'b0 ;
  assign y11141 = n26227 ;
  assign y11142 = ~n26228 ;
  assign y11143 = n26230 ;
  assign y11144 = ~n26231 ;
  assign y11145 = ~n26243 ;
  assign y11146 = n12858 ;
  assign y11147 = ~1'b0 ;
  assign y11148 = ~n14269 ;
  assign y11149 = ~n26246 ;
  assign y11150 = ~1'b0 ;
  assign y11151 = n26248 ;
  assign y11152 = ~n26251 ;
  assign y11153 = ~n26252 ;
  assign y11154 = n26253 ;
  assign y11155 = n26254 ;
  assign y11156 = n26255 ;
  assign y11157 = ~1'b0 ;
  assign y11158 = n26257 ;
  assign y11159 = ~n26259 ;
  assign y11160 = n26260 ;
  assign y11161 = n26261 ;
  assign y11162 = ~n26264 ;
  assign y11163 = n26268 ;
  assign y11164 = ~n26272 ;
  assign y11165 = ~1'b0 ;
  assign y11166 = ~n26275 ;
  assign y11167 = n26277 ;
  assign y11168 = n26279 ;
  assign y11169 = ~n26285 ;
  assign y11170 = ~n26287 ;
  assign y11171 = n26288 ;
  assign y11172 = ~n26290 ;
  assign y11173 = n26292 ;
  assign y11174 = ~n26295 ;
  assign y11175 = 1'b0 ;
  assign y11176 = ~n26297 ;
  assign y11177 = ~n26301 ;
  assign y11178 = ~n26303 ;
  assign y11179 = ~1'b0 ;
  assign y11180 = n26304 ;
  assign y11181 = ~n26306 ;
  assign y11182 = ~n26308 ;
  assign y11183 = ~n26309 ;
  assign y11184 = n26310 ;
  assign y11185 = ~n26314 ;
  assign y11186 = n26318 ;
  assign y11187 = ~n26319 ;
  assign y11188 = ~n26325 ;
  assign y11189 = ~n26329 ;
  assign y11190 = ~n26331 ;
  assign y11191 = ~1'b0 ;
  assign y11192 = ~n26333 ;
  assign y11193 = ~n26335 ;
  assign y11194 = ~1'b0 ;
  assign y11195 = ~n26339 ;
  assign y11196 = n26340 ;
  assign y11197 = ~1'b0 ;
  assign y11198 = ~n26342 ;
  assign y11199 = n26346 ;
  assign y11200 = n26348 ;
  assign y11201 = ~n26353 ;
  assign y11202 = n26354 ;
  assign y11203 = n26356 ;
  assign y11204 = ~n26358 ;
  assign y11205 = n26360 ;
  assign y11206 = n26362 ;
  assign y11207 = ~1'b0 ;
  assign y11208 = ~n26365 ;
  assign y11209 = ~n26369 ;
  assign y11210 = ~1'b0 ;
  assign y11211 = n26370 ;
  assign y11212 = ~n26371 ;
  assign y11213 = ~n26373 ;
  assign y11214 = n8095 ;
  assign y11215 = ~n26378 ;
  assign y11216 = ~1'b0 ;
  assign y11217 = ~n26380 ;
  assign y11218 = ~1'b0 ;
  assign y11219 = ~n26385 ;
  assign y11220 = n26390 ;
  assign y11221 = n26393 ;
  assign y11222 = ~n26395 ;
  assign y11223 = n26396 ;
  assign y11224 = ~n26397 ;
  assign y11225 = ~n26401 ;
  assign y11226 = ~1'b0 ;
  assign y11227 = ~n26403 ;
  assign y11228 = ~n26405 ;
  assign y11229 = ~n26409 ;
  assign y11230 = ~1'b0 ;
  assign y11231 = ~n26410 ;
  assign y11232 = ~n26413 ;
  assign y11233 = n26415 ;
  assign y11234 = n26419 ;
  assign y11235 = ~n26420 ;
  assign y11236 = ~n26423 ;
  assign y11237 = ~n26425 ;
  assign y11238 = n26435 ;
  assign y11239 = 1'b0 ;
  assign y11240 = n26436 ;
  assign y11241 = ~n26438 ;
  assign y11242 = ~n18835 ;
  assign y11243 = n26440 ;
  assign y11244 = ~n26441 ;
  assign y11245 = ~n26442 ;
  assign y11246 = n8658 ;
  assign y11247 = n26446 ;
  assign y11248 = n26447 ;
  assign y11249 = ~n26450 ;
  assign y11250 = ~n26452 ;
  assign y11251 = ~1'b0 ;
  assign y11252 = ~n26457 ;
  assign y11253 = ~n26458 ;
  assign y11254 = n26460 ;
  assign y11255 = ~1'b0 ;
  assign y11256 = n26463 ;
  assign y11257 = ~n26466 ;
  assign y11258 = ~1'b0 ;
  assign y11259 = n26468 ;
  assign y11260 = n26469 ;
  assign y11261 = n26473 ;
  assign y11262 = ~n26476 ;
  assign y11263 = ~n26485 ;
  assign y11264 = ~n26487 ;
  assign y11265 = ~1'b0 ;
  assign y11266 = ~1'b0 ;
  assign y11267 = ~n26491 ;
  assign y11268 = ~n26495 ;
  assign y11269 = ~n26496 ;
  assign y11270 = n26500 ;
  assign y11271 = ~n26502 ;
  assign y11272 = ~n26504 ;
  assign y11273 = ~n26505 ;
  assign y11274 = ~n26508 ;
  assign y11275 = ~n26509 ;
  assign y11276 = ~n26510 ;
  assign y11277 = ~n26511 ;
  assign y11278 = n26513 ;
  assign y11279 = ~1'b0 ;
  assign y11280 = n26514 ;
  assign y11281 = ~1'b0 ;
  assign y11282 = ~1'b0 ;
  assign y11283 = ~n26520 ;
  assign y11284 = ~n26522 ;
  assign y11285 = n26523 ;
  assign y11286 = ~n26525 ;
  assign y11287 = n26530 ;
  assign y11288 = n26532 ;
  assign y11289 = ~n26537 ;
  assign y11290 = ~1'b0 ;
  assign y11291 = n26538 ;
  assign y11292 = ~1'b0 ;
  assign y11293 = ~n26540 ;
  assign y11294 = n26541 ;
  assign y11295 = ~n26543 ;
  assign y11296 = n26544 ;
  assign y11297 = ~n26547 ;
  assign y11298 = ~n26550 ;
  assign y11299 = n26552 ;
  assign y11300 = n26553 ;
  assign y11301 = 1'b0 ;
  assign y11302 = n26554 ;
  assign y11303 = ~n26559 ;
  assign y11304 = ~n26562 ;
  assign y11305 = n5935 ;
  assign y11306 = ~n26566 ;
  assign y11307 = n26568 ;
  assign y11308 = ~n26569 ;
  assign y11309 = n6137 ;
  assign y11310 = ~n26571 ;
  assign y11311 = n26576 ;
  assign y11312 = n26577 ;
  assign y11313 = n26578 ;
  assign y11314 = n26580 ;
  assign y11315 = ~n26582 ;
  assign y11316 = ~n26583 ;
  assign y11317 = ~1'b0 ;
  assign y11318 = n26586 ;
  assign y11319 = ~n26589 ;
  assign y11320 = ~1'b0 ;
  assign y11321 = ~n26591 ;
  assign y11322 = ~1'b0 ;
  assign y11323 = ~n26592 ;
  assign y11324 = 1'b0 ;
  assign y11325 = ~n26595 ;
  assign y11326 = ~1'b0 ;
  assign y11327 = ~n26597 ;
  assign y11328 = ~1'b0 ;
  assign y11329 = ~1'b0 ;
  assign y11330 = ~n26600 ;
  assign y11331 = n26602 ;
  assign y11332 = n26608 ;
  assign y11333 = ~n26609 ;
  assign y11334 = n26610 ;
  assign y11335 = n26611 ;
  assign y11336 = n26612 ;
  assign y11337 = ~1'b0 ;
  assign y11338 = ~n26614 ;
  assign y11339 = ~n26616 ;
  assign y11340 = ~n26617 ;
  assign y11341 = ~n26618 ;
  assign y11342 = n26619 ;
  assign y11343 = ~n26620 ;
  assign y11344 = n26621 ;
  assign y11345 = ~n26623 ;
  assign y11346 = ~1'b0 ;
  assign y11347 = ~1'b0 ;
  assign y11348 = n22792 ;
  assign y11349 = ~n26625 ;
  assign y11350 = ~n26627 ;
  assign y11351 = ~n26221 ;
  assign y11352 = ~n26630 ;
  assign y11353 = n26635 ;
  assign y11354 = n26636 ;
  assign y11355 = ~n26637 ;
  assign y11356 = ~1'b0 ;
  assign y11357 = ~1'b0 ;
  assign y11358 = n26641 ;
  assign y11359 = ~1'b0 ;
  assign y11360 = ~n26648 ;
  assign y11361 = n26652 ;
  assign y11362 = ~n26653 ;
  assign y11363 = ~n26654 ;
  assign y11364 = ~n26655 ;
  assign y11365 = ~n26657 ;
  assign y11366 = n26659 ;
  assign y11367 = ~1'b0 ;
  assign y11368 = ~n26661 ;
  assign y11369 = ~1'b0 ;
  assign y11370 = ~n26662 ;
  assign y11371 = ~n26663 ;
  assign y11372 = n26664 ;
  assign y11373 = n26665 ;
  assign y11374 = n26668 ;
  assign y11375 = ~n26672 ;
  assign y11376 = ~n26675 ;
  assign y11377 = ~1'b0 ;
  assign y11378 = ~1'b0 ;
  assign y11379 = ~n26676 ;
  assign y11380 = ~1'b0 ;
  assign y11381 = ~1'b0 ;
  assign y11382 = n26680 ;
  assign y11383 = n26681 ;
  assign y11384 = n26683 ;
  assign y11385 = ~n26686 ;
  assign y11386 = ~1'b0 ;
  assign y11387 = ~1'b0 ;
  assign y11388 = ~1'b0 ;
  assign y11389 = ~1'b0 ;
  assign y11390 = ~1'b0 ;
  assign y11391 = ~n26689 ;
  assign y11392 = n26692 ;
  assign y11393 = ~n26693 ;
  assign y11394 = ~n4610 ;
  assign y11395 = ~n26694 ;
  assign y11396 = ~n26695 ;
  assign y11397 = ~n26700 ;
  assign y11398 = ~1'b0 ;
  assign y11399 = ~1'b0 ;
  assign y11400 = ~n26701 ;
  assign y11401 = n26708 ;
  assign y11402 = ~n14413 ;
  assign y11403 = n26709 ;
  assign y11404 = ~n26712 ;
  assign y11405 = n26715 ;
  assign y11406 = ~n26717 ;
  assign y11407 = ~1'b0 ;
  assign y11408 = ~n26720 ;
  assign y11409 = n26722 ;
  assign y11410 = ~n26724 ;
  assign y11411 = ~n26726 ;
  assign y11412 = n26729 ;
  assign y11413 = n26730 ;
  assign y11414 = ~n26736 ;
  assign y11415 = ~n26739 ;
  assign y11416 = n26741 ;
  assign y11417 = ~1'b0 ;
  assign y11418 = ~1'b0 ;
  assign y11419 = n26742 ;
  assign y11420 = n26744 ;
  assign y11421 = ~n26750 ;
  assign y11422 = ~1'b0 ;
  assign y11423 = ~n26752 ;
  assign y11424 = ~n26753 ;
  assign y11425 = n26754 ;
  assign y11426 = n26758 ;
  assign y11427 = n26762 ;
  assign y11428 = ~n26764 ;
  assign y11429 = n26765 ;
  assign y11430 = ~n26768 ;
  assign y11431 = n26769 ;
  assign y11432 = ~n26770 ;
  assign y11433 = ~n26771 ;
  assign y11434 = ~n26772 ;
  assign y11435 = n26773 ;
  assign y11436 = ~n26776 ;
  assign y11437 = ~n26777 ;
  assign y11438 = n26778 ;
  assign y11439 = n26780 ;
  assign y11440 = ~n26782 ;
  assign y11441 = ~n26786 ;
  assign y11442 = ~n26787 ;
  assign y11443 = ~n26789 ;
  assign y11444 = ~1'b0 ;
  assign y11445 = n2434 ;
  assign y11446 = n26790 ;
  assign y11447 = n26792 ;
  assign y11448 = ~n26795 ;
  assign y11449 = ~1'b0 ;
  assign y11450 = ~1'b0 ;
  assign y11451 = ~n26797 ;
  assign y11452 = ~n26799 ;
  assign y11453 = n26801 ;
  assign y11454 = n26803 ;
  assign y11455 = ~n26804 ;
  assign y11456 = ~n26807 ;
  assign y11457 = ~n26809 ;
  assign y11458 = n26810 ;
  assign y11459 = n26814 ;
  assign y11460 = ~n26819 ;
  assign y11461 = n26821 ;
  assign y11462 = n26823 ;
  assign y11463 = ~1'b0 ;
  assign y11464 = n26824 ;
  assign y11465 = n26825 ;
  assign y11466 = ~n26827 ;
  assign y11467 = ~1'b0 ;
  assign y11468 = ~1'b0 ;
  assign y11469 = ~1'b0 ;
  assign y11470 = ~n26834 ;
  assign y11471 = ~n26837 ;
  assign y11472 = ~1'b0 ;
  assign y11473 = 1'b0 ;
  assign y11474 = n26840 ;
  assign y11475 = n26842 ;
  assign y11476 = n26844 ;
  assign y11477 = n26845 ;
  assign y11478 = ~n26847 ;
  assign y11479 = n26849 ;
  assign y11480 = ~1'b0 ;
  assign y11481 = n26850 ;
  assign y11482 = n26852 ;
  assign y11483 = ~n26856 ;
  assign y11484 = ~n26857 ;
  assign y11485 = n26860 ;
  assign y11486 = n26861 ;
  assign y11487 = n26862 ;
  assign y11488 = ~n21547 ;
  assign y11489 = n26865 ;
  assign y11490 = ~1'b0 ;
  assign y11491 = ~n26867 ;
  assign y11492 = ~1'b0 ;
  assign y11493 = ~n26869 ;
  assign y11494 = ~n26871 ;
  assign y11495 = ~n26876 ;
  assign y11496 = n26877 ;
  assign y11497 = n16001 ;
  assign y11498 = n26878 ;
  assign y11499 = ~n26879 ;
  assign y11500 = ~n26881 ;
  assign y11501 = ~1'b0 ;
  assign y11502 = n26883 ;
  assign y11503 = n26885 ;
  assign y11504 = ~n26886 ;
  assign y11505 = ~1'b0 ;
  assign y11506 = n26889 ;
  assign y11507 = n26892 ;
  assign y11508 = n26894 ;
  assign y11509 = ~n26895 ;
  assign y11510 = n26896 ;
  assign y11511 = n26898 ;
  assign y11512 = ~1'b0 ;
  assign y11513 = n26899 ;
  assign y11514 = ~1'b0 ;
  assign y11515 = n26901 ;
  assign y11516 = n26903 ;
  assign y11517 = n26904 ;
  assign y11518 = n26908 ;
  assign y11519 = ~n26909 ;
  assign y11520 = n26910 ;
  assign y11521 = n26912 ;
  assign y11522 = ~n26913 ;
  assign y11523 = ~n26917 ;
  assign y11524 = n26918 ;
  assign y11525 = ~n26920 ;
  assign y11526 = ~n26923 ;
  assign y11527 = ~1'b0 ;
  assign y11528 = ~n26925 ;
  assign y11529 = n26926 ;
  assign y11530 = ~n26933 ;
  assign y11531 = n26935 ;
  assign y11532 = ~1'b0 ;
  assign y11533 = ~1'b0 ;
  assign y11534 = ~n26936 ;
  assign y11535 = ~n26938 ;
  assign y11536 = n26940 ;
  assign y11537 = ~n26941 ;
  assign y11538 = n25639 ;
  assign y11539 = n26943 ;
  assign y11540 = n26949 ;
  assign y11541 = ~1'b0 ;
  assign y11542 = ~1'b0 ;
  assign y11543 = n26951 ;
  assign y11544 = n26953 ;
  assign y11545 = ~1'b0 ;
  assign y11546 = ~n26956 ;
  assign y11547 = ~n26960 ;
  assign y11548 = n26965 ;
  assign y11549 = ~1'b0 ;
  assign y11550 = n26967 ;
  assign y11551 = n26969 ;
  assign y11552 = n26971 ;
  assign y11553 = ~1'b0 ;
  assign y11554 = n26972 ;
  assign y11555 = n26973 ;
  assign y11556 = ~1'b0 ;
  assign y11557 = n26974 ;
  assign y11558 = ~n26976 ;
  assign y11559 = ~n26980 ;
  assign y11560 = n26982 ;
  assign y11561 = ~n26983 ;
  assign y11562 = ~1'b0 ;
  assign y11563 = n26985 ;
  assign y11564 = n26987 ;
  assign y11565 = n26989 ;
  assign y11566 = n26991 ;
  assign y11567 = n26992 ;
  assign y11568 = ~n850 ;
  assign y11569 = n26993 ;
  assign y11570 = n26994 ;
  assign y11571 = ~n26997 ;
  assign y11572 = n27001 ;
  assign y11573 = n27003 ;
  assign y11574 = ~n27004 ;
  assign y11575 = n27005 ;
  assign y11576 = n27006 ;
  assign y11577 = ~n27008 ;
  assign y11578 = n27009 ;
  assign y11579 = n27010 ;
  assign y11580 = n27016 ;
  assign y11581 = n27021 ;
  assign y11582 = ~n27023 ;
  assign y11583 = ~1'b0 ;
  assign y11584 = ~1'b0 ;
  assign y11585 = n27024 ;
  assign y11586 = ~n27027 ;
  assign y11587 = n27035 ;
  assign y11588 = n27037 ;
  assign y11589 = ~n27043 ;
  assign y11590 = ~n349 ;
  assign y11591 = ~n27044 ;
  assign y11592 = ~1'b0 ;
  assign y11593 = ~n27046 ;
  assign y11594 = n27047 ;
  assign y11595 = n27049 ;
  assign y11596 = ~1'b0 ;
  assign y11597 = ~n27051 ;
  assign y11598 = n27054 ;
  assign y11599 = ~n27055 ;
  assign y11600 = ~n14225 ;
  assign y11601 = n27057 ;
  assign y11602 = ~n27059 ;
  assign y11603 = ~n27061 ;
  assign y11604 = n27063 ;
  assign y11605 = ~1'b0 ;
  assign y11606 = ~1'b0 ;
  assign y11607 = ~n27066 ;
  assign y11608 = n27067 ;
  assign y11609 = ~n27068 ;
  assign y11610 = n27075 ;
  assign y11611 = ~n27079 ;
  assign y11612 = n27080 ;
  assign y11613 = ~n27084 ;
  assign y11614 = ~n27087 ;
  assign y11615 = ~1'b0 ;
  assign y11616 = ~1'b0 ;
  assign y11617 = n27088 ;
  assign y11618 = ~n27089 ;
  assign y11619 = n27092 ;
  assign y11620 = n27093 ;
  assign y11621 = ~1'b0 ;
  assign y11622 = ~n27094 ;
  assign y11623 = ~1'b0 ;
  assign y11624 = ~n27099 ;
  assign y11625 = ~n27102 ;
  assign y11626 = n27104 ;
  assign y11627 = n27109 ;
  assign y11628 = ~n27112 ;
  assign y11629 = ~n27114 ;
  assign y11630 = n27117 ;
  assign y11631 = ~1'b0 ;
  assign y11632 = ~1'b0 ;
  assign y11633 = ~1'b0 ;
  assign y11634 = n27120 ;
  assign y11635 = ~n27122 ;
  assign y11636 = n27124 ;
  assign y11637 = ~1'b0 ;
  assign y11638 = ~n27126 ;
  assign y11639 = ~n27127 ;
  assign y11640 = ~n27129 ;
  assign y11641 = ~1'b0 ;
  assign y11642 = ~n27130 ;
  assign y11643 = n27132 ;
  assign y11644 = n27136 ;
  assign y11645 = ~1'b0 ;
  assign y11646 = n27140 ;
  assign y11647 = n27144 ;
  assign y11648 = n27148 ;
  assign y11649 = ~n27149 ;
  assign y11650 = n23069 ;
  assign y11651 = n27151 ;
  assign y11652 = ~n27152 ;
  assign y11653 = ~n27154 ;
  assign y11654 = n27156 ;
  assign y11655 = ~1'b0 ;
  assign y11656 = ~n27158 ;
  assign y11657 = n27162 ;
  assign y11658 = ~n27164 ;
  assign y11659 = n27166 ;
  assign y11660 = n27167 ;
  assign y11661 = ~n27169 ;
  assign y11662 = ~n27171 ;
  assign y11663 = ~n27173 ;
  assign y11664 = ~n27174 ;
  assign y11665 = ~n27177 ;
  assign y11666 = ~n27179 ;
  assign y11667 = ~n27180 ;
  assign y11668 = ~1'b0 ;
  assign y11669 = 1'b0 ;
  assign y11670 = n27181 ;
  assign y11671 = ~n27182 ;
  assign y11672 = n27184 ;
  assign y11673 = n27192 ;
  assign y11674 = n27194 ;
  assign y11675 = ~n27198 ;
  assign y11676 = n27201 ;
  assign y11677 = ~1'b0 ;
  assign y11678 = ~1'b0 ;
  assign y11679 = ~n27202 ;
  assign y11680 = n27205 ;
  assign y11681 = n27210 ;
  assign y11682 = ~n27212 ;
  assign y11683 = ~n27215 ;
  assign y11684 = n27219 ;
  assign y11685 = n27220 ;
  assign y11686 = ~1'b0 ;
  assign y11687 = ~1'b0 ;
  assign y11688 = ~1'b0 ;
  assign y11689 = n27221 ;
  assign y11690 = ~n27222 ;
  assign y11691 = ~n27226 ;
  assign y11692 = n27228 ;
  assign y11693 = ~1'b0 ;
  assign y11694 = ~n27234 ;
  assign y11695 = ~1'b0 ;
  assign y11696 = ~1'b0 ;
  assign y11697 = ~n27239 ;
  assign y11698 = n27242 ;
  assign y11699 = ~1'b0 ;
  assign y11700 = ~n27244 ;
  assign y11701 = ~n27245 ;
  assign y11702 = ~n27246 ;
  assign y11703 = n27247 ;
  assign y11704 = n27249 ;
  assign y11705 = ~n27252 ;
  assign y11706 = n27257 ;
  assign y11707 = n27259 ;
  assign y11708 = ~n27261 ;
  assign y11709 = ~1'b0 ;
  assign y11710 = ~n27265 ;
  assign y11711 = ~n27269 ;
  assign y11712 = n27271 ;
  assign y11713 = ~n27272 ;
  assign y11714 = n27273 ;
  assign y11715 = ~n27275 ;
  assign y11716 = ~n27281 ;
  assign y11717 = ~1'b0 ;
  assign y11718 = ~1'b0 ;
  assign y11719 = ~n27285 ;
  assign y11720 = ~n27287 ;
  assign y11721 = ~1'b0 ;
  assign y11722 = ~n27288 ;
  assign y11723 = n27292 ;
  assign y11724 = ~n27293 ;
  assign y11725 = n27300 ;
  assign y11726 = n27301 ;
  assign y11727 = ~n27305 ;
  assign y11728 = ~1'b0 ;
  assign y11729 = n27307 ;
  assign y11730 = n27309 ;
  assign y11731 = ~n27310 ;
  assign y11732 = ~n27311 ;
  assign y11733 = ~n27312 ;
  assign y11734 = ~n27316 ;
  assign y11735 = ~n27318 ;
  assign y11736 = ~n27321 ;
  assign y11737 = ~n27322 ;
  assign y11738 = ~1'b0 ;
  assign y11739 = ~n27327 ;
  assign y11740 = n27329 ;
  assign y11741 = n27331 ;
  assign y11742 = n27333 ;
  assign y11743 = ~n27336 ;
  assign y11744 = ~n27337 ;
  assign y11745 = n13672 ;
  assign y11746 = ~n27338 ;
  assign y11747 = ~n27341 ;
  assign y11748 = ~n27343 ;
  assign y11749 = ~n27345 ;
  assign y11750 = n27347 ;
  assign y11751 = ~1'b0 ;
  assign y11752 = n27349 ;
  assign y11753 = ~n27352 ;
  assign y11754 = n27353 ;
  assign y11755 = n27354 ;
  assign y11756 = n5355 ;
  assign y11757 = n27358 ;
  assign y11758 = n27361 ;
  assign y11759 = ~n27362 ;
  assign y11760 = ~1'b0 ;
  assign y11761 = n27365 ;
  assign y11762 = ~1'b0 ;
  assign y11763 = n27367 ;
  assign y11764 = ~n27369 ;
  assign y11765 = ~n27372 ;
  assign y11766 = n27373 ;
  assign y11767 = 1'b0 ;
  assign y11768 = ~1'b0 ;
  assign y11769 = ~1'b0 ;
  assign y11770 = ~n27375 ;
  assign y11771 = ~1'b0 ;
  assign y11772 = ~1'b0 ;
  assign y11773 = ~1'b0 ;
  assign y11774 = ~1'b0 ;
  assign y11775 = ~n27376 ;
  assign y11776 = n27377 ;
  assign y11777 = n27378 ;
  assign y11778 = ~n27380 ;
  assign y11779 = ~1'b0 ;
  assign y11780 = n27382 ;
  assign y11781 = n27386 ;
  assign y11782 = ~1'b0 ;
  assign y11783 = ~1'b0 ;
  assign y11784 = ~n27388 ;
  assign y11785 = ~n10809 ;
  assign y11786 = ~n27389 ;
  assign y11787 = n27394 ;
  assign y11788 = ~n27395 ;
  assign y11789 = ~n27396 ;
  assign y11790 = ~1'b0 ;
  assign y11791 = n27398 ;
  assign y11792 = n27399 ;
  assign y11793 = ~1'b0 ;
  assign y11794 = n8860 ;
  assign y11795 = n27402 ;
  assign y11796 = n27403 ;
  assign y11797 = ~n27404 ;
  assign y11798 = ~n27407 ;
  assign y11799 = n27408 ;
  assign y11800 = ~n27409 ;
  assign y11801 = ~1'b0 ;
  assign y11802 = n27410 ;
  assign y11803 = ~n27411 ;
  assign y11804 = ~1'b0 ;
  assign y11805 = n27413 ;
  assign y11806 = ~n27415 ;
  assign y11807 = ~n27417 ;
  assign y11808 = ~n15647 ;
  assign y11809 = n19820 ;
  assign y11810 = n27418 ;
  assign y11811 = ~n27421 ;
  assign y11812 = n27422 ;
  assign y11813 = n13457 ;
  assign y11814 = ~1'b0 ;
  assign y11815 = ~n27424 ;
  assign y11816 = ~n27425 ;
  assign y11817 = ~n27426 ;
  assign y11818 = ~n27436 ;
  assign y11819 = ~n27437 ;
  assign y11820 = n12470 ;
  assign y11821 = n27439 ;
  assign y11822 = ~n27441 ;
  assign y11823 = ~n27443 ;
  assign y11824 = ~n27444 ;
  assign y11825 = ~1'b0 ;
  assign y11826 = ~n27447 ;
  assign y11827 = ~n27450 ;
  assign y11828 = ~n27453 ;
  assign y11829 = ~n27456 ;
  assign y11830 = ~n27458 ;
  assign y11831 = ~n27459 ;
  assign y11832 = ~1'b0 ;
  assign y11833 = ~n27463 ;
  assign y11834 = ~1'b0 ;
  assign y11835 = n27469 ;
  assign y11836 = n27473 ;
  assign y11837 = ~1'b0 ;
  assign y11838 = n27474 ;
  assign y11839 = n27477 ;
  assign y11840 = n27478 ;
  assign y11841 = ~n27479 ;
  assign y11842 = ~1'b0 ;
  assign y11843 = n27482 ;
  assign y11844 = n27487 ;
  assign y11845 = ~1'b0 ;
  assign y11846 = ~n27489 ;
  assign y11847 = n27495 ;
  assign y11848 = n27496 ;
  assign y11849 = ~n27497 ;
  assign y11850 = n27499 ;
  assign y11851 = n27500 ;
  assign y11852 = n27503 ;
  assign y11853 = ~n27506 ;
  assign y11854 = ~n27509 ;
  assign y11855 = ~n27515 ;
  assign y11856 = ~1'b0 ;
  assign y11857 = 1'b0 ;
  assign y11858 = ~n27516 ;
  assign y11859 = n27520 ;
  assign y11860 = n27521 ;
  assign y11861 = ~n27523 ;
  assign y11862 = ~n27525 ;
  assign y11863 = ~1'b0 ;
  assign y11864 = ~n27529 ;
  assign y11865 = n27530 ;
  assign y11866 = ~1'b0 ;
  assign y11867 = ~1'b0 ;
  assign y11868 = ~n27531 ;
  assign y11869 = ~n27532 ;
  assign y11870 = n27533 ;
  assign y11871 = ~n27538 ;
  assign y11872 = ~1'b0 ;
  assign y11873 = n27539 ;
  assign y11874 = ~n27541 ;
  assign y11875 = ~1'b0 ;
  assign y11876 = ~1'b0 ;
  assign y11877 = n27545 ;
  assign y11878 = ~n27548 ;
  assign y11879 = ~n27550 ;
  assign y11880 = ~n27553 ;
  assign y11881 = ~n27557 ;
  assign y11882 = ~n27561 ;
  assign y11883 = ~n27564 ;
  assign y11884 = ~n27566 ;
  assign y11885 = ~1'b0 ;
  assign y11886 = ~n27568 ;
  assign y11887 = ~1'b0 ;
  assign y11888 = ~n27571 ;
  assign y11889 = n27572 ;
  assign y11890 = ~1'b0 ;
  assign y11891 = ~n27577 ;
  assign y11892 = n27579 ;
  assign y11893 = n27583 ;
  assign y11894 = ~n27585 ;
  assign y11895 = ~n27587 ;
  assign y11896 = ~1'b0 ;
  assign y11897 = ~1'b0 ;
  assign y11898 = ~1'b0 ;
  assign y11899 = ~n27588 ;
  assign y11900 = n27591 ;
  assign y11901 = ~n9710 ;
  assign y11902 = n27597 ;
  assign y11903 = ~n27599 ;
  assign y11904 = n27601 ;
  assign y11905 = ~1'b0 ;
  assign y11906 = ~n27606 ;
  assign y11907 = ~n27607 ;
  assign y11908 = n27614 ;
  assign y11909 = ~n27615 ;
  assign y11910 = n27620 ;
  assign y11911 = n27621 ;
  assign y11912 = n27622 ;
  assign y11913 = n27624 ;
  assign y11914 = ~n27631 ;
  assign y11915 = ~1'b0 ;
  assign y11916 = ~n27635 ;
  assign y11917 = n27637 ;
  assign y11918 = ~n27643 ;
  assign y11919 = ~1'b0 ;
  assign y11920 = n27644 ;
  assign y11921 = ~n27645 ;
  assign y11922 = n27647 ;
  assign y11923 = ~n27648 ;
  assign y11924 = ~n27651 ;
  assign y11925 = ~n27653 ;
  assign y11926 = n27658 ;
  assign y11927 = ~n27662 ;
  assign y11928 = ~1'b0 ;
  assign y11929 = ~1'b0 ;
  assign y11930 = n27664 ;
  assign y11931 = ~n27666 ;
  assign y11932 = ~1'b0 ;
  assign y11933 = ~n27668 ;
  assign y11934 = n27671 ;
  assign y11935 = ~n27672 ;
  assign y11936 = n27675 ;
  assign y11937 = ~n27677 ;
  assign y11938 = n27678 ;
  assign y11939 = n27680 ;
  assign y11940 = ~n27682 ;
  assign y11941 = n27683 ;
  assign y11942 = n27685 ;
  assign y11943 = ~n27687 ;
  assign y11944 = ~n27689 ;
  assign y11945 = n27690 ;
  assign y11946 = n2193 ;
  assign y11947 = ~1'b0 ;
  assign y11948 = ~n27692 ;
  assign y11949 = n27693 ;
  assign y11950 = n27694 ;
  assign y11951 = ~n27695 ;
  assign y11952 = n27701 ;
  assign y11953 = n27702 ;
  assign y11954 = ~n27705 ;
  assign y11955 = n27706 ;
  assign y11956 = n27708 ;
  assign y11957 = 1'b0 ;
  assign y11958 = n27710 ;
  assign y11959 = ~n27711 ;
  assign y11960 = n27716 ;
  assign y11961 = n27718 ;
  assign y11962 = ~n27719 ;
  assign y11963 = n17794 ;
  assign y11964 = ~n27722 ;
  assign y11965 = n27730 ;
  assign y11966 = n27731 ;
  assign y11967 = ~1'b0 ;
  assign y11968 = ~n27733 ;
  assign y11969 = ~1'b0 ;
  assign y11970 = ~n27735 ;
  assign y11971 = n27738 ;
  assign y11972 = ~n27740 ;
  assign y11973 = ~n27742 ;
  assign y11974 = n27745 ;
  assign y11975 = n27749 ;
  assign y11976 = n27752 ;
  assign y11977 = n27756 ;
  assign y11978 = ~n27757 ;
  assign y11979 = ~n27759 ;
  assign y11980 = n27761 ;
  assign y11981 = ~1'b0 ;
  assign y11982 = ~1'b0 ;
  assign y11983 = ~n21949 ;
  assign y11984 = ~n27764 ;
  assign y11985 = n27765 ;
  assign y11986 = n27766 ;
  assign y11987 = n27767 ;
  assign y11988 = ~1'b0 ;
  assign y11989 = ~n27770 ;
  assign y11990 = ~n27772 ;
  assign y11991 = ~n27773 ;
  assign y11992 = n27775 ;
  assign y11993 = n27777 ;
  assign y11994 = n27778 ;
  assign y11995 = n27781 ;
  assign y11996 = ~n27783 ;
  assign y11997 = n27784 ;
  assign y11998 = ~n27786 ;
  assign y11999 = n27789 ;
  assign y12000 = ~n27790 ;
  assign y12001 = n27792 ;
  assign y12002 = ~n27794 ;
  assign y12003 = n27796 ;
  assign y12004 = n27797 ;
  assign y12005 = ~n27799 ;
  assign y12006 = ~n27800 ;
  assign y12007 = ~n27801 ;
  assign y12008 = n27805 ;
  assign y12009 = ~1'b0 ;
  assign y12010 = n27809 ;
  assign y12011 = ~n27810 ;
  assign y12012 = ~n14855 ;
  assign y12013 = ~1'b0 ;
  assign y12014 = n27082 ;
  assign y12015 = n27811 ;
  assign y12016 = ~n27812 ;
  assign y12017 = ~n27813 ;
  assign y12018 = ~n27814 ;
  assign y12019 = n27821 ;
  assign y12020 = ~n27827 ;
  assign y12021 = ~1'b0 ;
  assign y12022 = ~n27829 ;
  assign y12023 = ~n27831 ;
  assign y12024 = ~n27833 ;
  assign y12025 = 1'b0 ;
  assign y12026 = ~n27835 ;
  assign y12027 = ~n27836 ;
  assign y12028 = ~n27838 ;
  assign y12029 = ~n27840 ;
  assign y12030 = ~n27842 ;
  assign y12031 = ~n27718 ;
  assign y12032 = n26528 ;
  assign y12033 = ~n27844 ;
  assign y12034 = ~n27848 ;
  assign y12035 = ~1'b0 ;
  assign y12036 = ~n27849 ;
  assign y12037 = n27852 ;
  assign y12038 = n27860 ;
  assign y12039 = n27861 ;
  assign y12040 = n27863 ;
  assign y12041 = ~n27865 ;
  assign y12042 = ~n27869 ;
  assign y12043 = n27870 ;
  assign y12044 = ~1'b0 ;
  assign y12045 = ~1'b0 ;
  assign y12046 = n27871 ;
  assign y12047 = ~n7795 ;
  assign y12048 = ~n27872 ;
  assign y12049 = ~n27875 ;
  assign y12050 = n27876 ;
  assign y12051 = n27877 ;
  assign y12052 = ~n27879 ;
  assign y12053 = n27882 ;
  assign y12054 = ~1'b0 ;
  assign y12055 = n27883 ;
  assign y12056 = ~n27887 ;
  assign y12057 = ~n27888 ;
  assign y12058 = ~1'b0 ;
  assign y12059 = n27889 ;
  assign y12060 = n27890 ;
  assign y12061 = ~n27892 ;
  assign y12062 = n27896 ;
  assign y12063 = ~n12841 ;
  assign y12064 = ~1'b0 ;
  assign y12065 = ~n27900 ;
  assign y12066 = ~1'b0 ;
  assign y12067 = ~n27901 ;
  assign y12068 = n27902 ;
  assign y12069 = ~n27904 ;
  assign y12070 = n27905 ;
  assign y12071 = n27906 ;
  assign y12072 = ~n27909 ;
  assign y12073 = n27911 ;
  assign y12074 = ~1'b0 ;
  assign y12075 = ~1'b0 ;
  assign y12076 = n27913 ;
  assign y12077 = ~n16219 ;
  assign y12078 = ~1'b0 ;
  assign y12079 = ~n27915 ;
  assign y12080 = n27916 ;
  assign y12081 = n27917 ;
  assign y12082 = ~1'b0 ;
  assign y12083 = n27919 ;
  assign y12084 = ~n27926 ;
  assign y12085 = n27928 ;
  assign y12086 = n27930 ;
  assign y12087 = ~n27931 ;
  assign y12088 = ~n27932 ;
  assign y12089 = n27934 ;
  assign y12090 = ~n20184 ;
  assign y12091 = n19005 ;
  assign y12092 = n27941 ;
  assign y12093 = n27944 ;
  assign y12094 = ~n27947 ;
  assign y12095 = ~n27951 ;
  assign y12096 = ~1'b0 ;
  assign y12097 = ~n27954 ;
  assign y12098 = n27959 ;
  assign y12099 = ~n5061 ;
  assign y12100 = ~n27963 ;
  assign y12101 = ~n27964 ;
  assign y12102 = ~n27967 ;
  assign y12103 = ~n27970 ;
  assign y12104 = n27975 ;
  assign y12105 = ~n27976 ;
  assign y12106 = n26168 ;
  assign y12107 = ~n27978 ;
  assign y12108 = n27980 ;
  assign y12109 = ~n27981 ;
  assign y12110 = ~n27984 ;
  assign y12111 = ~1'b0 ;
  assign y12112 = ~n27986 ;
  assign y12113 = ~n27987 ;
  assign y12114 = ~n27988 ;
  assign y12115 = n27989 ;
  assign y12116 = n28006 ;
  assign y12117 = n28007 ;
  assign y12118 = n28008 ;
  assign y12119 = ~1'b0 ;
  assign y12120 = ~n28010 ;
  assign y12121 = 1'b0 ;
  assign y12122 = n28013 ;
  assign y12123 = n28015 ;
  assign y12124 = ~n28018 ;
  assign y12125 = ~n28026 ;
  assign y12126 = n28028 ;
  assign y12127 = ~n28032 ;
  assign y12128 = ~1'b0 ;
  assign y12129 = ~n28037 ;
  assign y12130 = ~1'b0 ;
  assign y12131 = n28038 ;
  assign y12132 = n28039 ;
  assign y12133 = ~1'b0 ;
  assign y12134 = n28040 ;
  assign y12135 = n28042 ;
  assign y12136 = ~n28043 ;
  assign y12137 = n28045 ;
  assign y12138 = n28046 ;
  assign y12139 = n28048 ;
  assign y12140 = ~1'b0 ;
  assign y12141 = n28050 ;
  assign y12142 = ~n28053 ;
  assign y12143 = ~1'b0 ;
  assign y12144 = 1'b0 ;
  assign y12145 = ~1'b0 ;
  assign y12146 = n28055 ;
  assign y12147 = n28056 ;
  assign y12148 = ~n28057 ;
  assign y12149 = ~n28061 ;
  assign y12150 = ~n28062 ;
  assign y12151 = n28063 ;
  assign y12152 = n28065 ;
  assign y12153 = ~n28066 ;
  assign y12154 = ~n28078 ;
  assign y12155 = n28080 ;
  assign y12156 = n15784 ;
  assign y12157 = ~n28085 ;
  assign y12158 = ~n28086 ;
  assign y12159 = n28089 ;
  assign y12160 = n28092 ;
  assign y12161 = ~1'b0 ;
  assign y12162 = n28094 ;
  assign y12163 = ~1'b0 ;
  assign y12164 = n28095 ;
  assign y12165 = ~1'b0 ;
  assign y12166 = ~1'b0 ;
  assign y12167 = ~1'b0 ;
  assign y12168 = ~n28100 ;
  assign y12169 = ~n28102 ;
  assign y12170 = n28106 ;
  assign y12171 = ~n28109 ;
  assign y12172 = n28111 ;
  assign y12173 = n28112 ;
  assign y12174 = n28122 ;
  assign y12175 = ~n28124 ;
  assign y12176 = ~n28125 ;
  assign y12177 = n28126 ;
  assign y12178 = ~n18227 ;
  assign y12179 = n28128 ;
  assign y12180 = ~n28129 ;
  assign y12181 = n28130 ;
  assign y12182 = n28131 ;
  assign y12183 = ~n28135 ;
  assign y12184 = ~n28136 ;
  assign y12185 = n28138 ;
  assign y12186 = ~n14925 ;
  assign y12187 = ~1'b0 ;
  assign y12188 = ~1'b0 ;
  assign y12189 = n28139 ;
  assign y12190 = n28140 ;
  assign y12191 = n28142 ;
  assign y12192 = ~1'b0 ;
  assign y12193 = n28145 ;
  assign y12194 = ~n28147 ;
  assign y12195 = n28149 ;
  assign y12196 = ~1'b0 ;
  assign y12197 = n28151 ;
  assign y12198 = ~1'b0 ;
  assign y12199 = ~n28152 ;
  assign y12200 = ~n28154 ;
  assign y12201 = ~n1756 ;
  assign y12202 = n28156 ;
  assign y12203 = ~n28158 ;
  assign y12204 = ~n28159 ;
  assign y12205 = ~1'b0 ;
  assign y12206 = ~n28162 ;
  assign y12207 = n28163 ;
  assign y12208 = n28168 ;
  assign y12209 = ~n28172 ;
  assign y12210 = ~1'b0 ;
  assign y12211 = ~n28175 ;
  assign y12212 = ~n28176 ;
  assign y12213 = ~n28177 ;
  assign y12214 = n22540 ;
  assign y12215 = ~n28179 ;
  assign y12216 = ~1'b0 ;
  assign y12217 = ~n28181 ;
  assign y12218 = ~n28182 ;
  assign y12219 = ~1'b0 ;
  assign y12220 = ~n28187 ;
  assign y12221 = n28191 ;
  assign y12222 = n28194 ;
  assign y12223 = n28196 ;
  assign y12224 = n1952 ;
  assign y12225 = ~n28198 ;
  assign y12226 = n28199 ;
  assign y12227 = ~n28203 ;
  assign y12228 = ~1'b0 ;
  assign y12229 = ~n28206 ;
  assign y12230 = ~1'b0 ;
  assign y12231 = ~n28212 ;
  assign y12232 = ~1'b0 ;
  assign y12233 = ~1'b0 ;
  assign y12234 = ~n28214 ;
  assign y12235 = ~n28216 ;
  assign y12236 = n28219 ;
  assign y12237 = ~n28222 ;
  assign y12238 = n28223 ;
  assign y12239 = ~1'b0 ;
  assign y12240 = ~1'b0 ;
  assign y12241 = n28224 ;
  assign y12242 = ~1'b0 ;
  assign y12243 = ~n28226 ;
  assign y12244 = n28227 ;
  assign y12245 = ~n28230 ;
  assign y12246 = ~n28231 ;
  assign y12247 = n28237 ;
  assign y12248 = ~n28240 ;
  assign y12249 = n28242 ;
  assign y12250 = n28246 ;
  assign y12251 = ~n28250 ;
  assign y12252 = ~n28254 ;
  assign y12253 = ~1'b0 ;
  assign y12254 = n28255 ;
  assign y12255 = n28257 ;
  assign y12256 = ~n28259 ;
  assign y12257 = ~n28263 ;
  assign y12258 = ~n28264 ;
  assign y12259 = ~n28265 ;
  assign y12260 = ~1'b0 ;
  assign y12261 = ~1'b0 ;
  assign y12262 = ~n28267 ;
  assign y12263 = ~1'b0 ;
  assign y12264 = ~n28268 ;
  assign y12265 = ~n28269 ;
  assign y12266 = ~n28271 ;
  assign y12267 = n28273 ;
  assign y12268 = n28275 ;
  assign y12269 = ~n28277 ;
  assign y12270 = ~n28280 ;
  assign y12271 = ~n28281 ;
  assign y12272 = ~1'b0 ;
  assign y12273 = ~1'b0 ;
  assign y12274 = ~1'b0 ;
  assign y12275 = ~1'b0 ;
  assign y12276 = n28283 ;
  assign y12277 = n28284 ;
  assign y12278 = ~1'b0 ;
  assign y12279 = n28285 ;
  assign y12280 = n28287 ;
  assign y12281 = ~n28288 ;
  assign y12282 = n28289 ;
  assign y12283 = ~n28292 ;
  assign y12284 = n28300 ;
  assign y12285 = ~1'b0 ;
  assign y12286 = ~n28302 ;
  assign y12287 = ~1'b0 ;
  assign y12288 = ~n28304 ;
  assign y12289 = ~n28305 ;
  assign y12290 = n28306 ;
  assign y12291 = n28307 ;
  assign y12292 = n28308 ;
  assign y12293 = ~1'b0 ;
  assign y12294 = n28309 ;
  assign y12295 = ~n28312 ;
  assign y12296 = n28314 ;
  assign y12297 = ~n28317 ;
  assign y12298 = ~n28319 ;
  assign y12299 = n28326 ;
  assign y12300 = n28330 ;
  assign y12301 = n28334 ;
  assign y12302 = ~n28336 ;
  assign y12303 = ~n28337 ;
  assign y12304 = n8345 ;
  assign y12305 = ~1'b0 ;
  assign y12306 = ~1'b0 ;
  assign y12307 = n28339 ;
  assign y12308 = ~1'b0 ;
  assign y12309 = ~n28342 ;
  assign y12310 = ~1'b0 ;
  assign y12311 = n28348 ;
  assign y12312 = ~n28349 ;
  assign y12313 = ~n28351 ;
  assign y12314 = ~n28352 ;
  assign y12315 = ~n28355 ;
  assign y12316 = ~1'b0 ;
  assign y12317 = n28360 ;
  assign y12318 = n28362 ;
  assign y12319 = n28364 ;
  assign y12320 = ~1'b0 ;
  assign y12321 = n28366 ;
  assign y12322 = n28369 ;
  assign y12323 = ~n28370 ;
  assign y12324 = n28373 ;
  assign y12325 = ~n28374 ;
  assign y12326 = ~1'b0 ;
  assign y12327 = n28375 ;
  assign y12328 = ~1'b0 ;
  assign y12329 = ~1'b0 ;
  assign y12330 = ~1'b0 ;
  assign y12331 = n28376 ;
  assign y12332 = ~n28378 ;
  assign y12333 = n28384 ;
  assign y12334 = n28386 ;
  assign y12335 = n28387 ;
  assign y12336 = ~n28388 ;
  assign y12337 = ~n28391 ;
  assign y12338 = ~n28393 ;
  assign y12339 = n28394 ;
  assign y12340 = ~n28396 ;
  assign y12341 = n28399 ;
  assign y12342 = ~1'b0 ;
  assign y12343 = ~1'b0 ;
  assign y12344 = n28402 ;
  assign y12345 = ~n28403 ;
  assign y12346 = ~1'b0 ;
  assign y12347 = ~n28405 ;
  assign y12348 = n28407 ;
  assign y12349 = n28408 ;
  assign y12350 = ~n28409 ;
  assign y12351 = ~1'b0 ;
  assign y12352 = ~n28416 ;
  assign y12353 = ~n28417 ;
  assign y12354 = ~n28418 ;
  assign y12355 = n28420 ;
  assign y12356 = n28422 ;
  assign y12357 = n28423 ;
  assign y12358 = n28424 ;
  assign y12359 = ~1'b0 ;
  assign y12360 = n28426 ;
  assign y12361 = n28427 ;
  assign y12362 = ~1'b0 ;
  assign y12363 = ~n28431 ;
  assign y12364 = n28433 ;
  assign y12365 = ~n28437 ;
endmodule
