module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 ;
  wire n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6342 , n6343 , n6344 , n6346 , n6347 , n6348 ;
  assign n513 = x375 & ~x503 ;
  assign n514 = ~x375 & x503 ;
  assign n515 = ~x374 & x502 ;
  assign n516 = ~n514 & ~n515 ;
  assign n517 = ~x373 & x501 ;
  assign n518 = x372 & ~x500 ;
  assign n519 = ~n517 & n518 ;
  assign n520 = x373 & ~x501 ;
  assign n521 = ~n519 & ~n520 ;
  assign n522 = n516 & ~n521 ;
  assign n523 = ~x502 & ~n514 ;
  assign n524 = x374 & n523 ;
  assign n525 = ~x368 & x496 ;
  assign n526 = ~x371 & x499 ;
  assign n527 = ~x370 & x498 ;
  assign n528 = ~n526 & ~n527 ;
  assign n529 = ~x369 & x497 ;
  assign n530 = x367 & ~x495 ;
  assign n531 = ~x367 & x495 ;
  assign n532 = ~x366 & x494 ;
  assign n533 = ~n531 & ~n532 ;
  assign n534 = ~x365 & x493 ;
  assign n535 = x364 & ~x492 ;
  assign n536 = ~n534 & n535 ;
  assign n537 = x365 & ~x493 ;
  assign n538 = ~n536 & ~n537 ;
  assign n539 = n533 & ~n538 ;
  assign n540 = ~x494 & ~n531 ;
  assign n541 = x366 & n540 ;
  assign n542 = x359 & ~x487 ;
  assign n543 = ~x359 & x487 ;
  assign n544 = ~x358 & x486 ;
  assign n545 = ~n543 & ~n544 ;
  assign n546 = ~x357 & x485 ;
  assign n547 = x356 & ~x484 ;
  assign n548 = ~n546 & n547 ;
  assign n549 = x357 & ~x485 ;
  assign n550 = ~n548 & ~n549 ;
  assign n551 = n545 & ~n550 ;
  assign n552 = ~x486 & ~n543 ;
  assign n553 = x358 & n552 ;
  assign n554 = ~x352 & x480 ;
  assign n555 = ~x355 & x483 ;
  assign n556 = ~x354 & x482 ;
  assign n557 = ~n555 & ~n556 ;
  assign n558 = ~x353 & x481 ;
  assign n559 = x351 & ~x479 ;
  assign n560 = ~x351 & x479 ;
  assign n561 = ~x350 & x478 ;
  assign n562 = ~n560 & ~n561 ;
  assign n563 = ~x349 & x477 ;
  assign n564 = x348 & ~x476 ;
  assign n565 = ~n563 & n564 ;
  assign n566 = x349 & ~x477 ;
  assign n567 = ~n565 & ~n566 ;
  assign n568 = n562 & ~n567 ;
  assign n569 = ~x478 & ~n560 ;
  assign n570 = x350 & n569 ;
  assign n571 = x343 & ~x471 ;
  assign n572 = ~x343 & x471 ;
  assign n573 = ~x342 & x470 ;
  assign n574 = ~n572 & ~n573 ;
  assign n575 = ~x341 & x469 ;
  assign n576 = x340 & ~x468 ;
  assign n577 = ~n575 & n576 ;
  assign n578 = x341 & ~x469 ;
  assign n579 = ~n577 & ~n578 ;
  assign n580 = n574 & ~n579 ;
  assign n581 = ~x470 & ~n572 ;
  assign n582 = x342 & n581 ;
  assign n583 = ~x336 & x464 ;
  assign n584 = ~x339 & x467 ;
  assign n585 = ~x338 & x466 ;
  assign n586 = ~n584 & ~n585 ;
  assign n587 = ~x337 & x465 ;
  assign n588 = x335 & ~x463 ;
  assign n589 = ~x335 & x463 ;
  assign n590 = ~x334 & x462 ;
  assign n591 = ~n589 & ~n590 ;
  assign n592 = ~x333 & x461 ;
  assign n593 = x332 & ~x460 ;
  assign n594 = ~n592 & n593 ;
  assign n595 = x333 & ~x461 ;
  assign n596 = ~n594 & ~n595 ;
  assign n597 = n591 & ~n596 ;
  assign n598 = ~x462 & ~n589 ;
  assign n599 = x334 & n598 ;
  assign n600 = x327 & ~x455 ;
  assign n601 = ~x327 & x455 ;
  assign n602 = ~x326 & x454 ;
  assign n603 = ~n601 & ~n602 ;
  assign n604 = ~x325 & x453 ;
  assign n605 = x324 & ~x452 ;
  assign n606 = ~n604 & n605 ;
  assign n607 = x325 & ~x453 ;
  assign n608 = ~n606 & ~n607 ;
  assign n609 = n603 & ~n608 ;
  assign n610 = ~x454 & ~n601 ;
  assign n611 = x326 & n610 ;
  assign n612 = ~x323 & x451 ;
  assign n613 = ~x322 & x450 ;
  assign n614 = ~n612 & ~n613 ;
  assign n615 = ~x321 & x449 ;
  assign n616 = x319 & ~x447 ;
  assign n617 = ~x319 & x447 ;
  assign n618 = ~x318 & x446 ;
  assign n619 = ~n617 & ~n618 ;
  assign n620 = ~x316 & x444 ;
  assign n621 = ~x317 & x445 ;
  assign n622 = ~n620 & ~n621 ;
  assign n623 = n619 & n622 ;
  assign n624 = x315 & ~x443 ;
  assign n625 = ~x315 & x443 ;
  assign n626 = ~x314 & x442 ;
  assign n627 = ~n625 & ~n626 ;
  assign n628 = ~x313 & x441 ;
  assign n629 = x312 & ~x440 ;
  assign n630 = ~n628 & n629 ;
  assign n631 = x313 & ~x441 ;
  assign n632 = ~n630 & ~n631 ;
  assign n633 = x314 & ~x442 ;
  assign n634 = n632 & ~n633 ;
  assign n635 = n627 & ~n634 ;
  assign n636 = ~n624 & ~n635 ;
  assign n637 = n623 & ~n636 ;
  assign n638 = x316 & ~x444 ;
  assign n639 = ~n621 & n638 ;
  assign n640 = x317 & ~x445 ;
  assign n641 = ~n639 & ~n640 ;
  assign n642 = n619 & ~n641 ;
  assign n643 = ~x446 & ~n617 ;
  assign n644 = x318 & n643 ;
  assign n645 = x303 & ~x431 ;
  assign n646 = ~x303 & x431 ;
  assign n647 = ~x302 & x430 ;
  assign n648 = ~n646 & ~n647 ;
  assign n649 = ~x300 & x428 ;
  assign n650 = ~x301 & x429 ;
  assign n651 = ~n649 & ~n650 ;
  assign n652 = n648 & n651 ;
  assign n653 = x299 & ~x427 ;
  assign n654 = ~x299 & x427 ;
  assign n655 = ~x298 & x426 ;
  assign n656 = ~n654 & ~n655 ;
  assign n657 = ~x297 & x425 ;
  assign n658 = x296 & ~x424 ;
  assign n659 = ~n657 & n658 ;
  assign n660 = x297 & ~x425 ;
  assign n661 = ~n659 & ~n660 ;
  assign n662 = x298 & ~x426 ;
  assign n663 = n661 & ~n662 ;
  assign n664 = n656 & ~n663 ;
  assign n665 = ~n653 & ~n664 ;
  assign n666 = n652 & ~n665 ;
  assign n667 = x300 & ~x428 ;
  assign n668 = ~n650 & n667 ;
  assign n669 = x301 & ~x429 ;
  assign n670 = ~n668 & ~n669 ;
  assign n671 = n648 & ~n670 ;
  assign n672 = ~x430 & ~n646 ;
  assign n673 = x302 & n672 ;
  assign n674 = ~x288 & x416 ;
  assign n675 = ~x287 & x415 ;
  assign n676 = ~x286 & x414 ;
  assign n677 = ~x285 & x413 ;
  assign n678 = ~x284 & x412 ;
  assign n679 = ~x283 & x411 ;
  assign n680 = ~x282 & x410 ;
  assign n681 = ~x279 & x407 ;
  assign n682 = ~x278 & x406 ;
  assign n683 = ~x277 & x405 ;
  assign n684 = ~x276 & x404 ;
  assign n685 = ~x275 & x403 ;
  assign n686 = ~x274 & x402 ;
  assign n687 = ~x271 & x399 ;
  assign n688 = ~x270 & x398 ;
  assign n689 = ~x269 & x397 ;
  assign n690 = ~x268 & x396 ;
  assign n691 = ~x267 & x395 ;
  assign n692 = ~x266 & x394 ;
  assign n693 = ~x263 & x391 ;
  assign n694 = ~x262 & x390 ;
  assign n695 = ~x259 & x387 ;
  assign n696 = x256 & ~x384 ;
  assign n697 = x257 & n696 ;
  assign n698 = x385 & ~n697 ;
  assign n699 = ~x258 & x386 ;
  assign n700 = ~x257 & ~n696 ;
  assign n701 = ~n699 & ~n700 ;
  assign n702 = ~n698 & n701 ;
  assign n703 = x258 & ~x386 ;
  assign n704 = ~n702 & ~n703 ;
  assign n705 = ~n695 & ~n704 ;
  assign n706 = x259 & ~x387 ;
  assign n707 = ~n705 & ~n706 ;
  assign n708 = ~x260 & n707 ;
  assign n709 = ~x388 & ~n708 ;
  assign n710 = x260 & ~n707 ;
  assign n711 = ~n709 & ~n710 ;
  assign n712 = ~x261 & n711 ;
  assign n713 = ~x389 & ~n712 ;
  assign n714 = x261 & ~n711 ;
  assign n715 = ~n713 & ~n714 ;
  assign n716 = ~n694 & ~n715 ;
  assign n717 = x262 & ~x390 ;
  assign n718 = ~n716 & ~n717 ;
  assign n719 = ~n693 & ~n718 ;
  assign n720 = x263 & ~x391 ;
  assign n721 = ~n719 & ~n720 ;
  assign n722 = ~x264 & n721 ;
  assign n723 = ~x392 & ~n722 ;
  assign n724 = x264 & ~n721 ;
  assign n725 = ~n723 & ~n724 ;
  assign n726 = ~x265 & n725 ;
  assign n727 = ~x393 & ~n726 ;
  assign n728 = x265 & ~n725 ;
  assign n729 = ~n727 & ~n728 ;
  assign n730 = ~n692 & ~n729 ;
  assign n731 = x266 & ~x394 ;
  assign n732 = ~n730 & ~n731 ;
  assign n733 = ~n691 & ~n732 ;
  assign n734 = x267 & ~x395 ;
  assign n735 = ~n733 & ~n734 ;
  assign n736 = ~n690 & ~n735 ;
  assign n737 = x268 & ~x396 ;
  assign n738 = ~n736 & ~n737 ;
  assign n739 = ~n689 & ~n738 ;
  assign n740 = x269 & ~x397 ;
  assign n741 = ~n739 & ~n740 ;
  assign n742 = ~n688 & ~n741 ;
  assign n743 = x270 & ~x398 ;
  assign n744 = ~n742 & ~n743 ;
  assign n745 = ~n687 & ~n744 ;
  assign n746 = x271 & ~x399 ;
  assign n747 = ~n745 & ~n746 ;
  assign n748 = ~x272 & n747 ;
  assign n749 = ~x400 & ~n748 ;
  assign n750 = x272 & ~n747 ;
  assign n751 = ~n749 & ~n750 ;
  assign n752 = ~x273 & n751 ;
  assign n753 = ~x401 & ~n752 ;
  assign n754 = x273 & ~n751 ;
  assign n755 = ~n753 & ~n754 ;
  assign n756 = ~n686 & ~n755 ;
  assign n757 = x274 & ~x402 ;
  assign n758 = ~n756 & ~n757 ;
  assign n759 = ~n685 & ~n758 ;
  assign n760 = x275 & ~x403 ;
  assign n761 = ~n759 & ~n760 ;
  assign n762 = ~n684 & ~n761 ;
  assign n763 = x276 & ~x404 ;
  assign n764 = ~n762 & ~n763 ;
  assign n765 = ~n683 & ~n764 ;
  assign n766 = x277 & ~x405 ;
  assign n767 = ~n765 & ~n766 ;
  assign n768 = ~n682 & ~n767 ;
  assign n769 = x278 & ~x406 ;
  assign n770 = ~n768 & ~n769 ;
  assign n771 = ~n681 & ~n770 ;
  assign n772 = x279 & ~x407 ;
  assign n773 = ~n771 & ~n772 ;
  assign n774 = ~x280 & n773 ;
  assign n775 = ~x408 & ~n774 ;
  assign n776 = x280 & ~n773 ;
  assign n777 = ~n775 & ~n776 ;
  assign n778 = ~x281 & n777 ;
  assign n779 = ~x409 & ~n778 ;
  assign n780 = x281 & ~n777 ;
  assign n781 = ~n779 & ~n780 ;
  assign n782 = ~n680 & ~n781 ;
  assign n783 = x282 & ~x410 ;
  assign n784 = ~n782 & ~n783 ;
  assign n785 = ~n679 & ~n784 ;
  assign n786 = x283 & ~x411 ;
  assign n787 = ~n785 & ~n786 ;
  assign n788 = ~n678 & ~n787 ;
  assign n789 = x284 & ~x412 ;
  assign n790 = ~n788 & ~n789 ;
  assign n791 = ~n677 & ~n790 ;
  assign n792 = x285 & ~x413 ;
  assign n793 = ~n791 & ~n792 ;
  assign n794 = ~n676 & ~n793 ;
  assign n795 = x286 & ~x414 ;
  assign n796 = ~n794 & ~n795 ;
  assign n797 = ~n675 & ~n796 ;
  assign n798 = x287 & ~x415 ;
  assign n799 = ~n797 & ~n798 ;
  assign n800 = ~x295 & x423 ;
  assign n801 = ~x294 & x422 ;
  assign n802 = ~n800 & ~n801 ;
  assign n803 = ~x292 & x420 ;
  assign n804 = ~x293 & x421 ;
  assign n805 = ~n803 & ~n804 ;
  assign n806 = n802 & n805 ;
  assign n807 = ~x289 & x417 ;
  assign n808 = ~x291 & x419 ;
  assign n809 = ~x290 & x418 ;
  assign n810 = ~n808 & ~n809 ;
  assign n811 = ~n807 & n810 ;
  assign n812 = n806 & n811 ;
  assign n813 = ~n799 & n812 ;
  assign n814 = ~n674 & n813 ;
  assign n815 = x295 & ~x423 ;
  assign n816 = x292 & ~x420 ;
  assign n817 = ~n804 & n816 ;
  assign n818 = x293 & ~x421 ;
  assign n819 = ~n817 & ~n818 ;
  assign n820 = n802 & ~n819 ;
  assign n821 = ~x422 & ~n800 ;
  assign n822 = x294 & n821 ;
  assign n823 = x291 & ~x419 ;
  assign n824 = ~x416 & ~n807 ;
  assign n825 = x288 & n824 ;
  assign n826 = x289 & ~x417 ;
  assign n827 = ~n825 & ~n826 ;
  assign n828 = x290 & ~x418 ;
  assign n829 = n827 & ~n828 ;
  assign n830 = n810 & ~n829 ;
  assign n831 = ~n823 & ~n830 ;
  assign n832 = n806 & ~n831 ;
  assign n833 = ~n822 & ~n832 ;
  assign n834 = ~n820 & n833 ;
  assign n835 = ~n815 & n834 ;
  assign n836 = ~n814 & n835 ;
  assign n837 = ~x296 & x424 ;
  assign n838 = ~n657 & ~n837 ;
  assign n839 = n656 & n838 ;
  assign n840 = n652 & n839 ;
  assign n841 = ~n836 & n840 ;
  assign n842 = ~n673 & ~n841 ;
  assign n843 = ~n671 & n842 ;
  assign n844 = ~n666 & n843 ;
  assign n845 = ~n645 & n844 ;
  assign n846 = ~x304 & x432 ;
  assign n847 = ~x311 & x439 ;
  assign n848 = ~x310 & x438 ;
  assign n849 = ~n847 & ~n848 ;
  assign n850 = ~x309 & x437 ;
  assign n851 = ~x308 & x436 ;
  assign n852 = ~n850 & ~n851 ;
  assign n853 = n849 & n852 ;
  assign n854 = ~x305 & x433 ;
  assign n855 = ~x307 & x435 ;
  assign n856 = ~x306 & x434 ;
  assign n857 = ~n855 & ~n856 ;
  assign n858 = ~n854 & n857 ;
  assign n859 = n853 & n858 ;
  assign n860 = ~n846 & n859 ;
  assign n861 = ~n845 & n860 ;
  assign n862 = x311 & ~x439 ;
  assign n863 = x307 & ~x435 ;
  assign n864 = ~x432 & ~n854 ;
  assign n865 = x304 & n864 ;
  assign n866 = x305 & ~x433 ;
  assign n867 = ~n865 & ~n866 ;
  assign n868 = x306 & ~x434 ;
  assign n869 = n867 & ~n868 ;
  assign n870 = n857 & ~n869 ;
  assign n871 = ~n863 & ~n870 ;
  assign n872 = n853 & ~n871 ;
  assign n873 = x308 & ~x436 ;
  assign n874 = ~n850 & n873 ;
  assign n875 = x309 & ~x437 ;
  assign n876 = ~n874 & ~n875 ;
  assign n877 = x310 & ~x438 ;
  assign n878 = n876 & ~n877 ;
  assign n879 = n849 & ~n878 ;
  assign n880 = ~n872 & ~n879 ;
  assign n881 = ~n862 & n880 ;
  assign n882 = ~n861 & n881 ;
  assign n883 = ~x312 & x440 ;
  assign n884 = ~n628 & ~n883 ;
  assign n885 = n623 & n884 ;
  assign n886 = n627 & n885 ;
  assign n887 = ~n882 & n886 ;
  assign n888 = ~n644 & ~n887 ;
  assign n889 = ~n642 & n888 ;
  assign n890 = ~n637 & n889 ;
  assign n891 = ~n616 & n890 ;
  assign n892 = ~x320 & x448 ;
  assign n893 = ~n891 & ~n892 ;
  assign n894 = ~n615 & n893 ;
  assign n895 = n614 & n894 ;
  assign n896 = x323 & ~x451 ;
  assign n897 = x320 & ~x448 ;
  assign n898 = ~n615 & n897 ;
  assign n899 = x321 & ~x449 ;
  assign n900 = ~n898 & ~n899 ;
  assign n901 = x322 & ~x450 ;
  assign n902 = n900 & ~n901 ;
  assign n903 = n614 & ~n902 ;
  assign n904 = ~n896 & ~n903 ;
  assign n905 = ~n895 & n904 ;
  assign n906 = ~x324 & x452 ;
  assign n907 = ~n604 & ~n906 ;
  assign n908 = n603 & n907 ;
  assign n909 = ~n905 & n908 ;
  assign n910 = ~n611 & ~n909 ;
  assign n911 = ~n609 & n910 ;
  assign n912 = ~n600 & n911 ;
  assign n913 = ~x331 & x459 ;
  assign n914 = ~x330 & x458 ;
  assign n915 = ~n913 & ~n914 ;
  assign n916 = ~x329 & x457 ;
  assign n917 = ~x328 & x456 ;
  assign n918 = ~n916 & ~n917 ;
  assign n919 = n915 & n918 ;
  assign n920 = ~n912 & n919 ;
  assign n921 = x331 & ~x459 ;
  assign n922 = x328 & ~x456 ;
  assign n923 = ~n916 & n922 ;
  assign n924 = x329 & ~x457 ;
  assign n925 = ~n923 & ~n924 ;
  assign n926 = x330 & ~x458 ;
  assign n927 = n925 & ~n926 ;
  assign n928 = n915 & ~n927 ;
  assign n929 = ~n921 & ~n928 ;
  assign n930 = ~n920 & n929 ;
  assign n931 = ~x332 & x460 ;
  assign n932 = ~n592 & ~n931 ;
  assign n933 = n591 & n932 ;
  assign n934 = ~n930 & n933 ;
  assign n935 = ~n599 & ~n934 ;
  assign n936 = ~n597 & n935 ;
  assign n937 = ~n588 & n936 ;
  assign n938 = ~n587 & ~n937 ;
  assign n939 = n586 & n938 ;
  assign n940 = ~n583 & n939 ;
  assign n941 = x339 & ~x467 ;
  assign n942 = ~x464 & ~n587 ;
  assign n943 = x336 & n942 ;
  assign n944 = x337 & ~x465 ;
  assign n945 = ~n943 & ~n944 ;
  assign n946 = x338 & ~x466 ;
  assign n947 = n945 & ~n946 ;
  assign n948 = n586 & ~n947 ;
  assign n949 = ~n941 & ~n948 ;
  assign n950 = ~n940 & n949 ;
  assign n951 = ~x340 & x468 ;
  assign n952 = ~n575 & ~n951 ;
  assign n953 = n574 & n952 ;
  assign n954 = ~n950 & n953 ;
  assign n955 = ~n582 & ~n954 ;
  assign n956 = ~n580 & n955 ;
  assign n957 = ~n571 & n956 ;
  assign n958 = ~x347 & x475 ;
  assign n959 = ~x346 & x474 ;
  assign n960 = ~n958 & ~n959 ;
  assign n961 = ~x345 & x473 ;
  assign n962 = ~x344 & x472 ;
  assign n963 = ~n961 & ~n962 ;
  assign n964 = n960 & n963 ;
  assign n965 = ~n957 & n964 ;
  assign n966 = x347 & ~x475 ;
  assign n967 = x344 & ~x472 ;
  assign n968 = ~n961 & n967 ;
  assign n969 = x345 & ~x473 ;
  assign n970 = ~n968 & ~n969 ;
  assign n971 = x346 & ~x474 ;
  assign n972 = n970 & ~n971 ;
  assign n973 = n960 & ~n972 ;
  assign n974 = ~n966 & ~n973 ;
  assign n975 = ~n965 & n974 ;
  assign n976 = ~x348 & x476 ;
  assign n977 = ~n563 & ~n976 ;
  assign n978 = n562 & n977 ;
  assign n979 = ~n975 & n978 ;
  assign n980 = ~n570 & ~n979 ;
  assign n981 = ~n568 & n980 ;
  assign n982 = ~n559 & n981 ;
  assign n983 = ~n558 & ~n982 ;
  assign n984 = n557 & n983 ;
  assign n985 = ~n554 & n984 ;
  assign n986 = x355 & ~x483 ;
  assign n987 = ~x480 & ~n558 ;
  assign n988 = x352 & n987 ;
  assign n989 = x353 & ~x481 ;
  assign n990 = ~n988 & ~n989 ;
  assign n991 = x354 & ~x482 ;
  assign n992 = n990 & ~n991 ;
  assign n993 = n557 & ~n992 ;
  assign n994 = ~n986 & ~n993 ;
  assign n995 = ~n985 & n994 ;
  assign n996 = ~x356 & x484 ;
  assign n997 = ~n546 & ~n996 ;
  assign n998 = n545 & n997 ;
  assign n999 = ~n995 & n998 ;
  assign n1000 = ~n553 & ~n999 ;
  assign n1001 = ~n551 & n1000 ;
  assign n1002 = ~n542 & n1001 ;
  assign n1003 = ~x363 & x491 ;
  assign n1004 = ~x362 & x490 ;
  assign n1005 = ~n1003 & ~n1004 ;
  assign n1006 = ~x361 & x489 ;
  assign n1007 = ~x360 & x488 ;
  assign n1008 = ~n1006 & ~n1007 ;
  assign n1009 = n1005 & n1008 ;
  assign n1010 = ~n1002 & n1009 ;
  assign n1011 = x363 & ~x491 ;
  assign n1012 = x360 & ~x488 ;
  assign n1013 = ~n1006 & n1012 ;
  assign n1014 = x361 & ~x489 ;
  assign n1015 = ~n1013 & ~n1014 ;
  assign n1016 = x362 & ~x490 ;
  assign n1017 = n1015 & ~n1016 ;
  assign n1018 = n1005 & ~n1017 ;
  assign n1019 = ~n1011 & ~n1018 ;
  assign n1020 = ~n1010 & n1019 ;
  assign n1021 = ~x364 & x492 ;
  assign n1022 = ~n534 & ~n1021 ;
  assign n1023 = n533 & n1022 ;
  assign n1024 = ~n1020 & n1023 ;
  assign n1025 = ~n541 & ~n1024 ;
  assign n1026 = ~n539 & n1025 ;
  assign n1027 = ~n530 & n1026 ;
  assign n1028 = ~n529 & ~n1027 ;
  assign n1029 = n528 & n1028 ;
  assign n1030 = ~n525 & n1029 ;
  assign n1031 = x371 & ~x499 ;
  assign n1032 = ~x496 & ~n529 ;
  assign n1033 = x368 & n1032 ;
  assign n1034 = x369 & ~x497 ;
  assign n1035 = ~n1033 & ~n1034 ;
  assign n1036 = x370 & ~x498 ;
  assign n1037 = n1035 & ~n1036 ;
  assign n1038 = n528 & ~n1037 ;
  assign n1039 = ~n1031 & ~n1038 ;
  assign n1040 = ~n1030 & n1039 ;
  assign n1041 = ~x372 & x500 ;
  assign n1042 = ~n517 & ~n1041 ;
  assign n1043 = n516 & n1042 ;
  assign n1044 = ~n1040 & n1043 ;
  assign n1045 = ~n524 & ~n1044 ;
  assign n1046 = ~n522 & n1045 ;
  assign n1047 = ~n513 & n1046 ;
  assign n1048 = ~x379 & x507 ;
  assign n1049 = ~x378 & x506 ;
  assign n1050 = ~n1048 & ~n1049 ;
  assign n1051 = ~x377 & x505 ;
  assign n1052 = ~x376 & x504 ;
  assign n1053 = ~n1051 & ~n1052 ;
  assign n1054 = n1050 & n1053 ;
  assign n1055 = ~n1047 & n1054 ;
  assign n1056 = x379 & ~x507 ;
  assign n1057 = x376 & ~x504 ;
  assign n1058 = ~n1051 & n1057 ;
  assign n1059 = x377 & ~x505 ;
  assign n1060 = ~n1058 & ~n1059 ;
  assign n1061 = x378 & ~x506 ;
  assign n1062 = n1060 & ~n1061 ;
  assign n1063 = n1050 & ~n1062 ;
  assign n1064 = ~n1056 & ~n1063 ;
  assign n1065 = ~n1055 & n1064 ;
  assign n1066 = ~x380 & x508 ;
  assign n1067 = x383 & ~x511 ;
  assign n1068 = ~x382 & x510 ;
  assign n1069 = ~x381 & x509 ;
  assign n1070 = ~n1068 & ~n1069 ;
  assign n1071 = ~n1067 & n1070 ;
  assign n1072 = ~n1066 & n1071 ;
  assign n1073 = ~n1065 & n1072 ;
  assign n1074 = x380 & ~x508 ;
  assign n1075 = x381 & ~x509 ;
  assign n1076 = ~n1074 & ~n1075 ;
  assign n1077 = n1070 & ~n1076 ;
  assign n1078 = x382 & ~x510 ;
  assign n1079 = ~n1077 & ~n1078 ;
  assign n1080 = ~n1067 & ~n1079 ;
  assign n1081 = ~n1073 & ~n1080 ;
  assign n1082 = ~x383 & x511 ;
  assign n1083 = n1081 & ~n1082 ;
  assign n1084 = x384 & n1083 ;
  assign n1085 = x256 & ~n1083 ;
  assign n1086 = ~n1084 & ~n1085 ;
  assign n1087 = ~x511 & n1081 ;
  assign n1088 = x383 & ~n1087 ;
  assign n1089 = x119 & ~x247 ;
  assign n1090 = ~x119 & x247 ;
  assign n1091 = ~x118 & x246 ;
  assign n1092 = ~n1090 & ~n1091 ;
  assign n1093 = ~x117 & x245 ;
  assign n1094 = x116 & ~x244 ;
  assign n1095 = ~n1093 & n1094 ;
  assign n1096 = x117 & ~x245 ;
  assign n1097 = ~n1095 & ~n1096 ;
  assign n1098 = n1092 & ~n1097 ;
  assign n1099 = ~x246 & ~n1090 ;
  assign n1100 = x118 & n1099 ;
  assign n1101 = ~x112 & x240 ;
  assign n1102 = ~x115 & x243 ;
  assign n1103 = ~x114 & x242 ;
  assign n1104 = ~n1102 & ~n1103 ;
  assign n1105 = ~x113 & x241 ;
  assign n1106 = x111 & ~x239 ;
  assign n1107 = ~x111 & x239 ;
  assign n1108 = ~x110 & x238 ;
  assign n1109 = ~n1107 & ~n1108 ;
  assign n1110 = ~x109 & x237 ;
  assign n1111 = x108 & ~x236 ;
  assign n1112 = ~n1110 & n1111 ;
  assign n1113 = x109 & ~x237 ;
  assign n1114 = ~n1112 & ~n1113 ;
  assign n1115 = n1109 & ~n1114 ;
  assign n1116 = ~x238 & ~n1107 ;
  assign n1117 = x110 & n1116 ;
  assign n1118 = x103 & ~x231 ;
  assign n1119 = ~x103 & x231 ;
  assign n1120 = ~x102 & x230 ;
  assign n1121 = ~n1119 & ~n1120 ;
  assign n1122 = ~x101 & x229 ;
  assign n1123 = x100 & ~x228 ;
  assign n1124 = ~n1122 & n1123 ;
  assign n1125 = x101 & ~x229 ;
  assign n1126 = ~n1124 & ~n1125 ;
  assign n1127 = n1121 & ~n1126 ;
  assign n1128 = ~x230 & ~n1119 ;
  assign n1129 = x102 & n1128 ;
  assign n1130 = ~x96 & x224 ;
  assign n1131 = ~x99 & x227 ;
  assign n1132 = ~x98 & x226 ;
  assign n1133 = ~n1131 & ~n1132 ;
  assign n1134 = ~x97 & x225 ;
  assign n1135 = x95 & ~x223 ;
  assign n1136 = ~x95 & x223 ;
  assign n1137 = ~x94 & x222 ;
  assign n1138 = ~n1136 & ~n1137 ;
  assign n1139 = ~x93 & x221 ;
  assign n1140 = x92 & ~x220 ;
  assign n1141 = ~n1139 & n1140 ;
  assign n1142 = x93 & ~x221 ;
  assign n1143 = ~n1141 & ~n1142 ;
  assign n1144 = n1138 & ~n1143 ;
  assign n1145 = ~x222 & ~n1136 ;
  assign n1146 = x94 & n1145 ;
  assign n1147 = x87 & ~x215 ;
  assign n1148 = ~x87 & x215 ;
  assign n1149 = ~x86 & x214 ;
  assign n1150 = ~n1148 & ~n1149 ;
  assign n1151 = ~x85 & x213 ;
  assign n1152 = x84 & ~x212 ;
  assign n1153 = ~n1151 & n1152 ;
  assign n1154 = x85 & ~x213 ;
  assign n1155 = ~n1153 & ~n1154 ;
  assign n1156 = n1150 & ~n1155 ;
  assign n1157 = ~x214 & ~n1148 ;
  assign n1158 = x86 & n1157 ;
  assign n1159 = ~x80 & x208 ;
  assign n1160 = ~x83 & x211 ;
  assign n1161 = ~x82 & x210 ;
  assign n1162 = ~n1160 & ~n1161 ;
  assign n1163 = ~x81 & x209 ;
  assign n1164 = x79 & ~x207 ;
  assign n1165 = ~x79 & x207 ;
  assign n1166 = ~x78 & x206 ;
  assign n1167 = ~n1165 & ~n1166 ;
  assign n1168 = ~x77 & x205 ;
  assign n1169 = x76 & ~x204 ;
  assign n1170 = ~n1168 & n1169 ;
  assign n1171 = x77 & ~x205 ;
  assign n1172 = ~n1170 & ~n1171 ;
  assign n1173 = n1167 & ~n1172 ;
  assign n1174 = ~x206 & ~n1165 ;
  assign n1175 = x78 & n1174 ;
  assign n1176 = x71 & ~x199 ;
  assign n1177 = ~x71 & x199 ;
  assign n1178 = ~x70 & x198 ;
  assign n1179 = ~n1177 & ~n1178 ;
  assign n1180 = ~x69 & x197 ;
  assign n1181 = x68 & ~x196 ;
  assign n1182 = ~n1180 & n1181 ;
  assign n1183 = x69 & ~x197 ;
  assign n1184 = ~n1182 & ~n1183 ;
  assign n1185 = n1179 & ~n1184 ;
  assign n1186 = ~x198 & ~n1177 ;
  assign n1187 = x70 & n1186 ;
  assign n1188 = ~x67 & x195 ;
  assign n1189 = ~x66 & x194 ;
  assign n1190 = ~n1188 & ~n1189 ;
  assign n1191 = ~x65 & x193 ;
  assign n1192 = x63 & ~x191 ;
  assign n1193 = ~x63 & x191 ;
  assign n1194 = ~x62 & x190 ;
  assign n1195 = ~n1193 & ~n1194 ;
  assign n1196 = ~x60 & x188 ;
  assign n1197 = ~x61 & x189 ;
  assign n1198 = ~n1196 & ~n1197 ;
  assign n1199 = n1195 & n1198 ;
  assign n1200 = x59 & ~x187 ;
  assign n1201 = ~x59 & x187 ;
  assign n1202 = ~x58 & x186 ;
  assign n1203 = ~n1201 & ~n1202 ;
  assign n1204 = ~x57 & x185 ;
  assign n1205 = x56 & ~x184 ;
  assign n1206 = ~n1204 & n1205 ;
  assign n1207 = x57 & ~x185 ;
  assign n1208 = ~n1206 & ~n1207 ;
  assign n1209 = x58 & ~x186 ;
  assign n1210 = n1208 & ~n1209 ;
  assign n1211 = n1203 & ~n1210 ;
  assign n1212 = ~n1200 & ~n1211 ;
  assign n1213 = n1199 & ~n1212 ;
  assign n1214 = x60 & ~x188 ;
  assign n1215 = ~n1197 & n1214 ;
  assign n1216 = x61 & ~x189 ;
  assign n1217 = ~n1215 & ~n1216 ;
  assign n1218 = n1195 & ~n1217 ;
  assign n1219 = ~x190 & ~n1193 ;
  assign n1220 = x62 & n1219 ;
  assign n1221 = x47 & ~x175 ;
  assign n1222 = ~x47 & x175 ;
  assign n1223 = ~x46 & x174 ;
  assign n1224 = ~n1222 & ~n1223 ;
  assign n1225 = ~x44 & x172 ;
  assign n1226 = ~x45 & x173 ;
  assign n1227 = ~n1225 & ~n1226 ;
  assign n1228 = n1224 & n1227 ;
  assign n1229 = x43 & ~x171 ;
  assign n1230 = ~x43 & x171 ;
  assign n1231 = ~x42 & x170 ;
  assign n1232 = ~n1230 & ~n1231 ;
  assign n1233 = ~x41 & x169 ;
  assign n1234 = x40 & ~x168 ;
  assign n1235 = ~n1233 & n1234 ;
  assign n1236 = x41 & ~x169 ;
  assign n1237 = ~n1235 & ~n1236 ;
  assign n1238 = x42 & ~x170 ;
  assign n1239 = n1237 & ~n1238 ;
  assign n1240 = n1232 & ~n1239 ;
  assign n1241 = ~n1229 & ~n1240 ;
  assign n1242 = n1228 & ~n1241 ;
  assign n1243 = x44 & ~x172 ;
  assign n1244 = ~n1226 & n1243 ;
  assign n1245 = x45 & ~x173 ;
  assign n1246 = ~n1244 & ~n1245 ;
  assign n1247 = n1224 & ~n1246 ;
  assign n1248 = ~x174 & ~n1222 ;
  assign n1249 = x46 & n1248 ;
  assign n1250 = ~x32 & x160 ;
  assign n1251 = ~x31 & x159 ;
  assign n1252 = ~x30 & x158 ;
  assign n1253 = ~x29 & x157 ;
  assign n1254 = ~x28 & x156 ;
  assign n1255 = ~x27 & x155 ;
  assign n1256 = ~x26 & x154 ;
  assign n1257 = ~x23 & x151 ;
  assign n1258 = ~x22 & x150 ;
  assign n1259 = ~x21 & x149 ;
  assign n1260 = ~x20 & x148 ;
  assign n1261 = ~x19 & x147 ;
  assign n1262 = ~x18 & x146 ;
  assign n1263 = ~x15 & x143 ;
  assign n1264 = ~x14 & x142 ;
  assign n1265 = ~x13 & x141 ;
  assign n1266 = ~x12 & x140 ;
  assign n1267 = ~x11 & x139 ;
  assign n1268 = ~x10 & x138 ;
  assign n1269 = ~x7 & x135 ;
  assign n1270 = ~x6 & x134 ;
  assign n1271 = ~x3 & x131 ;
  assign n1272 = x0 & ~x128 ;
  assign n1273 = x1 & ~x129 ;
  assign n1274 = ~n1272 & ~n1273 ;
  assign n1275 = ~x2 & x130 ;
  assign n1276 = ~x1 & x129 ;
  assign n1277 = ~n1275 & ~n1276 ;
  assign n1278 = ~n1274 & n1277 ;
  assign n1279 = x2 & ~x130 ;
  assign n1280 = ~n1278 & ~n1279 ;
  assign n1281 = ~n1271 & ~n1280 ;
  assign n1282 = x3 & ~x131 ;
  assign n1283 = ~n1281 & ~n1282 ;
  assign n1284 = ~x4 & n1283 ;
  assign n1285 = ~x132 & ~n1284 ;
  assign n1286 = x4 & ~n1283 ;
  assign n1287 = ~n1285 & ~n1286 ;
  assign n1288 = ~x5 & n1287 ;
  assign n1289 = ~x133 & ~n1288 ;
  assign n1290 = x5 & ~n1287 ;
  assign n1291 = ~n1289 & ~n1290 ;
  assign n1292 = ~n1270 & ~n1291 ;
  assign n1293 = x6 & ~x134 ;
  assign n1294 = ~n1292 & ~n1293 ;
  assign n1295 = ~n1269 & ~n1294 ;
  assign n1296 = x7 & ~x135 ;
  assign n1297 = ~n1295 & ~n1296 ;
  assign n1298 = ~x8 & n1297 ;
  assign n1299 = ~x136 & ~n1298 ;
  assign n1300 = x8 & ~n1297 ;
  assign n1301 = ~n1299 & ~n1300 ;
  assign n1302 = ~x9 & n1301 ;
  assign n1303 = ~x137 & ~n1302 ;
  assign n1304 = x9 & ~n1301 ;
  assign n1305 = ~n1303 & ~n1304 ;
  assign n1306 = ~n1268 & ~n1305 ;
  assign n1307 = x10 & ~x138 ;
  assign n1308 = ~n1306 & ~n1307 ;
  assign n1309 = ~n1267 & ~n1308 ;
  assign n1310 = x11 & ~x139 ;
  assign n1311 = ~n1309 & ~n1310 ;
  assign n1312 = ~n1266 & ~n1311 ;
  assign n1313 = x12 & ~x140 ;
  assign n1314 = ~n1312 & ~n1313 ;
  assign n1315 = ~n1265 & ~n1314 ;
  assign n1316 = x13 & ~x141 ;
  assign n1317 = ~n1315 & ~n1316 ;
  assign n1318 = ~n1264 & ~n1317 ;
  assign n1319 = x14 & ~x142 ;
  assign n1320 = ~n1318 & ~n1319 ;
  assign n1321 = ~n1263 & ~n1320 ;
  assign n1322 = x15 & ~x143 ;
  assign n1323 = ~n1321 & ~n1322 ;
  assign n1324 = ~x16 & n1323 ;
  assign n1325 = ~x144 & ~n1324 ;
  assign n1326 = x16 & ~n1323 ;
  assign n1327 = ~n1325 & ~n1326 ;
  assign n1328 = ~x17 & n1327 ;
  assign n1329 = ~x145 & ~n1328 ;
  assign n1330 = x17 & ~n1327 ;
  assign n1331 = ~n1329 & ~n1330 ;
  assign n1332 = ~n1262 & ~n1331 ;
  assign n1333 = x18 & ~x146 ;
  assign n1334 = ~n1332 & ~n1333 ;
  assign n1335 = ~n1261 & ~n1334 ;
  assign n1336 = x19 & ~x147 ;
  assign n1337 = ~n1335 & ~n1336 ;
  assign n1338 = ~n1260 & ~n1337 ;
  assign n1339 = x20 & ~x148 ;
  assign n1340 = ~n1338 & ~n1339 ;
  assign n1341 = ~n1259 & ~n1340 ;
  assign n1342 = x21 & ~x149 ;
  assign n1343 = ~n1341 & ~n1342 ;
  assign n1344 = ~n1258 & ~n1343 ;
  assign n1345 = x22 & ~x150 ;
  assign n1346 = ~n1344 & ~n1345 ;
  assign n1347 = ~n1257 & ~n1346 ;
  assign n1348 = x23 & ~x151 ;
  assign n1349 = ~n1347 & ~n1348 ;
  assign n1350 = ~x24 & n1349 ;
  assign n1351 = ~x152 & ~n1350 ;
  assign n1352 = x24 & ~n1349 ;
  assign n1353 = ~n1351 & ~n1352 ;
  assign n1354 = ~x25 & n1353 ;
  assign n1355 = ~x153 & ~n1354 ;
  assign n1356 = x25 & ~n1353 ;
  assign n1357 = ~n1355 & ~n1356 ;
  assign n1358 = ~n1256 & ~n1357 ;
  assign n1359 = x26 & ~x154 ;
  assign n1360 = ~n1358 & ~n1359 ;
  assign n1361 = ~n1255 & ~n1360 ;
  assign n1362 = x27 & ~x155 ;
  assign n1363 = ~n1361 & ~n1362 ;
  assign n1364 = ~n1254 & ~n1363 ;
  assign n1365 = x28 & ~x156 ;
  assign n1366 = ~n1364 & ~n1365 ;
  assign n1367 = ~n1253 & ~n1366 ;
  assign n1368 = x29 & ~x157 ;
  assign n1369 = ~n1367 & ~n1368 ;
  assign n1370 = ~n1252 & ~n1369 ;
  assign n1371 = x30 & ~x158 ;
  assign n1372 = ~n1370 & ~n1371 ;
  assign n1373 = ~n1251 & ~n1372 ;
  assign n1374 = x31 & ~x159 ;
  assign n1375 = ~n1373 & ~n1374 ;
  assign n1376 = ~x39 & x167 ;
  assign n1377 = ~x38 & x166 ;
  assign n1378 = ~n1376 & ~n1377 ;
  assign n1379 = ~x36 & x164 ;
  assign n1380 = ~x37 & x165 ;
  assign n1381 = ~n1379 & ~n1380 ;
  assign n1382 = n1378 & n1381 ;
  assign n1383 = ~x33 & x161 ;
  assign n1384 = ~x35 & x163 ;
  assign n1385 = ~x34 & x162 ;
  assign n1386 = ~n1384 & ~n1385 ;
  assign n1387 = ~n1383 & n1386 ;
  assign n1388 = n1382 & n1387 ;
  assign n1389 = ~n1375 & n1388 ;
  assign n1390 = ~n1250 & n1389 ;
  assign n1391 = x39 & ~x167 ;
  assign n1392 = x36 & ~x164 ;
  assign n1393 = ~n1380 & n1392 ;
  assign n1394 = x37 & ~x165 ;
  assign n1395 = ~n1393 & ~n1394 ;
  assign n1396 = n1378 & ~n1395 ;
  assign n1397 = ~x166 & ~n1376 ;
  assign n1398 = x38 & n1397 ;
  assign n1399 = x35 & ~x163 ;
  assign n1400 = ~x160 & ~n1383 ;
  assign n1401 = x32 & n1400 ;
  assign n1402 = x33 & ~x161 ;
  assign n1403 = ~n1401 & ~n1402 ;
  assign n1404 = x34 & ~x162 ;
  assign n1405 = n1403 & ~n1404 ;
  assign n1406 = n1386 & ~n1405 ;
  assign n1407 = ~n1399 & ~n1406 ;
  assign n1408 = n1382 & ~n1407 ;
  assign n1409 = ~n1398 & ~n1408 ;
  assign n1410 = ~n1396 & n1409 ;
  assign n1411 = ~n1391 & n1410 ;
  assign n1412 = ~n1390 & n1411 ;
  assign n1413 = ~x40 & x168 ;
  assign n1414 = ~n1233 & ~n1413 ;
  assign n1415 = n1232 & n1414 ;
  assign n1416 = n1228 & n1415 ;
  assign n1417 = ~n1412 & n1416 ;
  assign n1418 = ~n1249 & ~n1417 ;
  assign n1419 = ~n1247 & n1418 ;
  assign n1420 = ~n1242 & n1419 ;
  assign n1421 = ~n1221 & n1420 ;
  assign n1422 = ~x48 & x176 ;
  assign n1423 = ~x55 & x183 ;
  assign n1424 = ~x54 & x182 ;
  assign n1425 = ~n1423 & ~n1424 ;
  assign n1426 = ~x53 & x181 ;
  assign n1427 = ~x52 & x180 ;
  assign n1428 = ~n1426 & ~n1427 ;
  assign n1429 = n1425 & n1428 ;
  assign n1430 = ~x49 & x177 ;
  assign n1431 = ~x51 & x179 ;
  assign n1432 = ~x50 & x178 ;
  assign n1433 = ~n1431 & ~n1432 ;
  assign n1434 = ~n1430 & n1433 ;
  assign n1435 = n1429 & n1434 ;
  assign n1436 = ~n1422 & n1435 ;
  assign n1437 = ~n1421 & n1436 ;
  assign n1438 = x55 & ~x183 ;
  assign n1439 = x51 & ~x179 ;
  assign n1440 = ~x176 & ~n1430 ;
  assign n1441 = x48 & n1440 ;
  assign n1442 = x49 & ~x177 ;
  assign n1443 = ~n1441 & ~n1442 ;
  assign n1444 = x50 & ~x178 ;
  assign n1445 = n1443 & ~n1444 ;
  assign n1446 = n1433 & ~n1445 ;
  assign n1447 = ~n1439 & ~n1446 ;
  assign n1448 = n1429 & ~n1447 ;
  assign n1449 = x52 & ~x180 ;
  assign n1450 = ~n1426 & n1449 ;
  assign n1451 = x53 & ~x181 ;
  assign n1452 = ~n1450 & ~n1451 ;
  assign n1453 = x54 & ~x182 ;
  assign n1454 = n1452 & ~n1453 ;
  assign n1455 = n1425 & ~n1454 ;
  assign n1456 = ~n1448 & ~n1455 ;
  assign n1457 = ~n1438 & n1456 ;
  assign n1458 = ~n1437 & n1457 ;
  assign n1459 = ~x56 & x184 ;
  assign n1460 = ~n1204 & ~n1459 ;
  assign n1461 = n1199 & n1460 ;
  assign n1462 = n1203 & n1461 ;
  assign n1463 = ~n1458 & n1462 ;
  assign n1464 = ~n1220 & ~n1463 ;
  assign n1465 = ~n1218 & n1464 ;
  assign n1466 = ~n1213 & n1465 ;
  assign n1467 = ~n1192 & n1466 ;
  assign n1468 = ~x64 & x192 ;
  assign n1469 = ~n1467 & ~n1468 ;
  assign n1470 = ~n1191 & n1469 ;
  assign n1471 = n1190 & n1470 ;
  assign n1472 = x67 & ~x195 ;
  assign n1473 = x64 & ~x192 ;
  assign n1474 = ~n1191 & n1473 ;
  assign n1475 = x65 & ~x193 ;
  assign n1476 = ~n1474 & ~n1475 ;
  assign n1477 = x66 & ~x194 ;
  assign n1478 = n1476 & ~n1477 ;
  assign n1479 = n1190 & ~n1478 ;
  assign n1480 = ~n1472 & ~n1479 ;
  assign n1481 = ~n1471 & n1480 ;
  assign n1482 = ~x68 & x196 ;
  assign n1483 = ~n1180 & ~n1482 ;
  assign n1484 = n1179 & n1483 ;
  assign n1485 = ~n1481 & n1484 ;
  assign n1486 = ~n1187 & ~n1485 ;
  assign n1487 = ~n1185 & n1486 ;
  assign n1488 = ~n1176 & n1487 ;
  assign n1489 = ~x75 & x203 ;
  assign n1490 = ~x74 & x202 ;
  assign n1491 = ~n1489 & ~n1490 ;
  assign n1492 = ~x73 & x201 ;
  assign n1493 = ~x72 & x200 ;
  assign n1494 = ~n1492 & ~n1493 ;
  assign n1495 = n1491 & n1494 ;
  assign n1496 = ~n1488 & n1495 ;
  assign n1497 = x75 & ~x203 ;
  assign n1498 = x72 & ~x200 ;
  assign n1499 = ~n1492 & n1498 ;
  assign n1500 = x73 & ~x201 ;
  assign n1501 = ~n1499 & ~n1500 ;
  assign n1502 = x74 & ~x202 ;
  assign n1503 = n1501 & ~n1502 ;
  assign n1504 = n1491 & ~n1503 ;
  assign n1505 = ~n1497 & ~n1504 ;
  assign n1506 = ~n1496 & n1505 ;
  assign n1507 = ~x76 & x204 ;
  assign n1508 = ~n1168 & ~n1507 ;
  assign n1509 = n1167 & n1508 ;
  assign n1510 = ~n1506 & n1509 ;
  assign n1511 = ~n1175 & ~n1510 ;
  assign n1512 = ~n1173 & n1511 ;
  assign n1513 = ~n1164 & n1512 ;
  assign n1514 = ~n1163 & ~n1513 ;
  assign n1515 = n1162 & n1514 ;
  assign n1516 = ~n1159 & n1515 ;
  assign n1517 = x83 & ~x211 ;
  assign n1518 = ~x208 & ~n1163 ;
  assign n1519 = x80 & n1518 ;
  assign n1520 = x81 & ~x209 ;
  assign n1521 = ~n1519 & ~n1520 ;
  assign n1522 = x82 & ~x210 ;
  assign n1523 = n1521 & ~n1522 ;
  assign n1524 = n1162 & ~n1523 ;
  assign n1525 = ~n1517 & ~n1524 ;
  assign n1526 = ~n1516 & n1525 ;
  assign n1527 = ~x84 & x212 ;
  assign n1528 = ~n1151 & ~n1527 ;
  assign n1529 = n1150 & n1528 ;
  assign n1530 = ~n1526 & n1529 ;
  assign n1531 = ~n1158 & ~n1530 ;
  assign n1532 = ~n1156 & n1531 ;
  assign n1533 = ~n1147 & n1532 ;
  assign n1534 = ~x91 & x219 ;
  assign n1535 = ~x90 & x218 ;
  assign n1536 = ~n1534 & ~n1535 ;
  assign n1537 = ~x89 & x217 ;
  assign n1538 = ~x88 & x216 ;
  assign n1539 = ~n1537 & ~n1538 ;
  assign n1540 = n1536 & n1539 ;
  assign n1541 = ~n1533 & n1540 ;
  assign n1542 = x91 & ~x219 ;
  assign n1543 = x88 & ~x216 ;
  assign n1544 = ~n1537 & n1543 ;
  assign n1545 = x89 & ~x217 ;
  assign n1546 = ~n1544 & ~n1545 ;
  assign n1547 = x90 & ~x218 ;
  assign n1548 = n1546 & ~n1547 ;
  assign n1549 = n1536 & ~n1548 ;
  assign n1550 = ~n1542 & ~n1549 ;
  assign n1551 = ~n1541 & n1550 ;
  assign n1552 = ~x92 & x220 ;
  assign n1553 = ~n1139 & ~n1552 ;
  assign n1554 = n1138 & n1553 ;
  assign n1555 = ~n1551 & n1554 ;
  assign n1556 = ~n1146 & ~n1555 ;
  assign n1557 = ~n1144 & n1556 ;
  assign n1558 = ~n1135 & n1557 ;
  assign n1559 = ~n1134 & ~n1558 ;
  assign n1560 = n1133 & n1559 ;
  assign n1561 = ~n1130 & n1560 ;
  assign n1562 = x99 & ~x227 ;
  assign n1563 = ~x224 & ~n1134 ;
  assign n1564 = x96 & n1563 ;
  assign n1565 = x97 & ~x225 ;
  assign n1566 = ~n1564 & ~n1565 ;
  assign n1567 = x98 & ~x226 ;
  assign n1568 = n1566 & ~n1567 ;
  assign n1569 = n1133 & ~n1568 ;
  assign n1570 = ~n1562 & ~n1569 ;
  assign n1571 = ~n1561 & n1570 ;
  assign n1572 = ~x100 & x228 ;
  assign n1573 = ~n1122 & ~n1572 ;
  assign n1574 = n1121 & n1573 ;
  assign n1575 = ~n1571 & n1574 ;
  assign n1576 = ~n1129 & ~n1575 ;
  assign n1577 = ~n1127 & n1576 ;
  assign n1578 = ~n1118 & n1577 ;
  assign n1579 = ~x107 & x235 ;
  assign n1580 = ~x106 & x234 ;
  assign n1581 = ~n1579 & ~n1580 ;
  assign n1582 = ~x105 & x233 ;
  assign n1583 = ~x104 & x232 ;
  assign n1584 = ~n1582 & ~n1583 ;
  assign n1585 = n1581 & n1584 ;
  assign n1586 = ~n1578 & n1585 ;
  assign n1587 = x107 & ~x235 ;
  assign n1588 = x104 & ~x232 ;
  assign n1589 = ~n1582 & n1588 ;
  assign n1590 = x105 & ~x233 ;
  assign n1591 = ~n1589 & ~n1590 ;
  assign n1592 = x106 & ~x234 ;
  assign n1593 = n1591 & ~n1592 ;
  assign n1594 = n1581 & ~n1593 ;
  assign n1595 = ~n1587 & ~n1594 ;
  assign n1596 = ~n1586 & n1595 ;
  assign n1597 = ~x108 & x236 ;
  assign n1598 = ~n1110 & ~n1597 ;
  assign n1599 = n1109 & n1598 ;
  assign n1600 = ~n1596 & n1599 ;
  assign n1601 = ~n1117 & ~n1600 ;
  assign n1602 = ~n1115 & n1601 ;
  assign n1603 = ~n1106 & n1602 ;
  assign n1604 = ~n1105 & ~n1603 ;
  assign n1605 = n1104 & n1604 ;
  assign n1606 = ~n1101 & n1605 ;
  assign n1607 = x115 & ~x243 ;
  assign n1608 = ~x240 & ~n1105 ;
  assign n1609 = x112 & n1608 ;
  assign n1610 = x113 & ~x241 ;
  assign n1611 = ~n1609 & ~n1610 ;
  assign n1612 = x114 & ~x242 ;
  assign n1613 = n1611 & ~n1612 ;
  assign n1614 = n1104 & ~n1613 ;
  assign n1615 = ~n1607 & ~n1614 ;
  assign n1616 = ~n1606 & n1615 ;
  assign n1617 = ~x116 & x244 ;
  assign n1618 = ~n1093 & ~n1617 ;
  assign n1619 = n1092 & n1618 ;
  assign n1620 = ~n1616 & n1619 ;
  assign n1621 = ~n1100 & ~n1620 ;
  assign n1622 = ~n1098 & n1621 ;
  assign n1623 = ~n1089 & n1622 ;
  assign n1624 = ~x123 & x251 ;
  assign n1625 = ~x122 & x250 ;
  assign n1626 = ~n1624 & ~n1625 ;
  assign n1627 = ~x121 & x249 ;
  assign n1628 = ~x120 & x248 ;
  assign n1629 = ~n1627 & ~n1628 ;
  assign n1630 = n1626 & n1629 ;
  assign n1631 = ~n1623 & n1630 ;
  assign n1632 = x123 & ~x251 ;
  assign n1633 = x120 & ~x248 ;
  assign n1634 = ~n1627 & n1633 ;
  assign n1635 = x121 & ~x249 ;
  assign n1636 = ~n1634 & ~n1635 ;
  assign n1637 = x122 & ~x250 ;
  assign n1638 = n1636 & ~n1637 ;
  assign n1639 = n1626 & ~n1638 ;
  assign n1640 = ~n1632 & ~n1639 ;
  assign n1641 = ~n1631 & n1640 ;
  assign n1642 = ~x124 & x252 ;
  assign n1643 = x127 & ~x255 ;
  assign n1644 = ~x126 & x254 ;
  assign n1645 = ~x125 & x253 ;
  assign n1646 = ~n1644 & ~n1645 ;
  assign n1647 = ~n1643 & n1646 ;
  assign n1648 = ~n1642 & n1647 ;
  assign n1649 = ~n1641 & n1648 ;
  assign n1650 = x124 & ~x252 ;
  assign n1651 = x125 & ~x253 ;
  assign n1652 = ~n1650 & ~n1651 ;
  assign n1653 = n1646 & ~n1652 ;
  assign n1654 = x126 & ~x254 ;
  assign n1655 = ~n1653 & ~n1654 ;
  assign n1656 = ~n1643 & ~n1655 ;
  assign n1657 = ~n1649 & ~n1656 ;
  assign n1658 = ~x255 & n1657 ;
  assign n1659 = x127 & ~n1658 ;
  assign n1660 = n1088 & ~n1659 ;
  assign n1661 = ~x127 & x255 ;
  assign n1662 = n1657 & ~n1661 ;
  assign n1663 = x247 & n1662 ;
  assign n1664 = x119 & ~n1662 ;
  assign n1665 = ~n1663 & ~n1664 ;
  assign n1666 = x503 & n1083 ;
  assign n1667 = x375 & ~n1083 ;
  assign n1668 = ~n1666 & ~n1667 ;
  assign n1669 = ~n1665 & n1668 ;
  assign n1670 = n1665 & ~n1668 ;
  assign n1671 = x502 & n1083 ;
  assign n1672 = x374 & ~n1083 ;
  assign n1673 = ~n1671 & ~n1672 ;
  assign n1674 = x246 & n1662 ;
  assign n1675 = x118 & ~n1662 ;
  assign n1676 = ~n1674 & ~n1675 ;
  assign n1677 = ~n1673 & n1676 ;
  assign n1678 = ~n1670 & ~n1677 ;
  assign n1679 = x244 & n1662 ;
  assign n1680 = x116 & ~n1662 ;
  assign n1681 = ~n1679 & ~n1680 ;
  assign n1682 = x245 & n1662 ;
  assign n1683 = x117 & ~n1662 ;
  assign n1684 = ~n1682 & ~n1683 ;
  assign n1685 = x501 & n1083 ;
  assign n1686 = x373 & ~n1083 ;
  assign n1687 = ~n1685 & ~n1686 ;
  assign n1688 = n1684 & ~n1687 ;
  assign n1689 = x500 & n1083 ;
  assign n1690 = x372 & ~n1083 ;
  assign n1691 = ~n1689 & ~n1690 ;
  assign n1692 = ~n1688 & n1691 ;
  assign n1693 = ~n1681 & n1692 ;
  assign n1694 = ~n1684 & n1687 ;
  assign n1695 = ~n1693 & ~n1694 ;
  assign n1696 = n1678 & ~n1695 ;
  assign n1697 = n1673 & ~n1676 ;
  assign n1698 = ~n1670 & n1697 ;
  assign n1699 = x496 & n1083 ;
  assign n1700 = x368 & ~n1083 ;
  assign n1701 = ~n1699 & ~n1700 ;
  assign n1702 = x240 & n1662 ;
  assign n1703 = x112 & ~n1662 ;
  assign n1704 = ~n1702 & ~n1703 ;
  assign n1705 = ~n1701 & n1704 ;
  assign n1706 = x243 & n1662 ;
  assign n1707 = x115 & ~n1662 ;
  assign n1708 = ~n1706 & ~n1707 ;
  assign n1709 = x499 & n1083 ;
  assign n1710 = x371 & ~n1083 ;
  assign n1711 = ~n1709 & ~n1710 ;
  assign n1712 = n1708 & ~n1711 ;
  assign n1713 = x498 & n1083 ;
  assign n1714 = x370 & ~n1083 ;
  assign n1715 = ~n1713 & ~n1714 ;
  assign n1716 = x242 & n1662 ;
  assign n1717 = x114 & ~n1662 ;
  assign n1718 = ~n1716 & ~n1717 ;
  assign n1719 = ~n1715 & n1718 ;
  assign n1720 = ~n1712 & ~n1719 ;
  assign n1721 = x241 & n1662 ;
  assign n1722 = x113 & ~n1662 ;
  assign n1723 = ~n1721 & ~n1722 ;
  assign n1724 = x497 & n1083 ;
  assign n1725 = x369 & ~n1083 ;
  assign n1726 = ~n1724 & ~n1725 ;
  assign n1727 = n1723 & ~n1726 ;
  assign n1728 = x239 & n1662 ;
  assign n1729 = x111 & ~n1662 ;
  assign n1730 = ~n1728 & ~n1729 ;
  assign n1731 = x495 & n1083 ;
  assign n1732 = x367 & ~n1083 ;
  assign n1733 = ~n1731 & ~n1732 ;
  assign n1734 = ~n1730 & n1733 ;
  assign n1735 = n1730 & ~n1733 ;
  assign n1736 = x494 & n1083 ;
  assign n1737 = x366 & ~n1083 ;
  assign n1738 = ~n1736 & ~n1737 ;
  assign n1739 = x238 & n1662 ;
  assign n1740 = x110 & ~n1662 ;
  assign n1741 = ~n1739 & ~n1740 ;
  assign n1742 = ~n1738 & n1741 ;
  assign n1743 = ~n1735 & ~n1742 ;
  assign n1744 = x237 & n1662 ;
  assign n1745 = x109 & ~n1662 ;
  assign n1746 = ~n1744 & ~n1745 ;
  assign n1747 = x493 & n1083 ;
  assign n1748 = x365 & ~n1083 ;
  assign n1749 = ~n1747 & ~n1748 ;
  assign n1750 = n1746 & ~n1749 ;
  assign n1751 = x236 & n1662 ;
  assign n1752 = x108 & ~n1662 ;
  assign n1753 = ~n1751 & ~n1752 ;
  assign n1754 = x492 & n1083 ;
  assign n1755 = x364 & ~n1083 ;
  assign n1756 = ~n1754 & ~n1755 ;
  assign n1757 = ~n1753 & n1756 ;
  assign n1758 = ~n1750 & n1757 ;
  assign n1759 = ~n1746 & n1749 ;
  assign n1760 = ~n1758 & ~n1759 ;
  assign n1761 = n1743 & ~n1760 ;
  assign n1762 = n1738 & ~n1741 ;
  assign n1763 = ~n1735 & n1762 ;
  assign n1764 = x231 & n1662 ;
  assign n1765 = x103 & ~n1662 ;
  assign n1766 = ~n1764 & ~n1765 ;
  assign n1767 = x487 & n1083 ;
  assign n1768 = x359 & ~n1083 ;
  assign n1769 = ~n1767 & ~n1768 ;
  assign n1770 = ~n1766 & n1769 ;
  assign n1771 = n1766 & ~n1769 ;
  assign n1772 = x486 & n1083 ;
  assign n1773 = x358 & ~n1083 ;
  assign n1774 = ~n1772 & ~n1773 ;
  assign n1775 = x230 & n1662 ;
  assign n1776 = x102 & ~n1662 ;
  assign n1777 = ~n1775 & ~n1776 ;
  assign n1778 = ~n1774 & n1777 ;
  assign n1779 = ~n1771 & ~n1778 ;
  assign n1780 = x229 & n1662 ;
  assign n1781 = x101 & ~n1662 ;
  assign n1782 = ~n1780 & ~n1781 ;
  assign n1783 = x485 & n1083 ;
  assign n1784 = x357 & ~n1083 ;
  assign n1785 = ~n1783 & ~n1784 ;
  assign n1786 = n1782 & ~n1785 ;
  assign n1787 = x228 & n1662 ;
  assign n1788 = x100 & ~n1662 ;
  assign n1789 = ~n1787 & ~n1788 ;
  assign n1790 = x484 & n1083 ;
  assign n1791 = x356 & ~n1083 ;
  assign n1792 = ~n1790 & ~n1791 ;
  assign n1793 = ~n1789 & n1792 ;
  assign n1794 = ~n1786 & n1793 ;
  assign n1795 = ~n1782 & n1785 ;
  assign n1796 = ~n1794 & ~n1795 ;
  assign n1797 = n1779 & ~n1796 ;
  assign n1798 = n1774 & ~n1777 ;
  assign n1799 = ~n1771 & n1798 ;
  assign n1800 = x480 & n1083 ;
  assign n1801 = x352 & ~n1083 ;
  assign n1802 = ~n1800 & ~n1801 ;
  assign n1803 = x224 & n1662 ;
  assign n1804 = x96 & ~n1662 ;
  assign n1805 = ~n1803 & ~n1804 ;
  assign n1806 = ~n1802 & n1805 ;
  assign n1807 = x227 & n1662 ;
  assign n1808 = x99 & ~n1662 ;
  assign n1809 = ~n1807 & ~n1808 ;
  assign n1810 = x483 & n1083 ;
  assign n1811 = x355 & ~n1083 ;
  assign n1812 = ~n1810 & ~n1811 ;
  assign n1813 = n1809 & ~n1812 ;
  assign n1814 = x482 & n1083 ;
  assign n1815 = x354 & ~n1083 ;
  assign n1816 = ~n1814 & ~n1815 ;
  assign n1817 = x226 & n1662 ;
  assign n1818 = x98 & ~n1662 ;
  assign n1819 = ~n1817 & ~n1818 ;
  assign n1820 = ~n1816 & n1819 ;
  assign n1821 = ~n1813 & ~n1820 ;
  assign n1822 = x225 & n1662 ;
  assign n1823 = x97 & ~n1662 ;
  assign n1824 = ~n1822 & ~n1823 ;
  assign n1825 = x481 & n1083 ;
  assign n1826 = x353 & ~n1083 ;
  assign n1827 = ~n1825 & ~n1826 ;
  assign n1828 = n1824 & ~n1827 ;
  assign n1829 = x223 & n1662 ;
  assign n1830 = x95 & ~n1662 ;
  assign n1831 = ~n1829 & ~n1830 ;
  assign n1832 = x479 & n1083 ;
  assign n1833 = x351 & ~n1083 ;
  assign n1834 = ~n1832 & ~n1833 ;
  assign n1835 = ~n1831 & n1834 ;
  assign n1836 = n1831 & ~n1834 ;
  assign n1837 = x478 & n1083 ;
  assign n1838 = x350 & ~n1083 ;
  assign n1839 = ~n1837 & ~n1838 ;
  assign n1840 = x222 & n1662 ;
  assign n1841 = x94 & ~n1662 ;
  assign n1842 = ~n1840 & ~n1841 ;
  assign n1843 = ~n1839 & n1842 ;
  assign n1844 = ~n1836 & ~n1843 ;
  assign n1845 = x221 & n1662 ;
  assign n1846 = x93 & ~n1662 ;
  assign n1847 = ~n1845 & ~n1846 ;
  assign n1848 = x477 & n1083 ;
  assign n1849 = x349 & ~n1083 ;
  assign n1850 = ~n1848 & ~n1849 ;
  assign n1851 = n1847 & ~n1850 ;
  assign n1852 = x220 & n1662 ;
  assign n1853 = x92 & ~n1662 ;
  assign n1854 = ~n1852 & ~n1853 ;
  assign n1855 = x476 & n1083 ;
  assign n1856 = x348 & ~n1083 ;
  assign n1857 = ~n1855 & ~n1856 ;
  assign n1858 = ~n1854 & n1857 ;
  assign n1859 = ~n1851 & n1858 ;
  assign n1860 = ~n1847 & n1850 ;
  assign n1861 = ~n1859 & ~n1860 ;
  assign n1862 = n1844 & ~n1861 ;
  assign n1863 = n1839 & ~n1842 ;
  assign n1864 = ~n1836 & n1863 ;
  assign n1865 = x215 & n1662 ;
  assign n1866 = x87 & ~n1662 ;
  assign n1867 = ~n1865 & ~n1866 ;
  assign n1868 = x471 & n1083 ;
  assign n1869 = x343 & ~n1083 ;
  assign n1870 = ~n1868 & ~n1869 ;
  assign n1871 = ~n1867 & n1870 ;
  assign n1872 = n1867 & ~n1870 ;
  assign n1873 = x470 & n1083 ;
  assign n1874 = x342 & ~n1083 ;
  assign n1875 = ~n1873 & ~n1874 ;
  assign n1876 = x214 & n1662 ;
  assign n1877 = x86 & ~n1662 ;
  assign n1878 = ~n1876 & ~n1877 ;
  assign n1879 = ~n1875 & n1878 ;
  assign n1880 = ~n1872 & ~n1879 ;
  assign n1881 = x213 & n1662 ;
  assign n1882 = x85 & ~n1662 ;
  assign n1883 = ~n1881 & ~n1882 ;
  assign n1884 = x469 & n1083 ;
  assign n1885 = x341 & ~n1083 ;
  assign n1886 = ~n1884 & ~n1885 ;
  assign n1887 = n1883 & ~n1886 ;
  assign n1888 = x212 & n1662 ;
  assign n1889 = x84 & ~n1662 ;
  assign n1890 = ~n1888 & ~n1889 ;
  assign n1891 = x468 & n1083 ;
  assign n1892 = x340 & ~n1083 ;
  assign n1893 = ~n1891 & ~n1892 ;
  assign n1894 = ~n1890 & n1893 ;
  assign n1895 = ~n1887 & n1894 ;
  assign n1896 = ~n1883 & n1886 ;
  assign n1897 = ~n1895 & ~n1896 ;
  assign n1898 = n1880 & ~n1897 ;
  assign n1899 = n1875 & ~n1878 ;
  assign n1900 = ~n1872 & n1899 ;
  assign n1901 = x464 & n1083 ;
  assign n1902 = x336 & ~n1083 ;
  assign n1903 = ~n1901 & ~n1902 ;
  assign n1904 = x208 & n1662 ;
  assign n1905 = x80 & ~n1662 ;
  assign n1906 = ~n1904 & ~n1905 ;
  assign n1907 = ~n1903 & n1906 ;
  assign n1908 = x211 & n1662 ;
  assign n1909 = x83 & ~n1662 ;
  assign n1910 = ~n1908 & ~n1909 ;
  assign n1911 = x467 & n1083 ;
  assign n1912 = x339 & ~n1083 ;
  assign n1913 = ~n1911 & ~n1912 ;
  assign n1914 = n1910 & ~n1913 ;
  assign n1915 = x466 & n1083 ;
  assign n1916 = x338 & ~n1083 ;
  assign n1917 = ~n1915 & ~n1916 ;
  assign n1918 = x210 & n1662 ;
  assign n1919 = x82 & ~n1662 ;
  assign n1920 = ~n1918 & ~n1919 ;
  assign n1921 = ~n1917 & n1920 ;
  assign n1922 = ~n1914 & ~n1921 ;
  assign n1923 = x209 & n1662 ;
  assign n1924 = x81 & ~n1662 ;
  assign n1925 = ~n1923 & ~n1924 ;
  assign n1926 = x465 & n1083 ;
  assign n1927 = x337 & ~n1083 ;
  assign n1928 = ~n1926 & ~n1927 ;
  assign n1929 = n1925 & ~n1928 ;
  assign n1930 = x207 & n1662 ;
  assign n1931 = x79 & ~n1662 ;
  assign n1932 = ~n1930 & ~n1931 ;
  assign n1933 = x463 & n1083 ;
  assign n1934 = x335 & ~n1083 ;
  assign n1935 = ~n1933 & ~n1934 ;
  assign n1936 = ~n1932 & n1935 ;
  assign n1937 = n1932 & ~n1935 ;
  assign n1938 = x462 & n1083 ;
  assign n1939 = x334 & ~n1083 ;
  assign n1940 = ~n1938 & ~n1939 ;
  assign n1941 = x206 & n1662 ;
  assign n1942 = x78 & ~n1662 ;
  assign n1943 = ~n1941 & ~n1942 ;
  assign n1944 = ~n1940 & n1943 ;
  assign n1945 = ~n1937 & ~n1944 ;
  assign n1946 = x205 & n1662 ;
  assign n1947 = x77 & ~n1662 ;
  assign n1948 = ~n1946 & ~n1947 ;
  assign n1949 = x461 & n1083 ;
  assign n1950 = x333 & ~n1083 ;
  assign n1951 = ~n1949 & ~n1950 ;
  assign n1952 = n1948 & ~n1951 ;
  assign n1953 = x204 & n1662 ;
  assign n1954 = x76 & ~n1662 ;
  assign n1955 = ~n1953 & ~n1954 ;
  assign n1956 = x460 & n1083 ;
  assign n1957 = x332 & ~n1083 ;
  assign n1958 = ~n1956 & ~n1957 ;
  assign n1959 = ~n1955 & n1958 ;
  assign n1960 = ~n1952 & n1959 ;
  assign n1961 = ~n1948 & n1951 ;
  assign n1962 = ~n1960 & ~n1961 ;
  assign n1963 = n1945 & ~n1962 ;
  assign n1964 = n1940 & ~n1943 ;
  assign n1965 = ~n1937 & n1964 ;
  assign n1966 = x199 & n1662 ;
  assign n1967 = x71 & ~n1662 ;
  assign n1968 = ~n1966 & ~n1967 ;
  assign n1969 = x455 & n1083 ;
  assign n1970 = x327 & ~n1083 ;
  assign n1971 = ~n1969 & ~n1970 ;
  assign n1972 = ~n1968 & n1971 ;
  assign n1973 = n1968 & ~n1971 ;
  assign n1974 = x454 & n1083 ;
  assign n1975 = x326 & ~n1083 ;
  assign n1976 = ~n1974 & ~n1975 ;
  assign n1977 = x198 & n1662 ;
  assign n1978 = x70 & ~n1662 ;
  assign n1979 = ~n1977 & ~n1978 ;
  assign n1980 = ~n1976 & n1979 ;
  assign n1981 = ~n1973 & ~n1980 ;
  assign n1982 = x197 & n1662 ;
  assign n1983 = x69 & ~n1662 ;
  assign n1984 = ~n1982 & ~n1983 ;
  assign n1985 = x453 & n1083 ;
  assign n1986 = x325 & ~n1083 ;
  assign n1987 = ~n1985 & ~n1986 ;
  assign n1988 = n1984 & ~n1987 ;
  assign n1989 = x196 & n1662 ;
  assign n1990 = x68 & ~n1662 ;
  assign n1991 = ~n1989 & ~n1990 ;
  assign n1992 = x452 & n1083 ;
  assign n1993 = x324 & ~n1083 ;
  assign n1994 = ~n1992 & ~n1993 ;
  assign n1995 = ~n1991 & n1994 ;
  assign n1996 = ~n1988 & n1995 ;
  assign n1997 = ~n1984 & n1987 ;
  assign n1998 = ~n1996 & ~n1997 ;
  assign n1999 = n1981 & ~n1998 ;
  assign n2000 = n1976 & ~n1979 ;
  assign n2001 = ~n1973 & n2000 ;
  assign n2002 = x195 & n1662 ;
  assign n2003 = x67 & ~n1662 ;
  assign n2004 = ~n2002 & ~n2003 ;
  assign n2005 = x451 & n1083 ;
  assign n2006 = x323 & ~n1083 ;
  assign n2007 = ~n2005 & ~n2006 ;
  assign n2008 = n2004 & ~n2007 ;
  assign n2009 = x450 & n1083 ;
  assign n2010 = x322 & ~n1083 ;
  assign n2011 = ~n2009 & ~n2010 ;
  assign n2012 = x194 & n1662 ;
  assign n2013 = x66 & ~n1662 ;
  assign n2014 = ~n2012 & ~n2013 ;
  assign n2015 = ~n2011 & n2014 ;
  assign n2016 = ~n2008 & ~n2015 ;
  assign n2017 = x448 & n1083 ;
  assign n2018 = x320 & ~n1083 ;
  assign n2019 = ~n2017 & ~n2018 ;
  assign n2020 = x192 & n1662 ;
  assign n2021 = x64 & ~n1662 ;
  assign n2022 = ~n2020 & ~n2021 ;
  assign n2023 = ~n2019 & n2022 ;
  assign n2024 = x193 & n1662 ;
  assign n2025 = x65 & ~n1662 ;
  assign n2026 = ~n2024 & ~n2025 ;
  assign n2027 = x449 & n1083 ;
  assign n2028 = x321 & ~n1083 ;
  assign n2029 = ~n2027 & ~n2028 ;
  assign n2030 = n2026 & ~n2029 ;
  assign n2031 = x191 & n1662 ;
  assign n2032 = x63 & ~n1662 ;
  assign n2033 = ~n2031 & ~n2032 ;
  assign n2034 = x447 & n1083 ;
  assign n2035 = x319 & ~n1083 ;
  assign n2036 = ~n2034 & ~n2035 ;
  assign n2037 = ~n2033 & n2036 ;
  assign n2038 = n2033 & ~n2036 ;
  assign n2039 = x446 & n1083 ;
  assign n2040 = x318 & ~n1083 ;
  assign n2041 = ~n2039 & ~n2040 ;
  assign n2042 = x190 & n1662 ;
  assign n2043 = x62 & ~n1662 ;
  assign n2044 = ~n2042 & ~n2043 ;
  assign n2045 = ~n2041 & n2044 ;
  assign n2046 = ~n2038 & ~n2045 ;
  assign n2047 = x188 & n1662 ;
  assign n2048 = x60 & ~n1662 ;
  assign n2049 = ~n2047 & ~n2048 ;
  assign n2050 = x444 & n1083 ;
  assign n2051 = x316 & ~n1083 ;
  assign n2052 = ~n2050 & ~n2051 ;
  assign n2053 = n2049 & ~n2052 ;
  assign n2054 = x189 & n1662 ;
  assign n2055 = x61 & ~n1662 ;
  assign n2056 = ~n2054 & ~n2055 ;
  assign n2057 = x445 & n1083 ;
  assign n2058 = x317 & ~n1083 ;
  assign n2059 = ~n2057 & ~n2058 ;
  assign n2060 = n2056 & ~n2059 ;
  assign n2061 = ~n2053 & ~n2060 ;
  assign n2062 = n2046 & n2061 ;
  assign n2063 = x187 & n1662 ;
  assign n2064 = x59 & ~n1662 ;
  assign n2065 = ~n2063 & ~n2064 ;
  assign n2066 = x443 & n1083 ;
  assign n2067 = x315 & ~n1083 ;
  assign n2068 = ~n2066 & ~n2067 ;
  assign n2069 = ~n2065 & n2068 ;
  assign n2070 = n2065 & ~n2068 ;
  assign n2071 = x186 & n1662 ;
  assign n2072 = x58 & ~n1662 ;
  assign n2073 = ~n2071 & ~n2072 ;
  assign n2074 = x442 & n1083 ;
  assign n2075 = x314 & ~n1083 ;
  assign n2076 = ~n2074 & ~n2075 ;
  assign n2077 = n2073 & ~n2076 ;
  assign n2078 = ~n2070 & ~n2077 ;
  assign n2079 = x185 & n1662 ;
  assign n2080 = x57 & ~n1662 ;
  assign n2081 = ~n2079 & ~n2080 ;
  assign n2082 = x441 & n1083 ;
  assign n2083 = x313 & ~n1083 ;
  assign n2084 = ~n2082 & ~n2083 ;
  assign n2085 = n2081 & ~n2084 ;
  assign n2086 = x184 & n1662 ;
  assign n2087 = x56 & ~n1662 ;
  assign n2088 = ~n2086 & ~n2087 ;
  assign n2089 = x440 & n1083 ;
  assign n2090 = x312 & ~n1083 ;
  assign n2091 = ~n2089 & ~n2090 ;
  assign n2092 = ~n2088 & n2091 ;
  assign n2093 = ~n2085 & n2092 ;
  assign n2094 = ~n2081 & n2084 ;
  assign n2095 = ~n2093 & ~n2094 ;
  assign n2096 = ~n2073 & n2076 ;
  assign n2097 = n2095 & ~n2096 ;
  assign n2098 = n2078 & ~n2097 ;
  assign n2099 = ~n2069 & ~n2098 ;
  assign n2100 = n2062 & ~n2099 ;
  assign n2101 = ~n2049 & n2052 ;
  assign n2102 = ~n2060 & n2101 ;
  assign n2103 = ~n2056 & n2059 ;
  assign n2104 = ~n2102 & ~n2103 ;
  assign n2105 = n2046 & ~n2104 ;
  assign n2106 = n2041 & ~n2044 ;
  assign n2107 = ~n2038 & n2106 ;
  assign n2108 = x175 & n1662 ;
  assign n2109 = x47 & ~n1662 ;
  assign n2110 = ~n2108 & ~n2109 ;
  assign n2111 = x431 & n1083 ;
  assign n2112 = x303 & ~n1083 ;
  assign n2113 = ~n2111 & ~n2112 ;
  assign n2114 = ~n2110 & n2113 ;
  assign n2115 = n2110 & ~n2113 ;
  assign n2116 = x430 & n1083 ;
  assign n2117 = x302 & ~n1083 ;
  assign n2118 = ~n2116 & ~n2117 ;
  assign n2119 = x174 & n1662 ;
  assign n2120 = x46 & ~n1662 ;
  assign n2121 = ~n2119 & ~n2120 ;
  assign n2122 = ~n2118 & n2121 ;
  assign n2123 = ~n2115 & ~n2122 ;
  assign n2124 = x172 & n1662 ;
  assign n2125 = x44 & ~n1662 ;
  assign n2126 = ~n2124 & ~n2125 ;
  assign n2127 = x428 & n1083 ;
  assign n2128 = x300 & ~n1083 ;
  assign n2129 = ~n2127 & ~n2128 ;
  assign n2130 = n2126 & ~n2129 ;
  assign n2131 = x173 & n1662 ;
  assign n2132 = x45 & ~n1662 ;
  assign n2133 = ~n2131 & ~n2132 ;
  assign n2134 = x429 & n1083 ;
  assign n2135 = x301 & ~n1083 ;
  assign n2136 = ~n2134 & ~n2135 ;
  assign n2137 = n2133 & ~n2136 ;
  assign n2138 = ~n2130 & ~n2137 ;
  assign n2139 = n2123 & n2138 ;
  assign n2140 = x171 & n1662 ;
  assign n2141 = x43 & ~n1662 ;
  assign n2142 = ~n2140 & ~n2141 ;
  assign n2143 = x427 & n1083 ;
  assign n2144 = x299 & ~n1083 ;
  assign n2145 = ~n2143 & ~n2144 ;
  assign n2146 = ~n2142 & n2145 ;
  assign n2147 = n2142 & ~n2145 ;
  assign n2148 = x170 & n1662 ;
  assign n2149 = x42 & ~n1662 ;
  assign n2150 = ~n2148 & ~n2149 ;
  assign n2151 = x426 & n1083 ;
  assign n2152 = x298 & ~n1083 ;
  assign n2153 = ~n2151 & ~n2152 ;
  assign n2154 = n2150 & ~n2153 ;
  assign n2155 = ~n2147 & ~n2154 ;
  assign n2156 = x169 & n1662 ;
  assign n2157 = x41 & ~n1662 ;
  assign n2158 = ~n2156 & ~n2157 ;
  assign n2159 = x425 & n1083 ;
  assign n2160 = x297 & ~n1083 ;
  assign n2161 = ~n2159 & ~n2160 ;
  assign n2162 = n2158 & ~n2161 ;
  assign n2163 = x168 & n1662 ;
  assign n2164 = x40 & ~n1662 ;
  assign n2165 = ~n2163 & ~n2164 ;
  assign n2166 = x424 & n1083 ;
  assign n2167 = x296 & ~n1083 ;
  assign n2168 = ~n2166 & ~n2167 ;
  assign n2169 = ~n2165 & n2168 ;
  assign n2170 = ~n2162 & n2169 ;
  assign n2171 = ~n2158 & n2161 ;
  assign n2172 = ~n2170 & ~n2171 ;
  assign n2173 = ~n2150 & n2153 ;
  assign n2174 = n2172 & ~n2173 ;
  assign n2175 = n2155 & ~n2174 ;
  assign n2176 = ~n2146 & ~n2175 ;
  assign n2177 = n2139 & ~n2176 ;
  assign n2178 = ~n2126 & n2129 ;
  assign n2179 = ~n2137 & n2178 ;
  assign n2180 = ~n2133 & n2136 ;
  assign n2181 = ~n2179 & ~n2180 ;
  assign n2182 = n2123 & ~n2181 ;
  assign n2183 = n2118 & ~n2121 ;
  assign n2184 = ~n2115 & n2183 ;
  assign n2185 = x416 & n1083 ;
  assign n2186 = x288 & ~n1083 ;
  assign n2187 = ~n2185 & ~n2186 ;
  assign n2188 = x160 & n1662 ;
  assign n2189 = x32 & ~n1662 ;
  assign n2190 = ~n2188 & ~n2189 ;
  assign n2191 = ~n2187 & n2190 ;
  assign n2192 = x159 & n1662 ;
  assign n2193 = x31 & ~n1662 ;
  assign n2194 = ~n2192 & ~n2193 ;
  assign n2195 = x415 & n1083 ;
  assign n2196 = x287 & ~n1083 ;
  assign n2197 = ~n2195 & ~n2196 ;
  assign n2198 = n2194 & ~n2197 ;
  assign n2199 = x158 & n1662 ;
  assign n2200 = x30 & ~n1662 ;
  assign n2201 = ~n2199 & ~n2200 ;
  assign n2202 = x414 & n1083 ;
  assign n2203 = x286 & ~n1083 ;
  assign n2204 = ~n2202 & ~n2203 ;
  assign n2205 = n2201 & ~n2204 ;
  assign n2206 = x157 & n1662 ;
  assign n2207 = x29 & ~n1662 ;
  assign n2208 = ~n2206 & ~n2207 ;
  assign n2209 = x413 & n1083 ;
  assign n2210 = x285 & ~n1083 ;
  assign n2211 = ~n2209 & ~n2210 ;
  assign n2212 = n2208 & ~n2211 ;
  assign n2213 = x156 & n1662 ;
  assign n2214 = x28 & ~n1662 ;
  assign n2215 = ~n2213 & ~n2214 ;
  assign n2216 = x412 & n1083 ;
  assign n2217 = x284 & ~n1083 ;
  assign n2218 = ~n2216 & ~n2217 ;
  assign n2219 = n2215 & ~n2218 ;
  assign n2220 = x155 & n1662 ;
  assign n2221 = x27 & ~n1662 ;
  assign n2222 = ~n2220 & ~n2221 ;
  assign n2223 = x411 & n1083 ;
  assign n2224 = x283 & ~n1083 ;
  assign n2225 = ~n2223 & ~n2224 ;
  assign n2226 = n2222 & ~n2225 ;
  assign n2227 = x154 & n1662 ;
  assign n2228 = x26 & ~n1662 ;
  assign n2229 = ~n2227 & ~n2228 ;
  assign n2230 = x410 & n1083 ;
  assign n2231 = x282 & ~n1083 ;
  assign n2232 = ~n2230 & ~n2231 ;
  assign n2233 = n2229 & ~n2232 ;
  assign n2234 = x409 & n1083 ;
  assign n2235 = x281 & ~n1083 ;
  assign n2236 = ~n2234 & ~n2235 ;
  assign n2237 = x408 & n1083 ;
  assign n2238 = x280 & ~n1083 ;
  assign n2239 = ~n2237 & ~n2238 ;
  assign n2240 = x151 & n1662 ;
  assign n2241 = x23 & ~n1662 ;
  assign n2242 = ~n2240 & ~n2241 ;
  assign n2243 = x407 & n1083 ;
  assign n2244 = x279 & ~n1083 ;
  assign n2245 = ~n2243 & ~n2244 ;
  assign n2246 = n2242 & ~n2245 ;
  assign n2247 = x150 & n1662 ;
  assign n2248 = x22 & ~n1662 ;
  assign n2249 = ~n2247 & ~n2248 ;
  assign n2250 = x406 & n1083 ;
  assign n2251 = x278 & ~n1083 ;
  assign n2252 = ~n2250 & ~n2251 ;
  assign n2253 = n2249 & ~n2252 ;
  assign n2254 = x149 & n1662 ;
  assign n2255 = x21 & ~n1662 ;
  assign n2256 = ~n2254 & ~n2255 ;
  assign n2257 = x405 & n1083 ;
  assign n2258 = x277 & ~n1083 ;
  assign n2259 = ~n2257 & ~n2258 ;
  assign n2260 = n2256 & ~n2259 ;
  assign n2261 = x148 & n1662 ;
  assign n2262 = x20 & ~n1662 ;
  assign n2263 = ~n2261 & ~n2262 ;
  assign n2264 = x404 & n1083 ;
  assign n2265 = x276 & ~n1083 ;
  assign n2266 = ~n2264 & ~n2265 ;
  assign n2267 = n2263 & ~n2266 ;
  assign n2268 = x147 & n1662 ;
  assign n2269 = x19 & ~n1662 ;
  assign n2270 = ~n2268 & ~n2269 ;
  assign n2271 = x403 & n1083 ;
  assign n2272 = x275 & ~n1083 ;
  assign n2273 = ~n2271 & ~n2272 ;
  assign n2274 = n2270 & ~n2273 ;
  assign n2275 = x146 & n1662 ;
  assign n2276 = x18 & ~n1662 ;
  assign n2277 = ~n2275 & ~n2276 ;
  assign n2278 = x402 & n1083 ;
  assign n2279 = x274 & ~n1083 ;
  assign n2280 = ~n2278 & ~n2279 ;
  assign n2281 = n2277 & ~n2280 ;
  assign n2282 = x401 & n1083 ;
  assign n2283 = x273 & ~n1083 ;
  assign n2284 = ~n2282 & ~n2283 ;
  assign n2285 = x400 & n1083 ;
  assign n2286 = x272 & ~n1083 ;
  assign n2287 = ~n2285 & ~n2286 ;
  assign n2288 = x143 & n1662 ;
  assign n2289 = x15 & ~n1662 ;
  assign n2290 = ~n2288 & ~n2289 ;
  assign n2291 = x399 & n1083 ;
  assign n2292 = x271 & ~n1083 ;
  assign n2293 = ~n2291 & ~n2292 ;
  assign n2294 = n2290 & ~n2293 ;
  assign n2295 = x142 & n1662 ;
  assign n2296 = x14 & ~n1662 ;
  assign n2297 = ~n2295 & ~n2296 ;
  assign n2298 = x398 & n1083 ;
  assign n2299 = x270 & ~n1083 ;
  assign n2300 = ~n2298 & ~n2299 ;
  assign n2301 = n2297 & ~n2300 ;
  assign n2302 = x141 & n1662 ;
  assign n2303 = x13 & ~n1662 ;
  assign n2304 = ~n2302 & ~n2303 ;
  assign n2305 = x397 & n1083 ;
  assign n2306 = x269 & ~n1083 ;
  assign n2307 = ~n2305 & ~n2306 ;
  assign n2308 = n2304 & ~n2307 ;
  assign n2309 = x140 & n1662 ;
  assign n2310 = x12 & ~n1662 ;
  assign n2311 = ~n2309 & ~n2310 ;
  assign n2312 = x396 & n1083 ;
  assign n2313 = x268 & ~n1083 ;
  assign n2314 = ~n2312 & ~n2313 ;
  assign n2315 = n2311 & ~n2314 ;
  assign n2316 = x139 & n1662 ;
  assign n2317 = x11 & ~n1662 ;
  assign n2318 = ~n2316 & ~n2317 ;
  assign n2319 = x395 & n1083 ;
  assign n2320 = x267 & ~n1083 ;
  assign n2321 = ~n2319 & ~n2320 ;
  assign n2322 = n2318 & ~n2321 ;
  assign n2323 = x138 & n1662 ;
  assign n2324 = x10 & ~n1662 ;
  assign n2325 = ~n2323 & ~n2324 ;
  assign n2326 = x394 & n1083 ;
  assign n2327 = x266 & ~n1083 ;
  assign n2328 = ~n2326 & ~n2327 ;
  assign n2329 = n2325 & ~n2328 ;
  assign n2330 = x393 & n1083 ;
  assign n2331 = x265 & ~n1083 ;
  assign n2332 = ~n2330 & ~n2331 ;
  assign n2333 = x392 & n1083 ;
  assign n2334 = x264 & ~n1083 ;
  assign n2335 = ~n2333 & ~n2334 ;
  assign n2336 = x135 & n1662 ;
  assign n2337 = x7 & ~n1662 ;
  assign n2338 = ~n2336 & ~n2337 ;
  assign n2339 = x391 & n1083 ;
  assign n2340 = x263 & ~n1083 ;
  assign n2341 = ~n2339 & ~n2340 ;
  assign n2342 = n2338 & ~n2341 ;
  assign n2343 = x390 & n1083 ;
  assign n2344 = x262 & ~n1083 ;
  assign n2345 = ~n2343 & ~n2344 ;
  assign n2346 = x134 & n1662 ;
  assign n2347 = x6 & ~n1662 ;
  assign n2348 = ~n2346 & ~n2347 ;
  assign n2349 = x389 & n1083 ;
  assign n2350 = x261 & ~n1083 ;
  assign n2351 = ~n2349 & ~n2350 ;
  assign n2352 = x133 & n1662 ;
  assign n2353 = x5 & ~n1662 ;
  assign n2354 = ~n2352 & ~n2353 ;
  assign n2355 = x388 & n1083 ;
  assign n2356 = x260 & ~n1083 ;
  assign n2357 = ~n2355 & ~n2356 ;
  assign n2358 = x132 & n1662 ;
  assign n2359 = x4 & ~n1662 ;
  assign n2360 = ~n2358 & ~n2359 ;
  assign n2361 = x131 & n1662 ;
  assign n2362 = x3 & ~n1662 ;
  assign n2363 = ~n2361 & ~n2362 ;
  assign n2364 = x387 & n1083 ;
  assign n2365 = x259 & ~n1083 ;
  assign n2366 = ~n2364 & ~n2365 ;
  assign n2367 = n2363 & ~n2366 ;
  assign n2368 = x385 & n1083 ;
  assign n2369 = x257 & ~n1083 ;
  assign n2370 = ~n2368 & ~n2369 ;
  assign n2371 = x128 & n1662 ;
  assign n2372 = x0 & ~n1662 ;
  assign n2373 = ~n2371 & ~n2372 ;
  assign n2374 = n1086 & ~n2373 ;
  assign n2375 = n2370 & n2374 ;
  assign n2376 = x129 & n1662 ;
  assign n2377 = x1 & ~n1662 ;
  assign n2378 = ~n2376 & ~n2377 ;
  assign n2379 = ~n2375 & n2378 ;
  assign n2380 = x130 & n1662 ;
  assign n2381 = x2 & ~n1662 ;
  assign n2382 = ~n2380 & ~n2381 ;
  assign n2383 = x386 & n1083 ;
  assign n2384 = x258 & ~n1083 ;
  assign n2385 = ~n2383 & ~n2384 ;
  assign n2386 = n2382 & ~n2385 ;
  assign n2387 = ~n2370 & ~n2374 ;
  assign n2388 = ~n2386 & ~n2387 ;
  assign n2389 = ~n2379 & n2388 ;
  assign n2390 = ~n2382 & n2385 ;
  assign n2391 = ~n2389 & ~n2390 ;
  assign n2392 = ~n2367 & ~n2391 ;
  assign n2393 = ~n2363 & n2366 ;
  assign n2394 = ~n2392 & ~n2393 ;
  assign n2395 = n2360 & n2394 ;
  assign n2396 = n2357 & ~n2395 ;
  assign n2397 = ~n2360 & ~n2394 ;
  assign n2398 = ~n2396 & ~n2397 ;
  assign n2399 = n2354 & n2398 ;
  assign n2400 = n2351 & ~n2399 ;
  assign n2401 = ~n2354 & ~n2398 ;
  assign n2402 = ~n2400 & ~n2401 ;
  assign n2403 = n2348 & n2402 ;
  assign n2404 = n2345 & ~n2403 ;
  assign n2405 = ~n2348 & ~n2402 ;
  assign n2406 = ~n2404 & ~n2405 ;
  assign n2407 = ~n2342 & ~n2406 ;
  assign n2408 = ~n2338 & n2341 ;
  assign n2409 = ~n2407 & ~n2408 ;
  assign n2410 = x136 & n1662 ;
  assign n2411 = x8 & ~n1662 ;
  assign n2412 = ~n2410 & ~n2411 ;
  assign n2413 = n2409 & n2412 ;
  assign n2414 = n2335 & ~n2413 ;
  assign n2415 = ~n2409 & ~n2412 ;
  assign n2416 = ~n2414 & ~n2415 ;
  assign n2417 = x137 & n1662 ;
  assign n2418 = x9 & ~n1662 ;
  assign n2419 = ~n2417 & ~n2418 ;
  assign n2420 = n2416 & n2419 ;
  assign n2421 = n2332 & ~n2420 ;
  assign n2422 = ~n2416 & ~n2419 ;
  assign n2423 = ~n2421 & ~n2422 ;
  assign n2424 = ~n2329 & ~n2423 ;
  assign n2425 = ~n2325 & n2328 ;
  assign n2426 = ~n2424 & ~n2425 ;
  assign n2427 = ~n2322 & ~n2426 ;
  assign n2428 = ~n2318 & n2321 ;
  assign n2429 = ~n2427 & ~n2428 ;
  assign n2430 = ~n2315 & ~n2429 ;
  assign n2431 = ~n2311 & n2314 ;
  assign n2432 = ~n2430 & ~n2431 ;
  assign n2433 = ~n2308 & ~n2432 ;
  assign n2434 = ~n2304 & n2307 ;
  assign n2435 = ~n2433 & ~n2434 ;
  assign n2436 = ~n2301 & ~n2435 ;
  assign n2437 = ~n2297 & n2300 ;
  assign n2438 = ~n2436 & ~n2437 ;
  assign n2439 = ~n2294 & ~n2438 ;
  assign n2440 = ~n2290 & n2293 ;
  assign n2441 = ~n2439 & ~n2440 ;
  assign n2442 = x144 & n1662 ;
  assign n2443 = x16 & ~n1662 ;
  assign n2444 = ~n2442 & ~n2443 ;
  assign n2445 = n2441 & n2444 ;
  assign n2446 = n2287 & ~n2445 ;
  assign n2447 = ~n2441 & ~n2444 ;
  assign n2448 = ~n2446 & ~n2447 ;
  assign n2449 = x145 & n1662 ;
  assign n2450 = x17 & ~n1662 ;
  assign n2451 = ~n2449 & ~n2450 ;
  assign n2452 = n2448 & n2451 ;
  assign n2453 = n2284 & ~n2452 ;
  assign n2454 = ~n2448 & ~n2451 ;
  assign n2455 = ~n2453 & ~n2454 ;
  assign n2456 = ~n2281 & ~n2455 ;
  assign n2457 = ~n2277 & n2280 ;
  assign n2458 = ~n2456 & ~n2457 ;
  assign n2459 = ~n2274 & ~n2458 ;
  assign n2460 = ~n2270 & n2273 ;
  assign n2461 = ~n2459 & ~n2460 ;
  assign n2462 = ~n2267 & ~n2461 ;
  assign n2463 = ~n2263 & n2266 ;
  assign n2464 = ~n2462 & ~n2463 ;
  assign n2465 = ~n2260 & ~n2464 ;
  assign n2466 = ~n2256 & n2259 ;
  assign n2467 = ~n2465 & ~n2466 ;
  assign n2468 = ~n2253 & ~n2467 ;
  assign n2469 = ~n2249 & n2252 ;
  assign n2470 = ~n2468 & ~n2469 ;
  assign n2471 = ~n2246 & ~n2470 ;
  assign n2472 = ~n2242 & n2245 ;
  assign n2473 = ~n2471 & ~n2472 ;
  assign n2474 = x152 & n1662 ;
  assign n2475 = x24 & ~n1662 ;
  assign n2476 = ~n2474 & ~n2475 ;
  assign n2477 = n2473 & n2476 ;
  assign n2478 = n2239 & ~n2477 ;
  assign n2479 = ~n2473 & ~n2476 ;
  assign n2480 = ~n2478 & ~n2479 ;
  assign n2481 = x153 & n1662 ;
  assign n2482 = x25 & ~n1662 ;
  assign n2483 = ~n2481 & ~n2482 ;
  assign n2484 = n2480 & n2483 ;
  assign n2485 = n2236 & ~n2484 ;
  assign n2486 = ~n2480 & ~n2483 ;
  assign n2487 = ~n2485 & ~n2486 ;
  assign n2488 = ~n2233 & ~n2487 ;
  assign n2489 = ~n2229 & n2232 ;
  assign n2490 = ~n2488 & ~n2489 ;
  assign n2491 = ~n2226 & ~n2490 ;
  assign n2492 = ~n2222 & n2225 ;
  assign n2493 = ~n2491 & ~n2492 ;
  assign n2494 = ~n2219 & ~n2493 ;
  assign n2495 = ~n2215 & n2218 ;
  assign n2496 = ~n2494 & ~n2495 ;
  assign n2497 = ~n2212 & ~n2496 ;
  assign n2498 = ~n2208 & n2211 ;
  assign n2499 = ~n2497 & ~n2498 ;
  assign n2500 = ~n2205 & ~n2499 ;
  assign n2501 = ~n2201 & n2204 ;
  assign n2502 = ~n2500 & ~n2501 ;
  assign n2503 = ~n2198 & ~n2502 ;
  assign n2504 = ~n2194 & n2197 ;
  assign n2505 = ~n2503 & ~n2504 ;
  assign n2506 = x167 & n1662 ;
  assign n2507 = x39 & ~n1662 ;
  assign n2508 = ~n2506 & ~n2507 ;
  assign n2509 = x423 & n1083 ;
  assign n2510 = x295 & ~n1083 ;
  assign n2511 = ~n2509 & ~n2510 ;
  assign n2512 = n2508 & ~n2511 ;
  assign n2513 = x422 & n1083 ;
  assign n2514 = x294 & ~n1083 ;
  assign n2515 = ~n2513 & ~n2514 ;
  assign n2516 = x166 & n1662 ;
  assign n2517 = x38 & ~n1662 ;
  assign n2518 = ~n2516 & ~n2517 ;
  assign n2519 = ~n2515 & n2518 ;
  assign n2520 = ~n2512 & ~n2519 ;
  assign n2521 = x164 & n1662 ;
  assign n2522 = x36 & ~n1662 ;
  assign n2523 = ~n2521 & ~n2522 ;
  assign n2524 = x420 & n1083 ;
  assign n2525 = x292 & ~n1083 ;
  assign n2526 = ~n2524 & ~n2525 ;
  assign n2527 = n2523 & ~n2526 ;
  assign n2528 = x165 & n1662 ;
  assign n2529 = x37 & ~n1662 ;
  assign n2530 = ~n2528 & ~n2529 ;
  assign n2531 = x421 & n1083 ;
  assign n2532 = x293 & ~n1083 ;
  assign n2533 = ~n2531 & ~n2532 ;
  assign n2534 = n2530 & ~n2533 ;
  assign n2535 = ~n2527 & ~n2534 ;
  assign n2536 = n2520 & n2535 ;
  assign n2537 = x161 & n1662 ;
  assign n2538 = x33 & ~n1662 ;
  assign n2539 = ~n2537 & ~n2538 ;
  assign n2540 = x417 & n1083 ;
  assign n2541 = x289 & ~n1083 ;
  assign n2542 = ~n2540 & ~n2541 ;
  assign n2543 = n2539 & ~n2542 ;
  assign n2544 = x163 & n1662 ;
  assign n2545 = x35 & ~n1662 ;
  assign n2546 = ~n2544 & ~n2545 ;
  assign n2547 = x419 & n1083 ;
  assign n2548 = x291 & ~n1083 ;
  assign n2549 = ~n2547 & ~n2548 ;
  assign n2550 = n2546 & ~n2549 ;
  assign n2551 = x418 & n1083 ;
  assign n2552 = x290 & ~n1083 ;
  assign n2553 = ~n2551 & ~n2552 ;
  assign n2554 = x162 & n1662 ;
  assign n2555 = x34 & ~n1662 ;
  assign n2556 = ~n2554 & ~n2555 ;
  assign n2557 = ~n2553 & n2556 ;
  assign n2558 = ~n2550 & ~n2557 ;
  assign n2559 = ~n2543 & n2558 ;
  assign n2560 = n2536 & n2559 ;
  assign n2561 = ~n2505 & n2560 ;
  assign n2562 = ~n2191 & n2561 ;
  assign n2563 = ~n2508 & n2511 ;
  assign n2564 = ~n2523 & n2526 ;
  assign n2565 = ~n2534 & n2564 ;
  assign n2566 = ~n2530 & n2533 ;
  assign n2567 = ~n2565 & ~n2566 ;
  assign n2568 = n2520 & ~n2567 ;
  assign n2569 = ~n2512 & n2515 ;
  assign n2570 = ~n2518 & n2569 ;
  assign n2571 = ~n2546 & n2549 ;
  assign n2572 = ~n2550 & n2553 ;
  assign n2573 = ~n2556 & n2572 ;
  assign n2574 = n2187 & ~n2190 ;
  assign n2575 = ~n2539 & n2542 ;
  assign n2576 = ~n2574 & ~n2575 ;
  assign n2577 = n2559 & ~n2576 ;
  assign n2578 = ~n2573 & ~n2577 ;
  assign n2579 = ~n2571 & n2578 ;
  assign n2580 = n2536 & ~n2579 ;
  assign n2581 = ~n2570 & ~n2580 ;
  assign n2582 = ~n2568 & n2581 ;
  assign n2583 = ~n2563 & n2582 ;
  assign n2584 = ~n2562 & n2583 ;
  assign n2585 = n2165 & ~n2168 ;
  assign n2586 = ~n2162 & ~n2585 ;
  assign n2587 = n2155 & n2586 ;
  assign n2588 = n2139 & n2587 ;
  assign n2589 = ~n2584 & n2588 ;
  assign n2590 = ~n2184 & ~n2589 ;
  assign n2591 = ~n2182 & n2590 ;
  assign n2592 = ~n2177 & n2591 ;
  assign n2593 = ~n2114 & n2592 ;
  assign n2594 = x432 & n1083 ;
  assign n2595 = x304 & ~n1083 ;
  assign n2596 = ~n2594 & ~n2595 ;
  assign n2597 = x176 & n1662 ;
  assign n2598 = x48 & ~n1662 ;
  assign n2599 = ~n2597 & ~n2598 ;
  assign n2600 = ~n2596 & n2599 ;
  assign n2601 = x183 & n1662 ;
  assign n2602 = x55 & ~n1662 ;
  assign n2603 = ~n2601 & ~n2602 ;
  assign n2604 = x439 & n1083 ;
  assign n2605 = x311 & ~n1083 ;
  assign n2606 = ~n2604 & ~n2605 ;
  assign n2607 = n2603 & ~n2606 ;
  assign n2608 = x438 & n1083 ;
  assign n2609 = x310 & ~n1083 ;
  assign n2610 = ~n2608 & ~n2609 ;
  assign n2611 = x182 & n1662 ;
  assign n2612 = x54 & ~n1662 ;
  assign n2613 = ~n2611 & ~n2612 ;
  assign n2614 = ~n2610 & n2613 ;
  assign n2615 = ~n2607 & ~n2614 ;
  assign n2616 = x181 & n1662 ;
  assign n2617 = x53 & ~n1662 ;
  assign n2618 = ~n2616 & ~n2617 ;
  assign n2619 = x437 & n1083 ;
  assign n2620 = x309 & ~n1083 ;
  assign n2621 = ~n2619 & ~n2620 ;
  assign n2622 = n2618 & ~n2621 ;
  assign n2623 = x436 & n1083 ;
  assign n2624 = x308 & ~n1083 ;
  assign n2625 = ~n2623 & ~n2624 ;
  assign n2626 = x180 & n1662 ;
  assign n2627 = x52 & ~n1662 ;
  assign n2628 = ~n2626 & ~n2627 ;
  assign n2629 = ~n2625 & n2628 ;
  assign n2630 = ~n2622 & ~n2629 ;
  assign n2631 = n2615 & n2630 ;
  assign n2632 = x177 & n1662 ;
  assign n2633 = x49 & ~n1662 ;
  assign n2634 = ~n2632 & ~n2633 ;
  assign n2635 = x433 & n1083 ;
  assign n2636 = x305 & ~n1083 ;
  assign n2637 = ~n2635 & ~n2636 ;
  assign n2638 = n2634 & ~n2637 ;
  assign n2639 = x179 & n1662 ;
  assign n2640 = x51 & ~n1662 ;
  assign n2641 = ~n2639 & ~n2640 ;
  assign n2642 = x435 & n1083 ;
  assign n2643 = x307 & ~n1083 ;
  assign n2644 = ~n2642 & ~n2643 ;
  assign n2645 = n2641 & ~n2644 ;
  assign n2646 = x434 & n1083 ;
  assign n2647 = x306 & ~n1083 ;
  assign n2648 = ~n2646 & ~n2647 ;
  assign n2649 = x178 & n1662 ;
  assign n2650 = x50 & ~n1662 ;
  assign n2651 = ~n2649 & ~n2650 ;
  assign n2652 = ~n2648 & n2651 ;
  assign n2653 = ~n2645 & ~n2652 ;
  assign n2654 = ~n2638 & n2653 ;
  assign n2655 = n2631 & n2654 ;
  assign n2656 = ~n2600 & n2655 ;
  assign n2657 = ~n2593 & n2656 ;
  assign n2658 = ~n2603 & n2606 ;
  assign n2659 = ~n2641 & n2644 ;
  assign n2660 = ~n2645 & n2648 ;
  assign n2661 = ~n2651 & n2660 ;
  assign n2662 = n2596 & ~n2599 ;
  assign n2663 = ~n2634 & n2637 ;
  assign n2664 = ~n2662 & ~n2663 ;
  assign n2665 = n2654 & ~n2664 ;
  assign n2666 = ~n2661 & ~n2665 ;
  assign n2667 = ~n2659 & n2666 ;
  assign n2668 = n2631 & ~n2667 ;
  assign n2669 = n2625 & ~n2628 ;
  assign n2670 = ~n2622 & n2669 ;
  assign n2671 = ~n2618 & n2621 ;
  assign n2672 = ~n2670 & ~n2671 ;
  assign n2673 = n2610 & ~n2613 ;
  assign n2674 = n2672 & ~n2673 ;
  assign n2675 = n2615 & ~n2674 ;
  assign n2676 = ~n2668 & ~n2675 ;
  assign n2677 = ~n2658 & n2676 ;
  assign n2678 = ~n2657 & n2677 ;
  assign n2679 = n2088 & ~n2091 ;
  assign n2680 = ~n2085 & ~n2679 ;
  assign n2681 = n2062 & n2680 ;
  assign n2682 = n2078 & n2681 ;
  assign n2683 = ~n2678 & n2682 ;
  assign n2684 = ~n2107 & ~n2683 ;
  assign n2685 = ~n2105 & n2684 ;
  assign n2686 = ~n2100 & n2685 ;
  assign n2687 = ~n2037 & n2686 ;
  assign n2688 = ~n2030 & ~n2687 ;
  assign n2689 = ~n2023 & n2688 ;
  assign n2690 = n2016 & n2689 ;
  assign n2691 = ~n2004 & n2007 ;
  assign n2692 = n2019 & ~n2030 ;
  assign n2693 = ~n2022 & n2692 ;
  assign n2694 = ~n2026 & n2029 ;
  assign n2695 = ~n2693 & ~n2694 ;
  assign n2696 = n2011 & ~n2014 ;
  assign n2697 = n2695 & ~n2696 ;
  assign n2698 = n2016 & ~n2697 ;
  assign n2699 = ~n2691 & ~n2698 ;
  assign n2700 = ~n2690 & n2699 ;
  assign n2701 = n1991 & ~n1994 ;
  assign n2702 = ~n1988 & ~n2701 ;
  assign n2703 = n1981 & n2702 ;
  assign n2704 = ~n2700 & n2703 ;
  assign n2705 = ~n2001 & ~n2704 ;
  assign n2706 = ~n1999 & n2705 ;
  assign n2707 = ~n1972 & n2706 ;
  assign n2708 = x203 & n1662 ;
  assign n2709 = x75 & ~n1662 ;
  assign n2710 = ~n2708 & ~n2709 ;
  assign n2711 = x459 & n1083 ;
  assign n2712 = x331 & ~n1083 ;
  assign n2713 = ~n2711 & ~n2712 ;
  assign n2714 = n2710 & ~n2713 ;
  assign n2715 = x458 & n1083 ;
  assign n2716 = x330 & ~n1083 ;
  assign n2717 = ~n2715 & ~n2716 ;
  assign n2718 = x202 & n1662 ;
  assign n2719 = x74 & ~n1662 ;
  assign n2720 = ~n2718 & ~n2719 ;
  assign n2721 = ~n2717 & n2720 ;
  assign n2722 = ~n2714 & ~n2721 ;
  assign n2723 = x201 & n1662 ;
  assign n2724 = x73 & ~n1662 ;
  assign n2725 = ~n2723 & ~n2724 ;
  assign n2726 = x457 & n1083 ;
  assign n2727 = x329 & ~n1083 ;
  assign n2728 = ~n2726 & ~n2727 ;
  assign n2729 = n2725 & ~n2728 ;
  assign n2730 = x456 & n1083 ;
  assign n2731 = x328 & ~n1083 ;
  assign n2732 = ~n2730 & ~n2731 ;
  assign n2733 = x200 & n1662 ;
  assign n2734 = x72 & ~n1662 ;
  assign n2735 = ~n2733 & ~n2734 ;
  assign n2736 = ~n2732 & n2735 ;
  assign n2737 = ~n2729 & ~n2736 ;
  assign n2738 = n2722 & n2737 ;
  assign n2739 = ~n2707 & n2738 ;
  assign n2740 = ~n2710 & n2713 ;
  assign n2741 = n2732 & ~n2735 ;
  assign n2742 = ~n2729 & n2741 ;
  assign n2743 = ~n2725 & n2728 ;
  assign n2744 = ~n2742 & ~n2743 ;
  assign n2745 = n2717 & ~n2720 ;
  assign n2746 = n2744 & ~n2745 ;
  assign n2747 = n2722 & ~n2746 ;
  assign n2748 = ~n2740 & ~n2747 ;
  assign n2749 = ~n2739 & n2748 ;
  assign n2750 = n1955 & ~n1958 ;
  assign n2751 = ~n1952 & ~n2750 ;
  assign n2752 = n1945 & n2751 ;
  assign n2753 = ~n2749 & n2752 ;
  assign n2754 = ~n1965 & ~n2753 ;
  assign n2755 = ~n1963 & n2754 ;
  assign n2756 = ~n1936 & n2755 ;
  assign n2757 = ~n1929 & ~n2756 ;
  assign n2758 = n1922 & n2757 ;
  assign n2759 = ~n1907 & n2758 ;
  assign n2760 = ~n1910 & n1913 ;
  assign n2761 = n1903 & ~n1929 ;
  assign n2762 = ~n1906 & n2761 ;
  assign n2763 = ~n1925 & n1928 ;
  assign n2764 = ~n2762 & ~n2763 ;
  assign n2765 = n1917 & ~n1920 ;
  assign n2766 = n2764 & ~n2765 ;
  assign n2767 = n1922 & ~n2766 ;
  assign n2768 = ~n2760 & ~n2767 ;
  assign n2769 = ~n2759 & n2768 ;
  assign n2770 = n1890 & ~n1893 ;
  assign n2771 = ~n1887 & ~n2770 ;
  assign n2772 = n1880 & n2771 ;
  assign n2773 = ~n2769 & n2772 ;
  assign n2774 = ~n1900 & ~n2773 ;
  assign n2775 = ~n1898 & n2774 ;
  assign n2776 = ~n1871 & n2775 ;
  assign n2777 = x219 & n1662 ;
  assign n2778 = x91 & ~n1662 ;
  assign n2779 = ~n2777 & ~n2778 ;
  assign n2780 = x475 & n1083 ;
  assign n2781 = x347 & ~n1083 ;
  assign n2782 = ~n2780 & ~n2781 ;
  assign n2783 = n2779 & ~n2782 ;
  assign n2784 = x474 & n1083 ;
  assign n2785 = x346 & ~n1083 ;
  assign n2786 = ~n2784 & ~n2785 ;
  assign n2787 = x218 & n1662 ;
  assign n2788 = x90 & ~n1662 ;
  assign n2789 = ~n2787 & ~n2788 ;
  assign n2790 = ~n2786 & n2789 ;
  assign n2791 = ~n2783 & ~n2790 ;
  assign n2792 = x217 & n1662 ;
  assign n2793 = x89 & ~n1662 ;
  assign n2794 = ~n2792 & ~n2793 ;
  assign n2795 = x473 & n1083 ;
  assign n2796 = x345 & ~n1083 ;
  assign n2797 = ~n2795 & ~n2796 ;
  assign n2798 = n2794 & ~n2797 ;
  assign n2799 = x472 & n1083 ;
  assign n2800 = x344 & ~n1083 ;
  assign n2801 = ~n2799 & ~n2800 ;
  assign n2802 = x216 & n1662 ;
  assign n2803 = x88 & ~n1662 ;
  assign n2804 = ~n2802 & ~n2803 ;
  assign n2805 = ~n2801 & n2804 ;
  assign n2806 = ~n2798 & ~n2805 ;
  assign n2807 = n2791 & n2806 ;
  assign n2808 = ~n2776 & n2807 ;
  assign n2809 = ~n2779 & n2782 ;
  assign n2810 = n2801 & ~n2804 ;
  assign n2811 = ~n2798 & n2810 ;
  assign n2812 = ~n2794 & n2797 ;
  assign n2813 = ~n2811 & ~n2812 ;
  assign n2814 = n2786 & ~n2789 ;
  assign n2815 = n2813 & ~n2814 ;
  assign n2816 = n2791 & ~n2815 ;
  assign n2817 = ~n2809 & ~n2816 ;
  assign n2818 = ~n2808 & n2817 ;
  assign n2819 = n1854 & ~n1857 ;
  assign n2820 = ~n1851 & ~n2819 ;
  assign n2821 = n1844 & n2820 ;
  assign n2822 = ~n2818 & n2821 ;
  assign n2823 = ~n1864 & ~n2822 ;
  assign n2824 = ~n1862 & n2823 ;
  assign n2825 = ~n1835 & n2824 ;
  assign n2826 = ~n1828 & ~n2825 ;
  assign n2827 = n1821 & n2826 ;
  assign n2828 = ~n1806 & n2827 ;
  assign n2829 = ~n1809 & n1812 ;
  assign n2830 = n1802 & ~n1828 ;
  assign n2831 = ~n1805 & n2830 ;
  assign n2832 = ~n1824 & n1827 ;
  assign n2833 = ~n2831 & ~n2832 ;
  assign n2834 = n1816 & ~n1819 ;
  assign n2835 = n2833 & ~n2834 ;
  assign n2836 = n1821 & ~n2835 ;
  assign n2837 = ~n2829 & ~n2836 ;
  assign n2838 = ~n2828 & n2837 ;
  assign n2839 = n1789 & ~n1792 ;
  assign n2840 = ~n1786 & ~n2839 ;
  assign n2841 = n1779 & n2840 ;
  assign n2842 = ~n2838 & n2841 ;
  assign n2843 = ~n1799 & ~n2842 ;
  assign n2844 = ~n1797 & n2843 ;
  assign n2845 = ~n1770 & n2844 ;
  assign n2846 = x235 & n1662 ;
  assign n2847 = x107 & ~n1662 ;
  assign n2848 = ~n2846 & ~n2847 ;
  assign n2849 = x491 & n1083 ;
  assign n2850 = x363 & ~n1083 ;
  assign n2851 = ~n2849 & ~n2850 ;
  assign n2852 = n2848 & ~n2851 ;
  assign n2853 = x490 & n1083 ;
  assign n2854 = x362 & ~n1083 ;
  assign n2855 = ~n2853 & ~n2854 ;
  assign n2856 = x234 & n1662 ;
  assign n2857 = x106 & ~n1662 ;
  assign n2858 = ~n2856 & ~n2857 ;
  assign n2859 = ~n2855 & n2858 ;
  assign n2860 = ~n2852 & ~n2859 ;
  assign n2861 = x233 & n1662 ;
  assign n2862 = x105 & ~n1662 ;
  assign n2863 = ~n2861 & ~n2862 ;
  assign n2864 = x489 & n1083 ;
  assign n2865 = x361 & ~n1083 ;
  assign n2866 = ~n2864 & ~n2865 ;
  assign n2867 = n2863 & ~n2866 ;
  assign n2868 = x488 & n1083 ;
  assign n2869 = x360 & ~n1083 ;
  assign n2870 = ~n2868 & ~n2869 ;
  assign n2871 = x232 & n1662 ;
  assign n2872 = x104 & ~n1662 ;
  assign n2873 = ~n2871 & ~n2872 ;
  assign n2874 = ~n2870 & n2873 ;
  assign n2875 = ~n2867 & ~n2874 ;
  assign n2876 = n2860 & n2875 ;
  assign n2877 = ~n2845 & n2876 ;
  assign n2878 = ~n2848 & n2851 ;
  assign n2879 = n2870 & ~n2873 ;
  assign n2880 = ~n2867 & n2879 ;
  assign n2881 = ~n2863 & n2866 ;
  assign n2882 = ~n2880 & ~n2881 ;
  assign n2883 = n2855 & ~n2858 ;
  assign n2884 = n2882 & ~n2883 ;
  assign n2885 = n2860 & ~n2884 ;
  assign n2886 = ~n2878 & ~n2885 ;
  assign n2887 = ~n2877 & n2886 ;
  assign n2888 = n1753 & ~n1756 ;
  assign n2889 = ~n1750 & ~n2888 ;
  assign n2890 = n1743 & n2889 ;
  assign n2891 = ~n2887 & n2890 ;
  assign n2892 = ~n1763 & ~n2891 ;
  assign n2893 = ~n1761 & n2892 ;
  assign n2894 = ~n1734 & n2893 ;
  assign n2895 = ~n1727 & ~n2894 ;
  assign n2896 = n1720 & n2895 ;
  assign n2897 = ~n1705 & n2896 ;
  assign n2898 = ~n1708 & n1711 ;
  assign n2899 = n1701 & ~n1727 ;
  assign n2900 = ~n1704 & n2899 ;
  assign n2901 = ~n1723 & n1726 ;
  assign n2902 = ~n2900 & ~n2901 ;
  assign n2903 = n1715 & ~n1718 ;
  assign n2904 = n2902 & ~n2903 ;
  assign n2905 = n1720 & ~n2904 ;
  assign n2906 = ~n2898 & ~n2905 ;
  assign n2907 = ~n2897 & n2906 ;
  assign n2908 = n1681 & ~n1691 ;
  assign n2909 = ~n1688 & ~n2908 ;
  assign n2910 = n1678 & n2909 ;
  assign n2911 = ~n2907 & n2910 ;
  assign n2912 = ~n1698 & ~n2911 ;
  assign n2913 = ~n1696 & n2912 ;
  assign n2914 = ~n1669 & n2913 ;
  assign n2915 = x251 & n1662 ;
  assign n2916 = x123 & ~n1662 ;
  assign n2917 = ~n2915 & ~n2916 ;
  assign n2918 = x507 & n1083 ;
  assign n2919 = x379 & ~n1083 ;
  assign n2920 = ~n2918 & ~n2919 ;
  assign n2921 = n2917 & ~n2920 ;
  assign n2922 = x506 & n1083 ;
  assign n2923 = x378 & ~n1083 ;
  assign n2924 = ~n2922 & ~n2923 ;
  assign n2925 = x250 & n1662 ;
  assign n2926 = x122 & ~n1662 ;
  assign n2927 = ~n2925 & ~n2926 ;
  assign n2928 = ~n2924 & n2927 ;
  assign n2929 = ~n2921 & ~n2928 ;
  assign n2930 = x249 & n1662 ;
  assign n2931 = x121 & ~n1662 ;
  assign n2932 = ~n2930 & ~n2931 ;
  assign n2933 = x505 & n1083 ;
  assign n2934 = x377 & ~n1083 ;
  assign n2935 = ~n2933 & ~n2934 ;
  assign n2936 = n2932 & ~n2935 ;
  assign n2937 = x504 & n1083 ;
  assign n2938 = x376 & ~n1083 ;
  assign n2939 = ~n2937 & ~n2938 ;
  assign n2940 = x248 & n1662 ;
  assign n2941 = x120 & ~n1662 ;
  assign n2942 = ~n2940 & ~n2941 ;
  assign n2943 = ~n2939 & n2942 ;
  assign n2944 = ~n2936 & ~n2943 ;
  assign n2945 = n2929 & n2944 ;
  assign n2946 = ~n2914 & n2945 ;
  assign n2947 = ~n2917 & n2920 ;
  assign n2948 = ~n2936 & n2939 ;
  assign n2949 = ~n2942 & n2948 ;
  assign n2950 = ~n2932 & n2935 ;
  assign n2951 = ~n2949 & ~n2950 ;
  assign n2952 = n2924 & ~n2927 ;
  assign n2953 = n2951 & ~n2952 ;
  assign n2954 = n2929 & ~n2953 ;
  assign n2955 = ~n2947 & ~n2954 ;
  assign n2956 = ~n2946 & n2955 ;
  assign n2957 = x252 & n1662 ;
  assign n2958 = x124 & ~n1662 ;
  assign n2959 = ~n2957 & ~n2958 ;
  assign n2960 = x508 & n1083 ;
  assign n2961 = x380 & ~n1083 ;
  assign n2962 = ~n2960 & ~n2961 ;
  assign n2963 = n2959 & ~n2962 ;
  assign n2964 = ~n1088 & n1659 ;
  assign n2965 = x254 & n1662 ;
  assign n2966 = x126 & ~n1662 ;
  assign n2967 = ~n2965 & ~n2966 ;
  assign n2968 = x510 & n1083 ;
  assign n2969 = x382 & ~n1083 ;
  assign n2970 = ~n2968 & ~n2969 ;
  assign n2971 = n2967 & ~n2970 ;
  assign n2972 = x253 & n1662 ;
  assign n2973 = x125 & ~n1662 ;
  assign n2974 = ~n2972 & ~n2973 ;
  assign n2975 = x509 & n1083 ;
  assign n2976 = x381 & ~n1083 ;
  assign n2977 = ~n2975 & ~n2976 ;
  assign n2978 = n2974 & ~n2977 ;
  assign n2979 = ~n2971 & ~n2978 ;
  assign n2980 = ~n2964 & n2979 ;
  assign n2981 = ~n2963 & n2980 ;
  assign n2982 = ~n2956 & n2981 ;
  assign n2983 = ~n2959 & n2962 ;
  assign n2984 = ~n2974 & n2977 ;
  assign n2985 = ~n2983 & ~n2984 ;
  assign n2986 = n2979 & ~n2985 ;
  assign n2987 = ~n2967 & n2970 ;
  assign n2988 = ~n2986 & ~n2987 ;
  assign n2989 = ~n2964 & ~n2988 ;
  assign n2990 = ~n2982 & ~n2989 ;
  assign n2991 = ~n1660 & n2990 ;
  assign n2992 = ~n1086 & n2991 ;
  assign n2993 = ~n2373 & ~n2991 ;
  assign n2994 = ~n2992 & ~n2993 ;
  assign n5064 = ~n2994 & x512 ;
  assign n2995 = x374 & ~x502 ;
  assign n2996 = ~n513 & ~n2995 ;
  assign n2997 = ~n520 & n1041 ;
  assign n2998 = ~n517 & ~n2997 ;
  assign n2999 = n2996 & ~n2998 ;
  assign n3000 = x502 & ~n513 ;
  assign n3001 = ~x374 & n3000 ;
  assign n3002 = x368 & ~x496 ;
  assign n3003 = ~n1031 & ~n1036 ;
  assign n3004 = x366 & ~x494 ;
  assign n3005 = ~n530 & ~n3004 ;
  assign n3006 = ~n537 & n1021 ;
  assign n3007 = ~n534 & ~n3006 ;
  assign n3008 = n3005 & ~n3007 ;
  assign n3009 = x494 & ~n530 ;
  assign n3010 = ~x366 & n3009 ;
  assign n3011 = x358 & ~x486 ;
  assign n3012 = ~n542 & ~n3011 ;
  assign n3013 = ~n549 & n996 ;
  assign n3014 = ~n546 & ~n3013 ;
  assign n3015 = n3012 & ~n3014 ;
  assign n3016 = x486 & ~n542 ;
  assign n3017 = ~x358 & n3016 ;
  assign n3018 = x352 & ~x480 ;
  assign n3019 = ~n986 & ~n991 ;
  assign n3020 = x350 & ~x478 ;
  assign n3021 = ~n559 & ~n3020 ;
  assign n3022 = ~n566 & n976 ;
  assign n3023 = ~n563 & ~n3022 ;
  assign n3024 = n3021 & ~n3023 ;
  assign n3025 = x478 & ~n559 ;
  assign n3026 = ~x350 & n3025 ;
  assign n3027 = x342 & ~x470 ;
  assign n3028 = ~n571 & ~n3027 ;
  assign n3029 = ~n578 & n951 ;
  assign n3030 = ~n575 & ~n3029 ;
  assign n3031 = n3028 & ~n3030 ;
  assign n3032 = x470 & ~n571 ;
  assign n3033 = ~x342 & n3032 ;
  assign n3034 = x336 & ~x464 ;
  assign n3035 = ~n941 & ~n946 ;
  assign n3036 = x334 & ~x462 ;
  assign n3037 = ~n588 & ~n3036 ;
  assign n3038 = ~n595 & n931 ;
  assign n3039 = ~n592 & ~n3038 ;
  assign n3040 = n3037 & ~n3039 ;
  assign n3041 = x462 & ~n588 ;
  assign n3042 = ~x334 & n3041 ;
  assign n3043 = x326 & ~x454 ;
  assign n3044 = ~n600 & ~n3043 ;
  assign n3045 = ~n607 & n906 ;
  assign n3046 = ~n604 & ~n3045 ;
  assign n3047 = n3044 & ~n3046 ;
  assign n3048 = x454 & ~n600 ;
  assign n3049 = ~x326 & n3048 ;
  assign n3050 = ~n896 & ~n901 ;
  assign n3051 = x318 & ~x446 ;
  assign n3052 = ~n616 & ~n3051 ;
  assign n3053 = ~n638 & ~n640 ;
  assign n3054 = n3052 & n3053 ;
  assign n3055 = ~n624 & ~n633 ;
  assign n3056 = ~n631 & n883 ;
  assign n3057 = ~n628 & ~n3056 ;
  assign n3058 = ~n626 & n3057 ;
  assign n3059 = n3055 & ~n3058 ;
  assign n3060 = ~n625 & ~n3059 ;
  assign n3061 = n3054 & ~n3060 ;
  assign n3062 = n620 & ~n640 ;
  assign n3063 = ~n621 & ~n3062 ;
  assign n3064 = n3052 & ~n3063 ;
  assign n3065 = x446 & ~n616 ;
  assign n3066 = ~x318 & n3065 ;
  assign n3067 = x302 & ~x430 ;
  assign n3068 = ~n645 & ~n3067 ;
  assign n3069 = ~n667 & ~n669 ;
  assign n3070 = n3068 & n3069 ;
  assign n3071 = ~n653 & ~n662 ;
  assign n3072 = ~n660 & n837 ;
  assign n3073 = ~n657 & ~n3072 ;
  assign n3074 = ~n655 & n3073 ;
  assign n3075 = n3071 & ~n3074 ;
  assign n3076 = ~n654 & ~n3075 ;
  assign n3077 = n3070 & ~n3076 ;
  assign n3078 = n649 & ~n669 ;
  assign n3079 = ~n650 & ~n3078 ;
  assign n3080 = n3068 & ~n3079 ;
  assign n3081 = x430 & ~n645 ;
  assign n3082 = ~x302 & n3081 ;
  assign n3083 = x288 & ~x416 ;
  assign n3084 = ~x256 & x384 ;
  assign n3085 = ~x257 & n3084 ;
  assign n3086 = ~x385 & ~n3085 ;
  assign n3087 = x257 & ~n3084 ;
  assign n3088 = ~n703 & ~n3087 ;
  assign n3089 = ~n3086 & n3088 ;
  assign n3090 = ~n699 & ~n3089 ;
  assign n3091 = ~n706 & ~n3090 ;
  assign n3092 = ~n695 & ~n3091 ;
  assign n3093 = x260 & n3092 ;
  assign n3094 = x388 & ~n3093 ;
  assign n3095 = ~x260 & ~n3092 ;
  assign n3096 = ~n3094 & ~n3095 ;
  assign n3097 = x261 & n3096 ;
  assign n3098 = x389 & ~n3097 ;
  assign n3099 = ~x261 & ~n3096 ;
  assign n3100 = ~n3098 & ~n3099 ;
  assign n3101 = ~n717 & ~n3100 ;
  assign n3102 = ~n694 & ~n3101 ;
  assign n3103 = ~n720 & ~n3102 ;
  assign n3104 = ~n693 & ~n3103 ;
  assign n3105 = x264 & n3104 ;
  assign n3106 = x392 & ~n3105 ;
  assign n3107 = ~x264 & ~n3104 ;
  assign n3108 = ~n3106 & ~n3107 ;
  assign n3109 = x265 & n3108 ;
  assign n3110 = x393 & ~n3109 ;
  assign n3111 = ~x265 & ~n3108 ;
  assign n3112 = ~n3110 & ~n3111 ;
  assign n3113 = ~n731 & ~n3112 ;
  assign n3114 = ~n692 & ~n3113 ;
  assign n3115 = ~n734 & ~n3114 ;
  assign n3116 = ~n691 & ~n3115 ;
  assign n3117 = ~n737 & ~n3116 ;
  assign n3118 = ~n690 & ~n3117 ;
  assign n3119 = ~n740 & ~n3118 ;
  assign n3120 = ~n689 & ~n3119 ;
  assign n3121 = ~n743 & ~n3120 ;
  assign n3122 = ~n688 & ~n3121 ;
  assign n3123 = ~n746 & ~n3122 ;
  assign n3124 = ~n687 & ~n3123 ;
  assign n3125 = x272 & n3124 ;
  assign n3126 = x400 & ~n3125 ;
  assign n3127 = ~x272 & ~n3124 ;
  assign n3128 = ~n3126 & ~n3127 ;
  assign n3129 = x273 & n3128 ;
  assign n3130 = x401 & ~n3129 ;
  assign n3131 = ~x273 & ~n3128 ;
  assign n3132 = ~n3130 & ~n3131 ;
  assign n3133 = ~n757 & ~n3132 ;
  assign n3134 = ~n686 & ~n3133 ;
  assign n3135 = ~n760 & ~n3134 ;
  assign n3136 = ~n685 & ~n3135 ;
  assign n3137 = ~n763 & ~n3136 ;
  assign n3138 = ~n684 & ~n3137 ;
  assign n3139 = ~n766 & ~n3138 ;
  assign n3140 = ~n683 & ~n3139 ;
  assign n3141 = ~n769 & ~n3140 ;
  assign n3142 = ~n682 & ~n3141 ;
  assign n3143 = ~n772 & ~n3142 ;
  assign n3144 = ~n681 & ~n3143 ;
  assign n3145 = x280 & n3144 ;
  assign n3146 = x408 & ~n3145 ;
  assign n3147 = ~x280 & ~n3144 ;
  assign n3148 = ~n3146 & ~n3147 ;
  assign n3149 = x281 & n3148 ;
  assign n3150 = x409 & ~n3149 ;
  assign n3151 = ~x281 & ~n3148 ;
  assign n3152 = ~n3150 & ~n3151 ;
  assign n3153 = ~n783 & ~n3152 ;
  assign n3154 = ~n680 & ~n3153 ;
  assign n3155 = ~n786 & ~n3154 ;
  assign n3156 = ~n679 & ~n3155 ;
  assign n3157 = ~n789 & ~n3156 ;
  assign n3158 = ~n678 & ~n3157 ;
  assign n3159 = ~n792 & ~n3158 ;
  assign n3160 = ~n677 & ~n3159 ;
  assign n3161 = ~n795 & ~n3160 ;
  assign n3162 = ~n676 & ~n3161 ;
  assign n3163 = ~n798 & ~n3162 ;
  assign n3164 = ~n675 & ~n3163 ;
  assign n3165 = x294 & ~x422 ;
  assign n3166 = ~n815 & ~n3165 ;
  assign n3167 = ~n816 & ~n818 ;
  assign n3168 = n3166 & n3167 ;
  assign n3169 = ~n823 & ~n828 ;
  assign n3170 = ~n826 & n3169 ;
  assign n3171 = n3168 & n3170 ;
  assign n3172 = ~n3164 & n3171 ;
  assign n3173 = ~n3083 & n3172 ;
  assign n3174 = n803 & ~n818 ;
  assign n3175 = ~n804 & ~n3174 ;
  assign n3176 = n3166 & ~n3175 ;
  assign n3177 = x422 & ~n815 ;
  assign n3178 = ~x294 & n3177 ;
  assign n3179 = x416 & ~n826 ;
  assign n3180 = ~x288 & n3179 ;
  assign n3181 = ~n807 & ~n3180 ;
  assign n3182 = ~n809 & n3181 ;
  assign n3183 = n3169 & ~n3182 ;
  assign n3184 = ~n808 & ~n3183 ;
  assign n3185 = n3168 & ~n3184 ;
  assign n3186 = ~n3178 & ~n3185 ;
  assign n3187 = ~n3176 & n3186 ;
  assign n3188 = ~n800 & n3187 ;
  assign n3189 = ~n3173 & n3188 ;
  assign n3190 = ~n658 & ~n660 ;
  assign n3191 = n3071 & n3190 ;
  assign n3192 = n3070 & n3191 ;
  assign n3193 = ~n3189 & n3192 ;
  assign n3194 = ~n3082 & ~n3193 ;
  assign n3195 = ~n3080 & n3194 ;
  assign n3196 = ~n3077 & n3195 ;
  assign n3197 = ~n646 & n3196 ;
  assign n3198 = x304 & ~x432 ;
  assign n3199 = ~n862 & ~n877 ;
  assign n3200 = ~n873 & ~n875 ;
  assign n3201 = n3199 & n3200 ;
  assign n3202 = ~n863 & ~n868 ;
  assign n3203 = ~n866 & n3202 ;
  assign n3204 = n3201 & n3203 ;
  assign n3205 = ~n3198 & n3204 ;
  assign n3206 = ~n3197 & n3205 ;
  assign n3207 = x432 & ~n866 ;
  assign n3208 = ~x304 & n3207 ;
  assign n3209 = ~n854 & ~n3208 ;
  assign n3210 = ~n856 & n3209 ;
  assign n3211 = n3202 & ~n3210 ;
  assign n3212 = ~n855 & ~n3211 ;
  assign n3213 = n3201 & ~n3212 ;
  assign n3214 = n851 & ~n875 ;
  assign n3215 = ~n850 & ~n3214 ;
  assign n3216 = ~n848 & n3215 ;
  assign n3217 = n3199 & ~n3216 ;
  assign n3218 = ~n3213 & ~n3217 ;
  assign n3219 = ~n847 & n3218 ;
  assign n3220 = ~n3206 & n3219 ;
  assign n3221 = ~n629 & ~n631 ;
  assign n3222 = n3054 & n3221 ;
  assign n3223 = n3055 & n3222 ;
  assign n3224 = ~n3220 & n3223 ;
  assign n3225 = ~n3066 & ~n3224 ;
  assign n3226 = ~n3064 & n3225 ;
  assign n3227 = ~n3061 & n3226 ;
  assign n3228 = ~n617 & n3227 ;
  assign n3229 = ~n897 & ~n3228 ;
  assign n3230 = ~n899 & n3229 ;
  assign n3231 = n3050 & n3230 ;
  assign n3232 = n892 & ~n899 ;
  assign n3233 = ~n615 & ~n3232 ;
  assign n3234 = ~n613 & n3233 ;
  assign n3235 = n3050 & ~n3234 ;
  assign n3236 = ~n612 & ~n3235 ;
  assign n3237 = ~n3231 & n3236 ;
  assign n3238 = ~n605 & ~n607 ;
  assign n3239 = n3044 & n3238 ;
  assign n3240 = ~n3237 & n3239 ;
  assign n3241 = ~n3049 & ~n3240 ;
  assign n3242 = ~n3047 & n3241 ;
  assign n3243 = ~n601 & n3242 ;
  assign n3244 = ~n921 & ~n926 ;
  assign n3245 = ~n922 & ~n924 ;
  assign n3246 = n3244 & n3245 ;
  assign n3247 = ~n3243 & n3246 ;
  assign n3248 = n917 & ~n924 ;
  assign n3249 = ~n916 & ~n3248 ;
  assign n3250 = ~n914 & n3249 ;
  assign n3251 = n3244 & ~n3250 ;
  assign n3252 = ~n913 & ~n3251 ;
  assign n3253 = ~n3247 & n3252 ;
  assign n3254 = ~n593 & ~n595 ;
  assign n3255 = n3037 & n3254 ;
  assign n3256 = ~n3253 & n3255 ;
  assign n3257 = ~n3042 & ~n3256 ;
  assign n3258 = ~n3040 & n3257 ;
  assign n3259 = ~n589 & n3258 ;
  assign n3260 = ~n944 & ~n3259 ;
  assign n3261 = n3035 & n3260 ;
  assign n3262 = ~n3034 & n3261 ;
  assign n3263 = x464 & ~n944 ;
  assign n3264 = ~x336 & n3263 ;
  assign n3265 = ~n587 & ~n3264 ;
  assign n3266 = ~n585 & n3265 ;
  assign n3267 = n3035 & ~n3266 ;
  assign n3268 = ~n584 & ~n3267 ;
  assign n3269 = ~n3262 & n3268 ;
  assign n3270 = ~n576 & ~n578 ;
  assign n3271 = n3028 & n3270 ;
  assign n3272 = ~n3269 & n3271 ;
  assign n3273 = ~n3033 & ~n3272 ;
  assign n3274 = ~n3031 & n3273 ;
  assign n3275 = ~n572 & n3274 ;
  assign n3276 = ~n966 & ~n971 ;
  assign n3277 = ~n967 & ~n969 ;
  assign n3278 = n3276 & n3277 ;
  assign n3279 = ~n3275 & n3278 ;
  assign n3280 = n962 & ~n969 ;
  assign n3281 = ~n961 & ~n3280 ;
  assign n3282 = ~n959 & n3281 ;
  assign n3283 = n3276 & ~n3282 ;
  assign n3284 = ~n958 & ~n3283 ;
  assign n3285 = ~n3279 & n3284 ;
  assign n3286 = ~n564 & ~n566 ;
  assign n3287 = n3021 & n3286 ;
  assign n3288 = ~n3285 & n3287 ;
  assign n3289 = ~n3026 & ~n3288 ;
  assign n3290 = ~n3024 & n3289 ;
  assign n3291 = ~n560 & n3290 ;
  assign n3292 = ~n989 & ~n3291 ;
  assign n3293 = n3019 & n3292 ;
  assign n3294 = ~n3018 & n3293 ;
  assign n3295 = x480 & ~n989 ;
  assign n3296 = ~x352 & n3295 ;
  assign n3297 = ~n558 & ~n3296 ;
  assign n3298 = ~n556 & n3297 ;
  assign n3299 = n3019 & ~n3298 ;
  assign n3300 = ~n555 & ~n3299 ;
  assign n3301 = ~n3294 & n3300 ;
  assign n3302 = ~n547 & ~n549 ;
  assign n3303 = n3012 & n3302 ;
  assign n3304 = ~n3301 & n3303 ;
  assign n3305 = ~n3017 & ~n3304 ;
  assign n3306 = ~n3015 & n3305 ;
  assign n3307 = ~n543 & n3306 ;
  assign n3308 = ~n1011 & ~n1016 ;
  assign n3309 = ~n1012 & ~n1014 ;
  assign n3310 = n3308 & n3309 ;
  assign n3311 = ~n3307 & n3310 ;
  assign n3312 = n1007 & ~n1014 ;
  assign n3313 = ~n1006 & ~n3312 ;
  assign n3314 = ~n1004 & n3313 ;
  assign n3315 = n3308 & ~n3314 ;
  assign n3316 = ~n1003 & ~n3315 ;
  assign n3317 = ~n3311 & n3316 ;
  assign n3318 = ~n535 & ~n537 ;
  assign n3319 = n3005 & n3318 ;
  assign n3320 = ~n3317 & n3319 ;
  assign n3321 = ~n3010 & ~n3320 ;
  assign n3322 = ~n3008 & n3321 ;
  assign n3323 = ~n531 & n3322 ;
  assign n3324 = ~n1034 & ~n3323 ;
  assign n3325 = n3003 & n3324 ;
  assign n3326 = ~n3002 & n3325 ;
  assign n3327 = x496 & ~n1034 ;
  assign n3328 = ~x368 & n3327 ;
  assign n3329 = ~n529 & ~n3328 ;
  assign n3330 = ~n527 & n3329 ;
  assign n3331 = n3003 & ~n3330 ;
  assign n3332 = ~n526 & ~n3331 ;
  assign n3333 = ~n3326 & n3332 ;
  assign n3334 = ~n518 & ~n520 ;
  assign n3335 = n2996 & n3334 ;
  assign n3336 = ~n3333 & n3335 ;
  assign n3337 = ~n3001 & ~n3336 ;
  assign n3338 = ~n2999 & n3337 ;
  assign n3339 = ~n514 & n3338 ;
  assign n3340 = ~n1056 & ~n1061 ;
  assign n3341 = ~n1057 & ~n1059 ;
  assign n3342 = n3340 & n3341 ;
  assign n3343 = ~n3339 & n3342 ;
  assign n3344 = n1052 & ~n1059 ;
  assign n3345 = ~n1051 & ~n3344 ;
  assign n3346 = ~n1049 & n3345 ;
  assign n3347 = n3340 & ~n3346 ;
  assign n3348 = ~n1048 & ~n3347 ;
  assign n3349 = ~n3343 & n3348 ;
  assign n3350 = ~n1075 & ~n1078 ;
  assign n3351 = ~n1082 & n3350 ;
  assign n3352 = ~n1074 & n3351 ;
  assign n3353 = ~n3349 & n3352 ;
  assign n3354 = ~n1066 & ~n1069 ;
  assign n3355 = n3350 & ~n3354 ;
  assign n3356 = ~n1068 & ~n3355 ;
  assign n3357 = ~n1082 & ~n3356 ;
  assign n3358 = ~n3353 & ~n3357 ;
  assign n3359 = ~n1067 & n3358 ;
  assign n3360 = ~x384 & n3359 ;
  assign n3361 = ~x256 & ~n3359 ;
  assign n3362 = ~n3360 & ~n3361 ;
  assign n3363 = x511 & n3358 ;
  assign n3364 = ~x383 & ~n3363 ;
  assign n3365 = x118 & ~x246 ;
  assign n3366 = ~n1089 & ~n3365 ;
  assign n3367 = ~n1096 & n1617 ;
  assign n3368 = ~n1093 & ~n3367 ;
  assign n3369 = n3366 & ~n3368 ;
  assign n3370 = x246 & ~n1089 ;
  assign n3371 = ~x118 & n3370 ;
  assign n3372 = x112 & ~x240 ;
  assign n3373 = ~n1607 & ~n1612 ;
  assign n3374 = x110 & ~x238 ;
  assign n3375 = ~n1106 & ~n3374 ;
  assign n3376 = ~n1113 & n1597 ;
  assign n3377 = ~n1110 & ~n3376 ;
  assign n3378 = n3375 & ~n3377 ;
  assign n3379 = x238 & ~n1106 ;
  assign n3380 = ~x110 & n3379 ;
  assign n3381 = x102 & ~x230 ;
  assign n3382 = ~n1118 & ~n3381 ;
  assign n3383 = ~n1125 & n1572 ;
  assign n3384 = ~n1122 & ~n3383 ;
  assign n3385 = n3382 & ~n3384 ;
  assign n3386 = x230 & ~n1118 ;
  assign n3387 = ~x102 & n3386 ;
  assign n3388 = x96 & ~x224 ;
  assign n3389 = ~n1562 & ~n1567 ;
  assign n3390 = x94 & ~x222 ;
  assign n3391 = ~n1135 & ~n3390 ;
  assign n3392 = ~n1142 & n1552 ;
  assign n3393 = ~n1139 & ~n3392 ;
  assign n3394 = n3391 & ~n3393 ;
  assign n3395 = x222 & ~n1135 ;
  assign n3396 = ~x94 & n3395 ;
  assign n3397 = x86 & ~x214 ;
  assign n3398 = ~n1147 & ~n3397 ;
  assign n3399 = ~n1154 & n1527 ;
  assign n3400 = ~n1151 & ~n3399 ;
  assign n3401 = n3398 & ~n3400 ;
  assign n3402 = x214 & ~n1147 ;
  assign n3403 = ~x86 & n3402 ;
  assign n3404 = x80 & ~x208 ;
  assign n3405 = ~n1517 & ~n1522 ;
  assign n3406 = x78 & ~x206 ;
  assign n3407 = ~n1164 & ~n3406 ;
  assign n3408 = ~n1171 & n1507 ;
  assign n3409 = ~n1168 & ~n3408 ;
  assign n3410 = n3407 & ~n3409 ;
  assign n3411 = x206 & ~n1164 ;
  assign n3412 = ~x78 & n3411 ;
  assign n3413 = x70 & ~x198 ;
  assign n3414 = ~n1176 & ~n3413 ;
  assign n3415 = ~n1183 & n1482 ;
  assign n3416 = ~n1180 & ~n3415 ;
  assign n3417 = n3414 & ~n3416 ;
  assign n3418 = x198 & ~n1176 ;
  assign n3419 = ~x70 & n3418 ;
  assign n3420 = ~n1472 & ~n1477 ;
  assign n3421 = x62 & ~x190 ;
  assign n3422 = ~n1192 & ~n3421 ;
  assign n3423 = ~n1214 & ~n1216 ;
  assign n3424 = n3422 & n3423 ;
  assign n3425 = ~n1200 & ~n1209 ;
  assign n3426 = ~n1207 & n1459 ;
  assign n3427 = ~n1204 & ~n3426 ;
  assign n3428 = ~n1202 & n3427 ;
  assign n3429 = n3425 & ~n3428 ;
  assign n3430 = ~n1201 & ~n3429 ;
  assign n3431 = n3424 & ~n3430 ;
  assign n3432 = n1196 & ~n1216 ;
  assign n3433 = ~n1197 & ~n3432 ;
  assign n3434 = n3422 & ~n3433 ;
  assign n3435 = x190 & ~n1192 ;
  assign n3436 = ~x62 & n3435 ;
  assign n3437 = x46 & ~x174 ;
  assign n3438 = ~n1221 & ~n3437 ;
  assign n3439 = ~n1243 & ~n1245 ;
  assign n3440 = n3438 & n3439 ;
  assign n3441 = ~n1229 & ~n1238 ;
  assign n3442 = ~n1236 & n1413 ;
  assign n3443 = ~n1233 & ~n3442 ;
  assign n3444 = ~n1231 & n3443 ;
  assign n3445 = n3441 & ~n3444 ;
  assign n3446 = ~n1230 & ~n3445 ;
  assign n3447 = n3440 & ~n3446 ;
  assign n3448 = n1225 & ~n1245 ;
  assign n3449 = ~n1226 & ~n3448 ;
  assign n3450 = n3438 & ~n3449 ;
  assign n3451 = x174 & ~n1221 ;
  assign n3452 = ~x46 & n3451 ;
  assign n3453 = x32 & ~x160 ;
  assign n3454 = ~x0 & x128 ;
  assign n3455 = ~n1276 & ~n3454 ;
  assign n3456 = ~n1273 & ~n1279 ;
  assign n3457 = ~n3455 & n3456 ;
  assign n3458 = ~n1275 & ~n3457 ;
  assign n3459 = ~n1282 & ~n3458 ;
  assign n3460 = ~n1271 & ~n3459 ;
  assign n3461 = x4 & n3460 ;
  assign n3462 = x132 & ~n3461 ;
  assign n3463 = ~x4 & ~n3460 ;
  assign n3464 = ~n3462 & ~n3463 ;
  assign n3465 = x5 & n3464 ;
  assign n3466 = x133 & ~n3465 ;
  assign n3467 = ~x5 & ~n3464 ;
  assign n3468 = ~n3466 & ~n3467 ;
  assign n3469 = ~n1293 & ~n3468 ;
  assign n3470 = ~n1270 & ~n3469 ;
  assign n3471 = ~n1296 & ~n3470 ;
  assign n3472 = ~n1269 & ~n3471 ;
  assign n3473 = x8 & n3472 ;
  assign n3474 = x136 & ~n3473 ;
  assign n3475 = ~x8 & ~n3472 ;
  assign n3476 = ~n3474 & ~n3475 ;
  assign n3477 = x9 & n3476 ;
  assign n3478 = x137 & ~n3477 ;
  assign n3479 = ~x9 & ~n3476 ;
  assign n3480 = ~n3478 & ~n3479 ;
  assign n3481 = ~n1307 & ~n3480 ;
  assign n3482 = ~n1268 & ~n3481 ;
  assign n3483 = ~n1310 & ~n3482 ;
  assign n3484 = ~n1267 & ~n3483 ;
  assign n3485 = ~n1313 & ~n3484 ;
  assign n3486 = ~n1266 & ~n3485 ;
  assign n3487 = ~n1316 & ~n3486 ;
  assign n3488 = ~n1265 & ~n3487 ;
  assign n3489 = ~n1319 & ~n3488 ;
  assign n3490 = ~n1264 & ~n3489 ;
  assign n3491 = ~n1322 & ~n3490 ;
  assign n3492 = ~n1263 & ~n3491 ;
  assign n3493 = x16 & n3492 ;
  assign n3494 = x144 & ~n3493 ;
  assign n3495 = ~x16 & ~n3492 ;
  assign n3496 = ~n3494 & ~n3495 ;
  assign n3497 = x17 & n3496 ;
  assign n3498 = x145 & ~n3497 ;
  assign n3499 = ~x17 & ~n3496 ;
  assign n3500 = ~n3498 & ~n3499 ;
  assign n3501 = ~n1333 & ~n3500 ;
  assign n3502 = ~n1262 & ~n3501 ;
  assign n3503 = ~n1336 & ~n3502 ;
  assign n3504 = ~n1261 & ~n3503 ;
  assign n3505 = ~n1339 & ~n3504 ;
  assign n3506 = ~n1260 & ~n3505 ;
  assign n3507 = ~n1342 & ~n3506 ;
  assign n3508 = ~n1259 & ~n3507 ;
  assign n3509 = ~n1345 & ~n3508 ;
  assign n3510 = ~n1258 & ~n3509 ;
  assign n3511 = ~n1348 & ~n3510 ;
  assign n3512 = ~n1257 & ~n3511 ;
  assign n3513 = x24 & n3512 ;
  assign n3514 = x152 & ~n3513 ;
  assign n3515 = ~x24 & ~n3512 ;
  assign n3516 = ~n3514 & ~n3515 ;
  assign n3517 = x25 & n3516 ;
  assign n3518 = x153 & ~n3517 ;
  assign n3519 = ~x25 & ~n3516 ;
  assign n3520 = ~n3518 & ~n3519 ;
  assign n3521 = ~n1359 & ~n3520 ;
  assign n3522 = ~n1256 & ~n3521 ;
  assign n3523 = ~n1362 & ~n3522 ;
  assign n3524 = ~n1255 & ~n3523 ;
  assign n3525 = ~n1365 & ~n3524 ;
  assign n3526 = ~n1254 & ~n3525 ;
  assign n3527 = ~n1368 & ~n3526 ;
  assign n3528 = ~n1253 & ~n3527 ;
  assign n3529 = ~n1371 & ~n3528 ;
  assign n3530 = ~n1252 & ~n3529 ;
  assign n3531 = ~n1374 & ~n3530 ;
  assign n3532 = ~n1251 & ~n3531 ;
  assign n3533 = x38 & ~x166 ;
  assign n3534 = ~n1391 & ~n3533 ;
  assign n3535 = ~n1392 & ~n1394 ;
  assign n3536 = n3534 & n3535 ;
  assign n3537 = ~n1399 & ~n1404 ;
  assign n3538 = ~n1402 & n3537 ;
  assign n3539 = n3536 & n3538 ;
  assign n3540 = ~n3532 & n3539 ;
  assign n3541 = ~n3453 & n3540 ;
  assign n3542 = n1379 & ~n1394 ;
  assign n3543 = ~n1380 & ~n3542 ;
  assign n3544 = n3534 & ~n3543 ;
  assign n3545 = x166 & ~n1391 ;
  assign n3546 = ~x38 & n3545 ;
  assign n3547 = x160 & ~n1402 ;
  assign n3548 = ~x32 & n3547 ;
  assign n3549 = ~n1383 & ~n3548 ;
  assign n3550 = ~n1385 & n3549 ;
  assign n3551 = n3537 & ~n3550 ;
  assign n3552 = ~n1384 & ~n3551 ;
  assign n3553 = n3536 & ~n3552 ;
  assign n3554 = ~n3546 & ~n3553 ;
  assign n3555 = ~n3544 & n3554 ;
  assign n3556 = ~n1376 & n3555 ;
  assign n3557 = ~n3541 & n3556 ;
  assign n3558 = ~n1234 & ~n1236 ;
  assign n3559 = n3441 & n3558 ;
  assign n3560 = n3440 & n3559 ;
  assign n3561 = ~n3557 & n3560 ;
  assign n3562 = ~n3452 & ~n3561 ;
  assign n3563 = ~n3450 & n3562 ;
  assign n3564 = ~n3447 & n3563 ;
  assign n3565 = ~n1222 & n3564 ;
  assign n3566 = x48 & ~x176 ;
  assign n3567 = ~n1438 & ~n1453 ;
  assign n3568 = ~n1449 & ~n1451 ;
  assign n3569 = n3567 & n3568 ;
  assign n3570 = ~n1439 & ~n1444 ;
  assign n3571 = ~n1442 & n3570 ;
  assign n3572 = n3569 & n3571 ;
  assign n3573 = ~n3566 & n3572 ;
  assign n3574 = ~n3565 & n3573 ;
  assign n3575 = x176 & ~n1442 ;
  assign n3576 = ~x48 & n3575 ;
  assign n3577 = ~n1430 & ~n3576 ;
  assign n3578 = ~n1432 & n3577 ;
  assign n3579 = n3570 & ~n3578 ;
  assign n3580 = ~n1431 & ~n3579 ;
  assign n3581 = n3569 & ~n3580 ;
  assign n3582 = n1427 & ~n1451 ;
  assign n3583 = ~n1426 & ~n3582 ;
  assign n3584 = ~n1424 & n3583 ;
  assign n3585 = n3567 & ~n3584 ;
  assign n3586 = ~n3581 & ~n3585 ;
  assign n3587 = ~n1423 & n3586 ;
  assign n3588 = ~n3574 & n3587 ;
  assign n3589 = ~n1205 & ~n1207 ;
  assign n3590 = n3424 & n3589 ;
  assign n3591 = n3425 & n3590 ;
  assign n3592 = ~n3588 & n3591 ;
  assign n3593 = ~n3436 & ~n3592 ;
  assign n3594 = ~n3434 & n3593 ;
  assign n3595 = ~n3431 & n3594 ;
  assign n3596 = ~n1193 & n3595 ;
  assign n3597 = ~n1473 & ~n3596 ;
  assign n3598 = ~n1475 & n3597 ;
  assign n3599 = n3420 & n3598 ;
  assign n3600 = n1468 & ~n1475 ;
  assign n3601 = ~n1191 & ~n3600 ;
  assign n3602 = ~n1189 & n3601 ;
  assign n3603 = n3420 & ~n3602 ;
  assign n3604 = ~n1188 & ~n3603 ;
  assign n3605 = ~n3599 & n3604 ;
  assign n3606 = ~n1181 & ~n1183 ;
  assign n3607 = n3414 & n3606 ;
  assign n3608 = ~n3605 & n3607 ;
  assign n3609 = ~n3419 & ~n3608 ;
  assign n3610 = ~n3417 & n3609 ;
  assign n3611 = ~n1177 & n3610 ;
  assign n3612 = ~n1497 & ~n1502 ;
  assign n3613 = ~n1498 & ~n1500 ;
  assign n3614 = n3612 & n3613 ;
  assign n3615 = ~n3611 & n3614 ;
  assign n3616 = n1493 & ~n1500 ;
  assign n3617 = ~n1492 & ~n3616 ;
  assign n3618 = ~n1490 & n3617 ;
  assign n3619 = n3612 & ~n3618 ;
  assign n3620 = ~n1489 & ~n3619 ;
  assign n3621 = ~n3615 & n3620 ;
  assign n3622 = ~n1169 & ~n1171 ;
  assign n3623 = n3407 & n3622 ;
  assign n3624 = ~n3621 & n3623 ;
  assign n3625 = ~n3412 & ~n3624 ;
  assign n3626 = ~n3410 & n3625 ;
  assign n3627 = ~n1165 & n3626 ;
  assign n3628 = ~n1520 & ~n3627 ;
  assign n3629 = n3405 & n3628 ;
  assign n3630 = ~n3404 & n3629 ;
  assign n3631 = x208 & ~n1520 ;
  assign n3632 = ~x80 & n3631 ;
  assign n3633 = ~n1163 & ~n3632 ;
  assign n3634 = ~n1161 & n3633 ;
  assign n3635 = n3405 & ~n3634 ;
  assign n3636 = ~n1160 & ~n3635 ;
  assign n3637 = ~n3630 & n3636 ;
  assign n3638 = ~n1152 & ~n1154 ;
  assign n3639 = n3398 & n3638 ;
  assign n3640 = ~n3637 & n3639 ;
  assign n3641 = ~n3403 & ~n3640 ;
  assign n3642 = ~n3401 & n3641 ;
  assign n3643 = ~n1148 & n3642 ;
  assign n3644 = ~n1542 & ~n1547 ;
  assign n3645 = ~n1543 & ~n1545 ;
  assign n3646 = n3644 & n3645 ;
  assign n3647 = ~n3643 & n3646 ;
  assign n3648 = n1538 & ~n1545 ;
  assign n3649 = ~n1537 & ~n3648 ;
  assign n3650 = ~n1535 & n3649 ;
  assign n3651 = n3644 & ~n3650 ;
  assign n3652 = ~n1534 & ~n3651 ;
  assign n3653 = ~n3647 & n3652 ;
  assign n3654 = ~n1140 & ~n1142 ;
  assign n3655 = n3391 & n3654 ;
  assign n3656 = ~n3653 & n3655 ;
  assign n3657 = ~n3396 & ~n3656 ;
  assign n3658 = ~n3394 & n3657 ;
  assign n3659 = ~n1136 & n3658 ;
  assign n3660 = ~n1565 & ~n3659 ;
  assign n3661 = n3389 & n3660 ;
  assign n3662 = ~n3388 & n3661 ;
  assign n3663 = x224 & ~n1565 ;
  assign n3664 = ~x96 & n3663 ;
  assign n3665 = ~n1134 & ~n3664 ;
  assign n3666 = ~n1132 & n3665 ;
  assign n3667 = n3389 & ~n3666 ;
  assign n3668 = ~n1131 & ~n3667 ;
  assign n3669 = ~n3662 & n3668 ;
  assign n3670 = ~n1123 & ~n1125 ;
  assign n3671 = n3382 & n3670 ;
  assign n3672 = ~n3669 & n3671 ;
  assign n3673 = ~n3387 & ~n3672 ;
  assign n3674 = ~n3385 & n3673 ;
  assign n3675 = ~n1119 & n3674 ;
  assign n3676 = ~n1587 & ~n1592 ;
  assign n3677 = ~n1588 & ~n1590 ;
  assign n3678 = n3676 & n3677 ;
  assign n3679 = ~n3675 & n3678 ;
  assign n3680 = n1583 & ~n1590 ;
  assign n3681 = ~n1582 & ~n3680 ;
  assign n3682 = ~n1580 & n3681 ;
  assign n3683 = n3676 & ~n3682 ;
  assign n3684 = ~n1579 & ~n3683 ;
  assign n3685 = ~n3679 & n3684 ;
  assign n3686 = ~n1111 & ~n1113 ;
  assign n3687 = n3375 & n3686 ;
  assign n3688 = ~n3685 & n3687 ;
  assign n3689 = ~n3380 & ~n3688 ;
  assign n3690 = ~n3378 & n3689 ;
  assign n3691 = ~n1107 & n3690 ;
  assign n3692 = ~n1610 & ~n3691 ;
  assign n3693 = n3373 & n3692 ;
  assign n3694 = ~n3372 & n3693 ;
  assign n3695 = x240 & ~n1610 ;
  assign n3696 = ~x112 & n3695 ;
  assign n3697 = ~n1105 & ~n3696 ;
  assign n3698 = ~n1103 & n3697 ;
  assign n3699 = n3373 & ~n3698 ;
  assign n3700 = ~n1102 & ~n3699 ;
  assign n3701 = ~n3694 & n3700 ;
  assign n3702 = ~n1094 & ~n1096 ;
  assign n3703 = n3366 & n3702 ;
  assign n3704 = ~n3701 & n3703 ;
  assign n3705 = ~n3371 & ~n3704 ;
  assign n3706 = ~n3369 & n3705 ;
  assign n3707 = ~n1090 & n3706 ;
  assign n3708 = ~n1632 & ~n1637 ;
  assign n3709 = ~n1633 & ~n1635 ;
  assign n3710 = n3708 & n3709 ;
  assign n3711 = ~n3707 & n3710 ;
  assign n3712 = n1628 & ~n1635 ;
  assign n3713 = ~n1627 & ~n3712 ;
  assign n3714 = ~n1625 & n3713 ;
  assign n3715 = n3708 & ~n3714 ;
  assign n3716 = ~n1624 & ~n3715 ;
  assign n3717 = ~n3711 & n3716 ;
  assign n3718 = ~n1651 & ~n1654 ;
  assign n3719 = ~n1661 & n3718 ;
  assign n3720 = ~n1650 & n3719 ;
  assign n3721 = ~n3717 & n3720 ;
  assign n3722 = ~n1642 & ~n1645 ;
  assign n3723 = n3718 & ~n3722 ;
  assign n3724 = ~n1644 & ~n3723 ;
  assign n3725 = ~n1661 & ~n3724 ;
  assign n3726 = ~n3721 & ~n3725 ;
  assign n3727 = x255 & n3726 ;
  assign n3728 = ~x127 & ~n3727 ;
  assign n3729 = n3364 & ~n3728 ;
  assign n3730 = ~n1643 & n3726 ;
  assign n3731 = ~x247 & n3730 ;
  assign n3732 = ~x119 & ~n3730 ;
  assign n3733 = ~n3731 & ~n3732 ;
  assign n3734 = ~x503 & n3359 ;
  assign n3735 = ~x375 & ~n3359 ;
  assign n3736 = ~n3734 & ~n3735 ;
  assign n3737 = ~n3733 & n3736 ;
  assign n3738 = n3733 & ~n3736 ;
  assign n3739 = ~x502 & n3359 ;
  assign n3740 = ~x374 & ~n3359 ;
  assign n3741 = ~n3739 & ~n3740 ;
  assign n3742 = ~x246 & n3730 ;
  assign n3743 = ~x118 & ~n3730 ;
  assign n3744 = ~n3742 & ~n3743 ;
  assign n3745 = ~n3741 & n3744 ;
  assign n3746 = ~n3738 & ~n3745 ;
  assign n3747 = ~x244 & n3730 ;
  assign n3748 = ~x116 & ~n3730 ;
  assign n3749 = ~n3747 & ~n3748 ;
  assign n3750 = ~x245 & n3730 ;
  assign n3751 = ~x117 & ~n3730 ;
  assign n3752 = ~n3750 & ~n3751 ;
  assign n3753 = ~x501 & n3359 ;
  assign n3754 = ~x373 & ~n3359 ;
  assign n3755 = ~n3753 & ~n3754 ;
  assign n3756 = n3752 & ~n3755 ;
  assign n3757 = ~x500 & n3359 ;
  assign n3758 = ~x372 & ~n3359 ;
  assign n3759 = ~n3757 & ~n3758 ;
  assign n3760 = ~n3756 & n3759 ;
  assign n3761 = ~n3749 & n3760 ;
  assign n3762 = ~n3752 & n3755 ;
  assign n3763 = ~n3761 & ~n3762 ;
  assign n3764 = n3746 & ~n3763 ;
  assign n3765 = n3741 & ~n3744 ;
  assign n3766 = ~n3738 & n3765 ;
  assign n3767 = ~x496 & n3359 ;
  assign n3768 = ~x368 & ~n3359 ;
  assign n3769 = ~n3767 & ~n3768 ;
  assign n3770 = ~x240 & n3730 ;
  assign n3771 = ~x112 & ~n3730 ;
  assign n3772 = ~n3770 & ~n3771 ;
  assign n3773 = ~n3769 & n3772 ;
  assign n3774 = ~x243 & n3730 ;
  assign n3775 = ~x115 & ~n3730 ;
  assign n3776 = ~n3774 & ~n3775 ;
  assign n3777 = ~x499 & n3359 ;
  assign n3778 = ~x371 & ~n3359 ;
  assign n3779 = ~n3777 & ~n3778 ;
  assign n3780 = n3776 & ~n3779 ;
  assign n3781 = ~x498 & n3359 ;
  assign n3782 = ~x370 & ~n3359 ;
  assign n3783 = ~n3781 & ~n3782 ;
  assign n3784 = ~x242 & n3730 ;
  assign n3785 = ~x114 & ~n3730 ;
  assign n3786 = ~n3784 & ~n3785 ;
  assign n3787 = ~n3783 & n3786 ;
  assign n3788 = ~n3780 & ~n3787 ;
  assign n3789 = ~x241 & n3730 ;
  assign n3790 = ~x113 & ~n3730 ;
  assign n3791 = ~n3789 & ~n3790 ;
  assign n3792 = ~x497 & n3359 ;
  assign n3793 = ~x369 & ~n3359 ;
  assign n3794 = ~n3792 & ~n3793 ;
  assign n3795 = n3791 & ~n3794 ;
  assign n3796 = ~x239 & n3730 ;
  assign n3797 = ~x111 & ~n3730 ;
  assign n3798 = ~n3796 & ~n3797 ;
  assign n3799 = ~x495 & n3359 ;
  assign n3800 = ~x367 & ~n3359 ;
  assign n3801 = ~n3799 & ~n3800 ;
  assign n3802 = ~n3798 & n3801 ;
  assign n3803 = n3798 & ~n3801 ;
  assign n3804 = ~x494 & n3359 ;
  assign n3805 = ~x366 & ~n3359 ;
  assign n3806 = ~n3804 & ~n3805 ;
  assign n3807 = ~x238 & n3730 ;
  assign n3808 = ~x110 & ~n3730 ;
  assign n3809 = ~n3807 & ~n3808 ;
  assign n3810 = ~n3806 & n3809 ;
  assign n3811 = ~n3803 & ~n3810 ;
  assign n3812 = ~x237 & n3730 ;
  assign n3813 = ~x109 & ~n3730 ;
  assign n3814 = ~n3812 & ~n3813 ;
  assign n3815 = ~x493 & n3359 ;
  assign n3816 = ~x365 & ~n3359 ;
  assign n3817 = ~n3815 & ~n3816 ;
  assign n3818 = n3814 & ~n3817 ;
  assign n3819 = ~x236 & n3730 ;
  assign n3820 = ~x108 & ~n3730 ;
  assign n3821 = ~n3819 & ~n3820 ;
  assign n3822 = ~x492 & n3359 ;
  assign n3823 = ~x364 & ~n3359 ;
  assign n3824 = ~n3822 & ~n3823 ;
  assign n3825 = ~n3821 & n3824 ;
  assign n3826 = ~n3818 & n3825 ;
  assign n3827 = ~n3814 & n3817 ;
  assign n3828 = ~n3826 & ~n3827 ;
  assign n3829 = n3811 & ~n3828 ;
  assign n3830 = n3806 & ~n3809 ;
  assign n3831 = ~n3803 & n3830 ;
  assign n3832 = ~x231 & n3730 ;
  assign n3833 = ~x103 & ~n3730 ;
  assign n3834 = ~n3832 & ~n3833 ;
  assign n3835 = ~x487 & n3359 ;
  assign n3836 = ~x359 & ~n3359 ;
  assign n3837 = ~n3835 & ~n3836 ;
  assign n3838 = ~n3834 & n3837 ;
  assign n3839 = n3834 & ~n3837 ;
  assign n3840 = ~x486 & n3359 ;
  assign n3841 = ~x358 & ~n3359 ;
  assign n3842 = ~n3840 & ~n3841 ;
  assign n3843 = ~x230 & n3730 ;
  assign n3844 = ~x102 & ~n3730 ;
  assign n3845 = ~n3843 & ~n3844 ;
  assign n3846 = ~n3842 & n3845 ;
  assign n3847 = ~n3839 & ~n3846 ;
  assign n3848 = ~x229 & n3730 ;
  assign n3849 = ~x101 & ~n3730 ;
  assign n3850 = ~n3848 & ~n3849 ;
  assign n3851 = ~x485 & n3359 ;
  assign n3852 = ~x357 & ~n3359 ;
  assign n3853 = ~n3851 & ~n3852 ;
  assign n3854 = n3850 & ~n3853 ;
  assign n3855 = ~x228 & n3730 ;
  assign n3856 = ~x100 & ~n3730 ;
  assign n3857 = ~n3855 & ~n3856 ;
  assign n3858 = ~x484 & n3359 ;
  assign n3859 = ~x356 & ~n3359 ;
  assign n3860 = ~n3858 & ~n3859 ;
  assign n3861 = ~n3857 & n3860 ;
  assign n3862 = ~n3854 & n3861 ;
  assign n3863 = ~n3850 & n3853 ;
  assign n3864 = ~n3862 & ~n3863 ;
  assign n3865 = n3847 & ~n3864 ;
  assign n3866 = n3842 & ~n3845 ;
  assign n3867 = ~n3839 & n3866 ;
  assign n3868 = ~x480 & n3359 ;
  assign n3869 = ~x352 & ~n3359 ;
  assign n3870 = ~n3868 & ~n3869 ;
  assign n3871 = ~x224 & n3730 ;
  assign n3872 = ~x96 & ~n3730 ;
  assign n3873 = ~n3871 & ~n3872 ;
  assign n3874 = ~n3870 & n3873 ;
  assign n3875 = ~x227 & n3730 ;
  assign n3876 = ~x99 & ~n3730 ;
  assign n3877 = ~n3875 & ~n3876 ;
  assign n3878 = ~x483 & n3359 ;
  assign n3879 = ~x355 & ~n3359 ;
  assign n3880 = ~n3878 & ~n3879 ;
  assign n3881 = n3877 & ~n3880 ;
  assign n3882 = ~x482 & n3359 ;
  assign n3883 = ~x354 & ~n3359 ;
  assign n3884 = ~n3882 & ~n3883 ;
  assign n3885 = ~x226 & n3730 ;
  assign n3886 = ~x98 & ~n3730 ;
  assign n3887 = ~n3885 & ~n3886 ;
  assign n3888 = ~n3884 & n3887 ;
  assign n3889 = ~n3881 & ~n3888 ;
  assign n3890 = ~x225 & n3730 ;
  assign n3891 = ~x97 & ~n3730 ;
  assign n3892 = ~n3890 & ~n3891 ;
  assign n3893 = ~x481 & n3359 ;
  assign n3894 = ~x353 & ~n3359 ;
  assign n3895 = ~n3893 & ~n3894 ;
  assign n3896 = n3892 & ~n3895 ;
  assign n3897 = ~x223 & n3730 ;
  assign n3898 = ~x95 & ~n3730 ;
  assign n3899 = ~n3897 & ~n3898 ;
  assign n3900 = ~x479 & n3359 ;
  assign n3901 = ~x351 & ~n3359 ;
  assign n3902 = ~n3900 & ~n3901 ;
  assign n3903 = ~n3899 & n3902 ;
  assign n3904 = n3899 & ~n3902 ;
  assign n3905 = ~x478 & n3359 ;
  assign n3906 = ~x350 & ~n3359 ;
  assign n3907 = ~n3905 & ~n3906 ;
  assign n3908 = ~x222 & n3730 ;
  assign n3909 = ~x94 & ~n3730 ;
  assign n3910 = ~n3908 & ~n3909 ;
  assign n3911 = ~n3907 & n3910 ;
  assign n3912 = ~n3904 & ~n3911 ;
  assign n3913 = ~x221 & n3730 ;
  assign n3914 = ~x93 & ~n3730 ;
  assign n3915 = ~n3913 & ~n3914 ;
  assign n3916 = ~x477 & n3359 ;
  assign n3917 = ~x349 & ~n3359 ;
  assign n3918 = ~n3916 & ~n3917 ;
  assign n3919 = n3915 & ~n3918 ;
  assign n3920 = ~x220 & n3730 ;
  assign n3921 = ~x92 & ~n3730 ;
  assign n3922 = ~n3920 & ~n3921 ;
  assign n3923 = ~x476 & n3359 ;
  assign n3924 = ~x348 & ~n3359 ;
  assign n3925 = ~n3923 & ~n3924 ;
  assign n3926 = ~n3922 & n3925 ;
  assign n3927 = ~n3919 & n3926 ;
  assign n3928 = ~n3915 & n3918 ;
  assign n3929 = ~n3927 & ~n3928 ;
  assign n3930 = n3912 & ~n3929 ;
  assign n3931 = n3907 & ~n3910 ;
  assign n3932 = ~n3904 & n3931 ;
  assign n3933 = ~x215 & n3730 ;
  assign n3934 = ~x87 & ~n3730 ;
  assign n3935 = ~n3933 & ~n3934 ;
  assign n3936 = ~x471 & n3359 ;
  assign n3937 = ~x343 & ~n3359 ;
  assign n3938 = ~n3936 & ~n3937 ;
  assign n3939 = ~n3935 & n3938 ;
  assign n3940 = n3935 & ~n3938 ;
  assign n3941 = ~x470 & n3359 ;
  assign n3942 = ~x342 & ~n3359 ;
  assign n3943 = ~n3941 & ~n3942 ;
  assign n3944 = ~x214 & n3730 ;
  assign n3945 = ~x86 & ~n3730 ;
  assign n3946 = ~n3944 & ~n3945 ;
  assign n3947 = ~n3943 & n3946 ;
  assign n3948 = ~n3940 & ~n3947 ;
  assign n3949 = ~x213 & n3730 ;
  assign n3950 = ~x85 & ~n3730 ;
  assign n3951 = ~n3949 & ~n3950 ;
  assign n3952 = ~x469 & n3359 ;
  assign n3953 = ~x341 & ~n3359 ;
  assign n3954 = ~n3952 & ~n3953 ;
  assign n3955 = n3951 & ~n3954 ;
  assign n3956 = ~x212 & n3730 ;
  assign n3957 = ~x84 & ~n3730 ;
  assign n3958 = ~n3956 & ~n3957 ;
  assign n3959 = ~x468 & n3359 ;
  assign n3960 = ~x340 & ~n3359 ;
  assign n3961 = ~n3959 & ~n3960 ;
  assign n3962 = ~n3958 & n3961 ;
  assign n3963 = ~n3955 & n3962 ;
  assign n3964 = ~n3951 & n3954 ;
  assign n3965 = ~n3963 & ~n3964 ;
  assign n3966 = n3948 & ~n3965 ;
  assign n3967 = n3943 & ~n3946 ;
  assign n3968 = ~n3940 & n3967 ;
  assign n3969 = ~x464 & n3359 ;
  assign n3970 = ~x336 & ~n3359 ;
  assign n3971 = ~n3969 & ~n3970 ;
  assign n3972 = ~x208 & n3730 ;
  assign n3973 = ~x80 & ~n3730 ;
  assign n3974 = ~n3972 & ~n3973 ;
  assign n3975 = ~n3971 & n3974 ;
  assign n3976 = ~x211 & n3730 ;
  assign n3977 = ~x83 & ~n3730 ;
  assign n3978 = ~n3976 & ~n3977 ;
  assign n3979 = ~x467 & n3359 ;
  assign n3980 = ~x339 & ~n3359 ;
  assign n3981 = ~n3979 & ~n3980 ;
  assign n3982 = n3978 & ~n3981 ;
  assign n3983 = ~x466 & n3359 ;
  assign n3984 = ~x338 & ~n3359 ;
  assign n3985 = ~n3983 & ~n3984 ;
  assign n3986 = ~x210 & n3730 ;
  assign n3987 = ~x82 & ~n3730 ;
  assign n3988 = ~n3986 & ~n3987 ;
  assign n3989 = ~n3985 & n3988 ;
  assign n3990 = ~n3982 & ~n3989 ;
  assign n3991 = ~x209 & n3730 ;
  assign n3992 = ~x81 & ~n3730 ;
  assign n3993 = ~n3991 & ~n3992 ;
  assign n3994 = ~x465 & n3359 ;
  assign n3995 = ~x337 & ~n3359 ;
  assign n3996 = ~n3994 & ~n3995 ;
  assign n3997 = n3993 & ~n3996 ;
  assign n3998 = ~x207 & n3730 ;
  assign n3999 = ~x79 & ~n3730 ;
  assign n4000 = ~n3998 & ~n3999 ;
  assign n4001 = ~x463 & n3359 ;
  assign n4002 = ~x335 & ~n3359 ;
  assign n4003 = ~n4001 & ~n4002 ;
  assign n4004 = ~n4000 & n4003 ;
  assign n4005 = n4000 & ~n4003 ;
  assign n4006 = ~x462 & n3359 ;
  assign n4007 = ~x334 & ~n3359 ;
  assign n4008 = ~n4006 & ~n4007 ;
  assign n4009 = ~x206 & n3730 ;
  assign n4010 = ~x78 & ~n3730 ;
  assign n4011 = ~n4009 & ~n4010 ;
  assign n4012 = ~n4008 & n4011 ;
  assign n4013 = ~n4005 & ~n4012 ;
  assign n4014 = ~x205 & n3730 ;
  assign n4015 = ~x77 & ~n3730 ;
  assign n4016 = ~n4014 & ~n4015 ;
  assign n4017 = ~x461 & n3359 ;
  assign n4018 = ~x333 & ~n3359 ;
  assign n4019 = ~n4017 & ~n4018 ;
  assign n4020 = n4016 & ~n4019 ;
  assign n4021 = ~x204 & n3730 ;
  assign n4022 = ~x76 & ~n3730 ;
  assign n4023 = ~n4021 & ~n4022 ;
  assign n4024 = ~x460 & n3359 ;
  assign n4025 = ~x332 & ~n3359 ;
  assign n4026 = ~n4024 & ~n4025 ;
  assign n4027 = ~n4023 & n4026 ;
  assign n4028 = ~n4020 & n4027 ;
  assign n4029 = ~n4016 & n4019 ;
  assign n4030 = ~n4028 & ~n4029 ;
  assign n4031 = n4013 & ~n4030 ;
  assign n4032 = n4008 & ~n4011 ;
  assign n4033 = ~n4005 & n4032 ;
  assign n4034 = ~x199 & n3730 ;
  assign n4035 = ~x71 & ~n3730 ;
  assign n4036 = ~n4034 & ~n4035 ;
  assign n4037 = ~x455 & n3359 ;
  assign n4038 = ~x327 & ~n3359 ;
  assign n4039 = ~n4037 & ~n4038 ;
  assign n4040 = ~n4036 & n4039 ;
  assign n4041 = n4036 & ~n4039 ;
  assign n4042 = ~x454 & n3359 ;
  assign n4043 = ~x326 & ~n3359 ;
  assign n4044 = ~n4042 & ~n4043 ;
  assign n4045 = ~x198 & n3730 ;
  assign n4046 = ~x70 & ~n3730 ;
  assign n4047 = ~n4045 & ~n4046 ;
  assign n4048 = ~n4044 & n4047 ;
  assign n4049 = ~n4041 & ~n4048 ;
  assign n4050 = ~x197 & n3730 ;
  assign n4051 = ~x69 & ~n3730 ;
  assign n4052 = ~n4050 & ~n4051 ;
  assign n4053 = ~x453 & n3359 ;
  assign n4054 = ~x325 & ~n3359 ;
  assign n4055 = ~n4053 & ~n4054 ;
  assign n4056 = n4052 & ~n4055 ;
  assign n4057 = ~x196 & n3730 ;
  assign n4058 = ~x68 & ~n3730 ;
  assign n4059 = ~n4057 & ~n4058 ;
  assign n4060 = ~x452 & n3359 ;
  assign n4061 = ~x324 & ~n3359 ;
  assign n4062 = ~n4060 & ~n4061 ;
  assign n4063 = ~n4059 & n4062 ;
  assign n4064 = ~n4056 & n4063 ;
  assign n4065 = ~n4052 & n4055 ;
  assign n4066 = ~n4064 & ~n4065 ;
  assign n4067 = n4049 & ~n4066 ;
  assign n4068 = n4044 & ~n4047 ;
  assign n4069 = ~n4041 & n4068 ;
  assign n4070 = ~x195 & n3730 ;
  assign n4071 = ~x67 & ~n3730 ;
  assign n4072 = ~n4070 & ~n4071 ;
  assign n4073 = ~x451 & n3359 ;
  assign n4074 = ~x323 & ~n3359 ;
  assign n4075 = ~n4073 & ~n4074 ;
  assign n4076 = n4072 & ~n4075 ;
  assign n4077 = ~x450 & n3359 ;
  assign n4078 = ~x322 & ~n3359 ;
  assign n4079 = ~n4077 & ~n4078 ;
  assign n4080 = ~x194 & n3730 ;
  assign n4081 = ~x66 & ~n3730 ;
  assign n4082 = ~n4080 & ~n4081 ;
  assign n4083 = ~n4079 & n4082 ;
  assign n4084 = ~n4076 & ~n4083 ;
  assign n4085 = ~x448 & n3359 ;
  assign n4086 = ~x320 & ~n3359 ;
  assign n4087 = ~n4085 & ~n4086 ;
  assign n4088 = ~x192 & n3730 ;
  assign n4089 = ~x64 & ~n3730 ;
  assign n4090 = ~n4088 & ~n4089 ;
  assign n4091 = ~n4087 & n4090 ;
  assign n4092 = ~x193 & n3730 ;
  assign n4093 = ~x65 & ~n3730 ;
  assign n4094 = ~n4092 & ~n4093 ;
  assign n4095 = ~x449 & n3359 ;
  assign n4096 = ~x321 & ~n3359 ;
  assign n4097 = ~n4095 & ~n4096 ;
  assign n4098 = n4094 & ~n4097 ;
  assign n4099 = ~x191 & n3730 ;
  assign n4100 = ~x63 & ~n3730 ;
  assign n4101 = ~n4099 & ~n4100 ;
  assign n4102 = ~x447 & n3359 ;
  assign n4103 = ~x319 & ~n3359 ;
  assign n4104 = ~n4102 & ~n4103 ;
  assign n4105 = ~n4101 & n4104 ;
  assign n4106 = n4101 & ~n4104 ;
  assign n4107 = ~x446 & n3359 ;
  assign n4108 = ~x318 & ~n3359 ;
  assign n4109 = ~n4107 & ~n4108 ;
  assign n4110 = ~x190 & n3730 ;
  assign n4111 = ~x62 & ~n3730 ;
  assign n4112 = ~n4110 & ~n4111 ;
  assign n4113 = ~n4109 & n4112 ;
  assign n4114 = ~n4106 & ~n4113 ;
  assign n4115 = ~x188 & n3730 ;
  assign n4116 = ~x60 & ~n3730 ;
  assign n4117 = ~n4115 & ~n4116 ;
  assign n4118 = ~x444 & n3359 ;
  assign n4119 = ~x316 & ~n3359 ;
  assign n4120 = ~n4118 & ~n4119 ;
  assign n4121 = n4117 & ~n4120 ;
  assign n4122 = ~x189 & n3730 ;
  assign n4123 = ~x61 & ~n3730 ;
  assign n4124 = ~n4122 & ~n4123 ;
  assign n4125 = ~x445 & n3359 ;
  assign n4126 = ~x317 & ~n3359 ;
  assign n4127 = ~n4125 & ~n4126 ;
  assign n4128 = n4124 & ~n4127 ;
  assign n4129 = ~n4121 & ~n4128 ;
  assign n4130 = n4114 & n4129 ;
  assign n4131 = ~x187 & n3730 ;
  assign n4132 = ~x59 & ~n3730 ;
  assign n4133 = ~n4131 & ~n4132 ;
  assign n4134 = ~x443 & n3359 ;
  assign n4135 = ~x315 & ~n3359 ;
  assign n4136 = ~n4134 & ~n4135 ;
  assign n4137 = ~n4133 & n4136 ;
  assign n4138 = n4133 & ~n4136 ;
  assign n4139 = ~x186 & n3730 ;
  assign n4140 = ~x58 & ~n3730 ;
  assign n4141 = ~n4139 & ~n4140 ;
  assign n4142 = ~x442 & n3359 ;
  assign n4143 = ~x314 & ~n3359 ;
  assign n4144 = ~n4142 & ~n4143 ;
  assign n4145 = n4141 & ~n4144 ;
  assign n4146 = ~n4138 & ~n4145 ;
  assign n4147 = ~x185 & n3730 ;
  assign n4148 = ~x57 & ~n3730 ;
  assign n4149 = ~n4147 & ~n4148 ;
  assign n4150 = ~x441 & n3359 ;
  assign n4151 = ~x313 & ~n3359 ;
  assign n4152 = ~n4150 & ~n4151 ;
  assign n4153 = n4149 & ~n4152 ;
  assign n4154 = ~x184 & n3730 ;
  assign n4155 = ~x56 & ~n3730 ;
  assign n4156 = ~n4154 & ~n4155 ;
  assign n4157 = ~x440 & n3359 ;
  assign n4158 = ~x312 & ~n3359 ;
  assign n4159 = ~n4157 & ~n4158 ;
  assign n4160 = ~n4156 & n4159 ;
  assign n4161 = ~n4153 & n4160 ;
  assign n4162 = ~n4149 & n4152 ;
  assign n4163 = ~n4161 & ~n4162 ;
  assign n4164 = ~n4141 & n4144 ;
  assign n4165 = n4163 & ~n4164 ;
  assign n4166 = n4146 & ~n4165 ;
  assign n4167 = ~n4137 & ~n4166 ;
  assign n4168 = n4130 & ~n4167 ;
  assign n4169 = ~n4117 & n4120 ;
  assign n4170 = ~n4128 & n4169 ;
  assign n4171 = ~n4124 & n4127 ;
  assign n4172 = ~n4170 & ~n4171 ;
  assign n4173 = n4114 & ~n4172 ;
  assign n4174 = n4109 & ~n4112 ;
  assign n4175 = ~n4106 & n4174 ;
  assign n4176 = ~x175 & n3730 ;
  assign n4177 = ~x47 & ~n3730 ;
  assign n4178 = ~n4176 & ~n4177 ;
  assign n4179 = ~x431 & n3359 ;
  assign n4180 = ~x303 & ~n3359 ;
  assign n4181 = ~n4179 & ~n4180 ;
  assign n4182 = ~n4178 & n4181 ;
  assign n4183 = n4178 & ~n4181 ;
  assign n4184 = ~x430 & n3359 ;
  assign n4185 = ~x302 & ~n3359 ;
  assign n4186 = ~n4184 & ~n4185 ;
  assign n4187 = ~x174 & n3730 ;
  assign n4188 = ~x46 & ~n3730 ;
  assign n4189 = ~n4187 & ~n4188 ;
  assign n4190 = ~n4186 & n4189 ;
  assign n4191 = ~n4183 & ~n4190 ;
  assign n4192 = ~x172 & n3730 ;
  assign n4193 = ~x44 & ~n3730 ;
  assign n4194 = ~n4192 & ~n4193 ;
  assign n4195 = ~x428 & n3359 ;
  assign n4196 = ~x300 & ~n3359 ;
  assign n4197 = ~n4195 & ~n4196 ;
  assign n4198 = n4194 & ~n4197 ;
  assign n4199 = ~x173 & n3730 ;
  assign n4200 = ~x45 & ~n3730 ;
  assign n4201 = ~n4199 & ~n4200 ;
  assign n4202 = ~x429 & n3359 ;
  assign n4203 = ~x301 & ~n3359 ;
  assign n4204 = ~n4202 & ~n4203 ;
  assign n4205 = n4201 & ~n4204 ;
  assign n4206 = ~n4198 & ~n4205 ;
  assign n4207 = n4191 & n4206 ;
  assign n4208 = ~x171 & n3730 ;
  assign n4209 = ~x43 & ~n3730 ;
  assign n4210 = ~n4208 & ~n4209 ;
  assign n4211 = ~x427 & n3359 ;
  assign n4212 = ~x299 & ~n3359 ;
  assign n4213 = ~n4211 & ~n4212 ;
  assign n4214 = ~n4210 & n4213 ;
  assign n4215 = n4210 & ~n4213 ;
  assign n4216 = ~x170 & n3730 ;
  assign n4217 = ~x42 & ~n3730 ;
  assign n4218 = ~n4216 & ~n4217 ;
  assign n4219 = ~x426 & n3359 ;
  assign n4220 = ~x298 & ~n3359 ;
  assign n4221 = ~n4219 & ~n4220 ;
  assign n4222 = n4218 & ~n4221 ;
  assign n4223 = ~n4215 & ~n4222 ;
  assign n4224 = ~x169 & n3730 ;
  assign n4225 = ~x41 & ~n3730 ;
  assign n4226 = ~n4224 & ~n4225 ;
  assign n4227 = ~x425 & n3359 ;
  assign n4228 = ~x297 & ~n3359 ;
  assign n4229 = ~n4227 & ~n4228 ;
  assign n4230 = n4226 & ~n4229 ;
  assign n4231 = ~x168 & n3730 ;
  assign n4232 = ~x40 & ~n3730 ;
  assign n4233 = ~n4231 & ~n4232 ;
  assign n4234 = ~x424 & n3359 ;
  assign n4235 = ~x296 & ~n3359 ;
  assign n4236 = ~n4234 & ~n4235 ;
  assign n4237 = ~n4233 & n4236 ;
  assign n4238 = ~n4230 & n4237 ;
  assign n4239 = ~n4226 & n4229 ;
  assign n4240 = ~n4238 & ~n4239 ;
  assign n4241 = ~n4218 & n4221 ;
  assign n4242 = n4240 & ~n4241 ;
  assign n4243 = n4223 & ~n4242 ;
  assign n4244 = ~n4214 & ~n4243 ;
  assign n4245 = n4207 & ~n4244 ;
  assign n4246 = ~n4194 & n4197 ;
  assign n4247 = ~n4205 & n4246 ;
  assign n4248 = ~n4201 & n4204 ;
  assign n4249 = ~n4247 & ~n4248 ;
  assign n4250 = n4191 & ~n4249 ;
  assign n4251 = n4186 & ~n4189 ;
  assign n4252 = ~n4183 & n4251 ;
  assign n4253 = ~x416 & n3359 ;
  assign n4254 = ~x288 & ~n3359 ;
  assign n4255 = ~n4253 & ~n4254 ;
  assign n4256 = ~x160 & n3730 ;
  assign n4257 = ~x32 & ~n3730 ;
  assign n4258 = ~n4256 & ~n4257 ;
  assign n4259 = ~n4255 & n4258 ;
  assign n4260 = ~x159 & n3730 ;
  assign n4261 = ~x31 & ~n3730 ;
  assign n4262 = ~n4260 & ~n4261 ;
  assign n4263 = ~x415 & n3359 ;
  assign n4264 = ~x287 & ~n3359 ;
  assign n4265 = ~n4263 & ~n4264 ;
  assign n4266 = n4262 & ~n4265 ;
  assign n4267 = ~x158 & n3730 ;
  assign n4268 = ~x30 & ~n3730 ;
  assign n4269 = ~n4267 & ~n4268 ;
  assign n4270 = ~x414 & n3359 ;
  assign n4271 = ~x286 & ~n3359 ;
  assign n4272 = ~n4270 & ~n4271 ;
  assign n4273 = n4269 & ~n4272 ;
  assign n4274 = ~x157 & n3730 ;
  assign n4275 = ~x29 & ~n3730 ;
  assign n4276 = ~n4274 & ~n4275 ;
  assign n4277 = ~x413 & n3359 ;
  assign n4278 = ~x285 & ~n3359 ;
  assign n4279 = ~n4277 & ~n4278 ;
  assign n4280 = n4276 & ~n4279 ;
  assign n4281 = ~x156 & n3730 ;
  assign n4282 = ~x28 & ~n3730 ;
  assign n4283 = ~n4281 & ~n4282 ;
  assign n4284 = ~x412 & n3359 ;
  assign n4285 = ~x284 & ~n3359 ;
  assign n4286 = ~n4284 & ~n4285 ;
  assign n4287 = n4283 & ~n4286 ;
  assign n4288 = ~x155 & n3730 ;
  assign n4289 = ~x27 & ~n3730 ;
  assign n4290 = ~n4288 & ~n4289 ;
  assign n4291 = ~x411 & n3359 ;
  assign n4292 = ~x283 & ~n3359 ;
  assign n4293 = ~n4291 & ~n4292 ;
  assign n4294 = n4290 & ~n4293 ;
  assign n4295 = ~x154 & n3730 ;
  assign n4296 = ~x26 & ~n3730 ;
  assign n4297 = ~n4295 & ~n4296 ;
  assign n4298 = ~x410 & n3359 ;
  assign n4299 = ~x282 & ~n3359 ;
  assign n4300 = ~n4298 & ~n4299 ;
  assign n4301 = n4297 & ~n4300 ;
  assign n4302 = ~x409 & n3359 ;
  assign n4303 = ~x281 & ~n3359 ;
  assign n4304 = ~n4302 & ~n4303 ;
  assign n4305 = ~x408 & n3359 ;
  assign n4306 = ~x280 & ~n3359 ;
  assign n4307 = ~n4305 & ~n4306 ;
  assign n4308 = ~x151 & n3730 ;
  assign n4309 = ~x23 & ~n3730 ;
  assign n4310 = ~n4308 & ~n4309 ;
  assign n4311 = ~x407 & n3359 ;
  assign n4312 = ~x279 & ~n3359 ;
  assign n4313 = ~n4311 & ~n4312 ;
  assign n4314 = n4310 & ~n4313 ;
  assign n4315 = ~x150 & n3730 ;
  assign n4316 = ~x22 & ~n3730 ;
  assign n4317 = ~n4315 & ~n4316 ;
  assign n4318 = ~x406 & n3359 ;
  assign n4319 = ~x278 & ~n3359 ;
  assign n4320 = ~n4318 & ~n4319 ;
  assign n4321 = n4317 & ~n4320 ;
  assign n4322 = ~x149 & n3730 ;
  assign n4323 = ~x21 & ~n3730 ;
  assign n4324 = ~n4322 & ~n4323 ;
  assign n4325 = ~x405 & n3359 ;
  assign n4326 = ~x277 & ~n3359 ;
  assign n4327 = ~n4325 & ~n4326 ;
  assign n4328 = n4324 & ~n4327 ;
  assign n4329 = ~x148 & n3730 ;
  assign n4330 = ~x20 & ~n3730 ;
  assign n4331 = ~n4329 & ~n4330 ;
  assign n4332 = ~x404 & n3359 ;
  assign n4333 = ~x276 & ~n3359 ;
  assign n4334 = ~n4332 & ~n4333 ;
  assign n4335 = n4331 & ~n4334 ;
  assign n4336 = ~x147 & n3730 ;
  assign n4337 = ~x19 & ~n3730 ;
  assign n4338 = ~n4336 & ~n4337 ;
  assign n4339 = ~x403 & n3359 ;
  assign n4340 = ~x275 & ~n3359 ;
  assign n4341 = ~n4339 & ~n4340 ;
  assign n4342 = n4338 & ~n4341 ;
  assign n4343 = ~x146 & n3730 ;
  assign n4344 = ~x18 & ~n3730 ;
  assign n4345 = ~n4343 & ~n4344 ;
  assign n4346 = ~x402 & n3359 ;
  assign n4347 = ~x274 & ~n3359 ;
  assign n4348 = ~n4346 & ~n4347 ;
  assign n4349 = n4345 & ~n4348 ;
  assign n4350 = ~x401 & n3359 ;
  assign n4351 = ~x273 & ~n3359 ;
  assign n4352 = ~n4350 & ~n4351 ;
  assign n4353 = ~x400 & n3359 ;
  assign n4354 = ~x272 & ~n3359 ;
  assign n4355 = ~n4353 & ~n4354 ;
  assign n4356 = ~x143 & n3730 ;
  assign n4357 = ~x15 & ~n3730 ;
  assign n4358 = ~n4356 & ~n4357 ;
  assign n4359 = ~x399 & n3359 ;
  assign n4360 = ~x271 & ~n3359 ;
  assign n4361 = ~n4359 & ~n4360 ;
  assign n4362 = n4358 & ~n4361 ;
  assign n4363 = ~x142 & n3730 ;
  assign n4364 = ~x14 & ~n3730 ;
  assign n4365 = ~n4363 & ~n4364 ;
  assign n4366 = ~x398 & n3359 ;
  assign n4367 = ~x270 & ~n3359 ;
  assign n4368 = ~n4366 & ~n4367 ;
  assign n4369 = n4365 & ~n4368 ;
  assign n4370 = ~x141 & n3730 ;
  assign n4371 = ~x13 & ~n3730 ;
  assign n4372 = ~n4370 & ~n4371 ;
  assign n4373 = ~x397 & n3359 ;
  assign n4374 = ~x269 & ~n3359 ;
  assign n4375 = ~n4373 & ~n4374 ;
  assign n4376 = n4372 & ~n4375 ;
  assign n4377 = ~x140 & n3730 ;
  assign n4378 = ~x12 & ~n3730 ;
  assign n4379 = ~n4377 & ~n4378 ;
  assign n4380 = ~x396 & n3359 ;
  assign n4381 = ~x268 & ~n3359 ;
  assign n4382 = ~n4380 & ~n4381 ;
  assign n4383 = n4379 & ~n4382 ;
  assign n4384 = ~x139 & n3730 ;
  assign n4385 = ~x11 & ~n3730 ;
  assign n4386 = ~n4384 & ~n4385 ;
  assign n4387 = ~x395 & n3359 ;
  assign n4388 = ~x267 & ~n3359 ;
  assign n4389 = ~n4387 & ~n4388 ;
  assign n4390 = n4386 & ~n4389 ;
  assign n4391 = ~x138 & n3730 ;
  assign n4392 = ~x10 & ~n3730 ;
  assign n4393 = ~n4391 & ~n4392 ;
  assign n4394 = ~x394 & n3359 ;
  assign n4395 = ~x266 & ~n3359 ;
  assign n4396 = ~n4394 & ~n4395 ;
  assign n4397 = n4393 & ~n4396 ;
  assign n4398 = ~x393 & n3359 ;
  assign n4399 = ~x265 & ~n3359 ;
  assign n4400 = ~n4398 & ~n4399 ;
  assign n4401 = ~x392 & n3359 ;
  assign n4402 = ~x264 & ~n3359 ;
  assign n4403 = ~n4401 & ~n4402 ;
  assign n4404 = ~x135 & n3730 ;
  assign n4405 = ~x7 & ~n3730 ;
  assign n4406 = ~n4404 & ~n4405 ;
  assign n4407 = ~x391 & n3359 ;
  assign n4408 = ~x263 & ~n3359 ;
  assign n4409 = ~n4407 & ~n4408 ;
  assign n4410 = n4406 & ~n4409 ;
  assign n4411 = ~x390 & n3359 ;
  assign n4412 = ~x262 & ~n3359 ;
  assign n4413 = ~n4411 & ~n4412 ;
  assign n4414 = ~x134 & n3730 ;
  assign n4415 = ~x6 & ~n3730 ;
  assign n4416 = ~n4414 & ~n4415 ;
  assign n4417 = ~x389 & n3359 ;
  assign n4418 = ~x261 & ~n3359 ;
  assign n4419 = ~n4417 & ~n4418 ;
  assign n4420 = ~x133 & n3730 ;
  assign n4421 = ~x5 & ~n3730 ;
  assign n4422 = ~n4420 & ~n4421 ;
  assign n4423 = ~x388 & n3359 ;
  assign n4424 = ~x260 & ~n3359 ;
  assign n4425 = ~n4423 & ~n4424 ;
  assign n4426 = ~x132 & n3730 ;
  assign n4427 = ~x4 & ~n3730 ;
  assign n4428 = ~n4426 & ~n4427 ;
  assign n4429 = ~x131 & n3730 ;
  assign n4430 = ~x3 & ~n3730 ;
  assign n4431 = ~n4429 & ~n4430 ;
  assign n4432 = ~x387 & n3359 ;
  assign n4433 = ~x259 & ~n3359 ;
  assign n4434 = ~n4432 & ~n4433 ;
  assign n4435 = n4431 & ~n4434 ;
  assign n4436 = ~x385 & n3359 ;
  assign n4437 = ~x257 & ~n3359 ;
  assign n4438 = ~n4436 & ~n4437 ;
  assign n4439 = ~x128 & n3730 ;
  assign n4440 = ~x0 & ~n3730 ;
  assign n4441 = ~n4439 & ~n4440 ;
  assign n4442 = n3362 & ~n4441 ;
  assign n4443 = n4438 & n4442 ;
  assign n4444 = ~x129 & n3730 ;
  assign n4445 = ~x1 & ~n3730 ;
  assign n4446 = ~n4444 & ~n4445 ;
  assign n4447 = ~n4443 & n4446 ;
  assign n4448 = ~x130 & n3730 ;
  assign n4449 = ~x2 & ~n3730 ;
  assign n4450 = ~n4448 & ~n4449 ;
  assign n4451 = ~x386 & n3359 ;
  assign n4452 = ~x258 & ~n3359 ;
  assign n4453 = ~n4451 & ~n4452 ;
  assign n4454 = n4450 & ~n4453 ;
  assign n4455 = ~n4438 & ~n4442 ;
  assign n4456 = ~n4454 & ~n4455 ;
  assign n4457 = ~n4447 & n4456 ;
  assign n4458 = ~n4450 & n4453 ;
  assign n4459 = ~n4457 & ~n4458 ;
  assign n4460 = ~n4435 & ~n4459 ;
  assign n4461 = ~n4431 & n4434 ;
  assign n4462 = ~n4460 & ~n4461 ;
  assign n4463 = n4428 & n4462 ;
  assign n4464 = n4425 & ~n4463 ;
  assign n4465 = ~n4428 & ~n4462 ;
  assign n4466 = ~n4464 & ~n4465 ;
  assign n4467 = n4422 & n4466 ;
  assign n4468 = n4419 & ~n4467 ;
  assign n4469 = ~n4422 & ~n4466 ;
  assign n4470 = ~n4468 & ~n4469 ;
  assign n4471 = n4416 & n4470 ;
  assign n4472 = n4413 & ~n4471 ;
  assign n4473 = ~n4416 & ~n4470 ;
  assign n4474 = ~n4472 & ~n4473 ;
  assign n4475 = ~n4410 & ~n4474 ;
  assign n4476 = ~n4406 & n4409 ;
  assign n4477 = ~n4475 & ~n4476 ;
  assign n4478 = ~x136 & n3730 ;
  assign n4479 = ~x8 & ~n3730 ;
  assign n4480 = ~n4478 & ~n4479 ;
  assign n4481 = n4477 & n4480 ;
  assign n4482 = n4403 & ~n4481 ;
  assign n4483 = ~n4477 & ~n4480 ;
  assign n4484 = ~n4482 & ~n4483 ;
  assign n4485 = ~x137 & n3730 ;
  assign n4486 = ~x9 & ~n3730 ;
  assign n4487 = ~n4485 & ~n4486 ;
  assign n4488 = n4484 & n4487 ;
  assign n4489 = n4400 & ~n4488 ;
  assign n4490 = ~n4484 & ~n4487 ;
  assign n4491 = ~n4489 & ~n4490 ;
  assign n4492 = ~n4397 & ~n4491 ;
  assign n4493 = ~n4393 & n4396 ;
  assign n4494 = ~n4492 & ~n4493 ;
  assign n4495 = ~n4390 & ~n4494 ;
  assign n4496 = ~n4386 & n4389 ;
  assign n4497 = ~n4495 & ~n4496 ;
  assign n4498 = ~n4383 & ~n4497 ;
  assign n4499 = ~n4379 & n4382 ;
  assign n4500 = ~n4498 & ~n4499 ;
  assign n4501 = ~n4376 & ~n4500 ;
  assign n4502 = ~n4372 & n4375 ;
  assign n4503 = ~n4501 & ~n4502 ;
  assign n4504 = ~n4369 & ~n4503 ;
  assign n4505 = ~n4365 & n4368 ;
  assign n4506 = ~n4504 & ~n4505 ;
  assign n4507 = ~n4362 & ~n4506 ;
  assign n4508 = ~n4358 & n4361 ;
  assign n4509 = ~n4507 & ~n4508 ;
  assign n4510 = ~x144 & n3730 ;
  assign n4511 = ~x16 & ~n3730 ;
  assign n4512 = ~n4510 & ~n4511 ;
  assign n4513 = n4509 & n4512 ;
  assign n4514 = n4355 & ~n4513 ;
  assign n4515 = ~n4509 & ~n4512 ;
  assign n4516 = ~n4514 & ~n4515 ;
  assign n4517 = ~x145 & n3730 ;
  assign n4518 = ~x17 & ~n3730 ;
  assign n4519 = ~n4517 & ~n4518 ;
  assign n4520 = n4516 & n4519 ;
  assign n4521 = n4352 & ~n4520 ;
  assign n4522 = ~n4516 & ~n4519 ;
  assign n4523 = ~n4521 & ~n4522 ;
  assign n4524 = ~n4349 & ~n4523 ;
  assign n4525 = ~n4345 & n4348 ;
  assign n4526 = ~n4524 & ~n4525 ;
  assign n4527 = ~n4342 & ~n4526 ;
  assign n4528 = ~n4338 & n4341 ;
  assign n4529 = ~n4527 & ~n4528 ;
  assign n4530 = ~n4335 & ~n4529 ;
  assign n4531 = ~n4331 & n4334 ;
  assign n4532 = ~n4530 & ~n4531 ;
  assign n4533 = ~n4328 & ~n4532 ;
  assign n4534 = ~n4324 & n4327 ;
  assign n4535 = ~n4533 & ~n4534 ;
  assign n4536 = ~n4321 & ~n4535 ;
  assign n4537 = ~n4317 & n4320 ;
  assign n4538 = ~n4536 & ~n4537 ;
  assign n4539 = ~n4314 & ~n4538 ;
  assign n4540 = ~n4310 & n4313 ;
  assign n4541 = ~n4539 & ~n4540 ;
  assign n4542 = ~x152 & n3730 ;
  assign n4543 = ~x24 & ~n3730 ;
  assign n4544 = ~n4542 & ~n4543 ;
  assign n4545 = n4541 & n4544 ;
  assign n4546 = n4307 & ~n4545 ;
  assign n4547 = ~n4541 & ~n4544 ;
  assign n4548 = ~n4546 & ~n4547 ;
  assign n4549 = ~x153 & n3730 ;
  assign n4550 = ~x25 & ~n3730 ;
  assign n4551 = ~n4549 & ~n4550 ;
  assign n4552 = n4548 & n4551 ;
  assign n4553 = n4304 & ~n4552 ;
  assign n4554 = ~n4548 & ~n4551 ;
  assign n4555 = ~n4553 & ~n4554 ;
  assign n4556 = ~n4301 & ~n4555 ;
  assign n4557 = ~n4297 & n4300 ;
  assign n4558 = ~n4556 & ~n4557 ;
  assign n4559 = ~n4294 & ~n4558 ;
  assign n4560 = ~n4290 & n4293 ;
  assign n4561 = ~n4559 & ~n4560 ;
  assign n4562 = ~n4287 & ~n4561 ;
  assign n4563 = ~n4283 & n4286 ;
  assign n4564 = ~n4562 & ~n4563 ;
  assign n4565 = ~n4280 & ~n4564 ;
  assign n4566 = ~n4276 & n4279 ;
  assign n4567 = ~n4565 & ~n4566 ;
  assign n4568 = ~n4273 & ~n4567 ;
  assign n4569 = ~n4269 & n4272 ;
  assign n4570 = ~n4568 & ~n4569 ;
  assign n4571 = ~n4266 & ~n4570 ;
  assign n4572 = ~n4262 & n4265 ;
  assign n4573 = ~n4571 & ~n4572 ;
  assign n4574 = ~x167 & n3730 ;
  assign n4575 = ~x39 & ~n3730 ;
  assign n4576 = ~n4574 & ~n4575 ;
  assign n4577 = ~x423 & n3359 ;
  assign n4578 = ~x295 & ~n3359 ;
  assign n4579 = ~n4577 & ~n4578 ;
  assign n4580 = n4576 & ~n4579 ;
  assign n4581 = ~x422 & n3359 ;
  assign n4582 = ~x294 & ~n3359 ;
  assign n4583 = ~n4581 & ~n4582 ;
  assign n4584 = ~x166 & n3730 ;
  assign n4585 = ~x38 & ~n3730 ;
  assign n4586 = ~n4584 & ~n4585 ;
  assign n4587 = ~n4583 & n4586 ;
  assign n4588 = ~n4580 & ~n4587 ;
  assign n4589 = ~x164 & n3730 ;
  assign n4590 = ~x36 & ~n3730 ;
  assign n4591 = ~n4589 & ~n4590 ;
  assign n4592 = ~x420 & n3359 ;
  assign n4593 = ~x292 & ~n3359 ;
  assign n4594 = ~n4592 & ~n4593 ;
  assign n4595 = n4591 & ~n4594 ;
  assign n4596 = ~x165 & n3730 ;
  assign n4597 = ~x37 & ~n3730 ;
  assign n4598 = ~n4596 & ~n4597 ;
  assign n4599 = ~x421 & n3359 ;
  assign n4600 = ~x293 & ~n3359 ;
  assign n4601 = ~n4599 & ~n4600 ;
  assign n4602 = n4598 & ~n4601 ;
  assign n4603 = ~n4595 & ~n4602 ;
  assign n4604 = n4588 & n4603 ;
  assign n4605 = ~x161 & n3730 ;
  assign n4606 = ~x33 & ~n3730 ;
  assign n4607 = ~n4605 & ~n4606 ;
  assign n4608 = ~x417 & n3359 ;
  assign n4609 = ~x289 & ~n3359 ;
  assign n4610 = ~n4608 & ~n4609 ;
  assign n4611 = n4607 & ~n4610 ;
  assign n4612 = ~x163 & n3730 ;
  assign n4613 = ~x35 & ~n3730 ;
  assign n4614 = ~n4612 & ~n4613 ;
  assign n4615 = ~x419 & n3359 ;
  assign n4616 = ~x291 & ~n3359 ;
  assign n4617 = ~n4615 & ~n4616 ;
  assign n4618 = n4614 & ~n4617 ;
  assign n4619 = ~x418 & n3359 ;
  assign n4620 = ~x290 & ~n3359 ;
  assign n4621 = ~n4619 & ~n4620 ;
  assign n4622 = ~x162 & n3730 ;
  assign n4623 = ~x34 & ~n3730 ;
  assign n4624 = ~n4622 & ~n4623 ;
  assign n4625 = ~n4621 & n4624 ;
  assign n4626 = ~n4618 & ~n4625 ;
  assign n4627 = ~n4611 & n4626 ;
  assign n4628 = n4604 & n4627 ;
  assign n4629 = ~n4573 & n4628 ;
  assign n4630 = ~n4259 & n4629 ;
  assign n4631 = ~n4576 & n4579 ;
  assign n4632 = ~n4591 & n4594 ;
  assign n4633 = ~n4602 & n4632 ;
  assign n4634 = ~n4598 & n4601 ;
  assign n4635 = ~n4633 & ~n4634 ;
  assign n4636 = n4588 & ~n4635 ;
  assign n4637 = ~n4580 & n4583 ;
  assign n4638 = ~n4586 & n4637 ;
  assign n4639 = ~n4614 & n4617 ;
  assign n4640 = ~n4618 & n4621 ;
  assign n4641 = ~n4624 & n4640 ;
  assign n4642 = n4255 & ~n4258 ;
  assign n4643 = ~n4607 & n4610 ;
  assign n4644 = ~n4642 & ~n4643 ;
  assign n4645 = n4627 & ~n4644 ;
  assign n4646 = ~n4641 & ~n4645 ;
  assign n4647 = ~n4639 & n4646 ;
  assign n4648 = n4604 & ~n4647 ;
  assign n4649 = ~n4638 & ~n4648 ;
  assign n4650 = ~n4636 & n4649 ;
  assign n4651 = ~n4631 & n4650 ;
  assign n4652 = ~n4630 & n4651 ;
  assign n4653 = n4233 & ~n4236 ;
  assign n4654 = ~n4230 & ~n4653 ;
  assign n4655 = n4223 & n4654 ;
  assign n4656 = n4207 & n4655 ;
  assign n4657 = ~n4652 & n4656 ;
  assign n4658 = ~n4252 & ~n4657 ;
  assign n4659 = ~n4250 & n4658 ;
  assign n4660 = ~n4245 & n4659 ;
  assign n4661 = ~n4182 & n4660 ;
  assign n4662 = ~x432 & n3359 ;
  assign n4663 = ~x304 & ~n3359 ;
  assign n4664 = ~n4662 & ~n4663 ;
  assign n4665 = ~x176 & n3730 ;
  assign n4666 = ~x48 & ~n3730 ;
  assign n4667 = ~n4665 & ~n4666 ;
  assign n4668 = ~n4664 & n4667 ;
  assign n4669 = ~x183 & n3730 ;
  assign n4670 = ~x55 & ~n3730 ;
  assign n4671 = ~n4669 & ~n4670 ;
  assign n4672 = ~x439 & n3359 ;
  assign n4673 = ~x311 & ~n3359 ;
  assign n4674 = ~n4672 & ~n4673 ;
  assign n4675 = n4671 & ~n4674 ;
  assign n4676 = ~x438 & n3359 ;
  assign n4677 = ~x310 & ~n3359 ;
  assign n4678 = ~n4676 & ~n4677 ;
  assign n4679 = ~x182 & n3730 ;
  assign n4680 = ~x54 & ~n3730 ;
  assign n4681 = ~n4679 & ~n4680 ;
  assign n4682 = ~n4678 & n4681 ;
  assign n4683 = ~n4675 & ~n4682 ;
  assign n4684 = ~x181 & n3730 ;
  assign n4685 = ~x53 & ~n3730 ;
  assign n4686 = ~n4684 & ~n4685 ;
  assign n4687 = ~x437 & n3359 ;
  assign n4688 = ~x309 & ~n3359 ;
  assign n4689 = ~n4687 & ~n4688 ;
  assign n4690 = n4686 & ~n4689 ;
  assign n4691 = ~x436 & n3359 ;
  assign n4692 = ~x308 & ~n3359 ;
  assign n4693 = ~n4691 & ~n4692 ;
  assign n4694 = ~x180 & n3730 ;
  assign n4695 = ~x52 & ~n3730 ;
  assign n4696 = ~n4694 & ~n4695 ;
  assign n4697 = ~n4693 & n4696 ;
  assign n4698 = ~n4690 & ~n4697 ;
  assign n4699 = n4683 & n4698 ;
  assign n4700 = ~x177 & n3730 ;
  assign n4701 = ~x49 & ~n3730 ;
  assign n4702 = ~n4700 & ~n4701 ;
  assign n4703 = ~x433 & n3359 ;
  assign n4704 = ~x305 & ~n3359 ;
  assign n4705 = ~n4703 & ~n4704 ;
  assign n4706 = n4702 & ~n4705 ;
  assign n4707 = ~x179 & n3730 ;
  assign n4708 = ~x51 & ~n3730 ;
  assign n4709 = ~n4707 & ~n4708 ;
  assign n4710 = ~x435 & n3359 ;
  assign n4711 = ~x307 & ~n3359 ;
  assign n4712 = ~n4710 & ~n4711 ;
  assign n4713 = n4709 & ~n4712 ;
  assign n4714 = ~x434 & n3359 ;
  assign n4715 = ~x306 & ~n3359 ;
  assign n4716 = ~n4714 & ~n4715 ;
  assign n4717 = ~x178 & n3730 ;
  assign n4718 = ~x50 & ~n3730 ;
  assign n4719 = ~n4717 & ~n4718 ;
  assign n4720 = ~n4716 & n4719 ;
  assign n4721 = ~n4713 & ~n4720 ;
  assign n4722 = ~n4706 & n4721 ;
  assign n4723 = n4699 & n4722 ;
  assign n4724 = ~n4668 & n4723 ;
  assign n4725 = ~n4661 & n4724 ;
  assign n4726 = ~n4671 & n4674 ;
  assign n4727 = ~n4709 & n4712 ;
  assign n4728 = ~n4713 & n4716 ;
  assign n4729 = ~n4719 & n4728 ;
  assign n4730 = n4664 & ~n4667 ;
  assign n4731 = ~n4702 & n4705 ;
  assign n4732 = ~n4730 & ~n4731 ;
  assign n4733 = n4722 & ~n4732 ;
  assign n4734 = ~n4729 & ~n4733 ;
  assign n4735 = ~n4727 & n4734 ;
  assign n4736 = n4699 & ~n4735 ;
  assign n4737 = n4693 & ~n4696 ;
  assign n4738 = ~n4690 & n4737 ;
  assign n4739 = ~n4686 & n4689 ;
  assign n4740 = ~n4738 & ~n4739 ;
  assign n4741 = n4678 & ~n4681 ;
  assign n4742 = n4740 & ~n4741 ;
  assign n4743 = n4683 & ~n4742 ;
  assign n4744 = ~n4736 & ~n4743 ;
  assign n4745 = ~n4726 & n4744 ;
  assign n4746 = ~n4725 & n4745 ;
  assign n4747 = n4156 & ~n4159 ;
  assign n4748 = ~n4153 & ~n4747 ;
  assign n4749 = n4130 & n4748 ;
  assign n4750 = n4146 & n4749 ;
  assign n4751 = ~n4746 & n4750 ;
  assign n4752 = ~n4175 & ~n4751 ;
  assign n4753 = ~n4173 & n4752 ;
  assign n4754 = ~n4168 & n4753 ;
  assign n4755 = ~n4105 & n4754 ;
  assign n4756 = ~n4098 & ~n4755 ;
  assign n4757 = ~n4091 & n4756 ;
  assign n4758 = n4084 & n4757 ;
  assign n4759 = ~n4072 & n4075 ;
  assign n4760 = n4087 & ~n4098 ;
  assign n4761 = ~n4090 & n4760 ;
  assign n4762 = ~n4094 & n4097 ;
  assign n4763 = ~n4761 & ~n4762 ;
  assign n4764 = n4079 & ~n4082 ;
  assign n4765 = n4763 & ~n4764 ;
  assign n4766 = n4084 & ~n4765 ;
  assign n4767 = ~n4759 & ~n4766 ;
  assign n4768 = ~n4758 & n4767 ;
  assign n4769 = n4059 & ~n4062 ;
  assign n4770 = ~n4056 & ~n4769 ;
  assign n4771 = n4049 & n4770 ;
  assign n4772 = ~n4768 & n4771 ;
  assign n4773 = ~n4069 & ~n4772 ;
  assign n4774 = ~n4067 & n4773 ;
  assign n4775 = ~n4040 & n4774 ;
  assign n4776 = ~x203 & n3730 ;
  assign n4777 = ~x75 & ~n3730 ;
  assign n4778 = ~n4776 & ~n4777 ;
  assign n4779 = ~x459 & n3359 ;
  assign n4780 = ~x331 & ~n3359 ;
  assign n4781 = ~n4779 & ~n4780 ;
  assign n4782 = n4778 & ~n4781 ;
  assign n4783 = ~x458 & n3359 ;
  assign n4784 = ~x330 & ~n3359 ;
  assign n4785 = ~n4783 & ~n4784 ;
  assign n4786 = ~x202 & n3730 ;
  assign n4787 = ~x74 & ~n3730 ;
  assign n4788 = ~n4786 & ~n4787 ;
  assign n4789 = ~n4785 & n4788 ;
  assign n4790 = ~n4782 & ~n4789 ;
  assign n4791 = ~x201 & n3730 ;
  assign n4792 = ~x73 & ~n3730 ;
  assign n4793 = ~n4791 & ~n4792 ;
  assign n4794 = ~x457 & n3359 ;
  assign n4795 = ~x329 & ~n3359 ;
  assign n4796 = ~n4794 & ~n4795 ;
  assign n4797 = n4793 & ~n4796 ;
  assign n4798 = ~x456 & n3359 ;
  assign n4799 = ~x328 & ~n3359 ;
  assign n4800 = ~n4798 & ~n4799 ;
  assign n4801 = ~x200 & n3730 ;
  assign n4802 = ~x72 & ~n3730 ;
  assign n4803 = ~n4801 & ~n4802 ;
  assign n4804 = ~n4800 & n4803 ;
  assign n4805 = ~n4797 & ~n4804 ;
  assign n4806 = n4790 & n4805 ;
  assign n4807 = ~n4775 & n4806 ;
  assign n4808 = ~n4778 & n4781 ;
  assign n4809 = n4800 & ~n4803 ;
  assign n4810 = ~n4797 & n4809 ;
  assign n4811 = ~n4793 & n4796 ;
  assign n4812 = ~n4810 & ~n4811 ;
  assign n4813 = n4785 & ~n4788 ;
  assign n4814 = n4812 & ~n4813 ;
  assign n4815 = n4790 & ~n4814 ;
  assign n4816 = ~n4808 & ~n4815 ;
  assign n4817 = ~n4807 & n4816 ;
  assign n4818 = n4023 & ~n4026 ;
  assign n4819 = ~n4020 & ~n4818 ;
  assign n4820 = n4013 & n4819 ;
  assign n4821 = ~n4817 & n4820 ;
  assign n4822 = ~n4033 & ~n4821 ;
  assign n4823 = ~n4031 & n4822 ;
  assign n4824 = ~n4004 & n4823 ;
  assign n4825 = ~n3997 & ~n4824 ;
  assign n4826 = n3990 & n4825 ;
  assign n4827 = ~n3975 & n4826 ;
  assign n4828 = ~n3978 & n3981 ;
  assign n4829 = n3971 & ~n3997 ;
  assign n4830 = ~n3974 & n4829 ;
  assign n4831 = ~n3993 & n3996 ;
  assign n4832 = ~n4830 & ~n4831 ;
  assign n4833 = n3985 & ~n3988 ;
  assign n4834 = n4832 & ~n4833 ;
  assign n4835 = n3990 & ~n4834 ;
  assign n4836 = ~n4828 & ~n4835 ;
  assign n4837 = ~n4827 & n4836 ;
  assign n4838 = n3958 & ~n3961 ;
  assign n4839 = ~n3955 & ~n4838 ;
  assign n4840 = n3948 & n4839 ;
  assign n4841 = ~n4837 & n4840 ;
  assign n4842 = ~n3968 & ~n4841 ;
  assign n4843 = ~n3966 & n4842 ;
  assign n4844 = ~n3939 & n4843 ;
  assign n4845 = ~x219 & n3730 ;
  assign n4846 = ~x91 & ~n3730 ;
  assign n4847 = ~n4845 & ~n4846 ;
  assign n4848 = ~x475 & n3359 ;
  assign n4849 = ~x347 & ~n3359 ;
  assign n4850 = ~n4848 & ~n4849 ;
  assign n4851 = n4847 & ~n4850 ;
  assign n4852 = ~x474 & n3359 ;
  assign n4853 = ~x346 & ~n3359 ;
  assign n4854 = ~n4852 & ~n4853 ;
  assign n4855 = ~x218 & n3730 ;
  assign n4856 = ~x90 & ~n3730 ;
  assign n4857 = ~n4855 & ~n4856 ;
  assign n4858 = ~n4854 & n4857 ;
  assign n4859 = ~n4851 & ~n4858 ;
  assign n4860 = ~x217 & n3730 ;
  assign n4861 = ~x89 & ~n3730 ;
  assign n4862 = ~n4860 & ~n4861 ;
  assign n4863 = ~x473 & n3359 ;
  assign n4864 = ~x345 & ~n3359 ;
  assign n4865 = ~n4863 & ~n4864 ;
  assign n4866 = n4862 & ~n4865 ;
  assign n4867 = ~x472 & n3359 ;
  assign n4868 = ~x344 & ~n3359 ;
  assign n4869 = ~n4867 & ~n4868 ;
  assign n4870 = ~x216 & n3730 ;
  assign n4871 = ~x88 & ~n3730 ;
  assign n4872 = ~n4870 & ~n4871 ;
  assign n4873 = ~n4869 & n4872 ;
  assign n4874 = ~n4866 & ~n4873 ;
  assign n4875 = n4859 & n4874 ;
  assign n4876 = ~n4844 & n4875 ;
  assign n4877 = ~n4847 & n4850 ;
  assign n4878 = n4869 & ~n4872 ;
  assign n4879 = ~n4866 & n4878 ;
  assign n4880 = ~n4862 & n4865 ;
  assign n4881 = ~n4879 & ~n4880 ;
  assign n4882 = n4854 & ~n4857 ;
  assign n4883 = n4881 & ~n4882 ;
  assign n4884 = n4859 & ~n4883 ;
  assign n4885 = ~n4877 & ~n4884 ;
  assign n4886 = ~n4876 & n4885 ;
  assign n4887 = n3922 & ~n3925 ;
  assign n4888 = ~n3919 & ~n4887 ;
  assign n4889 = n3912 & n4888 ;
  assign n4890 = ~n4886 & n4889 ;
  assign n4891 = ~n3932 & ~n4890 ;
  assign n4892 = ~n3930 & n4891 ;
  assign n4893 = ~n3903 & n4892 ;
  assign n4894 = ~n3896 & ~n4893 ;
  assign n4895 = n3889 & n4894 ;
  assign n4896 = ~n3874 & n4895 ;
  assign n4897 = ~n3877 & n3880 ;
  assign n4898 = n3870 & ~n3896 ;
  assign n4899 = ~n3873 & n4898 ;
  assign n4900 = ~n3892 & n3895 ;
  assign n4901 = ~n4899 & ~n4900 ;
  assign n4902 = n3884 & ~n3887 ;
  assign n4903 = n4901 & ~n4902 ;
  assign n4904 = n3889 & ~n4903 ;
  assign n4905 = ~n4897 & ~n4904 ;
  assign n4906 = ~n4896 & n4905 ;
  assign n4907 = n3857 & ~n3860 ;
  assign n4908 = ~n3854 & ~n4907 ;
  assign n4909 = n3847 & n4908 ;
  assign n4910 = ~n4906 & n4909 ;
  assign n4911 = ~n3867 & ~n4910 ;
  assign n4912 = ~n3865 & n4911 ;
  assign n4913 = ~n3838 & n4912 ;
  assign n4914 = ~x235 & n3730 ;
  assign n4915 = ~x107 & ~n3730 ;
  assign n4916 = ~n4914 & ~n4915 ;
  assign n4917 = ~x491 & n3359 ;
  assign n4918 = ~x363 & ~n3359 ;
  assign n4919 = ~n4917 & ~n4918 ;
  assign n4920 = n4916 & ~n4919 ;
  assign n4921 = ~x490 & n3359 ;
  assign n4922 = ~x362 & ~n3359 ;
  assign n4923 = ~n4921 & ~n4922 ;
  assign n4924 = ~x234 & n3730 ;
  assign n4925 = ~x106 & ~n3730 ;
  assign n4926 = ~n4924 & ~n4925 ;
  assign n4927 = ~n4923 & n4926 ;
  assign n4928 = ~n4920 & ~n4927 ;
  assign n4929 = ~x233 & n3730 ;
  assign n4930 = ~x105 & ~n3730 ;
  assign n4931 = ~n4929 & ~n4930 ;
  assign n4932 = ~x489 & n3359 ;
  assign n4933 = ~x361 & ~n3359 ;
  assign n4934 = ~n4932 & ~n4933 ;
  assign n4935 = n4931 & ~n4934 ;
  assign n4936 = ~x488 & n3359 ;
  assign n4937 = ~x360 & ~n3359 ;
  assign n4938 = ~n4936 & ~n4937 ;
  assign n4939 = ~x232 & n3730 ;
  assign n4940 = ~x104 & ~n3730 ;
  assign n4941 = ~n4939 & ~n4940 ;
  assign n4942 = ~n4938 & n4941 ;
  assign n4943 = ~n4935 & ~n4942 ;
  assign n4944 = n4928 & n4943 ;
  assign n4945 = ~n4913 & n4944 ;
  assign n4946 = ~n4916 & n4919 ;
  assign n4947 = n4938 & ~n4941 ;
  assign n4948 = ~n4935 & n4947 ;
  assign n4949 = ~n4931 & n4934 ;
  assign n4950 = ~n4948 & ~n4949 ;
  assign n4951 = n4923 & ~n4926 ;
  assign n4952 = n4950 & ~n4951 ;
  assign n4953 = n4928 & ~n4952 ;
  assign n4954 = ~n4946 & ~n4953 ;
  assign n4955 = ~n4945 & n4954 ;
  assign n4956 = n3821 & ~n3824 ;
  assign n4957 = ~n3818 & ~n4956 ;
  assign n4958 = n3811 & n4957 ;
  assign n4959 = ~n4955 & n4958 ;
  assign n4960 = ~n3831 & ~n4959 ;
  assign n4961 = ~n3829 & n4960 ;
  assign n4962 = ~n3802 & n4961 ;
  assign n4963 = ~n3795 & ~n4962 ;
  assign n4964 = n3788 & n4963 ;
  assign n4965 = ~n3773 & n4964 ;
  assign n4966 = ~n3776 & n3779 ;
  assign n4967 = n3769 & ~n3795 ;
  assign n4968 = ~n3772 & n4967 ;
  assign n4969 = ~n3791 & n3794 ;
  assign n4970 = ~n4968 & ~n4969 ;
  assign n4971 = n3783 & ~n3786 ;
  assign n4972 = n4970 & ~n4971 ;
  assign n4973 = n3788 & ~n4972 ;
  assign n4974 = ~n4966 & ~n4973 ;
  assign n4975 = ~n4965 & n4974 ;
  assign n4976 = n3749 & ~n3759 ;
  assign n4977 = ~n3756 & ~n4976 ;
  assign n4978 = n3746 & n4977 ;
  assign n4979 = ~n4975 & n4978 ;
  assign n4980 = ~n3766 & ~n4979 ;
  assign n4981 = ~n3764 & n4980 ;
  assign n4982 = ~n3737 & n4981 ;
  assign n4983 = ~x251 & n3730 ;
  assign n4984 = ~x123 & ~n3730 ;
  assign n4985 = ~n4983 & ~n4984 ;
  assign n4986 = ~x507 & n3359 ;
  assign n4987 = ~x379 & ~n3359 ;
  assign n4988 = ~n4986 & ~n4987 ;
  assign n4989 = n4985 & ~n4988 ;
  assign n4990 = ~x506 & n3359 ;
  assign n4991 = ~x378 & ~n3359 ;
  assign n4992 = ~n4990 & ~n4991 ;
  assign n4993 = ~x250 & n3730 ;
  assign n4994 = ~x122 & ~n3730 ;
  assign n4995 = ~n4993 & ~n4994 ;
  assign n4996 = ~n4992 & n4995 ;
  assign n4997 = ~n4989 & ~n4996 ;
  assign n4998 = ~x249 & n3730 ;
  assign n4999 = ~x121 & ~n3730 ;
  assign n5000 = ~n4998 & ~n4999 ;
  assign n5001 = ~x505 & n3359 ;
  assign n5002 = ~x377 & ~n3359 ;
  assign n5003 = ~n5001 & ~n5002 ;
  assign n5004 = n5000 & ~n5003 ;
  assign n5005 = ~x504 & n3359 ;
  assign n5006 = ~x376 & ~n3359 ;
  assign n5007 = ~n5005 & ~n5006 ;
  assign n5008 = ~x248 & n3730 ;
  assign n5009 = ~x120 & ~n3730 ;
  assign n5010 = ~n5008 & ~n5009 ;
  assign n5011 = ~n5007 & n5010 ;
  assign n5012 = ~n5004 & ~n5011 ;
  assign n5013 = n4997 & n5012 ;
  assign n5014 = ~n4982 & n5013 ;
  assign n5015 = ~n4985 & n4988 ;
  assign n5016 = ~n5004 & n5007 ;
  assign n5017 = ~n5010 & n5016 ;
  assign n5018 = ~n5000 & n5003 ;
  assign n5019 = ~n5017 & ~n5018 ;
  assign n5020 = n4992 & ~n4995 ;
  assign n5021 = n5019 & ~n5020 ;
  assign n5022 = n4997 & ~n5021 ;
  assign n5023 = ~n5015 & ~n5022 ;
  assign n5024 = ~n5014 & n5023 ;
  assign n5025 = ~x252 & n3730 ;
  assign n5026 = ~x124 & ~n3730 ;
  assign n5027 = ~n5025 & ~n5026 ;
  assign n5028 = ~x508 & n3359 ;
  assign n5029 = ~x380 & ~n3359 ;
  assign n5030 = ~n5028 & ~n5029 ;
  assign n5031 = n5027 & ~n5030 ;
  assign n5032 = ~n3364 & n3728 ;
  assign n5033 = ~x254 & n3730 ;
  assign n5034 = ~x126 & ~n3730 ;
  assign n5035 = ~n5033 & ~n5034 ;
  assign n5036 = ~x510 & n3359 ;
  assign n5037 = ~x382 & ~n3359 ;
  assign n5038 = ~n5036 & ~n5037 ;
  assign n5039 = n5035 & ~n5038 ;
  assign n5040 = ~x253 & n3730 ;
  assign n5041 = ~x125 & ~n3730 ;
  assign n5042 = ~n5040 & ~n5041 ;
  assign n5043 = ~x509 & n3359 ;
  assign n5044 = ~x381 & ~n3359 ;
  assign n5045 = ~n5043 & ~n5044 ;
  assign n5046 = n5042 & ~n5045 ;
  assign n5047 = ~n5039 & ~n5046 ;
  assign n5048 = ~n5032 & n5047 ;
  assign n5049 = ~n5031 & n5048 ;
  assign n5050 = ~n5024 & n5049 ;
  assign n5051 = ~n5027 & n5030 ;
  assign n5052 = ~n5042 & n5045 ;
  assign n5053 = ~n5051 & ~n5052 ;
  assign n5054 = n5047 & ~n5053 ;
  assign n5055 = ~n5035 & n5038 ;
  assign n5056 = ~n5054 & ~n5055 ;
  assign n5057 = ~n5032 & ~n5056 ;
  assign n5058 = ~n5050 & ~n5057 ;
  assign n5059 = ~n3729 & n5058 ;
  assign n5060 = ~n3362 & n5059 ;
  assign n5061 = ~n4441 & ~n5059 ;
  assign n5062 = ~n5060 & ~n5061 ;
  assign n5065 = n5062 & ~x512 ;
  assign n5066 = ~n5064 & ~n5065 ;
  assign n5067 = ~n2370 & n2991 ;
  assign n5068 = ~n2378 & ~n2991 ;
  assign n5069 = ~n5067 & ~n5068 ;
  assign n5074 = ~n5069 & x513 ;
  assign n5070 = ~n4438 & n5059 ;
  assign n5071 = ~n4446 & ~n5059 ;
  assign n5072 = ~n5070 & ~n5071 ;
  assign n5075 = n5072 & ~x513 ;
  assign n5076 = ~n5074 & ~n5075 ;
  assign n5077 = ~n2385 & n2991 ;
  assign n5078 = ~n2382 & ~n2991 ;
  assign n5079 = ~n5077 & ~n5078 ;
  assign n5084 = ~n5079 & x514 ;
  assign n5080 = ~n4453 & n5059 ;
  assign n5081 = ~n4450 & ~n5059 ;
  assign n5082 = ~n5080 & ~n5081 ;
  assign n5085 = n5082 & ~x514 ;
  assign n5086 = ~n5084 & ~n5085 ;
  assign n5087 = ~n2366 & n2991 ;
  assign n5088 = ~n2363 & ~n2991 ;
  assign n5089 = ~n5087 & ~n5088 ;
  assign n5094 = ~n5089 & x515 ;
  assign n5090 = ~n4434 & n5059 ;
  assign n5091 = ~n4431 & ~n5059 ;
  assign n5092 = ~n5090 & ~n5091 ;
  assign n5095 = n5092 & ~x515 ;
  assign n5096 = ~n5094 & ~n5095 ;
  assign n5097 = ~n2357 & n2991 ;
  assign n5098 = ~n2360 & ~n2991 ;
  assign n5099 = ~n5097 & ~n5098 ;
  assign n5104 = ~n5099 & x516 ;
  assign n5100 = ~n4425 & n5059 ;
  assign n5101 = ~n4428 & ~n5059 ;
  assign n5102 = ~n5100 & ~n5101 ;
  assign n5105 = n5102 & ~x516 ;
  assign n5106 = ~n5104 & ~n5105 ;
  assign n5107 = ~n2351 & n2991 ;
  assign n5108 = ~n2354 & ~n2991 ;
  assign n5109 = ~n5107 & ~n5108 ;
  assign n5114 = ~n5109 & x517 ;
  assign n5110 = ~n4419 & n5059 ;
  assign n5111 = ~n4422 & ~n5059 ;
  assign n5112 = ~n5110 & ~n5111 ;
  assign n5115 = n5112 & ~x517 ;
  assign n5116 = ~n5114 & ~n5115 ;
  assign n5117 = ~n2345 & n2991 ;
  assign n5118 = ~n2348 & ~n2991 ;
  assign n5119 = ~n5117 & ~n5118 ;
  assign n5124 = ~n5119 & x518 ;
  assign n5120 = ~n4413 & n5059 ;
  assign n5121 = ~n4416 & ~n5059 ;
  assign n5122 = ~n5120 & ~n5121 ;
  assign n5125 = n5122 & ~x518 ;
  assign n5126 = ~n5124 & ~n5125 ;
  assign n5127 = ~n2341 & n2991 ;
  assign n5128 = ~n2338 & ~n2991 ;
  assign n5129 = ~n5127 & ~n5128 ;
  assign n5134 = ~n5129 & x519 ;
  assign n5130 = ~n4409 & n5059 ;
  assign n5131 = ~n4406 & ~n5059 ;
  assign n5132 = ~n5130 & ~n5131 ;
  assign n5135 = n5132 & ~x519 ;
  assign n5136 = ~n5134 & ~n5135 ;
  assign n5137 = ~n2335 & n2991 ;
  assign n5138 = ~n2412 & ~n2991 ;
  assign n5139 = ~n5137 & ~n5138 ;
  assign n5144 = ~n5139 & x520 ;
  assign n5140 = ~n4403 & n5059 ;
  assign n5141 = ~n4480 & ~n5059 ;
  assign n5142 = ~n5140 & ~n5141 ;
  assign n5145 = n5142 & ~x520 ;
  assign n5146 = ~n5144 & ~n5145 ;
  assign n5147 = ~n2332 & n2991 ;
  assign n5148 = ~n2419 & ~n2991 ;
  assign n5149 = ~n5147 & ~n5148 ;
  assign n5154 = ~n5149 & x521 ;
  assign n5150 = ~n4400 & n5059 ;
  assign n5151 = ~n4487 & ~n5059 ;
  assign n5152 = ~n5150 & ~n5151 ;
  assign n5155 = n5152 & ~x521 ;
  assign n5156 = ~n5154 & ~n5155 ;
  assign n5157 = ~n2328 & n2991 ;
  assign n5158 = ~n2325 & ~n2991 ;
  assign n5159 = ~n5157 & ~n5158 ;
  assign n5164 = ~n5159 & x522 ;
  assign n5160 = ~n4396 & n5059 ;
  assign n5161 = ~n4393 & ~n5059 ;
  assign n5162 = ~n5160 & ~n5161 ;
  assign n5165 = n5162 & ~x522 ;
  assign n5166 = ~n5164 & ~n5165 ;
  assign n5167 = ~n2321 & n2991 ;
  assign n5168 = ~n2318 & ~n2991 ;
  assign n5169 = ~n5167 & ~n5168 ;
  assign n5174 = ~n5169 & x523 ;
  assign n5170 = ~n4389 & n5059 ;
  assign n5171 = ~n4386 & ~n5059 ;
  assign n5172 = ~n5170 & ~n5171 ;
  assign n5175 = n5172 & ~x523 ;
  assign n5176 = ~n5174 & ~n5175 ;
  assign n5177 = ~n2314 & n2991 ;
  assign n5178 = ~n2311 & ~n2991 ;
  assign n5179 = ~n5177 & ~n5178 ;
  assign n5184 = ~n5179 & x524 ;
  assign n5180 = ~n4382 & n5059 ;
  assign n5181 = ~n4379 & ~n5059 ;
  assign n5182 = ~n5180 & ~n5181 ;
  assign n5185 = n5182 & ~x524 ;
  assign n5186 = ~n5184 & ~n5185 ;
  assign n5187 = ~n2307 & n2991 ;
  assign n5188 = ~n2304 & ~n2991 ;
  assign n5189 = ~n5187 & ~n5188 ;
  assign n5194 = ~n5189 & x525 ;
  assign n5190 = ~n4375 & n5059 ;
  assign n5191 = ~n4372 & ~n5059 ;
  assign n5192 = ~n5190 & ~n5191 ;
  assign n5195 = n5192 & ~x525 ;
  assign n5196 = ~n5194 & ~n5195 ;
  assign n5197 = ~n2300 & n2991 ;
  assign n5198 = ~n2297 & ~n2991 ;
  assign n5199 = ~n5197 & ~n5198 ;
  assign n5204 = ~n5199 & x526 ;
  assign n5200 = ~n4368 & n5059 ;
  assign n5201 = ~n4365 & ~n5059 ;
  assign n5202 = ~n5200 & ~n5201 ;
  assign n5205 = n5202 & ~x526 ;
  assign n5206 = ~n5204 & ~n5205 ;
  assign n5207 = ~n2293 & n2991 ;
  assign n5208 = ~n2290 & ~n2991 ;
  assign n5209 = ~n5207 & ~n5208 ;
  assign n5214 = ~n5209 & x527 ;
  assign n5210 = ~n4361 & n5059 ;
  assign n5211 = ~n4358 & ~n5059 ;
  assign n5212 = ~n5210 & ~n5211 ;
  assign n5215 = n5212 & ~x527 ;
  assign n5216 = ~n5214 & ~n5215 ;
  assign n5217 = ~n2287 & n2991 ;
  assign n5218 = ~n2444 & ~n2991 ;
  assign n5219 = ~n5217 & ~n5218 ;
  assign n5224 = ~n5219 & x528 ;
  assign n5220 = ~n4355 & n5059 ;
  assign n5221 = ~n4512 & ~n5059 ;
  assign n5222 = ~n5220 & ~n5221 ;
  assign n5225 = n5222 & ~x528 ;
  assign n5226 = ~n5224 & ~n5225 ;
  assign n5227 = ~n2284 & n2991 ;
  assign n5228 = ~n2451 & ~n2991 ;
  assign n5229 = ~n5227 & ~n5228 ;
  assign n5234 = ~n5229 & x529 ;
  assign n5230 = ~n4352 & n5059 ;
  assign n5231 = ~n4519 & ~n5059 ;
  assign n5232 = ~n5230 & ~n5231 ;
  assign n5235 = n5232 & ~x529 ;
  assign n5236 = ~n5234 & ~n5235 ;
  assign n5237 = ~n2280 & n2991 ;
  assign n5238 = ~n2277 & ~n2991 ;
  assign n5239 = ~n5237 & ~n5238 ;
  assign n5244 = ~n5239 & x530 ;
  assign n5240 = ~n4348 & n5059 ;
  assign n5241 = ~n4345 & ~n5059 ;
  assign n5242 = ~n5240 & ~n5241 ;
  assign n5245 = n5242 & ~x530 ;
  assign n5246 = ~n5244 & ~n5245 ;
  assign n5247 = ~n2273 & n2991 ;
  assign n5248 = ~n2270 & ~n2991 ;
  assign n5249 = ~n5247 & ~n5248 ;
  assign n5254 = ~n5249 & x531 ;
  assign n5250 = ~n4341 & n5059 ;
  assign n5251 = ~n4338 & ~n5059 ;
  assign n5252 = ~n5250 & ~n5251 ;
  assign n5255 = n5252 & ~x531 ;
  assign n5256 = ~n5254 & ~n5255 ;
  assign n5257 = ~n2266 & n2991 ;
  assign n5258 = ~n2263 & ~n2991 ;
  assign n5259 = ~n5257 & ~n5258 ;
  assign n5264 = ~n5259 & x532 ;
  assign n5260 = ~n4334 & n5059 ;
  assign n5261 = ~n4331 & ~n5059 ;
  assign n5262 = ~n5260 & ~n5261 ;
  assign n5265 = n5262 & ~x532 ;
  assign n5266 = ~n5264 & ~n5265 ;
  assign n5267 = ~n2259 & n2991 ;
  assign n5268 = ~n2256 & ~n2991 ;
  assign n5269 = ~n5267 & ~n5268 ;
  assign n5274 = ~n5269 & x533 ;
  assign n5270 = ~n4327 & n5059 ;
  assign n5271 = ~n4324 & ~n5059 ;
  assign n5272 = ~n5270 & ~n5271 ;
  assign n5275 = n5272 & ~x533 ;
  assign n5276 = ~n5274 & ~n5275 ;
  assign n5277 = ~n2252 & n2991 ;
  assign n5278 = ~n2249 & ~n2991 ;
  assign n5279 = ~n5277 & ~n5278 ;
  assign n5284 = ~n5279 & x534 ;
  assign n5280 = ~n4320 & n5059 ;
  assign n5281 = ~n4317 & ~n5059 ;
  assign n5282 = ~n5280 & ~n5281 ;
  assign n5285 = n5282 & ~x534 ;
  assign n5286 = ~n5284 & ~n5285 ;
  assign n5287 = ~n2245 & n2991 ;
  assign n5288 = ~n2242 & ~n2991 ;
  assign n5289 = ~n5287 & ~n5288 ;
  assign n5294 = ~n5289 & x535 ;
  assign n5290 = ~n4313 & n5059 ;
  assign n5291 = ~n4310 & ~n5059 ;
  assign n5292 = ~n5290 & ~n5291 ;
  assign n5295 = n5292 & ~x535 ;
  assign n5296 = ~n5294 & ~n5295 ;
  assign n5297 = ~n2239 & n2991 ;
  assign n5298 = ~n2476 & ~n2991 ;
  assign n5299 = ~n5297 & ~n5298 ;
  assign n5304 = ~n5299 & x536 ;
  assign n5300 = ~n4307 & n5059 ;
  assign n5301 = ~n4544 & ~n5059 ;
  assign n5302 = ~n5300 & ~n5301 ;
  assign n5305 = n5302 & ~x536 ;
  assign n5306 = ~n5304 & ~n5305 ;
  assign n5307 = ~n2236 & n2991 ;
  assign n5308 = ~n2483 & ~n2991 ;
  assign n5309 = ~n5307 & ~n5308 ;
  assign n5314 = ~n5309 & x537 ;
  assign n5310 = ~n4304 & n5059 ;
  assign n5311 = ~n4551 & ~n5059 ;
  assign n5312 = ~n5310 & ~n5311 ;
  assign n5315 = n5312 & ~x537 ;
  assign n5316 = ~n5314 & ~n5315 ;
  assign n5317 = ~n2232 & n2991 ;
  assign n5318 = ~n2229 & ~n2991 ;
  assign n5319 = ~n5317 & ~n5318 ;
  assign n5324 = ~n5319 & x538 ;
  assign n5320 = ~n4300 & n5059 ;
  assign n5321 = ~n4297 & ~n5059 ;
  assign n5322 = ~n5320 & ~n5321 ;
  assign n5325 = n5322 & ~x538 ;
  assign n5326 = ~n5324 & ~n5325 ;
  assign n5327 = ~n2225 & n2991 ;
  assign n5328 = ~n2222 & ~n2991 ;
  assign n5329 = ~n5327 & ~n5328 ;
  assign n5334 = ~n5329 & x539 ;
  assign n5330 = ~n4293 & n5059 ;
  assign n5331 = ~n4290 & ~n5059 ;
  assign n5332 = ~n5330 & ~n5331 ;
  assign n5335 = n5332 & ~x539 ;
  assign n5336 = ~n5334 & ~n5335 ;
  assign n5337 = ~n2218 & n2991 ;
  assign n5338 = ~n2215 & ~n2991 ;
  assign n5339 = ~n5337 & ~n5338 ;
  assign n5344 = ~n5339 & x540 ;
  assign n5340 = ~n4286 & n5059 ;
  assign n5341 = ~n4283 & ~n5059 ;
  assign n5342 = ~n5340 & ~n5341 ;
  assign n5345 = n5342 & ~x540 ;
  assign n5346 = ~n5344 & ~n5345 ;
  assign n5347 = ~n2211 & n2991 ;
  assign n5348 = ~n2208 & ~n2991 ;
  assign n5349 = ~n5347 & ~n5348 ;
  assign n5354 = ~n5349 & x541 ;
  assign n5350 = ~n4279 & n5059 ;
  assign n5351 = ~n4276 & ~n5059 ;
  assign n5352 = ~n5350 & ~n5351 ;
  assign n5355 = n5352 & ~x541 ;
  assign n5356 = ~n5354 & ~n5355 ;
  assign n5357 = ~n2204 & n2991 ;
  assign n5358 = ~n2201 & ~n2991 ;
  assign n5359 = ~n5357 & ~n5358 ;
  assign n5364 = ~n5359 & x542 ;
  assign n5360 = ~n4272 & n5059 ;
  assign n5361 = ~n4269 & ~n5059 ;
  assign n5362 = ~n5360 & ~n5361 ;
  assign n5365 = n5362 & ~x542 ;
  assign n5366 = ~n5364 & ~n5365 ;
  assign n5367 = ~n2197 & n2991 ;
  assign n5368 = ~n2194 & ~n2991 ;
  assign n5369 = ~n5367 & ~n5368 ;
  assign n5374 = ~n5369 & x543 ;
  assign n5370 = ~n4265 & n5059 ;
  assign n5371 = ~n4262 & ~n5059 ;
  assign n5372 = ~n5370 & ~n5371 ;
  assign n5375 = n5372 & ~x543 ;
  assign n5376 = ~n5374 & ~n5375 ;
  assign n5377 = ~n2187 & n2991 ;
  assign n5378 = ~n2190 & ~n2991 ;
  assign n5379 = ~n5377 & ~n5378 ;
  assign n5384 = ~n5379 & x544 ;
  assign n5380 = ~n4255 & n5059 ;
  assign n5381 = ~n4258 & ~n5059 ;
  assign n5382 = ~n5380 & ~n5381 ;
  assign n5385 = n5382 & ~x544 ;
  assign n5386 = ~n5384 & ~n5385 ;
  assign n5387 = ~n2542 & n2991 ;
  assign n5388 = ~n2539 & ~n2991 ;
  assign n5389 = ~n5387 & ~n5388 ;
  assign n5394 = ~n5389 & x545 ;
  assign n5390 = ~n4610 & n5059 ;
  assign n5391 = ~n4607 & ~n5059 ;
  assign n5392 = ~n5390 & ~n5391 ;
  assign n5395 = n5392 & ~x545 ;
  assign n5396 = ~n5394 & ~n5395 ;
  assign n5397 = ~n2553 & n2991 ;
  assign n5398 = ~n2556 & ~n2991 ;
  assign n5399 = ~n5397 & ~n5398 ;
  assign n5404 = ~n5399 & x546 ;
  assign n5400 = ~n4621 & n5059 ;
  assign n5401 = ~n4624 & ~n5059 ;
  assign n5402 = ~n5400 & ~n5401 ;
  assign n5405 = n5402 & ~x546 ;
  assign n5406 = ~n5404 & ~n5405 ;
  assign n5407 = ~n2549 & n2991 ;
  assign n5408 = ~n2546 & ~n2991 ;
  assign n5409 = ~n5407 & ~n5408 ;
  assign n5414 = ~n5409 & x547 ;
  assign n5410 = ~n4617 & n5059 ;
  assign n5411 = ~n4614 & ~n5059 ;
  assign n5412 = ~n5410 & ~n5411 ;
  assign n5415 = n5412 & ~x547 ;
  assign n5416 = ~n5414 & ~n5415 ;
  assign n5417 = ~n2526 & n2991 ;
  assign n5418 = ~n2523 & ~n2991 ;
  assign n5419 = ~n5417 & ~n5418 ;
  assign n5424 = ~n5419 & x548 ;
  assign n5420 = ~n4594 & n5059 ;
  assign n5421 = ~n4591 & ~n5059 ;
  assign n5422 = ~n5420 & ~n5421 ;
  assign n5425 = n5422 & ~x548 ;
  assign n5426 = ~n5424 & ~n5425 ;
  assign n5427 = ~n2533 & n2991 ;
  assign n5428 = ~n2530 & ~n2991 ;
  assign n5429 = ~n5427 & ~n5428 ;
  assign n5434 = ~n5429 & x549 ;
  assign n5430 = ~n4601 & n5059 ;
  assign n5431 = ~n4598 & ~n5059 ;
  assign n5432 = ~n5430 & ~n5431 ;
  assign n5435 = n5432 & ~x549 ;
  assign n5436 = ~n5434 & ~n5435 ;
  assign n5437 = ~n2515 & n2991 ;
  assign n5438 = ~n2518 & ~n2991 ;
  assign n5439 = ~n5437 & ~n5438 ;
  assign n5444 = ~n5439 & x550 ;
  assign n5440 = ~n4583 & n5059 ;
  assign n5441 = ~n4586 & ~n5059 ;
  assign n5442 = ~n5440 & ~n5441 ;
  assign n5445 = n5442 & ~x550 ;
  assign n5446 = ~n5444 & ~n5445 ;
  assign n5447 = ~n2511 & n2991 ;
  assign n5448 = ~n2508 & ~n2991 ;
  assign n5449 = ~n5447 & ~n5448 ;
  assign n5454 = ~n5449 & x551 ;
  assign n5450 = ~n4579 & n5059 ;
  assign n5451 = ~n4576 & ~n5059 ;
  assign n5452 = ~n5450 & ~n5451 ;
  assign n5455 = n5452 & ~x551 ;
  assign n5456 = ~n5454 & ~n5455 ;
  assign n5457 = ~n2168 & n2991 ;
  assign n5458 = ~n2165 & ~n2991 ;
  assign n5459 = ~n5457 & ~n5458 ;
  assign n5464 = ~n5459 & x552 ;
  assign n5460 = ~n4236 & n5059 ;
  assign n5461 = ~n4233 & ~n5059 ;
  assign n5462 = ~n5460 & ~n5461 ;
  assign n5465 = n5462 & ~x552 ;
  assign n5466 = ~n5464 & ~n5465 ;
  assign n5467 = ~n2161 & n2991 ;
  assign n5468 = ~n2158 & ~n2991 ;
  assign n5469 = ~n5467 & ~n5468 ;
  assign n5474 = ~n5469 & x553 ;
  assign n5470 = ~n4229 & n5059 ;
  assign n5471 = ~n4226 & ~n5059 ;
  assign n5472 = ~n5470 & ~n5471 ;
  assign n5475 = n5472 & ~x553 ;
  assign n5476 = ~n5474 & ~n5475 ;
  assign n5477 = ~n2153 & n2991 ;
  assign n5478 = ~n2150 & ~n2991 ;
  assign n5479 = ~n5477 & ~n5478 ;
  assign n5484 = ~n5479 & x554 ;
  assign n5480 = ~n4221 & n5059 ;
  assign n5481 = ~n4218 & ~n5059 ;
  assign n5482 = ~n5480 & ~n5481 ;
  assign n5485 = n5482 & ~x554 ;
  assign n5486 = ~n5484 & ~n5485 ;
  assign n5487 = ~n2145 & n2991 ;
  assign n5488 = ~n2142 & ~n2991 ;
  assign n5489 = ~n5487 & ~n5488 ;
  assign n5494 = ~n5489 & x555 ;
  assign n5490 = ~n4213 & n5059 ;
  assign n5491 = ~n4210 & ~n5059 ;
  assign n5492 = ~n5490 & ~n5491 ;
  assign n5495 = n5492 & ~x555 ;
  assign n5496 = ~n5494 & ~n5495 ;
  assign n5497 = ~n2129 & n2991 ;
  assign n5498 = ~n2126 & ~n2991 ;
  assign n5499 = ~n5497 & ~n5498 ;
  assign n5504 = ~n5499 & x556 ;
  assign n5500 = ~n4197 & n5059 ;
  assign n5501 = ~n4194 & ~n5059 ;
  assign n5502 = ~n5500 & ~n5501 ;
  assign n5505 = n5502 & ~x556 ;
  assign n5506 = ~n5504 & ~n5505 ;
  assign n5507 = ~n2136 & n2991 ;
  assign n5508 = ~n2133 & ~n2991 ;
  assign n5509 = ~n5507 & ~n5508 ;
  assign n5514 = ~n5509 & x557 ;
  assign n5510 = ~n4204 & n5059 ;
  assign n5511 = ~n4201 & ~n5059 ;
  assign n5512 = ~n5510 & ~n5511 ;
  assign n5515 = n5512 & ~x557 ;
  assign n5516 = ~n5514 & ~n5515 ;
  assign n5517 = ~n2118 & n2991 ;
  assign n5518 = ~n2121 & ~n2991 ;
  assign n5519 = ~n5517 & ~n5518 ;
  assign n5524 = ~n5519 & x558 ;
  assign n5520 = ~n4186 & n5059 ;
  assign n5521 = ~n4189 & ~n5059 ;
  assign n5522 = ~n5520 & ~n5521 ;
  assign n5525 = n5522 & ~x558 ;
  assign n5526 = ~n5524 & ~n5525 ;
  assign n5527 = ~n2113 & n2991 ;
  assign n5528 = ~n2110 & ~n2991 ;
  assign n5529 = ~n5527 & ~n5528 ;
  assign n5534 = ~n5529 & x559 ;
  assign n5530 = ~n4181 & n5059 ;
  assign n5531 = ~n4178 & ~n5059 ;
  assign n5532 = ~n5530 & ~n5531 ;
  assign n5535 = n5532 & ~x559 ;
  assign n5536 = ~n5534 & ~n5535 ;
  assign n5537 = ~n2596 & n2991 ;
  assign n5538 = ~n2599 & ~n2991 ;
  assign n5539 = ~n5537 & ~n5538 ;
  assign n5544 = ~n5539 & x560 ;
  assign n5540 = ~n4664 & n5059 ;
  assign n5541 = ~n4667 & ~n5059 ;
  assign n5542 = ~n5540 & ~n5541 ;
  assign n5545 = n5542 & ~x560 ;
  assign n5546 = ~n5544 & ~n5545 ;
  assign n5547 = ~n2637 & n2991 ;
  assign n5548 = ~n2634 & ~n2991 ;
  assign n5549 = ~n5547 & ~n5548 ;
  assign n5554 = ~n5549 & x561 ;
  assign n5550 = ~n4705 & n5059 ;
  assign n5551 = ~n4702 & ~n5059 ;
  assign n5552 = ~n5550 & ~n5551 ;
  assign n5555 = n5552 & ~x561 ;
  assign n5556 = ~n5554 & ~n5555 ;
  assign n5557 = ~n2648 & n2991 ;
  assign n5558 = ~n2651 & ~n2991 ;
  assign n5559 = ~n5557 & ~n5558 ;
  assign n5564 = ~n5559 & x562 ;
  assign n5560 = ~n4716 & n5059 ;
  assign n5561 = ~n4719 & ~n5059 ;
  assign n5562 = ~n5560 & ~n5561 ;
  assign n5565 = n5562 & ~x562 ;
  assign n5566 = ~n5564 & ~n5565 ;
  assign n5567 = ~n2644 & n2991 ;
  assign n5568 = ~n2641 & ~n2991 ;
  assign n5569 = ~n5567 & ~n5568 ;
  assign n5574 = ~n5569 & x563 ;
  assign n5570 = ~n4712 & n5059 ;
  assign n5571 = ~n4709 & ~n5059 ;
  assign n5572 = ~n5570 & ~n5571 ;
  assign n5575 = n5572 & ~x563 ;
  assign n5576 = ~n5574 & ~n5575 ;
  assign n5577 = ~n2625 & n2991 ;
  assign n5578 = ~n2628 & ~n2991 ;
  assign n5579 = ~n5577 & ~n5578 ;
  assign n5584 = ~n5579 & x564 ;
  assign n5580 = ~n4693 & n5059 ;
  assign n5581 = ~n4696 & ~n5059 ;
  assign n5582 = ~n5580 & ~n5581 ;
  assign n5585 = n5582 & ~x564 ;
  assign n5586 = ~n5584 & ~n5585 ;
  assign n5587 = ~n2621 & n2991 ;
  assign n5588 = ~n2618 & ~n2991 ;
  assign n5589 = ~n5587 & ~n5588 ;
  assign n5594 = ~n5589 & x565 ;
  assign n5590 = ~n4689 & n5059 ;
  assign n5591 = ~n4686 & ~n5059 ;
  assign n5592 = ~n5590 & ~n5591 ;
  assign n5595 = n5592 & ~x565 ;
  assign n5596 = ~n5594 & ~n5595 ;
  assign n5597 = ~n2610 & n2991 ;
  assign n5598 = ~n2613 & ~n2991 ;
  assign n5599 = ~n5597 & ~n5598 ;
  assign n5604 = ~n5599 & x566 ;
  assign n5600 = ~n4678 & n5059 ;
  assign n5601 = ~n4681 & ~n5059 ;
  assign n5602 = ~n5600 & ~n5601 ;
  assign n5605 = n5602 & ~x566 ;
  assign n5606 = ~n5604 & ~n5605 ;
  assign n5607 = ~n2606 & n2991 ;
  assign n5608 = ~n2603 & ~n2991 ;
  assign n5609 = ~n5607 & ~n5608 ;
  assign n5614 = ~n5609 & x567 ;
  assign n5610 = ~n4674 & n5059 ;
  assign n5611 = ~n4671 & ~n5059 ;
  assign n5612 = ~n5610 & ~n5611 ;
  assign n5615 = n5612 & ~x567 ;
  assign n5616 = ~n5614 & ~n5615 ;
  assign n5617 = ~n2091 & n2991 ;
  assign n5618 = ~n2088 & ~n2991 ;
  assign n5619 = ~n5617 & ~n5618 ;
  assign n5624 = ~n5619 & x568 ;
  assign n5620 = ~n4159 & n5059 ;
  assign n5621 = ~n4156 & ~n5059 ;
  assign n5622 = ~n5620 & ~n5621 ;
  assign n5625 = n5622 & ~x568 ;
  assign n5626 = ~n5624 & ~n5625 ;
  assign n5627 = ~n2084 & n2991 ;
  assign n5628 = ~n2081 & ~n2991 ;
  assign n5629 = ~n5627 & ~n5628 ;
  assign n5634 = ~n5629 & x569 ;
  assign n5630 = ~n4152 & n5059 ;
  assign n5631 = ~n4149 & ~n5059 ;
  assign n5632 = ~n5630 & ~n5631 ;
  assign n5635 = n5632 & ~x569 ;
  assign n5636 = ~n5634 & ~n5635 ;
  assign n5637 = ~n2076 & n2991 ;
  assign n5638 = ~n2073 & ~n2991 ;
  assign n5639 = ~n5637 & ~n5638 ;
  assign n5644 = ~n5639 & x570 ;
  assign n5640 = ~n4144 & n5059 ;
  assign n5641 = ~n4141 & ~n5059 ;
  assign n5642 = ~n5640 & ~n5641 ;
  assign n5645 = n5642 & ~x570 ;
  assign n5646 = ~n5644 & ~n5645 ;
  assign n5647 = ~n2068 & n2991 ;
  assign n5648 = ~n2065 & ~n2991 ;
  assign n5649 = ~n5647 & ~n5648 ;
  assign n5654 = ~n5649 & x571 ;
  assign n5650 = ~n4136 & n5059 ;
  assign n5651 = ~n4133 & ~n5059 ;
  assign n5652 = ~n5650 & ~n5651 ;
  assign n5655 = n5652 & ~x571 ;
  assign n5656 = ~n5654 & ~n5655 ;
  assign n5657 = ~n2052 & n2991 ;
  assign n5658 = ~n2049 & ~n2991 ;
  assign n5659 = ~n5657 & ~n5658 ;
  assign n5664 = ~n5659 & x572 ;
  assign n5660 = ~n4120 & n5059 ;
  assign n5661 = ~n4117 & ~n5059 ;
  assign n5662 = ~n5660 & ~n5661 ;
  assign n5665 = n5662 & ~x572 ;
  assign n5666 = ~n5664 & ~n5665 ;
  assign n5667 = ~n2059 & n2991 ;
  assign n5668 = ~n2056 & ~n2991 ;
  assign n5669 = ~n5667 & ~n5668 ;
  assign n5674 = ~n5669 & x573 ;
  assign n5670 = ~n4127 & n5059 ;
  assign n5671 = ~n4124 & ~n5059 ;
  assign n5672 = ~n5670 & ~n5671 ;
  assign n5675 = n5672 & ~x573 ;
  assign n5676 = ~n5674 & ~n5675 ;
  assign n5677 = ~n2041 & n2991 ;
  assign n5678 = ~n2044 & ~n2991 ;
  assign n5679 = ~n5677 & ~n5678 ;
  assign n5684 = ~n5679 & x574 ;
  assign n5680 = ~n4109 & n5059 ;
  assign n5681 = ~n4112 & ~n5059 ;
  assign n5682 = ~n5680 & ~n5681 ;
  assign n5685 = n5682 & ~x574 ;
  assign n5686 = ~n5684 & ~n5685 ;
  assign n5687 = ~n2036 & n2991 ;
  assign n5688 = ~n2033 & ~n2991 ;
  assign n5689 = ~n5687 & ~n5688 ;
  assign n5694 = ~n5689 & x575 ;
  assign n5690 = ~n4104 & n5059 ;
  assign n5691 = ~n4101 & ~n5059 ;
  assign n5692 = ~n5690 & ~n5691 ;
  assign n5695 = n5692 & ~x575 ;
  assign n5696 = ~n5694 & ~n5695 ;
  assign n5697 = ~n2019 & n2991 ;
  assign n5698 = ~n2022 & ~n2991 ;
  assign n5699 = ~n5697 & ~n5698 ;
  assign n5704 = ~n5699 & x576 ;
  assign n5700 = ~n4087 & n5059 ;
  assign n5701 = ~n4090 & ~n5059 ;
  assign n5702 = ~n5700 & ~n5701 ;
  assign n5705 = n5702 & ~x576 ;
  assign n5706 = ~n5704 & ~n5705 ;
  assign n5707 = ~n2029 & n2991 ;
  assign n5708 = ~n2026 & ~n2991 ;
  assign n5709 = ~n5707 & ~n5708 ;
  assign n5714 = ~n5709 & x577 ;
  assign n5710 = ~n4097 & n5059 ;
  assign n5711 = ~n4094 & ~n5059 ;
  assign n5712 = ~n5710 & ~n5711 ;
  assign n5715 = n5712 & ~x577 ;
  assign n5716 = ~n5714 & ~n5715 ;
  assign n5717 = ~n2011 & n2991 ;
  assign n5718 = ~n2014 & ~n2991 ;
  assign n5719 = ~n5717 & ~n5718 ;
  assign n5724 = ~n5719 & x578 ;
  assign n5720 = ~n4079 & n5059 ;
  assign n5721 = ~n4082 & ~n5059 ;
  assign n5722 = ~n5720 & ~n5721 ;
  assign n5725 = n5722 & ~x578 ;
  assign n5726 = ~n5724 & ~n5725 ;
  assign n5727 = ~n2007 & n2991 ;
  assign n5728 = ~n2004 & ~n2991 ;
  assign n5729 = ~n5727 & ~n5728 ;
  assign n5734 = ~n5729 & x579 ;
  assign n5730 = ~n4075 & n5059 ;
  assign n5731 = ~n4072 & ~n5059 ;
  assign n5732 = ~n5730 & ~n5731 ;
  assign n5735 = n5732 & ~x579 ;
  assign n5736 = ~n5734 & ~n5735 ;
  assign n5737 = ~n1994 & n2991 ;
  assign n5738 = ~n1991 & ~n2991 ;
  assign n5739 = ~n5737 & ~n5738 ;
  assign n5744 = ~n5739 & x580 ;
  assign n5740 = ~n4062 & n5059 ;
  assign n5741 = ~n4059 & ~n5059 ;
  assign n5742 = ~n5740 & ~n5741 ;
  assign n5745 = n5742 & ~x580 ;
  assign n5746 = ~n5744 & ~n5745 ;
  assign n5747 = ~n1987 & n2991 ;
  assign n5748 = ~n1984 & ~n2991 ;
  assign n5749 = ~n5747 & ~n5748 ;
  assign n5754 = ~n5749 & x581 ;
  assign n5750 = ~n4055 & n5059 ;
  assign n5751 = ~n4052 & ~n5059 ;
  assign n5752 = ~n5750 & ~n5751 ;
  assign n5755 = n5752 & ~x581 ;
  assign n5756 = ~n5754 & ~n5755 ;
  assign n5757 = ~n1976 & n2991 ;
  assign n5758 = ~n1979 & ~n2991 ;
  assign n5759 = ~n5757 & ~n5758 ;
  assign n5764 = ~n5759 & x582 ;
  assign n5760 = ~n4044 & n5059 ;
  assign n5761 = ~n4047 & ~n5059 ;
  assign n5762 = ~n5760 & ~n5761 ;
  assign n5765 = n5762 & ~x582 ;
  assign n5766 = ~n5764 & ~n5765 ;
  assign n5767 = ~n1971 & n2991 ;
  assign n5768 = ~n1968 & ~n2991 ;
  assign n5769 = ~n5767 & ~n5768 ;
  assign n5774 = ~n5769 & x583 ;
  assign n5770 = ~n4039 & n5059 ;
  assign n5771 = ~n4036 & ~n5059 ;
  assign n5772 = ~n5770 & ~n5771 ;
  assign n5775 = n5772 & ~x583 ;
  assign n5776 = ~n5774 & ~n5775 ;
  assign n5777 = ~n2732 & n2991 ;
  assign n5778 = ~n2735 & ~n2991 ;
  assign n5779 = ~n5777 & ~n5778 ;
  assign n5784 = ~n5779 & x584 ;
  assign n5780 = ~n4800 & n5059 ;
  assign n5781 = ~n4803 & ~n5059 ;
  assign n5782 = ~n5780 & ~n5781 ;
  assign n5785 = n5782 & ~x584 ;
  assign n5786 = ~n5784 & ~n5785 ;
  assign n5787 = ~n2728 & n2991 ;
  assign n5788 = ~n2725 & ~n2991 ;
  assign n5789 = ~n5787 & ~n5788 ;
  assign n5794 = ~n5789 & x585 ;
  assign n5790 = ~n4796 & n5059 ;
  assign n5791 = ~n4793 & ~n5059 ;
  assign n5792 = ~n5790 & ~n5791 ;
  assign n5795 = n5792 & ~x585 ;
  assign n5796 = ~n5794 & ~n5795 ;
  assign n5797 = ~n2717 & n2991 ;
  assign n5798 = ~n2720 & ~n2991 ;
  assign n5799 = ~n5797 & ~n5798 ;
  assign n5804 = ~n5799 & x586 ;
  assign n5800 = ~n4785 & n5059 ;
  assign n5801 = ~n4788 & ~n5059 ;
  assign n5802 = ~n5800 & ~n5801 ;
  assign n5805 = n5802 & ~x586 ;
  assign n5806 = ~n5804 & ~n5805 ;
  assign n5807 = ~n2713 & n2991 ;
  assign n5808 = ~n2710 & ~n2991 ;
  assign n5809 = ~n5807 & ~n5808 ;
  assign n5814 = ~n5809 & x587 ;
  assign n5810 = ~n4781 & n5059 ;
  assign n5811 = ~n4778 & ~n5059 ;
  assign n5812 = ~n5810 & ~n5811 ;
  assign n5815 = n5812 & ~x587 ;
  assign n5816 = ~n5814 & ~n5815 ;
  assign n5817 = ~n1958 & n2991 ;
  assign n5818 = ~n1955 & ~n2991 ;
  assign n5819 = ~n5817 & ~n5818 ;
  assign n5824 = ~n5819 & x588 ;
  assign n5820 = ~n4026 & n5059 ;
  assign n5821 = ~n4023 & ~n5059 ;
  assign n5822 = ~n5820 & ~n5821 ;
  assign n5825 = n5822 & ~x588 ;
  assign n5826 = ~n5824 & ~n5825 ;
  assign n5827 = ~n1951 & n2991 ;
  assign n5828 = ~n1948 & ~n2991 ;
  assign n5829 = ~n5827 & ~n5828 ;
  assign n5834 = ~n5829 & x589 ;
  assign n5830 = ~n4019 & n5059 ;
  assign n5831 = ~n4016 & ~n5059 ;
  assign n5832 = ~n5830 & ~n5831 ;
  assign n5835 = n5832 & ~x589 ;
  assign n5836 = ~n5834 & ~n5835 ;
  assign n5837 = ~n1940 & n2991 ;
  assign n5838 = ~n1943 & ~n2991 ;
  assign n5839 = ~n5837 & ~n5838 ;
  assign n5844 = ~n5839 & x590 ;
  assign n5840 = ~n4008 & n5059 ;
  assign n5841 = ~n4011 & ~n5059 ;
  assign n5842 = ~n5840 & ~n5841 ;
  assign n5845 = n5842 & ~x590 ;
  assign n5846 = ~n5844 & ~n5845 ;
  assign n5847 = ~n1935 & n2991 ;
  assign n5848 = ~n1932 & ~n2991 ;
  assign n5849 = ~n5847 & ~n5848 ;
  assign n5854 = ~n5849 & x591 ;
  assign n5850 = ~n4003 & n5059 ;
  assign n5851 = ~n4000 & ~n5059 ;
  assign n5852 = ~n5850 & ~n5851 ;
  assign n5855 = n5852 & ~x591 ;
  assign n5856 = ~n5854 & ~n5855 ;
  assign n5857 = ~n1903 & n2991 ;
  assign n5858 = ~n1906 & ~n2991 ;
  assign n5859 = ~n5857 & ~n5858 ;
  assign n5864 = ~n5859 & x592 ;
  assign n5860 = ~n3971 & n5059 ;
  assign n5861 = ~n3974 & ~n5059 ;
  assign n5862 = ~n5860 & ~n5861 ;
  assign n5865 = n5862 & ~x592 ;
  assign n5866 = ~n5864 & ~n5865 ;
  assign n5867 = ~n1928 & n2991 ;
  assign n5868 = ~n1925 & ~n2991 ;
  assign n5869 = ~n5867 & ~n5868 ;
  assign n5874 = ~n5869 & x593 ;
  assign n5870 = ~n3996 & n5059 ;
  assign n5871 = ~n3993 & ~n5059 ;
  assign n5872 = ~n5870 & ~n5871 ;
  assign n5875 = n5872 & ~x593 ;
  assign n5876 = ~n5874 & ~n5875 ;
  assign n5877 = ~n1917 & n2991 ;
  assign n5878 = ~n1920 & ~n2991 ;
  assign n5879 = ~n5877 & ~n5878 ;
  assign n5884 = ~n5879 & x594 ;
  assign n5880 = ~n3985 & n5059 ;
  assign n5881 = ~n3988 & ~n5059 ;
  assign n5882 = ~n5880 & ~n5881 ;
  assign n5885 = n5882 & ~x594 ;
  assign n5886 = ~n5884 & ~n5885 ;
  assign n5887 = ~n1913 & n2991 ;
  assign n5888 = ~n1910 & ~n2991 ;
  assign n5889 = ~n5887 & ~n5888 ;
  assign n5894 = ~n5889 & x595 ;
  assign n5890 = ~n3981 & n5059 ;
  assign n5891 = ~n3978 & ~n5059 ;
  assign n5892 = ~n5890 & ~n5891 ;
  assign n5895 = n5892 & ~x595 ;
  assign n5896 = ~n5894 & ~n5895 ;
  assign n5897 = ~n1893 & n2991 ;
  assign n5898 = ~n1890 & ~n2991 ;
  assign n5899 = ~n5897 & ~n5898 ;
  assign n5904 = ~n5899 & x596 ;
  assign n5900 = ~n3961 & n5059 ;
  assign n5901 = ~n3958 & ~n5059 ;
  assign n5902 = ~n5900 & ~n5901 ;
  assign n5905 = n5902 & ~x596 ;
  assign n5906 = ~n5904 & ~n5905 ;
  assign n5907 = ~n1886 & n2991 ;
  assign n5908 = ~n1883 & ~n2991 ;
  assign n5909 = ~n5907 & ~n5908 ;
  assign n5914 = ~n5909 & x597 ;
  assign n5910 = ~n3954 & n5059 ;
  assign n5911 = ~n3951 & ~n5059 ;
  assign n5912 = ~n5910 & ~n5911 ;
  assign n5915 = n5912 & ~x597 ;
  assign n5916 = ~n5914 & ~n5915 ;
  assign n5917 = ~n1875 & n2991 ;
  assign n5918 = ~n1878 & ~n2991 ;
  assign n5919 = ~n5917 & ~n5918 ;
  assign n5924 = ~n5919 & x598 ;
  assign n5920 = ~n3943 & n5059 ;
  assign n5921 = ~n3946 & ~n5059 ;
  assign n5922 = ~n5920 & ~n5921 ;
  assign n5925 = n5922 & ~x598 ;
  assign n5926 = ~n5924 & ~n5925 ;
  assign n5927 = ~n1870 & n2991 ;
  assign n5928 = ~n1867 & ~n2991 ;
  assign n5929 = ~n5927 & ~n5928 ;
  assign n5934 = ~n5929 & x599 ;
  assign n5930 = ~n3938 & n5059 ;
  assign n5931 = ~n3935 & ~n5059 ;
  assign n5932 = ~n5930 & ~n5931 ;
  assign n5935 = n5932 & ~x599 ;
  assign n5936 = ~n5934 & ~n5935 ;
  assign n5937 = ~n2801 & n2991 ;
  assign n5938 = ~n2804 & ~n2991 ;
  assign n5939 = ~n5937 & ~n5938 ;
  assign n5944 = ~n5939 & x600 ;
  assign n5940 = ~n4869 & n5059 ;
  assign n5941 = ~n4872 & ~n5059 ;
  assign n5942 = ~n5940 & ~n5941 ;
  assign n5945 = n5942 & ~x600 ;
  assign n5946 = ~n5944 & ~n5945 ;
  assign n5947 = ~n2797 & n2991 ;
  assign n5948 = ~n2794 & ~n2991 ;
  assign n5949 = ~n5947 & ~n5948 ;
  assign n5954 = ~n5949 & x601 ;
  assign n5950 = ~n4865 & n5059 ;
  assign n5951 = ~n4862 & ~n5059 ;
  assign n5952 = ~n5950 & ~n5951 ;
  assign n5955 = n5952 & ~x601 ;
  assign n5956 = ~n5954 & ~n5955 ;
  assign n5957 = ~n2786 & n2991 ;
  assign n5958 = ~n2789 & ~n2991 ;
  assign n5959 = ~n5957 & ~n5958 ;
  assign n5964 = ~n5959 & x602 ;
  assign n5960 = ~n4854 & n5059 ;
  assign n5961 = ~n4857 & ~n5059 ;
  assign n5962 = ~n5960 & ~n5961 ;
  assign n5965 = n5962 & ~x602 ;
  assign n5966 = ~n5964 & ~n5965 ;
  assign n5967 = ~n2782 & n2991 ;
  assign n5968 = ~n2779 & ~n2991 ;
  assign n5969 = ~n5967 & ~n5968 ;
  assign n5974 = ~n5969 & x603 ;
  assign n5970 = ~n4850 & n5059 ;
  assign n5971 = ~n4847 & ~n5059 ;
  assign n5972 = ~n5970 & ~n5971 ;
  assign n5975 = n5972 & ~x603 ;
  assign n5976 = ~n5974 & ~n5975 ;
  assign n5977 = ~n1857 & n2991 ;
  assign n5978 = ~n1854 & ~n2991 ;
  assign n5979 = ~n5977 & ~n5978 ;
  assign n5984 = ~n5979 & x604 ;
  assign n5980 = ~n3925 & n5059 ;
  assign n5981 = ~n3922 & ~n5059 ;
  assign n5982 = ~n5980 & ~n5981 ;
  assign n5985 = n5982 & ~x604 ;
  assign n5986 = ~n5984 & ~n5985 ;
  assign n5987 = ~n1850 & n2991 ;
  assign n5988 = ~n1847 & ~n2991 ;
  assign n5989 = ~n5987 & ~n5988 ;
  assign n5994 = ~n5989 & x605 ;
  assign n5990 = ~n3918 & n5059 ;
  assign n5991 = ~n3915 & ~n5059 ;
  assign n5992 = ~n5990 & ~n5991 ;
  assign n5995 = n5992 & ~x605 ;
  assign n5996 = ~n5994 & ~n5995 ;
  assign n5997 = ~n1839 & n2991 ;
  assign n5998 = ~n1842 & ~n2991 ;
  assign n5999 = ~n5997 & ~n5998 ;
  assign n6004 = ~n5999 & x606 ;
  assign n6000 = ~n3907 & n5059 ;
  assign n6001 = ~n3910 & ~n5059 ;
  assign n6002 = ~n6000 & ~n6001 ;
  assign n6005 = n6002 & ~x606 ;
  assign n6006 = ~n6004 & ~n6005 ;
  assign n6007 = ~n1834 & n2991 ;
  assign n6008 = ~n1831 & ~n2991 ;
  assign n6009 = ~n6007 & ~n6008 ;
  assign n6014 = ~n6009 & x607 ;
  assign n6010 = ~n3902 & n5059 ;
  assign n6011 = ~n3899 & ~n5059 ;
  assign n6012 = ~n6010 & ~n6011 ;
  assign n6015 = n6012 & ~x607 ;
  assign n6016 = ~n6014 & ~n6015 ;
  assign n6017 = ~n1802 & n2991 ;
  assign n6018 = ~n1805 & ~n2991 ;
  assign n6019 = ~n6017 & ~n6018 ;
  assign n6024 = ~n6019 & x608 ;
  assign n6020 = ~n3870 & n5059 ;
  assign n6021 = ~n3873 & ~n5059 ;
  assign n6022 = ~n6020 & ~n6021 ;
  assign n6025 = n6022 & ~x608 ;
  assign n6026 = ~n6024 & ~n6025 ;
  assign n6027 = ~n1827 & n2991 ;
  assign n6028 = ~n1824 & ~n2991 ;
  assign n6029 = ~n6027 & ~n6028 ;
  assign n6034 = ~n6029 & x609 ;
  assign n6030 = ~n3895 & n5059 ;
  assign n6031 = ~n3892 & ~n5059 ;
  assign n6032 = ~n6030 & ~n6031 ;
  assign n6035 = n6032 & ~x609 ;
  assign n6036 = ~n6034 & ~n6035 ;
  assign n6037 = ~n1816 & n2991 ;
  assign n6038 = ~n1819 & ~n2991 ;
  assign n6039 = ~n6037 & ~n6038 ;
  assign n6044 = ~n6039 & x610 ;
  assign n6040 = ~n3884 & n5059 ;
  assign n6041 = ~n3887 & ~n5059 ;
  assign n6042 = ~n6040 & ~n6041 ;
  assign n6045 = n6042 & ~x610 ;
  assign n6046 = ~n6044 & ~n6045 ;
  assign n6047 = ~n1812 & n2991 ;
  assign n6048 = ~n1809 & ~n2991 ;
  assign n6049 = ~n6047 & ~n6048 ;
  assign n6054 = ~n6049 & x611 ;
  assign n6050 = ~n3880 & n5059 ;
  assign n6051 = ~n3877 & ~n5059 ;
  assign n6052 = ~n6050 & ~n6051 ;
  assign n6055 = n6052 & ~x611 ;
  assign n6056 = ~n6054 & ~n6055 ;
  assign n6057 = ~n1792 & n2991 ;
  assign n6058 = ~n1789 & ~n2991 ;
  assign n6059 = ~n6057 & ~n6058 ;
  assign n6064 = ~n6059 & x612 ;
  assign n6060 = ~n3860 & n5059 ;
  assign n6061 = ~n3857 & ~n5059 ;
  assign n6062 = ~n6060 & ~n6061 ;
  assign n6065 = n6062 & ~x612 ;
  assign n6066 = ~n6064 & ~n6065 ;
  assign n6067 = ~n1785 & n2991 ;
  assign n6068 = ~n1782 & ~n2991 ;
  assign n6069 = ~n6067 & ~n6068 ;
  assign n6074 = ~n6069 & x613 ;
  assign n6070 = ~n3853 & n5059 ;
  assign n6071 = ~n3850 & ~n5059 ;
  assign n6072 = ~n6070 & ~n6071 ;
  assign n6075 = n6072 & ~x613 ;
  assign n6076 = ~n6074 & ~n6075 ;
  assign n6077 = ~n1774 & n2991 ;
  assign n6078 = ~n1777 & ~n2991 ;
  assign n6079 = ~n6077 & ~n6078 ;
  assign n6084 = ~n6079 & x614 ;
  assign n6080 = ~n3842 & n5059 ;
  assign n6081 = ~n3845 & ~n5059 ;
  assign n6082 = ~n6080 & ~n6081 ;
  assign n6085 = n6082 & ~x614 ;
  assign n6086 = ~n6084 & ~n6085 ;
  assign n6087 = ~n1769 & n2991 ;
  assign n6088 = ~n1766 & ~n2991 ;
  assign n6089 = ~n6087 & ~n6088 ;
  assign n6094 = ~n6089 & x615 ;
  assign n6090 = ~n3837 & n5059 ;
  assign n6091 = ~n3834 & ~n5059 ;
  assign n6092 = ~n6090 & ~n6091 ;
  assign n6095 = n6092 & ~x615 ;
  assign n6096 = ~n6094 & ~n6095 ;
  assign n6097 = ~n2870 & n2991 ;
  assign n6098 = ~n2873 & ~n2991 ;
  assign n6099 = ~n6097 & ~n6098 ;
  assign n6104 = ~n6099 & x616 ;
  assign n6100 = ~n4938 & n5059 ;
  assign n6101 = ~n4941 & ~n5059 ;
  assign n6102 = ~n6100 & ~n6101 ;
  assign n6105 = n6102 & ~x616 ;
  assign n6106 = ~n6104 & ~n6105 ;
  assign n6107 = ~n2866 & n2991 ;
  assign n6108 = ~n2863 & ~n2991 ;
  assign n6109 = ~n6107 & ~n6108 ;
  assign n6114 = ~n6109 & x617 ;
  assign n6110 = ~n4934 & n5059 ;
  assign n6111 = ~n4931 & ~n5059 ;
  assign n6112 = ~n6110 & ~n6111 ;
  assign n6115 = n6112 & ~x617 ;
  assign n6116 = ~n6114 & ~n6115 ;
  assign n6117 = ~n2855 & n2991 ;
  assign n6118 = ~n2858 & ~n2991 ;
  assign n6119 = ~n6117 & ~n6118 ;
  assign n6124 = ~n6119 & x618 ;
  assign n6120 = ~n4923 & n5059 ;
  assign n6121 = ~n4926 & ~n5059 ;
  assign n6122 = ~n6120 & ~n6121 ;
  assign n6125 = n6122 & ~x618 ;
  assign n6126 = ~n6124 & ~n6125 ;
  assign n6127 = ~n2851 & n2991 ;
  assign n6128 = ~n2848 & ~n2991 ;
  assign n6129 = ~n6127 & ~n6128 ;
  assign n6134 = ~n6129 & x619 ;
  assign n6130 = ~n4919 & n5059 ;
  assign n6131 = ~n4916 & ~n5059 ;
  assign n6132 = ~n6130 & ~n6131 ;
  assign n6135 = n6132 & ~x619 ;
  assign n6136 = ~n6134 & ~n6135 ;
  assign n6137 = ~n1756 & n2991 ;
  assign n6138 = ~n1753 & ~n2991 ;
  assign n6139 = ~n6137 & ~n6138 ;
  assign n6144 = ~n6139 & x620 ;
  assign n6140 = ~n3824 & n5059 ;
  assign n6141 = ~n3821 & ~n5059 ;
  assign n6142 = ~n6140 & ~n6141 ;
  assign n6145 = n6142 & ~x620 ;
  assign n6146 = ~n6144 & ~n6145 ;
  assign n6147 = ~n1749 & n2991 ;
  assign n6148 = ~n1746 & ~n2991 ;
  assign n6149 = ~n6147 & ~n6148 ;
  assign n6154 = ~n6149 & x621 ;
  assign n6150 = ~n3817 & n5059 ;
  assign n6151 = ~n3814 & ~n5059 ;
  assign n6152 = ~n6150 & ~n6151 ;
  assign n6155 = n6152 & ~x621 ;
  assign n6156 = ~n6154 & ~n6155 ;
  assign n6157 = ~n1738 & n2991 ;
  assign n6158 = ~n1741 & ~n2991 ;
  assign n6159 = ~n6157 & ~n6158 ;
  assign n6164 = ~n6159 & x622 ;
  assign n6160 = ~n3806 & n5059 ;
  assign n6161 = ~n3809 & ~n5059 ;
  assign n6162 = ~n6160 & ~n6161 ;
  assign n6165 = n6162 & ~x622 ;
  assign n6166 = ~n6164 & ~n6165 ;
  assign n6167 = ~n1733 & n2991 ;
  assign n6168 = ~n1730 & ~n2991 ;
  assign n6169 = ~n6167 & ~n6168 ;
  assign n6174 = ~n6169 & x623 ;
  assign n6170 = ~n3801 & n5059 ;
  assign n6171 = ~n3798 & ~n5059 ;
  assign n6172 = ~n6170 & ~n6171 ;
  assign n6175 = n6172 & ~x623 ;
  assign n6176 = ~n6174 & ~n6175 ;
  assign n6177 = ~n1701 & n2991 ;
  assign n6178 = ~n1704 & ~n2991 ;
  assign n6179 = ~n6177 & ~n6178 ;
  assign n6184 = ~n6179 & x624 ;
  assign n6180 = ~n3769 & n5059 ;
  assign n6181 = ~n3772 & ~n5059 ;
  assign n6182 = ~n6180 & ~n6181 ;
  assign n6185 = n6182 & ~x624 ;
  assign n6186 = ~n6184 & ~n6185 ;
  assign n6187 = ~n1726 & n2991 ;
  assign n6188 = ~n1723 & ~n2991 ;
  assign n6189 = ~n6187 & ~n6188 ;
  assign n6194 = ~n6189 & x625 ;
  assign n6190 = ~n3794 & n5059 ;
  assign n6191 = ~n3791 & ~n5059 ;
  assign n6192 = ~n6190 & ~n6191 ;
  assign n6195 = n6192 & ~x625 ;
  assign n6196 = ~n6194 & ~n6195 ;
  assign n6197 = ~n1715 & n2991 ;
  assign n6198 = ~n1718 & ~n2991 ;
  assign n6199 = ~n6197 & ~n6198 ;
  assign n6204 = ~n6199 & x626 ;
  assign n6200 = ~n3783 & n5059 ;
  assign n6201 = ~n3786 & ~n5059 ;
  assign n6202 = ~n6200 & ~n6201 ;
  assign n6205 = n6202 & ~x626 ;
  assign n6206 = ~n6204 & ~n6205 ;
  assign n6207 = ~n1711 & n2991 ;
  assign n6208 = ~n1708 & ~n2991 ;
  assign n6209 = ~n6207 & ~n6208 ;
  assign n6214 = ~n6209 & x627 ;
  assign n6210 = ~n3779 & n5059 ;
  assign n6211 = ~n3776 & ~n5059 ;
  assign n6212 = ~n6210 & ~n6211 ;
  assign n6215 = n6212 & ~x627 ;
  assign n6216 = ~n6214 & ~n6215 ;
  assign n6217 = ~n1691 & n2991 ;
  assign n6218 = ~n1681 & ~n2991 ;
  assign n6219 = ~n6217 & ~n6218 ;
  assign n6224 = ~n6219 & x628 ;
  assign n6220 = ~n3759 & n5059 ;
  assign n6221 = ~n3749 & ~n5059 ;
  assign n6222 = ~n6220 & ~n6221 ;
  assign n6225 = n6222 & ~x628 ;
  assign n6226 = ~n6224 & ~n6225 ;
  assign n6227 = ~n1687 & n2991 ;
  assign n6228 = ~n1684 & ~n2991 ;
  assign n6229 = ~n6227 & ~n6228 ;
  assign n6234 = ~n6229 & x629 ;
  assign n6230 = ~n3755 & n5059 ;
  assign n6231 = ~n3752 & ~n5059 ;
  assign n6232 = ~n6230 & ~n6231 ;
  assign n6235 = n6232 & ~x629 ;
  assign n6236 = ~n6234 & ~n6235 ;
  assign n6237 = ~n1673 & n2991 ;
  assign n6238 = ~n1676 & ~n2991 ;
  assign n6239 = ~n6237 & ~n6238 ;
  assign n6244 = ~n6239 & x630 ;
  assign n6240 = ~n3741 & n5059 ;
  assign n6241 = ~n3744 & ~n5059 ;
  assign n6242 = ~n6240 & ~n6241 ;
  assign n6245 = n6242 & ~x630 ;
  assign n6246 = ~n6244 & ~n6245 ;
  assign n6247 = ~n1668 & n2991 ;
  assign n6248 = ~n1665 & ~n2991 ;
  assign n6249 = ~n6247 & ~n6248 ;
  assign n6254 = ~n6249 & x631 ;
  assign n6250 = ~n3736 & n5059 ;
  assign n6251 = ~n3733 & ~n5059 ;
  assign n6252 = ~n6250 & ~n6251 ;
  assign n6255 = n6252 & ~x631 ;
  assign n6256 = ~n6254 & ~n6255 ;
  assign n6257 = ~n2939 & n2991 ;
  assign n6258 = ~n2942 & ~n2991 ;
  assign n6259 = ~n6257 & ~n6258 ;
  assign n6264 = ~n6259 & x632 ;
  assign n6260 = ~n5007 & n5059 ;
  assign n6261 = ~n5010 & ~n5059 ;
  assign n6262 = ~n6260 & ~n6261 ;
  assign n6265 = n6262 & ~x632 ;
  assign n6266 = ~n6264 & ~n6265 ;
  assign n6267 = ~n2935 & n2991 ;
  assign n6268 = ~n2932 & ~n2991 ;
  assign n6269 = ~n6267 & ~n6268 ;
  assign n6274 = ~n6269 & x633 ;
  assign n6270 = ~n5003 & n5059 ;
  assign n6271 = ~n5000 & ~n5059 ;
  assign n6272 = ~n6270 & ~n6271 ;
  assign n6275 = n6272 & ~x633 ;
  assign n6276 = ~n6274 & ~n6275 ;
  assign n6277 = ~n2924 & n2991 ;
  assign n6278 = ~n2927 & ~n2991 ;
  assign n6279 = ~n6277 & ~n6278 ;
  assign n6284 = ~n6279 & x634 ;
  assign n6280 = ~n4992 & n5059 ;
  assign n6281 = ~n4995 & ~n5059 ;
  assign n6282 = ~n6280 & ~n6281 ;
  assign n6285 = n6282 & ~x634 ;
  assign n6286 = ~n6284 & ~n6285 ;
  assign n6287 = ~n2920 & n2991 ;
  assign n6288 = ~n2917 & ~n2991 ;
  assign n6289 = ~n6287 & ~n6288 ;
  assign n6294 = ~n6289 & x635 ;
  assign n6290 = ~n4988 & n5059 ;
  assign n6291 = ~n4985 & ~n5059 ;
  assign n6292 = ~n6290 & ~n6291 ;
  assign n6295 = n6292 & ~x635 ;
  assign n6296 = ~n6294 & ~n6295 ;
  assign n6297 = ~n2962 & n2991 ;
  assign n6298 = ~n2959 & ~n2991 ;
  assign n6299 = ~n6297 & ~n6298 ;
  assign n6304 = ~n6299 & x636 ;
  assign n6300 = ~n5030 & n5059 ;
  assign n6301 = ~n5027 & ~n5059 ;
  assign n6302 = ~n6300 & ~n6301 ;
  assign n6305 = n6302 & ~x636 ;
  assign n6306 = ~n6304 & ~n6305 ;
  assign n6307 = ~n2977 & n2991 ;
  assign n6308 = ~n2974 & ~n2991 ;
  assign n6309 = ~n6307 & ~n6308 ;
  assign n6314 = ~n6309 & x637 ;
  assign n6310 = ~n5045 & n5059 ;
  assign n6311 = ~n5042 & ~n5059 ;
  assign n6312 = ~n6310 & ~n6311 ;
  assign n6315 = n6312 & ~x637 ;
  assign n6316 = ~n6314 & ~n6315 ;
  assign n6317 = ~n2970 & n2991 ;
  assign n6318 = ~n2967 & ~n2991 ;
  assign n6319 = ~n6317 & ~n6318 ;
  assign n6324 = ~n6319 & x638 ;
  assign n6320 = ~n5038 & n5059 ;
  assign n6321 = ~n5035 & ~n5059 ;
  assign n6322 = ~n6320 & ~n6321 ;
  assign n6325 = n6322 & ~x638 ;
  assign n6326 = ~n6324 & ~n6325 ;
  assign n6327 = ~n1088 & n2990 ;
  assign n6328 = n1659 & ~n6327 ;
  assign n6332 = n6328 & x639 ;
  assign n6329 = ~n3364 & n5058 ;
  assign n6330 = n3728 & ~n6329 ;
  assign n6333 = ~n6330 & ~x639 ;
  assign n6334 = ~n6332 & ~n6333 ;
  assign n6335 = n1083 & n2991 ;
  assign n6336 = n1662 & ~n2991 ;
  assign n6337 = ~n6335 & ~n6336 ;
  assign n6342 = ~n6337 & x640 ;
  assign n6338 = n3359 & n5059 ;
  assign n6339 = n3730 & ~n5059 ;
  assign n6340 = ~n6338 & ~n6339 ;
  assign n6343 = n6340 & ~x640 ;
  assign n6344 = ~n6342 & ~n6343 ;
  assign n6346 = n2991 & x641 ;
  assign n6347 = ~n5059 & ~x641 ;
  assign n6348 = ~n6346 & ~n6347 ;
  assign y0 = ~n5066 ;
  assign y1 = ~n5076 ;
  assign y2 = ~n5086 ;
  assign y3 = ~n5096 ;
  assign y4 = ~n5106 ;
  assign y5 = ~n5116 ;
  assign y6 = ~n5126 ;
  assign y7 = ~n5136 ;
  assign y8 = ~n5146 ;
  assign y9 = ~n5156 ;
  assign y10 = ~n5166 ;
  assign y11 = ~n5176 ;
  assign y12 = ~n5186 ;
  assign y13 = ~n5196 ;
  assign y14 = ~n5206 ;
  assign y15 = ~n5216 ;
  assign y16 = ~n5226 ;
  assign y17 = ~n5236 ;
  assign y18 = ~n5246 ;
  assign y19 = ~n5256 ;
  assign y20 = ~n5266 ;
  assign y21 = ~n5276 ;
  assign y22 = ~n5286 ;
  assign y23 = ~n5296 ;
  assign y24 = ~n5306 ;
  assign y25 = ~n5316 ;
  assign y26 = ~n5326 ;
  assign y27 = ~n5336 ;
  assign y28 = ~n5346 ;
  assign y29 = ~n5356 ;
  assign y30 = ~n5366 ;
  assign y31 = ~n5376 ;
  assign y32 = ~n5386 ;
  assign y33 = ~n5396 ;
  assign y34 = ~n5406 ;
  assign y35 = ~n5416 ;
  assign y36 = ~n5426 ;
  assign y37 = ~n5436 ;
  assign y38 = ~n5446 ;
  assign y39 = ~n5456 ;
  assign y40 = ~n5466 ;
  assign y41 = ~n5476 ;
  assign y42 = ~n5486 ;
  assign y43 = ~n5496 ;
  assign y44 = ~n5506 ;
  assign y45 = ~n5516 ;
  assign y46 = ~n5526 ;
  assign y47 = ~n5536 ;
  assign y48 = ~n5546 ;
  assign y49 = ~n5556 ;
  assign y50 = ~n5566 ;
  assign y51 = ~n5576 ;
  assign y52 = ~n5586 ;
  assign y53 = ~n5596 ;
  assign y54 = ~n5606 ;
  assign y55 = ~n5616 ;
  assign y56 = ~n5626 ;
  assign y57 = ~n5636 ;
  assign y58 = ~n5646 ;
  assign y59 = ~n5656 ;
  assign y60 = ~n5666 ;
  assign y61 = ~n5676 ;
  assign y62 = ~n5686 ;
  assign y63 = ~n5696 ;
  assign y64 = ~n5706 ;
  assign y65 = ~n5716 ;
  assign y66 = ~n5726 ;
  assign y67 = ~n5736 ;
  assign y68 = ~n5746 ;
  assign y69 = ~n5756 ;
  assign y70 = ~n5766 ;
  assign y71 = ~n5776 ;
  assign y72 = ~n5786 ;
  assign y73 = ~n5796 ;
  assign y74 = ~n5806 ;
  assign y75 = ~n5816 ;
  assign y76 = ~n5826 ;
  assign y77 = ~n5836 ;
  assign y78 = ~n5846 ;
  assign y79 = ~n5856 ;
  assign y80 = ~n5866 ;
  assign y81 = ~n5876 ;
  assign y82 = ~n5886 ;
  assign y83 = ~n5896 ;
  assign y84 = ~n5906 ;
  assign y85 = ~n5916 ;
  assign y86 = ~n5926 ;
  assign y87 = ~n5936 ;
  assign y88 = ~n5946 ;
  assign y89 = ~n5956 ;
  assign y90 = ~n5966 ;
  assign y91 = ~n5976 ;
  assign y92 = ~n5986 ;
  assign y93 = ~n5996 ;
  assign y94 = ~n6006 ;
  assign y95 = ~n6016 ;
  assign y96 = ~n6026 ;
  assign y97 = ~n6036 ;
  assign y98 = ~n6046 ;
  assign y99 = ~n6056 ;
  assign y100 = ~n6066 ;
  assign y101 = ~n6076 ;
  assign y102 = ~n6086 ;
  assign y103 = ~n6096 ;
  assign y104 = ~n6106 ;
  assign y105 = ~n6116 ;
  assign y106 = ~n6126 ;
  assign y107 = ~n6136 ;
  assign y108 = ~n6146 ;
  assign y109 = ~n6156 ;
  assign y110 = ~n6166 ;
  assign y111 = ~n6176 ;
  assign y112 = ~n6186 ;
  assign y113 = ~n6196 ;
  assign y114 = ~n6206 ;
  assign y115 = ~n6216 ;
  assign y116 = ~n6226 ;
  assign y117 = ~n6236 ;
  assign y118 = ~n6246 ;
  assign y119 = ~n6256 ;
  assign y120 = ~n6266 ;
  assign y121 = ~n6276 ;
  assign y122 = ~n6286 ;
  assign y123 = ~n6296 ;
  assign y124 = ~n6306 ;
  assign y125 = ~n6316 ;
  assign y126 = ~n6326 ;
  assign y127 = ~n6334 ;
  assign y128 = ~n6344 ;
  assign y129 = ~n6348 ;
endmodule
