module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , n46236 , n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , n46643 , n46644 , n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , n46674 , n46675 , n46676 , n46677 , n46678 , n46680 , n46681 , n46682 , n46683 , n46684 , n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , n46711 , n46712 , n46713 , n46714 , n46715 , n46716 , n46717 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , n46725 , n46726 , n46727 , n46728 , n46729 , n46730 , n46731 , n46732 , n46733 , n46734 , n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , n46751 , n46752 , n46753 , n46754 , n46755 , n46756 , n46757 , n46758 , n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , n46765 , n46766 , n46767 , n46768 , n46769 , n46770 , n46771 , n46772 , n46773 , n46774 , n46775 , n46776 , n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , n46785 , n46786 , n46787 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , n46795 , n46796 , n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , n46805 , n46806 , n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , n46815 , n46816 , n46817 , n46818 , n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , n46835 , n46836 , n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , n46845 , n46846 , n46847 , n46848 , n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , n46855 , n46856 , n46857 , n46858 , n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , n46865 , n46866 , n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , n46895 , n46896 , n46897 , n46898 , n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , n46905 , n46906 , n46907 , n46908 , n46909 , n46910 , n46911 , n46912 , n46913 , n46914 , n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , n46924 , n46925 , n46926 , n46927 , n46928 , n46929 , n46930 , n46931 , n46932 , n46933 , n46934 , n46935 , n46936 , n46937 , n46938 , n46939 , n46940 , n46941 , n46942 , n46943 , n46944 , n46945 , n46946 , n46947 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , n46954 , n46955 , n46956 , n46957 , n46958 , n46959 , n46960 , n46961 , n46962 , n46963 , n46964 , n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , n46974 , n46975 , n46976 , n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , n46985 , n46986 , n46987 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , n46995 , n46996 , n46997 , n46998 , n46999 , n47000 , n47001 , n47002 , n47003 , n47004 , n47005 , n47006 , n47007 , n47008 , n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , n47015 , n47016 , n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , n47025 , n47026 , n47027 , n47028 , n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , n47035 , n47036 , n47037 , n47038 , n47039 , n47040 , n47041 , n47042 , n47043 , n47044 , n47045 , n47046 , n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n47053 , n47054 , n47055 , n47056 , n47057 , n47058 , n47059 , n47060 , n47061 , n47062 , n47063 , n47064 , n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , n47071 , n47072 , n47073 , n47074 , n47075 , n47076 , n47077 , n47078 , n47079 , n47080 , n47081 , n47082 , n47083 , n47084 , n47085 , n47086 , n47087 , n47088 , n47089 , n47090 , n47091 , n47092 , n47093 , n47094 , n47095 , n47096 , n47097 , n47098 , n47099 , n47100 , n47101 , n47102 , n47103 , n47104 , n47105 , n47106 , n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n47113 , n47114 , n47116 , n47117 , n47118 , n47119 , n47120 , n47121 , n47122 , n47123 , n47124 , n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , n47131 , n47132 , n47133 , n47134 , n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , n47141 , n47142 , n47143 , n47144 , n47145 , n47146 , n47147 , n47148 , n47149 , n47150 , n47151 , n47152 , n47153 , n47154 , n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n47163 , n47164 , n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , n47185 , n47186 , n47187 , n47188 , n47189 , n47190 , n47191 , n47192 , n47193 , n47194 , n47195 , n47196 , n47197 , n47198 , n47199 , n47200 , n47201 , n47202 , n47203 , n47204 , n47205 , n47206 , n47207 , n47208 , n47209 , n47210 , n47211 , n47212 , n47213 , n47214 , n47215 , n47216 , n47217 , n47218 , n47219 , n47220 , n47221 , n47222 , n47223 , n47224 , n47225 , n47226 , n47227 , n47228 , n47229 , n47230 , n47231 , n47232 , n47233 , n47234 , n47235 , n47236 , n47237 , n47238 , n47239 , n47240 , n47241 , n47242 , n47243 , n47244 , n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , n47251 , n47252 , n47253 , n47254 , n47255 , n47256 , n47257 , n47258 , n47259 , n47260 , n47261 , n47262 , n47263 , n47264 , n47265 , n47266 , n47267 , n47268 , n47269 , n47270 , n47271 , n47272 , n47273 , n47274 , n47275 , n47276 , n47277 , n47278 , n47279 , n47280 , n47281 , n47282 , n47283 , n47284 , n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , n47291 , n47292 , n47293 , n47294 , n47295 , n47296 , n47297 , n47298 , n47299 , n47300 , n47301 , n47302 , n47303 , n47304 , n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , n47325 , n47326 , n47327 , n47328 , n47329 , n47330 , n47331 , n47332 , n47333 , n47334 , n47335 , n47336 , n47337 , n47338 , n47339 , n47340 , n47341 , n47342 , n47343 , n47344 , n47345 , n47346 , n47347 , n47348 , n47349 , n47350 , n47351 , n47352 , n47353 , n47354 , n47355 , n47356 , n47357 , n47358 , n47359 , n47360 , n47361 , n47362 , n47363 , n47364 , n47365 , n47366 , n47367 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , n47375 , n47376 , n47377 , n47378 , n47379 , n47380 , n47381 , n47382 , n47383 , n47384 , n47385 , n47386 , n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n47393 , n47394 , n47395 , n47396 , n47397 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , n47404 , n47405 , n47406 , n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , n47414 , n47415 , n47416 , n47417 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , n47424 , n47425 , n47426 , n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , n47435 , n47436 , n47437 , n47438 , n47439 , n47440 , n47441 , n47442 , n47443 , n47444 , n47445 , n47446 , n47447 , n47448 , n47449 , n47450 , n47451 , n47452 , n47453 , n47454 , n47455 , n47456 , n47457 , n47458 , n47459 , n47460 , n47461 , n47462 , n47463 , n47464 , n47465 , n47466 , n47467 , n47468 , n47469 , n47470 , n47471 , n47472 , n47473 , n47474 , n47475 , n47476 , n47477 , n47478 , n47479 , n47480 , n47481 , n47482 , n47483 , n47484 , n47485 , n47486 , n47487 , n47488 , n47489 , n47490 , n47491 , n47492 , n47493 , n47494 , n47495 , n47496 , n47497 , n47498 , n47499 , n47500 , n47501 , n47502 , n47503 , n47504 , n47505 , n47506 , n47507 , n47508 , n47509 , n47510 , n47511 , n47512 , n47513 , n47514 , n47515 , n47516 , n47517 , n47518 , n47519 , n47520 , n47521 , n47522 , n47523 , n47524 , n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , n47536 , n47537 , n47538 , n47539 , n47540 , n47541 , n47542 , n47543 , n47544 , n47545 , n47546 , n47547 , n47548 , n47549 , n47550 , n47551 , n47552 , n47553 , n47554 , n47555 , n47556 , n47557 , n47558 , n47559 , n47560 , n47561 , n47562 , n47563 , n47564 , n47565 , n47566 , n47567 , n47568 , n47569 , n47570 , n47571 , n47572 , n47573 , n47574 , n47575 , n47576 , n47577 , n47578 , n47579 , n47580 , n47581 , n47582 , n47583 , n47584 , n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , n47591 , n47592 , n47593 , n47594 , n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , n47601 , n47602 , n47603 , n47604 , n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , n47611 , n47612 , n47613 , n47614 , n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , n47621 , n47622 , n47623 , n47624 , n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , n47641 , n47642 , n47643 , n47644 , n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , n47651 , n47652 , n47653 , n47654 , n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , n47661 , n47662 , n47663 , n47664 , n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , n47671 , n47672 , n47673 , n47674 , n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , n47691 , n47692 , n47693 , n47694 , n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , n47701 , n47702 , n47703 , n47704 , n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , n47711 , n47712 , n47713 , n47714 , n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , n47721 , n47722 , n47723 , n47724 , n47725 , n47726 , n47727 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , n47734 , n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , n47741 , n47742 , n47743 , n47744 , n47745 , n47746 , n47747 , n47748 , n47749 , n47750 , n47751 , n47752 , n47753 , n47754 , n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , n47765 , n47766 , n47767 , n47768 , n47769 , n47770 , n47771 , n47772 , n47773 , n47774 , n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , n47791 , n47792 , n47793 , n47794 , n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , n47801 , n47802 , n47803 , n47804 , n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , n47811 , n47812 , n47813 , n47814 , n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , n47821 , n47822 , n47823 , n47824 , n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , n47831 , n47832 , n47833 , n47834 , n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n47843 , n47844 , n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , n47861 , n47862 , n47863 , n47864 , n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , n47871 , n47872 , n47873 , n47874 , n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , n47881 , n47882 , n47883 , n47884 , n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , n47891 , n47892 , n47893 , n47894 , n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , n47901 , n47902 , n47903 , n47904 , n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , n47911 , n47912 , n47913 , n47914 , n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , n47921 , n47922 , n47923 , n47924 , n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , n47931 , n47932 , n47933 , n47934 , n47935 , n47936 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , n47944 , n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , n47951 , n47952 , n47953 , n47954 , n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , n47981 , n47982 , n47983 , n47984 , n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , n47991 , n47992 , n47993 , n47994 , n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , n48001 , n48002 , n48003 , n48004 , n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , n48011 , n48012 , n48013 , n48014 , n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , n48021 , n48022 , n48023 , n48024 , n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , n48031 , n48032 , n48033 , n48034 , n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n48043 , n48044 , n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , n48051 , n48052 , n48053 , n48054 , n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , n48061 , n48062 , n48063 , n48064 , n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , n48071 , n48072 , n48073 , n48074 , n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , n48081 , n48082 , n48083 , n48084 , n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , n48101 , n48102 , n48103 , n48104 , n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , n48111 , n48112 , n48113 , n48114 , n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , n48121 , n48122 , n48123 , n48124 , n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , n48134 , n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , n48141 , n48142 , n48143 , n48144 , n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , n48151 , n48152 , n48153 , n48154 , n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , n48161 , n48162 , n48163 , n48164 , n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , n48191 , n48192 , n48193 , n48194 , n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , n48204 , n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n48213 , n48214 , n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , n48221 , n48222 , n48223 , n48224 , n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , n48231 , n48232 , n48233 , n48234 , n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , n48241 , n48242 , n48243 , n48244 , n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , n48251 , n48252 , n48253 , n48254 , n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , n48261 , n48262 , n48263 , n48264 , n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , n48271 , n48272 , n48273 , n48274 , n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , n48281 , n48282 , n48283 , n48284 , n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , n48291 , n48292 , n48293 , n48294 , n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , n48301 , n48302 , n48303 , n48304 , n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n48313 , n48314 , n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n48323 , n48324 , n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , n48331 , n48332 , n48334 , n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , n48341 , n48342 , n48343 , n48344 , n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , n48351 , n48352 , n48353 , n48354 , n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , n48361 , n48362 , n48363 , n48364 , n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , n48371 , n48372 , n48373 , n48374 , n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , n48381 , n48382 , n48383 , n48384 , n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , n48394 , n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , n48401 , n48402 , n48403 , n48404 , n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , n48411 , n48412 , n48413 , n48414 , n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , n48421 , n48422 , n48423 , n48424 , n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n48433 , n48434 , n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , n48441 , n48442 , n48443 , n48444 , n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48453 , n48454 , n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , n48461 , n48462 , n48463 , n48464 , n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , n48471 , n48472 , n48473 , n48474 , n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n48493 , n48494 , n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , n48501 , n48502 , n48503 , n48504 , n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , n48511 , n48512 , n48513 , n48514 , n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , n48521 , n48522 , n48523 , n48524 , n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , n48531 , n48532 , n48533 , n48534 , n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , n48541 , n48542 , n48543 , n48544 , n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , n48551 , n48552 , n48553 , n48554 , n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , n48561 , n48562 , n48563 , n48564 , n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , n48571 , n48572 , n48573 , n48574 , n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , n48581 , n48582 , n48583 , n48584 , n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , n48591 , n48592 , n48593 , n48594 , n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , n48601 , n48602 , n48603 , n48604 , n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , n48611 , n48612 , n48613 , n48614 , n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , n48621 , n48622 , n48623 , n48624 , n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , n48651 , n48652 , n48653 , n48654 , n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n48663 , n48664 , n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , n48671 , n48672 , n48673 , n48674 , n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , n48681 , n48682 , n48683 , n48684 , n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n48693 , n48694 , n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , n48701 , n48702 , n48703 , n48704 , n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , n48712 , n48713 , n48714 , n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , n48731 , n48732 , n48733 , n48734 , n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48753 , n48754 , n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , n48761 , n48762 , n48763 , n48764 , n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , n48774 , n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , n48781 , n48782 , n48783 , n48784 , n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , n48791 , n48792 , n48793 , n48794 , n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , n48804 , n48805 , n48806 , n48807 , n48808 , n48809 , n48810 , n48811 , n48812 , n48813 , n48814 , n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , n48821 , n48822 , n48823 , n48824 , n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , n48834 , n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , n48841 , n48842 , n48843 , n48844 , n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , n48851 , n48852 , n48853 , n48854 , n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 , n48864 , n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , n48881 , n48882 , n48883 , n48884 , n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , n48901 , n48902 , n48903 , n48904 , n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , n48921 , n48922 , n48923 , n48924 , n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , n48941 , n48942 , n48943 , n48944 , n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , n48961 , n48962 , n48963 , n48964 , n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , n48981 , n48982 , n48983 , n48984 , n48985 , n48986 , n48987 , n48988 , n48989 , n48990 , n48991 , n48992 , n48993 , n48994 , n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , n49001 , n49002 , n49003 , n49004 , n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , n49011 , n49012 , n49013 , n49014 , n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , n49024 , n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , n49051 , n49052 , n49053 , n49054 , n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , n49061 , n49062 , n49063 , n49064 , n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n49073 , n49074 , n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , n49082 , n49083 , n49084 , n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , n49091 , n49092 , n49093 , n49094 , n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , n49101 , n49102 , n49103 , n49104 , n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , n49111 , n49112 , n49113 , n49114 , n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , n49124 , n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , n49131 , n49132 , n49133 , n49134 , n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , n49141 , n49142 , n49143 , n49144 , n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n49153 , n49154 , n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , n49161 , n49162 , n49163 , n49164 , n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , n49171 , n49172 , n49173 , n49174 , n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , n49194 , n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n49213 , n49214 , n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , n49221 , n49222 , n49223 , n49224 , n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , n49231 , n49232 , n49233 , n49234 , n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , n49241 , n49242 , n49243 , n49244 , n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , n49251 , n49252 , n49253 , n49254 , n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , n49261 , n49262 , n49263 , n49264 , n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , n49281 , n49282 , n49283 , n49284 , n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , n49294 , n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , n49301 , n49302 , n49303 , n49304 , n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , n49311 , n49312 , n49313 , n49314 , n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , n49321 , n49322 , n49323 , n49324 , n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , n49331 , n49332 , n49333 , n49334 , n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , n49351 , n49352 , n49353 , n49354 , n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , n49391 , n49392 , n49393 , n49394 , n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , n49411 , n49412 , n49413 , n49414 , n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , n49421 , n49422 , n49423 , n49424 , n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , n49431 , n49432 , n49433 , n49434 , n49435 , n49436 , n49437 , n49438 , n49440 , n49441 , n49442 , n49443 , n49444 , n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , n49451 , n49452 , n49453 , n49454 , n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , n49461 , n49462 , n49463 , n49464 , n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , n49471 , n49472 , n49473 , n49474 , n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , n49481 , n49482 , n49483 , n49484 , n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , n49491 , n49492 , n49493 , n49494 , n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , n49501 , n49502 , n49503 , n49504 , n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , n49511 , n49512 , n49513 , n49514 , n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , n49521 , n49522 , n49523 , n49524 , n49525 , n49526 , n49527 , n49528 , n49529 , n49530 , n49531 , n49532 , n49533 , n49534 , n49535 , n49536 , n49537 , n49538 , n49539 , n49540 , n49541 , n49542 , n49543 , n49544 , n49545 , n49546 , n49547 , n49548 , n49549 , n49550 , n49551 , n49552 , n49553 , n49554 , n49555 , n49556 , n49557 , n49558 , n49559 , n49560 , n49561 , n49562 , n49563 , n49564 , n49565 , n49566 , n49567 , n49568 , n49569 , n49570 , n49571 , n49572 , n49573 , n49574 , n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , n49581 , n49582 , n49583 , n49584 , n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , n49591 , n49592 , n49593 , n49594 , n49595 , n49596 , n49597 , n49598 , n49599 , n49600 , n49601 , n49602 , n49603 , n49604 , n49605 , n49606 , n49607 , n49608 , n49609 , n49610 , n49611 , n49612 , n49613 , n49614 , n49615 , n49616 , n49617 , n49618 , n49619 , n49620 , n49621 , n49622 , n49623 , n49624 , n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , n49631 , n49632 , n49633 , n49634 , n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , n49641 , n49642 , n49643 , n49644 , n49645 , n49646 , n49647 , n49648 , n49649 , n49650 , n49651 , n49652 , n49653 , n49654 , n49655 , n49656 , n49657 , n49658 , n49659 , n49660 , n49661 , n49662 , n49663 , n49664 , n49665 , n49666 , n49667 , n49668 , n49669 , n49670 , n49671 , n49672 , n49673 , n49674 , n49675 , n49676 , n49677 , n49678 , n49679 , n49680 , n49681 , n49682 , n49683 , n49684 , n49685 , n49686 , n49687 , n49688 , n49689 , n49690 , n49691 , n49692 , n49693 , n49694 , n49695 , n49696 , n49697 , n49698 , n49699 , n49700 , n49701 , n49702 , n49703 , n49704 , n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , n49711 , n49712 , n49713 , n49714 , n49715 , n49716 , n49717 , n49718 , n49719 , n49720 , n49721 , n49722 , n49723 , n49724 , n49725 , n49726 , n49727 , n49728 , n49729 , n49730 , n49731 , n49732 , n49733 , n49734 , n49735 , n49736 , n49737 , n49738 , n49739 , n49740 , n49741 , n49742 , n49743 , n49744 , n49745 , n49746 , n49747 , n49748 , n49749 , n49750 , n49751 , n49752 , n49753 , n49754 , n49755 , n49756 , n49757 , n49758 , n49759 , n49760 , n49761 , n49762 , n49763 , n49764 , n49765 , n49766 , n49767 , n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , n49774 , n49775 , n49776 , n49777 , n49778 , n49779 , n49780 , n49781 , n49782 , n49784 , n49785 , n49786 , n49787 , n49788 , n49789 , n49790 , n49791 , n49792 , n49793 , n49794 , n49795 , n49796 , n49797 , n49798 , n49799 , n49800 , n49801 , n49802 , n49803 , n49804 , n49805 , n49806 , n49807 , n49808 , n49809 , n49810 , n49811 , n49812 , n49813 , n49814 , n49815 , n49816 , n49817 , n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , n49824 , n49825 , n49826 , n49827 , n49828 , n49829 , n49830 , n49831 , n49832 , n49833 , n49834 , n49835 , n49836 , n49837 , n49838 , n49839 , n49840 , n49841 , n49842 , n49843 , n49844 , n49845 , n49846 , n49847 , n49848 , n49849 , n49850 , n49851 , n49852 , n49853 , n49854 , n49855 , n49856 , n49857 , n49858 , n49859 , n49860 , n49861 , n49862 , n49863 , n49864 , n49865 , n49866 , n49867 , n49868 , n49869 , n49870 , n49871 , n49872 , n49873 , n49874 , n49875 , n49876 , n49877 , n49878 , n49879 , n49880 , n49881 , n49882 , n49883 , n49884 , n49885 , n49886 , n49887 , n49888 , n49889 , n49890 , n49891 , n49892 , n49893 , n49894 , n49895 , n49896 , n49897 , n49898 , n49899 , n49900 , n49901 , n49902 , n49903 , n49904 , n49905 , n49906 , n49907 , n49908 , n49909 , n49910 , n49911 , n49912 , n49913 , n49914 , n49915 , n49916 , n49917 , n49918 , n49919 , n49920 , n49921 , n49922 , n49923 , n49924 , n49925 , n49926 , n49927 , n49928 , n49929 , n49930 , n49931 , n49932 , n49933 , n49934 , n49935 , n49936 , n49937 , n49938 , n49939 , n49940 , n49941 , n49942 , n49943 , n49944 , n49945 , n49946 , n49947 , n49948 , n49949 , n49950 , n49951 , n49952 , n49953 , n49954 , n49955 , n49956 , n49957 , n49958 , n49959 , n49960 , n49961 , n49962 , n49963 , n49964 , n49965 , n49966 , n49967 , n49968 , n49969 , n49970 , n49971 , n49972 , n49973 , n49974 , n49975 , n49976 , n49977 , n49978 , n49979 , n49980 , n49981 , n49982 , n49983 , n49984 , n49985 , n49986 , n49987 , n49988 , n49989 , n49990 , n49991 , n49992 , n49993 , n49994 , n49995 , n49996 , n49997 , n49998 , n49999 , n50000 , n50001 , n50002 , n50003 , n50004 , n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , n50011 , n50012 , n50013 , n50014 , n50015 , n50016 , n50017 , n50018 , n50019 , n50020 , n50021 , n50022 , n50023 , n50024 , n50025 , n50026 , n50027 , n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , n50034 , n50035 , n50036 , n50037 , n50038 , n50039 , n50040 , n50041 , n50042 , n50043 , n50044 , n50045 , n50046 , n50047 , n50048 , n50049 , n50050 , n50051 , n50052 , n50053 , n50054 , n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , n50061 , n50062 , n50063 , n50064 , n50065 , n50066 , n50067 , n50068 , n50069 , n50070 , n50071 , n50072 , n50073 , n50074 , n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , n50081 , n50082 , n50083 , n50084 , n50085 , n50086 , n50087 , n50088 , n50089 , n50090 , n50091 , n50092 , n50093 , n50094 , n50095 , n50096 , n50097 , n50098 , n50099 , n50100 , n50101 , n50102 , n50103 , n50104 , n50105 , n50106 , n50107 , n50108 , n50109 , n50110 , n50112 , n50113 , n50114 , n50115 , n50116 , n50117 , n50118 , n50119 , n50120 , n50121 , n50122 , n50123 , n50124 , n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , n50131 , n50132 , n50133 , n50134 , n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , n50141 , n50142 , n50143 , n50144 , n50145 , n50146 , n50147 , n50148 , n50149 , n50150 , n50151 , n50152 , n50153 , n50154 , n50155 , n50156 , n50157 , n50158 , n50159 , n50160 , n50161 , n50162 , n50163 , n50164 , n50165 , n50166 , n50167 , n50168 , n50169 , n50170 , n50171 , n50172 , n50173 , n50174 , n50175 , n50176 , n50177 , n50178 , n50179 , n50180 , n50181 , n50182 , n50183 , n50184 , n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , n50191 , n50192 , n50193 , n50194 , n50195 , n50196 , n50197 , n50198 , n50199 , n50200 , n50201 , n50202 , n50203 , n50204 , n50205 , n50206 , n50207 , n50208 , n50209 , n50210 , n50211 , n50212 , n50213 , n50214 , n50215 , n50216 , n50217 , n50218 , n50219 , n50220 , n50221 , n50222 , n50223 , n50224 , n50225 , n50226 , n50227 , n50228 , n50229 , n50230 , n50231 , n50232 , n50233 , n50234 , n50235 , n50236 , n50237 , n50238 , n50239 , n50240 , n50241 , n50242 , n50243 , n50244 , n50245 , n50246 , n50247 , n50248 , n50249 , n50250 , n50251 , n50252 , n50253 , n50254 , n50255 , n50256 , n50257 , n50258 , n50259 , n50260 , n50261 , n50262 , n50263 , n50264 , n50265 , n50266 , n50267 , n50268 , n50269 , n50270 , n50271 , n50272 , n50273 , n50274 , n50275 , n50276 , n50277 , n50278 , n50279 , n50280 , n50281 , n50282 , n50283 , n50284 , n50285 , n50286 , n50287 , n50288 , n50289 , n50290 , n50291 , n50292 , n50293 , n50294 , n50295 , n50296 , n50297 , n50298 , n50299 , n50300 , n50301 , n50302 , n50303 , n50304 , n50305 , n50306 , n50307 , n50308 , n50309 , n50310 , n50311 , n50312 , n50313 , n50314 , n50315 , n50316 , n50317 , n50318 , n50319 , n50320 , n50321 , n50322 , n50323 , n50324 , n50325 , n50326 , n50327 , n50328 , n50329 , n50330 , n50331 , n50332 , n50333 , n50334 , n50335 , n50336 , n50337 , n50338 , n50339 , n50340 , n50341 , n50342 , n50343 , n50344 , n50345 , n50346 , n50347 , n50348 , n50349 , n50350 , n50351 , n50352 , n50353 , n50354 , n50355 , n50356 , n50357 , n50358 , n50359 , n50360 , n50361 , n50362 , n50363 , n50364 , n50365 , n50366 , n50367 , n50368 , n50369 , n50370 , n50371 , n50372 , n50373 , n50374 , n50375 , n50376 , n50377 , n50378 , n50379 , n50380 , n50381 , n50382 , n50383 , n50384 , n50385 , n50386 , n50387 , n50388 , n50389 , n50390 , n50391 , n50392 , n50393 , n50394 , n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , n50401 , n50402 , n50403 , n50404 , n50405 , n50406 , n50407 , n50408 , n50409 , n50410 , n50411 , n50412 , n50413 , n50414 , n50415 , n50416 , n50417 , n50418 , n50419 , n50420 , n50421 , n50422 , n50423 , n50424 , n50425 , n50426 , n50427 , n50428 , n50429 , n50430 , n50431 , n50432 , n50434 , n50435 , n50436 , n50437 , n50438 , n50439 , n50440 , n50441 , n50442 , n50443 , n50444 , n50445 , n50446 , n50447 , n50448 , n50449 , n50450 , n50451 , n50452 , n50453 , n50454 , n50455 , n50456 , n50457 , n50458 , n50459 , n50460 , n50461 , n50462 , n50463 , n50464 , n50465 , n50466 , n50467 , n50468 , n50469 , n50470 , n50471 , n50472 , n50473 , n50474 , n50475 , n50476 , n50477 , n50478 , n50479 , n50480 , n50481 , n50482 , n50483 , n50484 , n50485 , n50486 , n50487 , n50488 , n50489 , n50490 , n50491 , n50492 , n50493 , n50494 , n50495 , n50496 , n50497 , n50498 , n50499 , n50500 , n50501 , n50502 , n50503 , n50504 , n50505 , n50506 , n50507 , n50508 , n50509 , n50510 , n50511 , n50512 , n50513 , n50514 , n50515 , n50516 , n50517 , n50518 , n50519 , n50520 , n50521 , n50522 , n50523 , n50524 , n50525 , n50526 , n50527 , n50528 , n50529 , n50530 , n50531 , n50532 , n50533 , n50534 , n50535 , n50536 , n50537 , n50538 , n50539 , n50540 , n50541 , n50542 , n50543 , n50544 , n50545 , n50546 , n50547 , n50548 , n50549 , n50550 , n50551 , n50552 , n50553 , n50554 , n50555 , n50556 , n50557 , n50558 , n50559 , n50560 , n50561 , n50562 , n50563 , n50564 , n50565 , n50566 , n50567 , n50568 , n50569 , n50570 , n50571 , n50572 , n50573 , n50574 , n50575 , n50576 , n50577 , n50578 , n50579 , n50580 , n50581 , n50582 , n50583 , n50584 , n50585 , n50586 , n50587 , n50588 , n50589 , n50590 , n50591 , n50592 , n50593 , n50594 , n50595 , n50596 , n50597 , n50598 , n50599 , n50600 , n50601 , n50602 , n50603 , n50604 , n50605 , n50606 , n50607 , n50608 , n50609 , n50610 , n50611 , n50612 , n50613 , n50614 , n50615 , n50616 , n50617 , n50618 , n50619 , n50620 , n50621 , n50622 , n50623 , n50624 , n50625 , n50626 , n50627 , n50628 , n50629 , n50630 , n50631 , n50632 , n50633 , n50634 , n50635 , n50636 , n50637 , n50638 , n50639 , n50640 , n50641 , n50642 , n50643 , n50644 , n50645 , n50646 , n50647 , n50648 , n50649 , n50650 , n50651 , n50652 , n50653 , n50654 , n50655 , n50656 , n50657 , n50658 , n50659 , n50660 , n50661 , n50662 , n50663 , n50664 , n50665 , n50666 , n50667 , n50668 , n50669 , n50670 , n50671 , n50672 , n50673 , n50674 , n50675 , n50676 , n50677 , n50678 , n50679 , n50680 , n50681 , n50682 , n50683 , n50684 , n50685 , n50686 , n50687 , n50688 , n50689 , n50690 , n50691 , n50692 , n50693 , n50694 , n50695 , n50696 , n50697 , n50698 , n50699 , n50700 , n50701 , n50702 , n50703 , n50704 , n50705 , n50706 , n50707 , n50708 , n50709 , n50710 , n50711 , n50712 , n50713 , n50714 , n50715 , n50716 , n50717 , n50718 , n50719 , n50720 , n50721 , n50722 , n50723 , n50724 , n50725 , n50726 , n50727 , n50728 , n50729 , n50730 , n50731 , n50732 , n50733 , n50734 , n50735 , n50736 , n50737 , n50738 , n50740 , n50741 , n50742 , n50743 , n50744 , n50745 , n50746 , n50747 , n50748 , n50749 , n50750 , n50751 , n50752 , n50753 , n50754 , n50755 , n50756 , n50757 , n50758 , n50759 , n50760 , n50761 , n50762 , n50763 , n50764 , n50765 , n50766 , n50767 , n50768 , n50769 , n50770 , n50771 , n50772 , n50773 , n50774 , n50775 , n50776 , n50777 , n50778 , n50779 , n50780 , n50781 , n50782 , n50783 , n50784 , n50785 , n50786 , n50787 , n50788 , n50789 , n50790 , n50791 , n50792 , n50793 , n50794 , n50795 , n50796 , n50797 , n50798 , n50799 , n50800 , n50801 , n50802 , n50803 , n50804 , n50805 , n50806 , n50807 , n50808 , n50809 , n50810 , n50811 , n50812 , n50813 , n50814 , n50815 , n50816 , n50817 , n50818 , n50819 , n50820 , n50821 , n50822 , n50823 , n50824 , n50825 , n50826 , n50827 , n50828 , n50829 , n50830 , n50831 , n50832 , n50833 , n50834 , n50835 , n50836 , n50837 , n50838 , n50839 , n50840 , n50841 , n50842 , n50843 , n50844 , n50845 , n50846 , n50847 , n50848 , n50849 , n50850 , n50851 , n50852 , n50853 , n50854 , n50855 , n50856 , n50857 , n50858 , n50859 , n50860 , n50861 , n50862 , n50863 , n50864 , n50865 , n50866 , n50867 , n50868 , n50869 , n50870 , n50871 , n50872 , n50873 , n50874 , n50875 , n50876 , n50877 , n50878 , n50879 , n50880 , n50881 , n50882 , n50883 , n50884 , n50885 , n50886 , n50887 , n50888 , n50889 , n50890 , n50891 , n50892 , n50893 , n50894 , n50895 , n50896 , n50897 , n50898 , n50899 , n50900 , n50901 , n50902 , n50903 , n50904 , n50905 , n50906 , n50907 , n50908 , n50909 , n50910 , n50911 , n50912 , n50913 , n50914 , n50915 , n50916 , n50917 , n50918 , n50919 , n50920 , n50921 , n50922 , n50923 , n50924 , n50925 , n50926 , n50927 , n50928 , n50929 , n50930 , n50931 , n50932 , n50933 , n50934 , n50935 , n50936 , n50937 , n50938 , n50939 , n50940 , n50941 , n50942 , n50943 , n50944 , n50945 , n50946 , n50947 , n50948 , n50949 , n50950 , n50951 , n50952 , n50953 , n50954 , n50955 , n50956 , n50957 , n50958 , n50959 , n50960 , n50961 , n50962 , n50963 , n50964 , n50965 , n50966 , n50967 , n50968 , n50969 , n50970 , n50971 , n50972 , n50973 , n50974 , n50975 , n50976 , n50977 , n50978 , n50979 , n50980 , n50981 , n50982 , n50983 , n50984 , n50985 , n50986 , n50987 , n50988 , n50989 , n50990 , n50991 , n50992 , n50993 , n50994 , n50995 , n50996 , n50997 , n50998 , n50999 , n51000 , n51001 , n51002 , n51003 , n51004 , n51005 , n51006 , n51007 , n51008 , n51009 , n51010 , n51011 , n51012 , n51013 , n51014 , n51015 , n51016 , n51017 , n51018 , n51019 , n51020 , n51021 , n51022 , n51023 , n51024 , n51025 , n51026 , n51027 , n51028 , n51030 , n51031 , n51032 , n51033 , n51034 , n51035 , n51036 , n51037 , n51038 , n51039 , n51040 , n51041 , n51042 , n51043 , n51044 , n51045 , n51046 , n51047 , n51048 , n51049 , n51050 , n51051 , n51052 , n51053 , n51054 , n51055 , n51056 , n51057 , n51058 , n51059 , n51060 , n51061 , n51062 , n51063 , n51064 , n51065 , n51066 , n51067 , n51068 , n51069 , n51070 , n51071 , n51072 , n51073 , n51074 , n51075 , n51076 , n51077 , n51078 , n51079 , n51080 , n51081 , n51082 , n51083 , n51084 , n51085 , n51086 , n51087 , n51088 , n51089 , n51090 , n51091 , n51092 , n51093 , n51094 , n51095 , n51096 , n51097 , n51098 , n51099 , n51100 , n51101 , n51102 , n51103 , n51104 , n51105 , n51106 , n51107 , n51108 , n51109 , n51110 , n51111 , n51112 , n51113 , n51114 , n51115 , n51116 , n51117 , n51118 , n51119 , n51120 , n51121 , n51122 , n51123 , n51124 , n51125 , n51126 , n51127 , n51128 , n51129 , n51130 , n51131 , n51132 , n51133 , n51134 , n51135 , n51136 , n51137 , n51138 , n51139 , n51140 , n51141 , n51142 , n51143 , n51144 , n51145 , n51146 , n51147 , n51148 , n51149 , n51150 , n51151 , n51152 , n51153 , n51154 , n51155 , n51156 , n51157 , n51158 , n51159 , n51160 , n51161 , n51162 , n51163 , n51164 , n51165 , n51166 , n51167 , n51168 , n51169 , n51170 , n51171 , n51172 , n51173 , n51174 , n51175 , n51176 , n51177 , n51178 , n51179 , n51180 , n51181 , n51182 , n51183 , n51184 , n51185 , n51186 , n51187 , n51188 , n51189 , n51190 , n51191 , n51192 , n51193 , n51194 , n51195 , n51196 , n51197 , n51198 , n51199 , n51200 , n51201 , n51202 , n51203 , n51204 , n51205 , n51206 , n51207 , n51208 , n51209 , n51210 , n51211 , n51212 , n51213 , n51214 , n51215 , n51216 , n51217 , n51218 , n51219 , n51220 , n51221 , n51222 , n51223 , n51224 , n51225 , n51226 , n51227 , n51228 , n51229 , n51230 , n51231 , n51232 , n51233 , n51234 , n51235 , n51236 , n51237 , n51238 , n51239 , n51240 , n51241 , n51242 , n51243 , n51244 , n51245 , n51246 , n51247 , n51248 , n51249 , n51250 , n51251 , n51252 , n51253 , n51254 , n51255 , n51256 , n51257 , n51258 , n51259 , n51260 , n51261 , n51262 , n51263 , n51264 , n51265 , n51266 , n51267 , n51268 , n51269 , n51270 , n51271 , n51272 , n51273 , n51274 , n51275 , n51276 , n51277 , n51278 , n51279 , n51280 , n51281 , n51282 , n51283 , n51284 , n51285 , n51286 , n51287 , n51288 , n51289 , n51290 , n51291 , n51292 , n51293 , n51294 , n51295 , n51296 , n51297 , n51298 , n51299 , n51300 , n51301 , n51302 , n51303 , n51304 , n51305 , n51306 , n51307 , n51308 , n51309 , n51310 , n51311 , n51312 , n51313 , n51314 , n51315 , n51316 , n51317 , n51318 , n51320 , n51321 , n51322 , n51323 , n51324 , n51325 , n51326 , n51327 , n51328 , n51329 , n51330 , n51331 , n51332 , n51333 , n51334 , n51335 , n51336 , n51337 , n51338 , n51339 , n51340 , n51341 , n51342 , n51343 , n51344 , n51345 , n51346 , n51347 , n51348 , n51349 , n51350 , n51351 , n51352 , n51353 , n51354 , n51355 , n51356 , n51357 , n51358 , n51359 , n51360 , n51361 , n51362 , n51363 , n51364 , n51365 , n51366 , n51367 , n51368 , n51369 , n51370 , n51371 , n51372 , n51373 , n51374 , n51375 , n51376 , n51377 , n51378 , n51379 , n51380 , n51381 , n51382 , n51383 , n51384 , n51385 , n51386 , n51387 , n51388 , n51389 , n51390 , n51391 , n51392 , n51393 , n51394 , n51395 , n51396 , n51397 , n51398 , n51399 , n51400 , n51401 , n51402 , n51403 , n51404 , n51405 , n51406 , n51407 , n51408 , n51409 , n51410 , n51411 , n51412 , n51413 , n51414 , n51415 , n51416 , n51417 , n51418 , n51419 , n51420 , n51421 , n51422 , n51423 , n51424 , n51425 , n51426 , n51427 , n51428 , n51429 , n51430 , n51431 , n51432 , n51433 , n51434 , n51435 , n51436 , n51437 , n51438 , n51439 , n51440 , n51441 , n51442 , n51443 , n51444 , n51445 , n51446 , n51447 , n51448 , n51449 , n51450 , n51451 , n51452 , n51453 , n51454 , n51455 , n51456 , n51457 , n51458 , n51459 , n51460 , n51461 , n51462 , n51463 , n51464 , n51465 , n51466 , n51467 , n51468 , n51469 , n51470 , n51471 , n51472 , n51473 , n51474 , n51475 , n51476 , n51477 , n51478 , n51479 , n51480 , n51481 , n51482 , n51483 , n51484 , n51485 , n51486 , n51487 , n51488 , n51489 , n51490 , n51491 , n51492 , n51493 , n51494 , n51495 , n51496 , n51497 , n51498 , n51499 , n51500 , n51501 , n51502 , n51503 , n51504 , n51505 , n51506 , n51507 , n51508 , n51509 , n51510 , n51511 , n51512 , n51513 , n51514 , n51515 , n51516 , n51517 , n51518 , n51519 , n51520 , n51521 , n51522 , n51523 , n51524 , n51525 , n51526 , n51527 , n51528 , n51529 , n51530 , n51531 , n51532 , n51533 , n51534 , n51535 , n51536 , n51537 , n51538 , n51539 , n51540 , n51541 , n51542 , n51543 , n51544 , n51545 , n51546 , n51547 , n51548 , n51549 , n51550 , n51551 , n51552 , n51553 , n51554 , n51555 , n51556 , n51557 , n51558 , n51559 , n51560 , n51561 , n51562 , n51563 , n51564 , n51565 , n51566 , n51567 , n51568 , n51569 , n51570 , n51571 , n51572 , n51573 , n51574 , n51575 , n51576 , n51577 , n51578 , n51579 , n51580 , n51581 , n51582 , n51584 , n51585 , n51586 , n51587 , n51588 , n51589 , n51590 , n51591 , n51592 , n51593 , n51594 , n51595 , n51596 , n51597 , n51598 , n51599 , n51600 , n51601 , n51602 , n51603 , n51604 , n51605 , n51606 , n51607 , n51608 , n51609 , n51610 , n51611 , n51612 , n51613 , n51614 , n51615 , n51616 , n51617 , n51618 , n51619 , n51620 , n51621 , n51622 , n51623 , n51624 , n51625 , n51626 , n51627 , n51628 , n51629 , n51630 , n51631 , n51632 , n51633 , n51634 , n51635 , n51636 , n51637 , n51638 , n51639 , n51640 , n51641 , n51642 , n51643 , n51644 , n51645 , n51646 , n51647 , n51648 , n51649 , n51650 , n51651 , n51652 , n51653 , n51654 , n51655 , n51656 , n51657 , n51658 , n51659 , n51660 , n51661 , n51662 , n51663 , n51664 , n51665 , n51666 , n51667 , n51668 , n51669 , n51670 , n51671 , n51672 , n51673 , n51674 , n51675 , n51676 , n51677 , n51678 , n51679 , n51680 , n51681 , n51682 , n51683 , n51684 , n51685 , n51686 , n51687 , n51688 , n51689 , n51690 , n51691 , n51692 , n51693 , n51694 , n51695 , n51696 , n51697 , n51698 , n51699 , n51700 , n51701 , n51702 , n51703 , n51704 , n51705 , n51706 , n51707 , n51708 , n51709 , n51710 , n51711 , n51712 , n51713 , n51714 , n51715 , n51716 , n51717 , n51718 , n51719 , n51720 , n51721 , n51722 , n51723 , n51724 , n51725 , n51726 , n51727 , n51728 , n51729 , n51730 , n51731 , n51732 , n51733 , n51734 , n51735 , n51736 , n51737 , n51738 , n51739 , n51740 , n51741 , n51742 , n51743 , n51744 , n51745 , n51746 , n51747 , n51748 , n51749 , n51750 , n51751 , n51752 , n51753 , n51754 , n51755 , n51756 , n51757 , n51758 , n51759 , n51760 , n51761 , n51762 , n51763 , n51764 , n51765 , n51766 , n51767 , n51768 , n51769 , n51770 , n51771 , n51772 , n51773 , n51774 , n51775 , n51776 , n51777 , n51778 , n51779 , n51780 , n51781 , n51782 , n51783 , n51784 , n51785 , n51786 , n51787 , n51788 , n51789 , n51790 , n51791 , n51792 , n51793 , n51794 , n51795 , n51796 , n51797 , n51798 , n51799 , n51800 , n51801 , n51802 , n51803 , n51804 , n51805 , n51806 , n51807 , n51808 , n51809 , n51810 , n51811 , n51812 , n51813 , n51814 , n51815 , n51816 , n51817 , n51818 , n51819 , n51820 , n51821 , n51822 , n51823 , n51824 , n51825 , n51826 , n51827 , n51828 , n51829 , n51830 , n51831 , n51832 , n51834 , n51835 , n51836 , n51837 , n51838 , n51839 , n51840 , n51841 , n51842 , n51843 , n51844 , n51845 , n51846 , n51847 , n51848 , n51849 , n51850 , n51851 , n51852 , n51853 , n51854 , n51855 , n51856 , n51857 , n51858 , n51859 , n51860 , n51861 , n51862 , n51863 , n51864 , n51865 , n51866 , n51867 , n51868 , n51869 , n51870 , n51871 , n51872 , n51873 , n51874 , n51875 , n51876 , n51877 , n51878 , n51879 , n51880 , n51881 , n51882 , n51883 , n51884 , n51885 , n51886 , n51887 , n51888 , n51889 , n51890 , n51891 , n51892 , n51893 , n51894 , n51895 , n51896 , n51897 , n51898 , n51899 , n51900 , n51901 , n51902 , n51903 , n51904 , n51905 , n51906 , n51907 , n51908 , n51909 , n51910 , n51911 , n51912 , n51913 , n51914 , n51915 , n51916 , n51917 , n51918 , n51919 , n51920 , n51921 , n51922 , n51923 , n51924 , n51925 , n51926 , n51927 , n51928 , n51929 , n51930 , n51931 , n51932 , n51933 , n51934 , n51935 , n51936 , n51937 , n51938 , n51939 , n51940 , n51941 , n51942 , n51943 , n51944 , n51945 , n51946 , n51947 , n51948 , n51949 , n51950 , n51951 , n51952 , n51953 , n51954 , n51955 , n51956 , n51957 , n51958 , n51959 , n51960 , n51961 , n51962 , n51963 , n51964 , n51965 , n51966 , n51967 , n51968 , n51969 , n51970 , n51971 , n51972 , n51973 , n51974 , n51975 , n51976 , n51977 , n51978 , n51979 , n51980 , n51981 , n51982 , n51983 , n51984 , n51985 , n51986 , n51987 , n51988 , n51989 , n51990 , n51991 , n51992 , n51993 , n51994 , n51995 , n51996 , n51997 , n51998 , n51999 , n52000 , n52001 , n52002 , n52003 , n52004 , n52005 , n52006 , n52007 , n52008 , n52009 , n52010 , n52011 , n52012 , n52013 , n52014 , n52015 , n52016 , n52017 , n52018 , n52019 , n52020 , n52021 , n52022 , n52023 , n52024 , n52025 , n52026 , n52027 , n52028 , n52029 , n52030 , n52031 , n52032 , n52033 , n52034 , n52035 , n52036 , n52037 , n52038 , n52039 , n52040 , n52041 , n52042 , n52043 , n52044 , n52045 , n52046 , n52047 , n52048 , n52049 , n52050 , n52051 , n52052 , n52053 , n52054 , n52055 , n52056 , n52057 , n52058 , n52059 , n52060 , n52061 , n52062 , n52063 , n52064 , n52065 , n52066 , n52067 , n52068 , n52069 , n52070 , n52071 , n52072 , n52073 , n52074 , n52075 , n52076 , n52077 , n52078 , n52079 , n52080 , n52081 , n52082 , n52084 , n52085 , n52086 , n52087 , n52088 , n52089 , n52090 , n52091 , n52092 , n52093 , n52094 , n52095 , n52096 , n52097 , n52098 , n52099 , n52100 , n52101 , n52102 , n52103 , n52104 , n52105 , n52106 , n52107 , n52108 , n52109 , n52110 , n52111 , n52112 , n52113 , n52114 , n52115 , n52116 , n52117 , n52118 , n52119 , n52120 , n52121 , n52122 , n52123 , n52124 , n52125 , n52126 , n52127 , n52128 , n52129 , n52130 , n52131 , n52132 , n52133 , n52134 , n52135 , n52136 , n52137 , n52138 , n52139 , n52140 , n52141 , n52142 , n52143 , n52144 , n52145 , n52146 , n52147 , n52148 , n52149 , n52150 , n52151 , n52152 , n52153 , n52154 , n52155 , n52156 , n52157 , n52158 , n52159 , n52160 , n52161 , n52162 , n52163 , n52164 , n52165 , n52166 , n52167 , n52168 , n52169 , n52170 , n52171 , n52172 , n52173 , n52174 , n52175 , n52176 , n52177 , n52178 , n52179 , n52180 , n52181 , n52182 , n52183 , n52184 , n52185 , n52186 , n52187 , n52188 , n52189 , n52190 , n52191 , n52192 , n52193 , n52194 , n52195 , n52196 , n52197 , n52198 , n52199 , n52200 , n52201 , n52202 , n52203 , n52204 , n52205 , n52206 , n52207 , n52208 , n52209 , n52210 , n52211 , n52212 , n52213 , n52214 , n52215 , n52216 , n52217 , n52218 , n52219 , n52220 , n52221 , n52222 , n52223 , n52224 , n52225 , n52226 , n52227 , n52228 , n52229 , n52230 , n52231 , n52232 , n52233 , n52234 , n52235 , n52236 , n52237 , n52238 , n52239 , n52240 , n52241 , n52242 , n52243 , n52244 , n52245 , n52246 , n52247 , n52248 , n52249 , n52250 , n52251 , n52252 , n52253 , n52254 , n52255 , n52256 , n52257 , n52258 , n52259 , n52260 , n52261 , n52262 , n52263 , n52264 , n52265 , n52266 , n52267 , n52268 , n52269 , n52270 , n52271 , n52272 , n52273 , n52274 , n52275 , n52276 , n52277 , n52278 , n52279 , n52280 , n52281 , n52282 , n52283 , n52284 , n52285 , n52286 , n52287 , n52288 , n52289 , n52290 , n52291 , n52292 , n52293 , n52294 , n52295 , n52296 , n52297 , n52298 , n52299 , n52300 , n52301 , n52302 , n52303 , n52304 , n52305 , n52306 , n52308 , n52309 , n52310 , n52311 , n52312 , n52313 , n52314 , n52315 , n52316 , n52317 , n52318 , n52319 , n52320 , n52321 , n52322 , n52323 , n52324 , n52325 , n52326 , n52327 , n52328 , n52329 , n52330 , n52331 , n52332 , n52333 , n52334 , n52335 , n52336 , n52337 , n52338 , n52339 , n52340 , n52341 , n52342 , n52343 , n52344 , n52345 , n52346 , n52347 , n52348 , n52349 , n52350 , n52351 , n52352 , n52353 , n52354 , n52355 , n52356 , n52357 , n52358 , n52359 , n52360 , n52361 , n52362 , n52363 , n52364 , n52365 , n52366 , n52367 , n52368 , n52369 , n52370 , n52371 , n52372 , n52373 , n52374 , n52375 , n52376 , n52377 , n52378 , n52379 , n52380 , n52381 , n52382 , n52383 , n52384 , n52385 , n52386 , n52387 , n52388 , n52389 , n52390 , n52391 , n52392 , n52393 , n52394 , n52395 , n52396 , n52397 , n52398 , n52399 , n52400 , n52401 , n52402 , n52403 , n52404 , n52405 , n52406 , n52407 , n52408 , n52409 , n52410 , n52411 , n52412 , n52413 , n52414 , n52415 , n52416 , n52417 , n52418 , n52419 , n52420 , n52421 , n52422 , n52423 , n52424 , n52425 , n52426 , n52427 , n52428 , n52429 , n52430 , n52431 , n52432 , n52433 , n52434 , n52435 , n52436 , n52437 , n52438 , n52439 , n52440 , n52441 , n52442 , n52443 , n52444 , n52445 , n52446 , n52447 , n52448 , n52449 , n52450 , n52451 , n52452 , n52453 , n52454 , n52455 , n52456 , n52457 , n52458 , n52459 , n52460 , n52461 , n52462 , n52463 , n52464 , n52465 , n52466 , n52467 , n52468 , n52469 , n52470 , n52471 , n52472 , n52473 , n52474 , n52475 , n52476 , n52477 , n52478 , n52479 , n52480 , n52481 , n52482 , n52483 , n52484 , n52485 , n52486 , n52487 , n52488 , n52489 , n52490 , n52491 , n52492 , n52493 , n52494 , n52495 , n52496 , n52497 , n52498 , n52499 , n52500 , n52501 , n52502 , n52503 , n52504 , n52505 , n52506 , n52507 , n52508 , n52509 , n52510 , n52511 , n52512 , n52513 , n52514 , n52515 , n52516 , n52517 , n52518 , n52519 , n52520 , n52522 , n52523 , n52524 , n52525 , n52526 , n52527 , n52528 , n52529 , n52530 , n52531 , n52532 , n52533 , n52534 , n52535 , n52536 , n52537 , n52538 , n52539 , n52540 , n52541 , n52542 , n52543 , n52544 , n52545 , n52546 , n52547 , n52548 , n52549 , n52550 , n52551 , n52552 , n52553 , n52554 , n52555 , n52556 , n52557 , n52558 , n52559 , n52560 , n52561 , n52562 , n52563 , n52564 , n52565 , n52566 , n52567 , n52568 , n52569 , n52570 , n52571 , n52572 , n52573 , n52574 , n52575 , n52576 , n52577 , n52578 , n52579 , n52580 , n52581 , n52582 , n52583 , n52584 , n52585 , n52586 , n52587 , n52588 , n52589 , n52590 , n52591 , n52592 , n52593 , n52594 , n52595 , n52596 , n52597 , n52598 , n52599 , n52600 , n52601 , n52602 , n52603 , n52604 , n52605 , n52606 , n52607 , n52608 , n52609 , n52610 , n52611 , n52612 , n52613 , n52614 , n52615 , n52616 , n52617 , n52618 , n52619 , n52620 , n52621 , n52622 , n52623 , n52624 , n52625 , n52626 , n52627 , n52628 , n52629 , n52630 , n52631 , n52632 , n52633 , n52634 , n52635 , n52636 , n52637 , n52638 , n52639 , n52640 , n52641 , n52642 , n52643 , n52644 , n52645 , n52646 , n52647 , n52648 , n52649 , n52650 , n52651 , n52652 , n52653 , n52654 , n52655 , n52656 , n52657 , n52658 , n52659 , n52660 , n52661 , n52662 , n52663 , n52664 , n52665 , n52666 , n52667 , n52668 , n52669 , n52670 , n52671 , n52672 , n52673 , n52674 , n52675 , n52676 , n52677 , n52678 , n52679 , n52680 , n52681 , n52682 , n52683 , n52684 , n52685 , n52686 , n52687 , n52688 , n52689 , n52690 , n52691 , n52692 , n52693 , n52694 , n52695 , n52696 , n52697 , n52698 , n52699 , n52700 , n52701 , n52702 , n52703 , n52704 , n52705 , n52706 , n52707 , n52708 , n52709 , n52710 , n52711 , n52712 , n52713 , n52714 , n52715 , n52716 , n52717 , n52718 , n52719 , n52720 , n52721 , n52722 , n52723 , n52724 , n52725 , n52726 , n52728 , n52729 , n52730 , n52731 , n52732 , n52733 , n52734 , n52735 , n52736 , n52737 , n52738 , n52739 , n52740 , n52741 , n52742 , n52743 , n52744 , n52745 , n52746 , n52747 , n52748 , n52749 , n52750 , n52751 , n52752 , n52753 , n52754 , n52755 , n52756 , n52757 , n52758 , n52759 , n52760 , n52761 , n52762 , n52763 , n52764 , n52765 , n52766 , n52767 , n52768 , n52769 , n52770 , n52771 , n52772 , n52773 , n52774 , n52775 , n52776 , n52777 , n52778 , n52779 , n52780 , n52781 , n52782 , n52783 , n52784 , n52785 , n52786 , n52787 , n52788 , n52789 , n52790 , n52791 , n52792 , n52793 , n52794 , n52795 , n52796 , n52797 , n52798 , n52799 , n52800 , n52801 , n52802 , n52803 , n52804 , n52805 , n52806 , n52807 , n52808 , n52809 , n52810 , n52811 , n52812 , n52813 , n52814 , n52815 , n52816 , n52817 , n52818 , n52819 , n52820 , n52821 , n52822 , n52823 , n52824 , n52825 , n52826 , n52827 , n52828 , n52829 , n52830 , n52831 , n52832 , n52833 , n52834 , n52835 , n52836 , n52837 , n52838 , n52839 , n52840 , n52841 , n52842 , n52843 , n52844 , n52845 , n52846 , n52847 , n52848 , n52849 , n52850 , n52851 , n52852 , n52853 , n52854 , n52855 , n52856 , n52857 , n52858 , n52859 , n52860 , n52861 , n52862 , n52863 , n52864 , n52865 , n52866 , n52867 , n52868 , n52869 , n52870 , n52871 , n52872 , n52873 , n52874 , n52875 , n52876 , n52877 , n52878 , n52879 , n52880 , n52881 , n52882 , n52883 , n52884 , n52885 , n52886 , n52887 , n52888 , n52889 , n52890 , n52891 , n52892 , n52893 , n52894 , n52895 , n52896 , n52897 , n52898 , n52899 , n52900 , n52901 , n52902 , n52903 , n52904 , n52905 , n52906 , n52907 , n52908 , n52909 , n52910 , n52911 , n52912 , n52913 , n52914 , n52915 , n52916 , n52917 , n52918 , n52920 , n52921 , n52922 , n52923 , n52924 , n52925 , n52926 , n52927 , n52928 , n52929 , n52930 , n52931 , n52932 , n52933 , n52934 , n52935 , n52936 , n52937 , n52938 , n52939 , n52940 , n52941 , n52942 , n52943 , n52944 , n52945 , n52946 , n52947 , n52948 , n52949 , n52950 , n52951 , n52952 , n52953 , n52954 , n52955 , n52956 , n52957 , n52958 , n52959 , n52960 , n52961 , n52962 , n52963 , n52964 , n52965 , n52966 , n52967 , n52968 , n52969 , n52970 , n52971 , n52972 , n52973 , n52974 , n52975 , n52976 , n52977 , n52978 , n52979 , n52980 , n52981 , n52982 , n52983 , n52984 , n52985 , n52986 , n52987 , n52988 , n52989 , n52990 , n52991 , n52992 , n52993 , n52994 , n52995 , n52996 , n52997 , n52998 , n52999 , n53000 , n53001 , n53002 , n53003 , n53004 , n53005 , n53006 , n53007 , n53008 , n53009 , n53010 , n53011 , n53012 , n53013 , n53014 , n53015 , n53016 , n53017 , n53018 , n53019 , n53020 , n53021 , n53022 , n53023 , n53024 , n53025 , n53026 , n53027 , n53028 , n53029 , n53030 , n53031 , n53032 , n53033 , n53034 , n53035 , n53036 , n53037 , n53038 , n53039 , n53040 , n53041 , n53042 , n53043 , n53044 , n53045 , n53046 , n53047 , n53048 , n53049 , n53050 , n53051 , n53052 , n53053 , n53054 , n53055 , n53056 , n53057 , n53058 , n53059 , n53060 , n53061 , n53062 , n53063 , n53064 , n53065 , n53066 , n53067 , n53068 , n53069 , n53070 , n53071 , n53072 , n53073 , n53074 , n53075 , n53076 , n53077 , n53078 , n53079 , n53080 , n53081 , n53082 , n53083 , n53084 , n53085 , n53086 , n53087 , n53088 , n53089 , n53090 , n53092 , n53093 , n53094 , n53095 , n53096 , n53097 , n53098 , n53099 , n53100 , n53101 , n53102 , n53103 , n53104 , n53105 , n53106 , n53107 , n53108 , n53109 , n53110 , n53111 , n53112 , n53113 , n53114 , n53115 , n53116 , n53117 , n53118 , n53119 , n53120 , n53121 , n53122 , n53123 , n53124 , n53125 , n53126 , n53127 , n53128 , n53129 , n53130 , n53131 , n53132 , n53133 , n53134 , n53135 , n53136 , n53137 , n53138 , n53139 , n53140 , n53141 , n53142 , n53143 , n53144 , n53145 , n53146 , n53147 , n53148 , n53149 , n53150 , n53151 , n53152 , n53153 , n53154 , n53155 , n53156 , n53157 , n53158 , n53159 , n53160 , n53161 , n53162 , n53163 , n53164 , n53165 , n53166 , n53167 , n53168 , n53169 , n53170 , n53171 , n53172 , n53173 , n53174 , n53175 , n53176 , n53177 , n53178 , n53179 , n53180 , n53181 , n53182 , n53183 , n53184 , n53185 , n53186 , n53187 , n53188 , n53189 , n53190 , n53191 , n53192 , n53193 , n53194 , n53195 , n53196 , n53197 , n53198 , n53199 , n53200 , n53201 , n53202 , n53203 , n53204 , n53205 , n53206 , n53207 , n53208 , n53209 , n53210 , n53211 , n53212 , n53213 , n53214 , n53215 , n53216 , n53217 , n53218 , n53219 , n53220 , n53221 , n53222 , n53223 , n53224 , n53225 , n53226 , n53227 , n53228 , n53229 , n53230 , n53231 , n53232 , n53233 , n53234 , n53235 , n53236 , n53237 , n53238 , n53239 , n53240 , n53241 , n53242 , n53243 , n53244 , n53245 , n53246 , n53247 , n53248 , n53249 , n53250 , n53251 , n53252 , n53253 , n53254 , n53255 , n53256 , n53257 , n53258 , n53260 , n53261 , n53262 , n53263 , n53264 , n53265 , n53266 , n53267 , n53268 , n53269 , n53270 , n53271 , n53272 , n53273 , n53274 , n53275 , n53276 , n53277 , n53278 , n53279 , n53280 , n53281 , n53282 , n53283 , n53284 , n53285 , n53286 , n53287 , n53288 , n53289 , n53290 , n53291 , n53292 , n53293 , n53294 , n53295 , n53296 , n53297 , n53298 , n53299 , n53300 , n53301 , n53302 , n53303 , n53304 , n53305 , n53306 , n53307 , n53308 , n53309 , n53310 , n53311 , n53312 , n53313 , n53314 , n53315 , n53316 , n53317 , n53318 , n53319 , n53320 , n53321 , n53322 , n53323 , n53324 , n53325 , n53326 , n53327 , n53328 , n53329 , n53330 , n53331 , n53332 , n53333 , n53334 , n53335 , n53336 , n53337 , n53338 , n53339 , n53340 , n53341 , n53342 , n53343 , n53344 , n53345 , n53346 , n53347 , n53348 , n53349 , n53350 , n53351 , n53352 , n53353 , n53354 , n53355 , n53356 , n53357 , n53358 , n53359 , n53360 , n53361 , n53362 , n53363 , n53364 , n53365 , n53366 , n53367 , n53368 , n53369 , n53370 , n53371 , n53372 , n53373 , n53374 , n53375 , n53376 , n53377 , n53378 , n53379 , n53380 , n53381 , n53382 , n53383 , n53384 , n53385 , n53386 , n53387 , n53388 , n53389 , n53390 , n53391 , n53392 , n53393 , n53394 , n53395 , n53396 , n53397 , n53398 , n53399 , n53400 , n53401 , n53402 , n53403 , n53404 , n53405 , n53406 , n53407 , n53408 , n53409 , n53410 , n53411 , n53412 , n53414 , n53415 , n53416 , n53417 , n53418 , n53419 , n53420 , n53421 , n53422 , n53423 , n53424 , n53425 , n53426 , n53427 , n53428 , n53429 , n53430 , n53431 , n53432 , n53433 , n53434 , n53435 , n53436 , n53437 , n53438 , n53439 , n53440 , n53441 , n53442 , n53443 , n53444 , n53445 , n53446 , n53447 , n53448 , n53449 , n53450 , n53451 , n53452 , n53453 , n53454 , n53455 , n53456 , n53457 , n53458 , n53459 , n53460 , n53461 , n53462 , n53463 , n53464 , n53465 , n53466 , n53467 , n53468 , n53469 , n53470 , n53471 , n53472 , n53473 , n53474 , n53475 , n53476 , n53477 , n53478 , n53479 , n53480 , n53481 , n53482 , n53483 , n53484 , n53485 , n53486 , n53487 , n53488 , n53489 , n53490 , n53491 , n53492 , n53493 , n53494 , n53495 , n53496 , n53497 , n53498 , n53499 , n53500 , n53501 , n53502 , n53503 , n53504 , n53505 , n53506 , n53507 , n53508 , n53509 , n53510 , n53511 , n53512 , n53513 , n53514 , n53515 , n53516 , n53517 , n53518 , n53519 , n53520 , n53521 , n53522 , n53523 , n53524 , n53525 , n53526 , n53527 , n53528 , n53529 , n53530 , n53531 , n53532 , n53533 , n53534 , n53535 , n53536 , n53537 , n53538 , n53539 , n53540 , n53541 , n53542 , n53543 , n53544 , n53545 , n53546 , n53547 , n53548 , n53549 , n53550 , n53551 , n53552 , n53553 , n53554 , n53556 , n53557 , n53558 , n53559 , n53560 , n53561 , n53562 , n53563 , n53564 , n53565 , n53566 , n53567 , n53568 , n53569 , n53570 , n53571 , n53572 , n53573 , n53574 , n53575 , n53576 , n53577 , n53578 , n53579 , n53580 , n53581 , n53582 , n53583 , n53584 , n53585 , n53586 , n53587 , n53588 , n53589 , n53590 , n53591 , n53592 , n53593 , n53594 , n53595 , n53596 , n53597 , n53598 , n53599 , n53600 , n53601 , n53602 , n53603 , n53604 , n53605 , n53606 , n53607 , n53608 , n53609 , n53610 , n53611 , n53612 , n53613 , n53614 , n53615 , n53616 , n53617 , n53618 , n53619 , n53620 , n53621 , n53622 , n53623 , n53624 , n53625 , n53626 , n53627 , n53628 , n53629 , n53630 , n53631 , n53632 , n53633 , n53634 , n53635 , n53636 , n53637 , n53638 , n53639 , n53640 , n53641 , n53642 , n53643 , n53644 , n53645 , n53646 , n53647 , n53648 , n53649 , n53650 , n53651 , n53652 , n53653 , n53654 , n53655 , n53656 , n53657 , n53658 , n53659 , n53660 , n53661 , n53662 , n53663 , n53664 , n53665 , n53666 , n53667 , n53668 , n53669 , n53670 , n53671 , n53672 , n53673 , n53674 , n53675 , n53676 , n53677 , n53678 , n53679 , n53680 , n53681 , n53682 , n53683 , n53684 , n53685 , n53686 , n53688 , n53689 , n53690 , n53691 , n53692 , n53693 , n53694 , n53695 , n53696 , n53697 , n53698 , n53699 , n53700 , n53701 , n53702 , n53703 , n53704 , n53705 , n53706 , n53707 , n53708 , n53709 , n53710 , n53711 , n53712 , n53713 , n53714 , n53715 , n53716 , n53717 , n53718 , n53719 , n53720 , n53721 , n53722 , n53723 , n53724 , n53725 , n53726 , n53727 , n53728 , n53729 , n53730 , n53731 , n53732 , n53733 , n53734 , n53735 , n53736 , n53737 , n53738 , n53739 , n53740 , n53741 , n53742 , n53743 , n53744 , n53745 , n53746 , n53747 , n53748 , n53749 , n53750 , n53751 , n53752 , n53753 , n53754 , n53755 , n53756 , n53757 , n53758 , n53759 , n53760 , n53761 , n53762 , n53763 , n53764 , n53765 , n53766 , n53767 , n53768 , n53769 , n53770 , n53771 , n53772 , n53773 , n53774 , n53775 , n53776 , n53777 , n53778 , n53779 , n53780 , n53781 , n53782 , n53783 , n53784 , n53785 , n53786 , n53787 , n53788 , n53789 , n53790 , n53791 , n53792 , n53793 , n53794 , n53795 , n53796 , n53797 , n53798 , n53799 , n53800 , n53801 , n53802 , n53803 , n53804 , n53805 , n53806 , n53808 , n53809 , n53810 , n53811 , n53812 , n53813 , n53814 , n53815 , n53816 , n53817 , n53818 , n53819 , n53820 , n53821 , n53822 , n53823 , n53824 , n53825 , n53826 , n53827 , n53828 , n53829 , n53830 , n53831 , n53832 , n53833 , n53834 , n53835 , n53836 , n53837 , n53838 , n53839 , n53840 , n53841 , n53842 , n53843 , n53844 , n53845 , n53846 , n53847 , n53848 , n53849 , n53850 , n53851 , n53852 , n53853 , n53854 , n53855 , n53856 , n53857 , n53858 , n53859 , n53860 , n53861 , n53862 , n53863 , n53864 , n53865 , n53866 , n53867 , n53868 , n53869 , n53870 , n53871 , n53872 , n53873 , n53874 , n53875 , n53876 , n53877 , n53878 , n53879 , n53880 , n53881 , n53882 , n53883 , n53884 , n53885 , n53886 , n53887 , n53888 , n53889 , n53890 , n53891 , n53892 , n53893 , n53894 , n53895 , n53896 , n53897 , n53898 , n53899 , n53900 , n53901 , n53902 , n53904 , n53905 , n53906 , n53907 , n53908 , n53909 , n53910 , n53911 , n53912 , n53913 , n53914 , n53915 , n53916 , n53917 , n53918 , n53919 , n53920 , n53921 , n53922 , n53923 , n53924 , n53925 , n53926 , n53927 , n53928 , n53929 , n53930 , n53931 , n53932 , n53933 , n53934 , n53935 , n53936 , n53937 , n53938 , n53939 , n53940 , n53941 , n53942 , n53943 , n53944 , n53945 , n53946 , n53947 , n53948 , n53949 , n53950 , n53951 , n53952 , n53953 , n53954 , n53955 , n53956 , n53957 , n53958 , n53959 , n53960 , n53961 , n53962 , n53963 , n53964 , n53965 , n53966 , n53967 , n53968 , n53969 , n53970 , n53971 , n53972 , n53973 , n53974 , n53975 , n53976 , n53977 , n53978 , n53979 , n53980 , n53981 , n53982 , n53983 , n53984 , n53985 , n53986 , n53987 , n53988 , n53989 , n53990 , n53991 , n53992 , n53993 , n53994 , n53995 , n53996 , n53997 , n53998 , n53999 , n54000 , n54002 , n54003 , n54004 , n54005 , n54006 , n54007 , n54008 , n54009 , n54010 , n54011 , n54012 , n54013 , n54014 , n54015 , n54016 , n54017 , n54018 , n54019 , n54020 , n54021 , n54022 , n54023 , n54024 , n54025 , n54026 , n54027 , n54028 , n54029 , n54030 , n54031 , n54032 , n54033 , n54034 , n54035 , n54036 , n54037 , n54038 , n54039 , n54040 , n54041 , n54042 , n54043 , n54044 , n54045 , n54046 , n54047 , n54048 , n54049 , n54050 , n54051 , n54052 , n54053 , n54054 , n54055 , n54056 , n54057 , n54058 , n54059 , n54060 , n54061 , n54062 , n54063 , n54064 , n54065 , n54066 , n54067 , n54068 , n54069 , n54070 , n54071 , n54072 , n54073 , n54074 , n54075 , n54076 , n54077 , n54078 , n54079 , n54080 , n54082 , n54083 , n54084 , n54085 , n54086 , n54087 , n54088 , n54089 , n54090 , n54091 , n54092 , n54093 , n54094 , n54095 , n54096 , n54097 , n54098 , n54099 , n54100 , n54101 , n54102 , n54103 , n54104 , n54105 , n54106 , n54107 , n54108 , n54109 , n54110 , n54111 , n54112 , n54113 , n54114 , n54115 , n54116 , n54117 , n54118 , n54119 , n54120 , n54121 , n54122 , n54123 , n54124 , n54125 , n54126 , n54127 , n54128 , n54129 , n54130 , n54131 , n54132 , n54133 , n54134 , n54135 , n54136 , n54137 , n54138 , n54139 , n54140 , n54141 , n54142 , n54143 , n54144 , n54146 , n54147 , n54148 , n54149 , n54150 , n54151 , n54152 , n54153 , n54154 , n54155 , n54156 , n54157 , n54158 , n54159 , n54160 , n54161 , n54162 , n54163 , n54164 , n54165 , n54166 , n54167 , n54168 , n54169 , n54170 , n54171 , n54172 , n54173 , n54174 , n54175 , n54176 , n54177 , n54178 , n54179 , n54180 , n54181 , n54182 , n54183 , n54184 , n54185 , n54186 , n54187 , n54188 , n54189 , n54190 , n54191 , n54192 , n54193 , n54194 , n54195 , n54196 , n54197 , n54198 , n54199 , n54200 , n54202 , n54203 , n54204 , n54205 , n54206 , n54207 , n54208 , n54209 , n54210 , n54211 , n54212 , n54213 , n54214 , n54215 , n54216 , n54217 , n54218 , n54219 , n54220 , n54221 , n54222 , n54223 , n54224 , n54225 , n54226 , n54227 , n54228 , n54229 , n54230 , n54231 , n54232 , n54233 , n54234 , n54235 , n54236 , n54237 , n54238 , n54240 , n54241 , n54242 , n54243 , n54244 , n54245 , n54246 , n54247 , n54248 , n54249 , n54250 , n54251 , n54252 , n54253 , n54254 , n54255 , n54256 , n54257 , n54258 , n54259 , n54260 , n54262 , n54263 , n54264 ;
  assign n129 = x0 & x64 ;
  assign n130 = x2 & ~n129 ;
  assign n131 = ~x2 & ~n129 ;
  assign n132 = ~n130 & ~n131 ;
  assign n138 = n132 & x128 ;
  assign n133 = ~x0 & ~x64 ;
  assign n134 = ~x2 & ~n133 ;
  assign n135 = x2 & ~n133 ;
  assign n136 = ~n134 & ~n135 ;
  assign n139 = ~n136 & ~x128 ;
  assign n140 = ~n138 & ~n139 ;
  assign n141 = ~x0 & x1 ;
  assign n142 = x64 & n141 ;
  assign n143 = ~x1 & x2 ;
  assign n144 = x1 & ~x2 ;
  assign n145 = ~n143 & ~n144 ;
  assign n146 = x0 & n145 ;
  assign n147 = x65 & n146 ;
  assign n148 = ~n142 & ~n147 ;
  assign n149 = x0 & ~n145 ;
  assign n150 = x64 & ~x65 ;
  assign n151 = ~x64 & x65 ;
  assign n152 = ~n150 & ~n151 ;
  assign n153 = n149 & ~n152 ;
  assign n154 = n148 & ~n153 ;
  assign n155 = x2 & ~n154 ;
  assign n156 = x2 & ~n155 ;
  assign n157 = ~n154 & ~n155 ;
  assign n158 = ~n156 & ~n157 ;
  assign n159 = n130 & ~n158 ;
  assign n160 = ~n130 & n158 ;
  assign n161 = ~n159 & ~n160 ;
  assign n178 = n161 & x129 ;
  assign n162 = x0 & ~x1 ;
  assign n163 = ~x64 & n162 ;
  assign n164 = ~x0 & n145 ;
  assign n165 = ~x65 & n164 ;
  assign n166 = ~n163 & ~n165 ;
  assign n167 = ~x0 & ~n145 ;
  assign n168 = ~n152 & n167 ;
  assign n169 = n166 & ~n168 ;
  assign n170 = ~x2 & ~n169 ;
  assign n171 = ~x2 & ~n170 ;
  assign n172 = ~n169 & ~n170 ;
  assign n173 = ~n171 & ~n172 ;
  assign n174 = n134 & ~n173 ;
  assign n175 = ~n134 & n173 ;
  assign n176 = ~n174 & ~n175 ;
  assign n179 = ~n176 & ~x129 ;
  assign n180 = ~n178 & ~n179 ;
  assign n181 = x66 & n146 ;
  assign n182 = ~x1 & n167 ;
  assign n183 = x64 & n182 ;
  assign n184 = x65 & n141 ;
  assign n185 = ~n183 & ~n184 ;
  assign n186 = ~n181 & n185 ;
  assign n187 = x64 & ~x66 ;
  assign n188 = x65 & n187 ;
  assign n189 = x65 & ~x66 ;
  assign n190 = ~x65 & x66 ;
  assign n191 = ~n189 & ~n190 ;
  assign n192 = x64 & x65 ;
  assign n193 = n191 & ~n192 ;
  assign n194 = ~n188 & ~n193 ;
  assign n195 = n149 & n194 ;
  assign n196 = n186 & ~n195 ;
  assign n197 = x2 & ~n196 ;
  assign n198 = x2 & ~n197 ;
  assign n199 = ~n196 & ~n197 ;
  assign n200 = ~n198 & ~n199 ;
  assign n201 = n159 & ~n200 ;
  assign n202 = ~n159 & n200 ;
  assign n203 = ~n201 & ~n202 ;
  assign n225 = n203 & x130 ;
  assign n204 = ~x66 & n164 ;
  assign n205 = x1 & n149 ;
  assign n206 = ~x64 & n205 ;
  assign n207 = ~x65 & n162 ;
  assign n208 = ~n206 & ~n207 ;
  assign n209 = ~n204 & n208 ;
  assign n210 = ~x64 & x66 ;
  assign n211 = ~x65 & n210 ;
  assign n212 = ~x64 & ~x65 ;
  assign n213 = n191 & ~n212 ;
  assign n214 = ~n211 & ~n213 ;
  assign n215 = n167 & n214 ;
  assign n216 = n209 & ~n215 ;
  assign n217 = ~x2 & ~n216 ;
  assign n218 = ~x2 & ~n217 ;
  assign n219 = ~n216 & ~n217 ;
  assign n220 = ~n218 & ~n219 ;
  assign n221 = n174 & ~n220 ;
  assign n222 = ~n174 & n220 ;
  assign n223 = ~n221 & ~n222 ;
  assign n226 = ~n223 & ~x130 ;
  assign n227 = ~n225 & ~n226 ;
  assign n228 = x67 & n146 ;
  assign n229 = x65 & n182 ;
  assign n230 = x66 & n141 ;
  assign n231 = ~n229 & ~n230 ;
  assign n232 = ~n228 & n231 ;
  assign n233 = x65 & x66 ;
  assign n234 = ~n188 & ~n233 ;
  assign n235 = ~x66 & ~x67 ;
  assign n236 = x66 & x67 ;
  assign n237 = ~n235 & ~n236 ;
  assign n238 = ~n234 & n237 ;
  assign n239 = n234 & ~n237 ;
  assign n240 = ~n238 & ~n239 ;
  assign n241 = n149 & n240 ;
  assign n242 = n232 & ~n241 ;
  assign n243 = x2 & ~n242 ;
  assign n244 = x2 & ~n243 ;
  assign n245 = ~n242 & ~n243 ;
  assign n246 = ~n244 & ~n245 ;
  assign n247 = x2 & ~x3 ;
  assign n248 = ~x2 & x3 ;
  assign n249 = ~n247 & ~n248 ;
  assign n250 = x64 & ~n249 ;
  assign n251 = ~n246 & n250 ;
  assign n252 = n246 & ~n250 ;
  assign n253 = ~n251 & ~n252 ;
  assign n254 = n201 & n253 ;
  assign n255 = ~n201 & ~n253 ;
  assign n256 = ~n254 & ~n255 ;
  assign n281 = n256 & x131 ;
  assign n257 = ~x67 & n164 ;
  assign n258 = ~x65 & n205 ;
  assign n259 = ~x66 & n162 ;
  assign n260 = ~n258 & ~n259 ;
  assign n261 = ~n257 & n260 ;
  assign n262 = ~x65 & ~x66 ;
  assign n263 = ~n211 & ~n262 ;
  assign n264 = n237 & ~n263 ;
  assign n265 = ~n237 & n263 ;
  assign n266 = ~n264 & ~n265 ;
  assign n267 = n167 & n266 ;
  assign n268 = n261 & ~n267 ;
  assign n269 = ~x2 & ~n268 ;
  assign n270 = ~x2 & ~n269 ;
  assign n271 = ~n268 & ~n269 ;
  assign n272 = ~n270 & ~n271 ;
  assign n273 = ~x64 & ~n249 ;
  assign n274 = ~n272 & n273 ;
  assign n275 = n272 & ~n273 ;
  assign n276 = ~n274 & ~n275 ;
  assign n277 = n221 & n276 ;
  assign n278 = ~n221 & ~n276 ;
  assign n279 = ~n277 & ~n278 ;
  assign n282 = ~n279 & ~x131 ;
  assign n283 = ~n281 & ~n282 ;
  assign n284 = x5 & ~n250 ;
  assign n285 = ~x3 & x4 ;
  assign n286 = x3 & ~x4 ;
  assign n287 = ~n285 & ~n286 ;
  assign n288 = n249 & ~n287 ;
  assign n289 = x64 & n288 ;
  assign n290 = ~x4 & x5 ;
  assign n291 = x4 & ~x5 ;
  assign n292 = ~n290 & ~n291 ;
  assign n293 = ~n249 & n292 ;
  assign n294 = x65 & n293 ;
  assign n295 = ~n289 & ~n294 ;
  assign n296 = ~n249 & ~n292 ;
  assign n297 = ~n152 & n296 ;
  assign n298 = n295 & ~n297 ;
  assign n299 = x5 & ~n298 ;
  assign n300 = x5 & ~n299 ;
  assign n301 = ~n298 & ~n299 ;
  assign n302 = ~n300 & ~n301 ;
  assign n303 = n284 & ~n302 ;
  assign n304 = ~n284 & n302 ;
  assign n305 = ~n303 & ~n304 ;
  assign n306 = x68 & n146 ;
  assign n307 = x66 & n182 ;
  assign n308 = x67 & n141 ;
  assign n309 = ~n307 & ~n308 ;
  assign n310 = ~n306 & n309 ;
  assign n311 = ~n236 & ~n238 ;
  assign n312 = ~x67 & ~x68 ;
  assign n313 = x67 & x68 ;
  assign n314 = ~n312 & ~n313 ;
  assign n315 = ~n311 & n314 ;
  assign n316 = n311 & ~n314 ;
  assign n317 = ~n315 & ~n316 ;
  assign n318 = n149 & n317 ;
  assign n319 = n310 & ~n318 ;
  assign n320 = x2 & ~n319 ;
  assign n321 = x2 & ~n320 ;
  assign n322 = ~n319 & ~n320 ;
  assign n323 = ~n321 & ~n322 ;
  assign n324 = n305 & ~n323 ;
  assign n325 = n305 & ~n324 ;
  assign n326 = ~n323 & ~n324 ;
  assign n327 = ~n325 & ~n326 ;
  assign n328 = ~n251 & ~n254 ;
  assign n329 = ~n327 & ~n328 ;
  assign n330 = n327 & n328 ;
  assign n331 = ~n329 & ~n330 ;
  assign n368 = n331 & x132 ;
  assign n332 = ~x5 & ~n273 ;
  assign n333 = ~x64 & n288 ;
  assign n334 = ~x65 & n293 ;
  assign n335 = ~n333 & ~n334 ;
  assign n336 = ~n297 & n335 ;
  assign n337 = ~x5 & ~n336 ;
  assign n338 = ~x5 & ~n337 ;
  assign n339 = ~n336 & ~n337 ;
  assign n340 = ~n338 & ~n339 ;
  assign n341 = n332 & ~n340 ;
  assign n342 = ~n332 & n340 ;
  assign n343 = ~n341 & ~n342 ;
  assign n344 = ~x68 & n164 ;
  assign n345 = ~x66 & n205 ;
  assign n346 = ~x67 & n162 ;
  assign n347 = ~n345 & ~n346 ;
  assign n348 = ~n344 & n347 ;
  assign n349 = ~n235 & ~n264 ;
  assign n350 = n314 & ~n349 ;
  assign n351 = ~n314 & n349 ;
  assign n352 = ~n350 & ~n351 ;
  assign n353 = n167 & n352 ;
  assign n354 = n348 & ~n353 ;
  assign n355 = ~x2 & ~n354 ;
  assign n356 = ~x2 & ~n355 ;
  assign n357 = ~n354 & ~n355 ;
  assign n358 = ~n356 & ~n357 ;
  assign n359 = n343 & ~n358 ;
  assign n360 = n343 & ~n359 ;
  assign n361 = ~n358 & ~n359 ;
  assign n362 = ~n360 & ~n361 ;
  assign n363 = ~n274 & ~n277 ;
  assign n364 = ~n362 & ~n363 ;
  assign n365 = n362 & n363 ;
  assign n366 = ~n364 & ~n365 ;
  assign n369 = ~n366 & ~x132 ;
  assign n370 = ~n368 & ~n369 ;
  assign n371 = x66 & n293 ;
  assign n372 = n249 & ~n292 ;
  assign n373 = n287 & n372 ;
  assign n374 = x64 & n373 ;
  assign n375 = x65 & n288 ;
  assign n376 = ~n374 & ~n375 ;
  assign n377 = ~n371 & n376 ;
  assign n378 = ~n296 & n377 ;
  assign n379 = ~n194 & n377 ;
  assign n380 = ~n378 & ~n379 ;
  assign n381 = x5 & ~n380 ;
  assign n382 = ~x5 & n380 ;
  assign n383 = ~n381 & ~n382 ;
  assign n384 = n303 & ~n383 ;
  assign n385 = ~n303 & n383 ;
  assign n386 = ~n384 & ~n385 ;
  assign n387 = x69 & n146 ;
  assign n388 = x67 & n182 ;
  assign n389 = x68 & n141 ;
  assign n390 = ~n388 & ~n389 ;
  assign n391 = ~n387 & n390 ;
  assign n392 = ~n313 & ~n315 ;
  assign n393 = ~x68 & ~x69 ;
  assign n394 = x68 & x69 ;
  assign n395 = ~n393 & ~n394 ;
  assign n396 = ~n392 & n395 ;
  assign n397 = n392 & ~n395 ;
  assign n398 = ~n396 & ~n397 ;
  assign n399 = n149 & n398 ;
  assign n400 = n391 & ~n399 ;
  assign n401 = x2 & ~n400 ;
  assign n402 = x2 & ~n401 ;
  assign n403 = ~n400 & ~n401 ;
  assign n404 = ~n402 & ~n403 ;
  assign n405 = n386 & ~n404 ;
  assign n406 = n386 & ~n405 ;
  assign n407 = ~n404 & ~n405 ;
  assign n408 = ~n406 & ~n407 ;
  assign n409 = ~n324 & ~n329 ;
  assign n410 = ~n408 & ~n409 ;
  assign n411 = n408 & n409 ;
  assign n412 = ~n410 & ~n411 ;
  assign n451 = n412 & x133 ;
  assign n413 = ~x66 & n293 ;
  assign n414 = ~x64 & n373 ;
  assign n415 = ~x65 & n288 ;
  assign n416 = ~n414 & ~n415 ;
  assign n417 = ~n413 & n416 ;
  assign n418 = ~n296 & n417 ;
  assign n419 = ~n214 & n417 ;
  assign n420 = ~n418 & ~n419 ;
  assign n421 = ~x5 & ~n420 ;
  assign n422 = x5 & n420 ;
  assign n423 = ~n421 & ~n422 ;
  assign n424 = n341 & ~n423 ;
  assign n425 = ~n341 & n423 ;
  assign n426 = ~n424 & ~n425 ;
  assign n427 = ~x69 & n164 ;
  assign n428 = ~x67 & n205 ;
  assign n429 = ~x68 & n162 ;
  assign n430 = ~n428 & ~n429 ;
  assign n431 = ~n427 & n430 ;
  assign n432 = ~n312 & ~n350 ;
  assign n433 = n395 & ~n432 ;
  assign n434 = ~n395 & n432 ;
  assign n435 = ~n433 & ~n434 ;
  assign n436 = n167 & n435 ;
  assign n437 = n431 & ~n436 ;
  assign n438 = ~x2 & ~n437 ;
  assign n439 = ~x2 & ~n438 ;
  assign n440 = ~n437 & ~n438 ;
  assign n441 = ~n439 & ~n440 ;
  assign n442 = n426 & ~n441 ;
  assign n443 = n426 & ~n442 ;
  assign n444 = ~n441 & ~n442 ;
  assign n445 = ~n443 & ~n444 ;
  assign n446 = ~n359 & ~n364 ;
  assign n447 = ~n445 & ~n446 ;
  assign n448 = n445 & n446 ;
  assign n449 = ~n447 & ~n448 ;
  assign n452 = ~n449 & ~x133 ;
  assign n453 = ~n451 & ~n452 ;
  assign n454 = ~n405 & ~n410 ;
  assign n455 = x5 & ~x6 ;
  assign n456 = ~x5 & x6 ;
  assign n457 = ~n455 & ~n456 ;
  assign n458 = x64 & ~n457 ;
  assign n459 = n384 & n458 ;
  assign n460 = n384 & ~n459 ;
  assign n461 = n458 & ~n459 ;
  assign n462 = ~n460 & ~n461 ;
  assign n463 = x67 & n293 ;
  assign n464 = x65 & n373 ;
  assign n465 = x66 & n288 ;
  assign n466 = ~n464 & ~n465 ;
  assign n467 = ~n463 & n466 ;
  assign n468 = n240 & n296 ;
  assign n469 = n467 & ~n468 ;
  assign n470 = x5 & ~n469 ;
  assign n471 = x5 & ~n470 ;
  assign n472 = ~n469 & ~n470 ;
  assign n473 = ~n471 & ~n472 ;
  assign n474 = ~n462 & n473 ;
  assign n475 = n462 & ~n473 ;
  assign n476 = ~n474 & ~n475 ;
  assign n477 = x70 & n146 ;
  assign n478 = x68 & n182 ;
  assign n479 = x69 & n141 ;
  assign n480 = ~n478 & ~n479 ;
  assign n481 = ~n477 & n480 ;
  assign n482 = ~n394 & ~n396 ;
  assign n483 = ~x69 & ~x70 ;
  assign n484 = x69 & x70 ;
  assign n485 = ~n483 & ~n484 ;
  assign n486 = ~n482 & n485 ;
  assign n487 = n482 & ~n485 ;
  assign n488 = ~n486 & ~n487 ;
  assign n489 = n149 & n488 ;
  assign n490 = n481 & ~n489 ;
  assign n491 = x2 & ~n490 ;
  assign n492 = x2 & ~n491 ;
  assign n493 = ~n490 & ~n491 ;
  assign n494 = ~n492 & ~n493 ;
  assign n495 = ~n476 & ~n494 ;
  assign n496 = n476 & n494 ;
  assign n497 = ~n495 & ~n496 ;
  assign n498 = ~n454 & n497 ;
  assign n499 = n454 & ~n497 ;
  assign n500 = ~n498 & ~n499 ;
  assign n543 = n500 & x134 ;
  assign n501 = ~n442 & ~n447 ;
  assign n502 = ~x64 & ~n457 ;
  assign n503 = n424 & n502 ;
  assign n504 = n424 & ~n503 ;
  assign n505 = n502 & ~n503 ;
  assign n506 = ~n504 & ~n505 ;
  assign n507 = ~x67 & n293 ;
  assign n508 = ~x65 & n373 ;
  assign n509 = ~x66 & n288 ;
  assign n510 = ~n508 & ~n509 ;
  assign n511 = ~n507 & n510 ;
  assign n512 = n266 & n296 ;
  assign n513 = n511 & ~n512 ;
  assign n514 = ~x5 & ~n513 ;
  assign n515 = ~x5 & ~n514 ;
  assign n516 = ~n513 & ~n514 ;
  assign n517 = ~n515 & ~n516 ;
  assign n518 = ~n506 & n517 ;
  assign n519 = n506 & ~n517 ;
  assign n520 = ~n518 & ~n519 ;
  assign n521 = ~x70 & n164 ;
  assign n522 = ~x68 & n205 ;
  assign n523 = ~x69 & n162 ;
  assign n524 = ~n522 & ~n523 ;
  assign n525 = ~n521 & n524 ;
  assign n526 = ~n393 & ~n433 ;
  assign n527 = n485 & ~n526 ;
  assign n528 = ~n485 & n526 ;
  assign n529 = ~n527 & ~n528 ;
  assign n530 = n167 & n529 ;
  assign n531 = n525 & ~n530 ;
  assign n532 = ~x2 & ~n531 ;
  assign n533 = ~x2 & ~n532 ;
  assign n534 = ~n531 & ~n532 ;
  assign n535 = ~n533 & ~n534 ;
  assign n536 = ~n520 & ~n535 ;
  assign n537 = n520 & n535 ;
  assign n538 = ~n536 & ~n537 ;
  assign n539 = ~n501 & n538 ;
  assign n540 = n501 & ~n538 ;
  assign n541 = ~n539 & ~n540 ;
  assign n544 = ~n541 & ~x134 ;
  assign n545 = ~n543 & ~n544 ;
  assign n546 = ~n495 & ~n498 ;
  assign n547 = x71 & n146 ;
  assign n548 = x69 & n182 ;
  assign n549 = x70 & n141 ;
  assign n550 = ~n548 & ~n549 ;
  assign n551 = ~n547 & n550 ;
  assign n552 = ~n484 & ~n486 ;
  assign n553 = ~x70 & ~x71 ;
  assign n554 = x70 & x71 ;
  assign n555 = ~n553 & ~n554 ;
  assign n556 = ~n552 & n555 ;
  assign n557 = n552 & ~n555 ;
  assign n558 = ~n556 & ~n557 ;
  assign n559 = n149 & n558 ;
  assign n560 = n551 & ~n559 ;
  assign n561 = x2 & ~n560 ;
  assign n562 = x2 & ~n561 ;
  assign n563 = ~n560 & ~n561 ;
  assign n564 = ~n562 & ~n563 ;
  assign n565 = x8 & ~n458 ;
  assign n566 = ~x6 & x7 ;
  assign n567 = x6 & ~x7 ;
  assign n568 = ~n566 & ~n567 ;
  assign n569 = n457 & ~n568 ;
  assign n570 = x64 & n569 ;
  assign n571 = ~x7 & x8 ;
  assign n572 = x7 & ~x8 ;
  assign n573 = ~n571 & ~n572 ;
  assign n574 = ~n457 & n573 ;
  assign n575 = x65 & n574 ;
  assign n576 = ~n570 & ~n575 ;
  assign n577 = ~n457 & ~n573 ;
  assign n578 = ~n152 & n577 ;
  assign n579 = n576 & ~n578 ;
  assign n580 = x8 & ~n579 ;
  assign n581 = x8 & ~n580 ;
  assign n582 = ~n579 & ~n580 ;
  assign n583 = ~n581 & ~n582 ;
  assign n584 = n565 & ~n583 ;
  assign n585 = ~n565 & n583 ;
  assign n586 = ~n584 & ~n585 ;
  assign n587 = x68 & n293 ;
  assign n588 = x66 & n373 ;
  assign n589 = x67 & n288 ;
  assign n590 = ~n588 & ~n589 ;
  assign n591 = ~n587 & n590 ;
  assign n592 = n296 & n317 ;
  assign n593 = n591 & ~n592 ;
  assign n594 = x5 & ~n593 ;
  assign n595 = x5 & ~n594 ;
  assign n596 = ~n593 & ~n594 ;
  assign n597 = ~n595 & ~n596 ;
  assign n598 = n586 & ~n597 ;
  assign n599 = n586 & ~n598 ;
  assign n600 = ~n597 & ~n598 ;
  assign n601 = ~n599 & ~n600 ;
  assign n602 = ~n462 & ~n473 ;
  assign n603 = ~n459 & ~n602 ;
  assign n604 = ~n601 & ~n603 ;
  assign n605 = n601 & n603 ;
  assign n606 = ~n604 & ~n605 ;
  assign n607 = ~n564 & n606 ;
  assign n608 = n564 & ~n606 ;
  assign n609 = ~n607 & ~n608 ;
  assign n610 = ~n546 & n609 ;
  assign n611 = n546 & ~n609 ;
  assign n612 = ~n610 & ~n611 ;
  assign n668 = n612 & x135 ;
  assign n613 = ~n536 & ~n539 ;
  assign n614 = ~x71 & n164 ;
  assign n615 = ~x69 & n205 ;
  assign n616 = ~x70 & n162 ;
  assign n617 = ~n615 & ~n616 ;
  assign n618 = ~n614 & n617 ;
  assign n619 = ~n483 & ~n527 ;
  assign n620 = n555 & ~n619 ;
  assign n621 = ~n555 & n619 ;
  assign n622 = ~n620 & ~n621 ;
  assign n623 = n167 & n622 ;
  assign n624 = n618 & ~n623 ;
  assign n625 = ~x2 & ~n624 ;
  assign n626 = ~x2 & ~n625 ;
  assign n627 = ~n624 & ~n625 ;
  assign n628 = ~n626 & ~n627 ;
  assign n629 = ~x8 & ~n502 ;
  assign n630 = ~x64 & n569 ;
  assign n631 = ~x65 & n574 ;
  assign n632 = ~n630 & ~n631 ;
  assign n633 = ~n578 & n632 ;
  assign n634 = ~x8 & ~n633 ;
  assign n635 = ~x8 & ~n634 ;
  assign n636 = ~n633 & ~n634 ;
  assign n637 = ~n635 & ~n636 ;
  assign n638 = n629 & ~n637 ;
  assign n639 = ~n629 & n637 ;
  assign n640 = ~n638 & ~n639 ;
  assign n641 = ~x68 & n293 ;
  assign n642 = ~x66 & n373 ;
  assign n643 = ~x67 & n288 ;
  assign n644 = ~n642 & ~n643 ;
  assign n645 = ~n641 & n644 ;
  assign n646 = n296 & n352 ;
  assign n647 = n645 & ~n646 ;
  assign n648 = ~x5 & ~n647 ;
  assign n649 = ~x5 & ~n648 ;
  assign n650 = ~n647 & ~n648 ;
  assign n651 = ~n649 & ~n650 ;
  assign n652 = n640 & ~n651 ;
  assign n653 = n640 & ~n652 ;
  assign n654 = ~n651 & ~n652 ;
  assign n655 = ~n653 & ~n654 ;
  assign n656 = ~n506 & ~n517 ;
  assign n657 = ~n503 & ~n656 ;
  assign n658 = ~n655 & ~n657 ;
  assign n659 = n655 & n657 ;
  assign n660 = ~n658 & ~n659 ;
  assign n661 = ~n628 & n660 ;
  assign n662 = n628 & ~n660 ;
  assign n663 = ~n661 & ~n662 ;
  assign n664 = ~n613 & n663 ;
  assign n665 = n613 & ~n663 ;
  assign n666 = ~n664 & ~n665 ;
  assign n669 = ~n666 & ~x135 ;
  assign n670 = ~n668 & ~n669 ;
  assign n671 = x66 & n574 ;
  assign n672 = n457 & ~n573 ;
  assign n673 = n568 & n672 ;
  assign n674 = x64 & n673 ;
  assign n675 = x65 & n569 ;
  assign n676 = ~n674 & ~n675 ;
  assign n677 = ~n671 & n676 ;
  assign n678 = n194 & n577 ;
  assign n679 = n677 & ~n678 ;
  assign n680 = x8 & ~n679 ;
  assign n681 = x8 & ~n680 ;
  assign n682 = ~n679 & ~n680 ;
  assign n683 = ~n681 & ~n682 ;
  assign n684 = ~n584 & n683 ;
  assign n685 = n584 & ~n683 ;
  assign n686 = ~n684 & ~n685 ;
  assign n687 = x69 & n293 ;
  assign n688 = x67 & n373 ;
  assign n689 = x68 & n288 ;
  assign n690 = ~n688 & ~n689 ;
  assign n691 = ~n687 & n690 ;
  assign n692 = n296 & n398 ;
  assign n693 = n691 & ~n692 ;
  assign n694 = x5 & ~n693 ;
  assign n695 = x5 & ~n694 ;
  assign n696 = ~n693 & ~n694 ;
  assign n697 = ~n695 & ~n696 ;
  assign n698 = n686 & ~n697 ;
  assign n699 = n686 & ~n698 ;
  assign n700 = ~n697 & ~n698 ;
  assign n701 = ~n699 & ~n700 ;
  assign n702 = ~n598 & ~n604 ;
  assign n703 = n701 & n702 ;
  assign n704 = ~n701 & ~n702 ;
  assign n705 = ~n703 & ~n704 ;
  assign n706 = x72 & n146 ;
  assign n707 = x70 & n182 ;
  assign n708 = x71 & n141 ;
  assign n709 = ~n707 & ~n708 ;
  assign n710 = ~n706 & n709 ;
  assign n711 = ~n554 & ~n556 ;
  assign n712 = ~x71 & ~x72 ;
  assign n713 = x71 & x72 ;
  assign n714 = ~n712 & ~n713 ;
  assign n715 = ~n711 & n714 ;
  assign n716 = n711 & ~n714 ;
  assign n717 = ~n715 & ~n716 ;
  assign n718 = n149 & n717 ;
  assign n719 = n710 & ~n718 ;
  assign n720 = x2 & ~n719 ;
  assign n721 = x2 & ~n720 ;
  assign n722 = ~n719 & ~n720 ;
  assign n723 = ~n721 & ~n722 ;
  assign n724 = n705 & ~n723 ;
  assign n725 = n705 & ~n724 ;
  assign n726 = ~n723 & ~n724 ;
  assign n727 = ~n725 & ~n726 ;
  assign n728 = ~n607 & ~n610 ;
  assign n729 = ~n727 & ~n728 ;
  assign n730 = n727 & n728 ;
  assign n731 = ~n729 & ~n730 ;
  assign n789 = n731 & x136 ;
  assign n732 = ~x66 & n574 ;
  assign n733 = ~x64 & n673 ;
  assign n734 = ~x65 & n569 ;
  assign n735 = ~n733 & ~n734 ;
  assign n736 = ~n732 & n735 ;
  assign n737 = n214 & n577 ;
  assign n738 = n736 & ~n737 ;
  assign n739 = ~x8 & ~n738 ;
  assign n740 = ~x8 & ~n739 ;
  assign n741 = ~n738 & ~n739 ;
  assign n742 = ~n740 & ~n741 ;
  assign n743 = ~n638 & n742 ;
  assign n744 = n638 & ~n742 ;
  assign n745 = ~n743 & ~n744 ;
  assign n746 = ~x69 & n293 ;
  assign n747 = ~x67 & n373 ;
  assign n748 = ~x68 & n288 ;
  assign n749 = ~n747 & ~n748 ;
  assign n750 = ~n746 & n749 ;
  assign n751 = n296 & n435 ;
  assign n752 = n750 & ~n751 ;
  assign n753 = ~x5 & ~n752 ;
  assign n754 = ~x5 & ~n753 ;
  assign n755 = ~n752 & ~n753 ;
  assign n756 = ~n754 & ~n755 ;
  assign n757 = n745 & ~n756 ;
  assign n758 = n745 & ~n757 ;
  assign n759 = ~n756 & ~n757 ;
  assign n760 = ~n758 & ~n759 ;
  assign n761 = ~n652 & ~n658 ;
  assign n762 = n760 & n761 ;
  assign n763 = ~n760 & ~n761 ;
  assign n764 = ~n762 & ~n763 ;
  assign n765 = ~x72 & n164 ;
  assign n766 = ~x70 & n205 ;
  assign n767 = ~x71 & n162 ;
  assign n768 = ~n766 & ~n767 ;
  assign n769 = ~n765 & n768 ;
  assign n770 = ~n553 & ~n620 ;
  assign n771 = n714 & ~n770 ;
  assign n772 = ~n714 & n770 ;
  assign n773 = ~n771 & ~n772 ;
  assign n774 = n167 & n773 ;
  assign n775 = n769 & ~n774 ;
  assign n776 = ~x2 & ~n775 ;
  assign n777 = ~x2 & ~n776 ;
  assign n778 = ~n775 & ~n776 ;
  assign n779 = ~n777 & ~n778 ;
  assign n780 = n764 & ~n779 ;
  assign n781 = n764 & ~n780 ;
  assign n782 = ~n779 & ~n780 ;
  assign n783 = ~n781 & ~n782 ;
  assign n784 = ~n661 & ~n664 ;
  assign n785 = ~n783 & ~n784 ;
  assign n786 = n783 & n784 ;
  assign n787 = ~n785 & ~n786 ;
  assign n790 = ~n787 & ~x136 ;
  assign n791 = ~n789 & ~n790 ;
  assign n792 = x8 & ~x9 ;
  assign n793 = ~x8 & x9 ;
  assign n794 = ~n792 & ~n793 ;
  assign n795 = x64 & ~n794 ;
  assign n796 = ~n685 & n795 ;
  assign n797 = n685 & ~n795 ;
  assign n798 = ~n796 & ~n797 ;
  assign n799 = x67 & n574 ;
  assign n800 = x65 & n673 ;
  assign n801 = x66 & n569 ;
  assign n802 = ~n800 & ~n801 ;
  assign n803 = ~n799 & n802 ;
  assign n804 = n240 & n577 ;
  assign n805 = n803 & ~n804 ;
  assign n806 = x8 & ~n805 ;
  assign n807 = x8 & ~n806 ;
  assign n808 = ~n805 & ~n806 ;
  assign n809 = ~n807 & ~n808 ;
  assign n810 = ~n798 & ~n809 ;
  assign n811 = n798 & n809 ;
  assign n812 = ~n810 & ~n811 ;
  assign n813 = x70 & n293 ;
  assign n814 = x68 & n373 ;
  assign n815 = x69 & n288 ;
  assign n816 = ~n814 & ~n815 ;
  assign n817 = ~n813 & n816 ;
  assign n818 = n296 & n488 ;
  assign n819 = n817 & ~n818 ;
  assign n820 = x5 & ~n819 ;
  assign n821 = x5 & ~n820 ;
  assign n822 = ~n819 & ~n820 ;
  assign n823 = ~n821 & ~n822 ;
  assign n824 = n812 & ~n823 ;
  assign n825 = n812 & ~n824 ;
  assign n826 = ~n823 & ~n824 ;
  assign n827 = ~n825 & ~n826 ;
  assign n828 = ~n698 & ~n704 ;
  assign n829 = n827 & n828 ;
  assign n830 = ~n827 & ~n828 ;
  assign n831 = ~n829 & ~n830 ;
  assign n832 = x73 & n146 ;
  assign n833 = x71 & n182 ;
  assign n834 = x72 & n141 ;
  assign n835 = ~n833 & ~n834 ;
  assign n836 = ~n832 & n835 ;
  assign n837 = ~n713 & ~n715 ;
  assign n838 = ~x72 & ~x73 ;
  assign n839 = x72 & x73 ;
  assign n840 = ~n838 & ~n839 ;
  assign n841 = ~n837 & n840 ;
  assign n842 = n837 & ~n840 ;
  assign n843 = ~n841 & ~n842 ;
  assign n844 = n149 & n843 ;
  assign n845 = n836 & ~n844 ;
  assign n846 = x2 & ~n845 ;
  assign n847 = x2 & ~n846 ;
  assign n848 = ~n845 & ~n846 ;
  assign n849 = ~n847 & ~n848 ;
  assign n850 = n831 & ~n849 ;
  assign n851 = n831 & ~n850 ;
  assign n852 = ~n849 & ~n850 ;
  assign n853 = ~n851 & ~n852 ;
  assign n854 = ~n724 & ~n729 ;
  assign n855 = ~n853 & ~n854 ;
  assign n856 = n853 & n854 ;
  assign n857 = ~n855 & ~n856 ;
  assign n919 = n857 & x137 ;
  assign n858 = ~x64 & ~n794 ;
  assign n859 = ~n744 & n858 ;
  assign n860 = n744 & ~n858 ;
  assign n861 = ~n859 & ~n860 ;
  assign n862 = ~x67 & n574 ;
  assign n863 = ~x65 & n673 ;
  assign n864 = ~x66 & n569 ;
  assign n865 = ~n863 & ~n864 ;
  assign n866 = ~n862 & n865 ;
  assign n867 = n266 & n577 ;
  assign n868 = n866 & ~n867 ;
  assign n869 = ~x8 & ~n868 ;
  assign n870 = ~x8 & ~n869 ;
  assign n871 = ~n868 & ~n869 ;
  assign n872 = ~n870 & ~n871 ;
  assign n873 = ~n861 & ~n872 ;
  assign n874 = n861 & n872 ;
  assign n875 = ~n873 & ~n874 ;
  assign n876 = ~x70 & n293 ;
  assign n877 = ~x68 & n373 ;
  assign n878 = ~x69 & n288 ;
  assign n879 = ~n877 & ~n878 ;
  assign n880 = ~n876 & n879 ;
  assign n881 = n296 & n529 ;
  assign n882 = n880 & ~n881 ;
  assign n883 = ~x5 & ~n882 ;
  assign n884 = ~x5 & ~n883 ;
  assign n885 = ~n882 & ~n883 ;
  assign n886 = ~n884 & ~n885 ;
  assign n887 = n875 & ~n886 ;
  assign n888 = n875 & ~n887 ;
  assign n889 = ~n886 & ~n887 ;
  assign n890 = ~n888 & ~n889 ;
  assign n891 = ~n757 & ~n763 ;
  assign n892 = n890 & n891 ;
  assign n893 = ~n890 & ~n891 ;
  assign n894 = ~n892 & ~n893 ;
  assign n895 = ~x73 & n164 ;
  assign n896 = ~x71 & n205 ;
  assign n897 = ~x72 & n162 ;
  assign n898 = ~n896 & ~n897 ;
  assign n899 = ~n895 & n898 ;
  assign n900 = ~n712 & ~n771 ;
  assign n901 = n840 & ~n900 ;
  assign n902 = ~n840 & n900 ;
  assign n903 = ~n901 & ~n902 ;
  assign n904 = n167 & n903 ;
  assign n905 = n899 & ~n904 ;
  assign n906 = ~x2 & ~n905 ;
  assign n907 = ~x2 & ~n906 ;
  assign n908 = ~n905 & ~n906 ;
  assign n909 = ~n907 & ~n908 ;
  assign n910 = n894 & ~n909 ;
  assign n911 = n894 & ~n910 ;
  assign n912 = ~n909 & ~n910 ;
  assign n913 = ~n911 & ~n912 ;
  assign n914 = ~n780 & ~n785 ;
  assign n915 = ~n913 & ~n914 ;
  assign n916 = n913 & n914 ;
  assign n917 = ~n915 & ~n916 ;
  assign n920 = ~n917 & ~x137 ;
  assign n921 = ~n919 & ~n920 ;
  assign n922 = ~n850 & ~n855 ;
  assign n923 = n685 & n795 ;
  assign n924 = ~n810 & ~n923 ;
  assign n925 = x68 & n574 ;
  assign n926 = x66 & n673 ;
  assign n927 = x67 & n569 ;
  assign n928 = ~n926 & ~n927 ;
  assign n929 = ~n925 & n928 ;
  assign n930 = n317 & n577 ;
  assign n931 = n929 & ~n930 ;
  assign n932 = x8 & ~n931 ;
  assign n933 = x8 & ~n932 ;
  assign n934 = ~n931 & ~n932 ;
  assign n935 = ~n933 & ~n934 ;
  assign n936 = x11 & ~n795 ;
  assign n937 = ~x9 & x10 ;
  assign n938 = x9 & ~x10 ;
  assign n939 = ~n937 & ~n938 ;
  assign n940 = n794 & ~n939 ;
  assign n941 = x64 & n940 ;
  assign n942 = ~x10 & x11 ;
  assign n943 = x10 & ~x11 ;
  assign n944 = ~n942 & ~n943 ;
  assign n945 = ~n794 & n944 ;
  assign n946 = x65 & n945 ;
  assign n947 = ~n941 & ~n946 ;
  assign n948 = ~n794 & ~n944 ;
  assign n949 = ~n152 & n948 ;
  assign n950 = n947 & ~n949 ;
  assign n951 = x11 & ~n950 ;
  assign n952 = x11 & ~n951 ;
  assign n953 = ~n950 & ~n951 ;
  assign n954 = ~n952 & ~n953 ;
  assign n955 = n936 & ~n954 ;
  assign n956 = ~n936 & n954 ;
  assign n957 = ~n955 & ~n956 ;
  assign n958 = n935 & ~n957 ;
  assign n959 = ~n935 & n957 ;
  assign n960 = ~n958 & ~n959 ;
  assign n961 = ~n924 & n960 ;
  assign n962 = n924 & ~n960 ;
  assign n963 = ~n961 & ~n962 ;
  assign n964 = x71 & n293 ;
  assign n965 = x69 & n373 ;
  assign n966 = x70 & n288 ;
  assign n967 = ~n965 & ~n966 ;
  assign n968 = ~n964 & n967 ;
  assign n969 = n296 & n558 ;
  assign n970 = n968 & ~n969 ;
  assign n971 = x5 & ~n970 ;
  assign n972 = x5 & ~n971 ;
  assign n973 = ~n970 & ~n971 ;
  assign n974 = ~n972 & ~n973 ;
  assign n975 = n963 & ~n974 ;
  assign n976 = n963 & ~n975 ;
  assign n977 = ~n974 & ~n975 ;
  assign n978 = ~n976 & ~n977 ;
  assign n979 = ~n824 & ~n830 ;
  assign n980 = n978 & n979 ;
  assign n981 = ~n978 & ~n979 ;
  assign n982 = ~n980 & ~n981 ;
  assign n983 = x74 & n146 ;
  assign n984 = x72 & n182 ;
  assign n985 = x73 & n141 ;
  assign n986 = ~n984 & ~n985 ;
  assign n987 = ~n983 & n986 ;
  assign n988 = ~n839 & ~n841 ;
  assign n989 = ~x73 & ~x74 ;
  assign n990 = x73 & x74 ;
  assign n991 = ~n989 & ~n990 ;
  assign n992 = ~n988 & n991 ;
  assign n993 = n988 & ~n991 ;
  assign n994 = ~n992 & ~n993 ;
  assign n995 = n149 & n994 ;
  assign n996 = n987 & ~n995 ;
  assign n997 = x2 & ~n996 ;
  assign n998 = x2 & ~n997 ;
  assign n999 = ~n996 & ~n997 ;
  assign n1000 = ~n998 & ~n999 ;
  assign n1001 = ~n982 & n1000 ;
  assign n1002 = n982 & ~n1000 ;
  assign n1003 = ~n1001 & ~n1002 ;
  assign n1004 = ~n922 & n1003 ;
  assign n1005 = n922 & ~n1003 ;
  assign n1006 = ~n1004 & ~n1005 ;
  assign n1080 = n1006 & x138 ;
  assign n1007 = ~n910 & ~n915 ;
  assign n1008 = n744 & n858 ;
  assign n1009 = ~n873 & ~n1008 ;
  assign n1010 = ~x68 & n574 ;
  assign n1011 = ~x66 & n673 ;
  assign n1012 = ~x67 & n569 ;
  assign n1013 = ~n1011 & ~n1012 ;
  assign n1014 = ~n1010 & n1013 ;
  assign n1015 = n352 & n577 ;
  assign n1016 = n1014 & ~n1015 ;
  assign n1017 = ~x8 & ~n1016 ;
  assign n1018 = ~x8 & ~n1017 ;
  assign n1019 = ~n1016 & ~n1017 ;
  assign n1020 = ~n1018 & ~n1019 ;
  assign n1021 = ~x11 & ~n858 ;
  assign n1022 = ~x64 & n940 ;
  assign n1023 = ~x65 & n945 ;
  assign n1024 = ~n1022 & ~n1023 ;
  assign n1025 = ~n949 & n1024 ;
  assign n1026 = ~x11 & ~n1025 ;
  assign n1027 = ~x11 & ~n1026 ;
  assign n1028 = ~n1025 & ~n1026 ;
  assign n1029 = ~n1027 & ~n1028 ;
  assign n1030 = n1021 & ~n1029 ;
  assign n1031 = ~n1021 & n1029 ;
  assign n1032 = ~n1030 & ~n1031 ;
  assign n1033 = n1020 & ~n1032 ;
  assign n1034 = ~n1020 & n1032 ;
  assign n1035 = ~n1033 & ~n1034 ;
  assign n1036 = ~n1009 & n1035 ;
  assign n1037 = n1009 & ~n1035 ;
  assign n1038 = ~n1036 & ~n1037 ;
  assign n1039 = ~x71 & n293 ;
  assign n1040 = ~x69 & n373 ;
  assign n1041 = ~x70 & n288 ;
  assign n1042 = ~n1040 & ~n1041 ;
  assign n1043 = ~n1039 & n1042 ;
  assign n1044 = n296 & n622 ;
  assign n1045 = n1043 & ~n1044 ;
  assign n1046 = ~x5 & ~n1045 ;
  assign n1047 = ~x5 & ~n1046 ;
  assign n1048 = ~n1045 & ~n1046 ;
  assign n1049 = ~n1047 & ~n1048 ;
  assign n1050 = n1038 & ~n1049 ;
  assign n1051 = n1038 & ~n1050 ;
  assign n1052 = ~n1049 & ~n1050 ;
  assign n1053 = ~n1051 & ~n1052 ;
  assign n1054 = ~n887 & ~n893 ;
  assign n1055 = n1053 & n1054 ;
  assign n1056 = ~n1053 & ~n1054 ;
  assign n1057 = ~n1055 & ~n1056 ;
  assign n1058 = ~x74 & n164 ;
  assign n1059 = ~x72 & n205 ;
  assign n1060 = ~x73 & n162 ;
  assign n1061 = ~n1059 & ~n1060 ;
  assign n1062 = ~n1058 & n1061 ;
  assign n1063 = ~n838 & ~n901 ;
  assign n1064 = n991 & ~n1063 ;
  assign n1065 = ~n991 & n1063 ;
  assign n1066 = ~n1064 & ~n1065 ;
  assign n1067 = n167 & n1066 ;
  assign n1068 = n1062 & ~n1067 ;
  assign n1069 = ~x2 & ~n1068 ;
  assign n1070 = ~x2 & ~n1069 ;
  assign n1071 = ~n1068 & ~n1069 ;
  assign n1072 = ~n1070 & ~n1071 ;
  assign n1073 = ~n1057 & n1072 ;
  assign n1074 = n1057 & ~n1072 ;
  assign n1075 = ~n1073 & ~n1074 ;
  assign n1076 = ~n1007 & n1075 ;
  assign n1077 = n1007 & ~n1075 ;
  assign n1078 = ~n1076 & ~n1077 ;
  assign n1081 = ~n1078 & ~x138 ;
  assign n1082 = ~n1080 & ~n1081 ;
  assign n1083 = ~n1002 & ~n1004 ;
  assign n1084 = ~n975 & ~n981 ;
  assign n1085 = x72 & n293 ;
  assign n1086 = x70 & n373 ;
  assign n1087 = x71 & n288 ;
  assign n1088 = ~n1086 & ~n1087 ;
  assign n1089 = ~n1085 & n1088 ;
  assign n1090 = n296 & n717 ;
  assign n1091 = n1089 & ~n1090 ;
  assign n1092 = x5 & ~n1091 ;
  assign n1093 = x5 & ~n1092 ;
  assign n1094 = ~n1091 & ~n1092 ;
  assign n1095 = ~n1093 & ~n1094 ;
  assign n1096 = ~n959 & ~n961 ;
  assign n1097 = x66 & n945 ;
  assign n1098 = n794 & ~n944 ;
  assign n1099 = n939 & n1098 ;
  assign n1100 = x64 & n1099 ;
  assign n1101 = x65 & n940 ;
  assign n1102 = ~n1100 & ~n1101 ;
  assign n1103 = ~n1097 & n1102 ;
  assign n1104 = n194 & n948 ;
  assign n1105 = n1103 & ~n1104 ;
  assign n1106 = x11 & ~n1105 ;
  assign n1107 = x11 & ~n1106 ;
  assign n1108 = ~n1105 & ~n1106 ;
  assign n1109 = ~n1107 & ~n1108 ;
  assign n1110 = ~n955 & n1109 ;
  assign n1111 = n955 & ~n1109 ;
  assign n1112 = ~n1110 & ~n1111 ;
  assign n1113 = x69 & n574 ;
  assign n1114 = x67 & n673 ;
  assign n1115 = x68 & n569 ;
  assign n1116 = ~n1114 & ~n1115 ;
  assign n1117 = ~n1113 & n1116 ;
  assign n1118 = n398 & n577 ;
  assign n1119 = n1117 & ~n1118 ;
  assign n1120 = x8 & ~n1119 ;
  assign n1121 = x8 & ~n1120 ;
  assign n1122 = ~n1119 & ~n1120 ;
  assign n1123 = ~n1121 & ~n1122 ;
  assign n1124 = n1112 & ~n1123 ;
  assign n1125 = n1112 & ~n1124 ;
  assign n1126 = ~n1123 & ~n1124 ;
  assign n1127 = ~n1125 & ~n1126 ;
  assign n1128 = ~n1096 & ~n1127 ;
  assign n1129 = n1096 & n1127 ;
  assign n1130 = ~n1128 & ~n1129 ;
  assign n1131 = ~n1095 & n1130 ;
  assign n1132 = ~n1095 & ~n1131 ;
  assign n1133 = n1130 & ~n1131 ;
  assign n1134 = ~n1132 & ~n1133 ;
  assign n1135 = ~n1084 & ~n1134 ;
  assign n1136 = ~n1084 & ~n1135 ;
  assign n1137 = ~n1134 & ~n1135 ;
  assign n1138 = ~n1136 & ~n1137 ;
  assign n1139 = x75 & n146 ;
  assign n1140 = x73 & n182 ;
  assign n1141 = x74 & n141 ;
  assign n1142 = ~n1140 & ~n1141 ;
  assign n1143 = ~n1139 & n1142 ;
  assign n1144 = ~n990 & ~n992 ;
  assign n1145 = ~x74 & ~x75 ;
  assign n1146 = x74 & x75 ;
  assign n1147 = ~n1145 & ~n1146 ;
  assign n1148 = ~n1144 & n1147 ;
  assign n1149 = n1144 & ~n1147 ;
  assign n1150 = ~n1148 & ~n1149 ;
  assign n1151 = n149 & n1150 ;
  assign n1152 = n1143 & ~n1151 ;
  assign n1153 = x2 & ~n1152 ;
  assign n1154 = x2 & ~n1153 ;
  assign n1155 = ~n1152 & ~n1153 ;
  assign n1156 = ~n1154 & ~n1155 ;
  assign n1157 = ~n1138 & n1156 ;
  assign n1158 = n1138 & ~n1156 ;
  assign n1159 = ~n1157 & ~n1158 ;
  assign n1160 = ~n1083 & ~n1159 ;
  assign n1161 = n1083 & n1159 ;
  assign n1162 = ~n1160 & ~n1161 ;
  assign n1239 = n1162 & x139 ;
  assign n1163 = ~n1074 & ~n1076 ;
  assign n1164 = ~n1050 & ~n1056 ;
  assign n1165 = ~x72 & n293 ;
  assign n1166 = ~x70 & n373 ;
  assign n1167 = ~x71 & n288 ;
  assign n1168 = ~n1166 & ~n1167 ;
  assign n1169 = ~n1165 & n1168 ;
  assign n1170 = n296 & n773 ;
  assign n1171 = n1169 & ~n1170 ;
  assign n1172 = ~x5 & ~n1171 ;
  assign n1173 = ~x5 & ~n1172 ;
  assign n1174 = ~n1171 & ~n1172 ;
  assign n1175 = ~n1173 & ~n1174 ;
  assign n1176 = ~n1034 & ~n1036 ;
  assign n1177 = ~x66 & n945 ;
  assign n1178 = ~x64 & n1099 ;
  assign n1179 = ~x65 & n940 ;
  assign n1180 = ~n1178 & ~n1179 ;
  assign n1181 = ~n1177 & n1180 ;
  assign n1182 = n214 & n948 ;
  assign n1183 = n1181 & ~n1182 ;
  assign n1184 = ~x11 & ~n1183 ;
  assign n1185 = ~x11 & ~n1184 ;
  assign n1186 = ~n1183 & ~n1184 ;
  assign n1187 = ~n1185 & ~n1186 ;
  assign n1188 = ~n1030 & n1187 ;
  assign n1189 = n1030 & ~n1187 ;
  assign n1190 = ~n1188 & ~n1189 ;
  assign n1191 = ~x69 & n574 ;
  assign n1192 = ~x67 & n673 ;
  assign n1193 = ~x68 & n569 ;
  assign n1194 = ~n1192 & ~n1193 ;
  assign n1195 = ~n1191 & n1194 ;
  assign n1196 = n435 & n577 ;
  assign n1197 = n1195 & ~n1196 ;
  assign n1198 = ~x8 & ~n1197 ;
  assign n1199 = ~x8 & ~n1198 ;
  assign n1200 = ~n1197 & ~n1198 ;
  assign n1201 = ~n1199 & ~n1200 ;
  assign n1202 = n1190 & ~n1201 ;
  assign n1203 = n1190 & ~n1202 ;
  assign n1204 = ~n1201 & ~n1202 ;
  assign n1205 = ~n1203 & ~n1204 ;
  assign n1206 = ~n1176 & ~n1205 ;
  assign n1207 = n1176 & n1205 ;
  assign n1208 = ~n1206 & ~n1207 ;
  assign n1209 = ~n1175 & n1208 ;
  assign n1210 = ~n1175 & ~n1209 ;
  assign n1211 = n1208 & ~n1209 ;
  assign n1212 = ~n1210 & ~n1211 ;
  assign n1213 = ~n1164 & ~n1212 ;
  assign n1214 = ~n1164 & ~n1213 ;
  assign n1215 = ~n1212 & ~n1213 ;
  assign n1216 = ~n1214 & ~n1215 ;
  assign n1217 = ~x75 & n164 ;
  assign n1218 = ~x73 & n205 ;
  assign n1219 = ~x74 & n162 ;
  assign n1220 = ~n1218 & ~n1219 ;
  assign n1221 = ~n1217 & n1220 ;
  assign n1222 = ~n989 & ~n1064 ;
  assign n1223 = n1147 & ~n1222 ;
  assign n1224 = ~n1147 & n1222 ;
  assign n1225 = ~n1223 & ~n1224 ;
  assign n1226 = n167 & n1225 ;
  assign n1227 = n1221 & ~n1226 ;
  assign n1228 = ~x2 & ~n1227 ;
  assign n1229 = ~x2 & ~n1228 ;
  assign n1230 = ~n1227 & ~n1228 ;
  assign n1231 = ~n1229 & ~n1230 ;
  assign n1232 = ~n1216 & n1231 ;
  assign n1233 = n1216 & ~n1231 ;
  assign n1234 = ~n1232 & ~n1233 ;
  assign n1235 = ~n1163 & ~n1234 ;
  assign n1236 = n1163 & n1234 ;
  assign n1237 = ~n1235 & ~n1236 ;
  assign n1240 = ~n1237 & ~x139 ;
  assign n1241 = ~n1239 & ~n1240 ;
  assign n1242 = x11 & ~x12 ;
  assign n1243 = ~x11 & x12 ;
  assign n1244 = ~n1242 & ~n1243 ;
  assign n1245 = x64 & ~n1244 ;
  assign n1246 = ~n1111 & n1245 ;
  assign n1247 = n1111 & ~n1245 ;
  assign n1248 = ~n1246 & ~n1247 ;
  assign n1249 = x67 & n945 ;
  assign n1250 = x65 & n1099 ;
  assign n1251 = x66 & n940 ;
  assign n1252 = ~n1250 & ~n1251 ;
  assign n1253 = ~n1249 & n1252 ;
  assign n1254 = n240 & n948 ;
  assign n1255 = n1253 & ~n1254 ;
  assign n1256 = x11 & ~n1255 ;
  assign n1257 = x11 & ~n1256 ;
  assign n1258 = ~n1255 & ~n1256 ;
  assign n1259 = ~n1257 & ~n1258 ;
  assign n1260 = ~n1248 & ~n1259 ;
  assign n1261 = n1248 & n1259 ;
  assign n1262 = ~n1260 & ~n1261 ;
  assign n1263 = x70 & n574 ;
  assign n1264 = x68 & n673 ;
  assign n1265 = x69 & n569 ;
  assign n1266 = ~n1264 & ~n1265 ;
  assign n1267 = ~n1263 & n1266 ;
  assign n1268 = n488 & n577 ;
  assign n1269 = n1267 & ~n1268 ;
  assign n1270 = x8 & ~n1269 ;
  assign n1271 = x8 & ~n1270 ;
  assign n1272 = ~n1269 & ~n1270 ;
  assign n1273 = ~n1271 & ~n1272 ;
  assign n1274 = n1262 & ~n1273 ;
  assign n1275 = n1262 & ~n1274 ;
  assign n1276 = ~n1273 & ~n1274 ;
  assign n1277 = ~n1275 & ~n1276 ;
  assign n1278 = ~n1124 & ~n1128 ;
  assign n1279 = n1277 & n1278 ;
  assign n1280 = ~n1277 & ~n1278 ;
  assign n1281 = ~n1279 & ~n1280 ;
  assign n1282 = x73 & n293 ;
  assign n1283 = x71 & n373 ;
  assign n1284 = x72 & n288 ;
  assign n1285 = ~n1283 & ~n1284 ;
  assign n1286 = ~n1282 & n1285 ;
  assign n1287 = n296 & n843 ;
  assign n1288 = n1286 & ~n1287 ;
  assign n1289 = x5 & ~n1288 ;
  assign n1290 = x5 & ~n1289 ;
  assign n1291 = ~n1288 & ~n1289 ;
  assign n1292 = ~n1290 & ~n1291 ;
  assign n1293 = ~n1281 & n1292 ;
  assign n1294 = n1281 & ~n1292 ;
  assign n1295 = ~n1293 & ~n1294 ;
  assign n1296 = ~n1131 & ~n1135 ;
  assign n1297 = n1295 & ~n1296 ;
  assign n1298 = ~n1295 & n1296 ;
  assign n1299 = ~n1297 & ~n1298 ;
  assign n1300 = x76 & n146 ;
  assign n1301 = x74 & n182 ;
  assign n1302 = x75 & n141 ;
  assign n1303 = ~n1301 & ~n1302 ;
  assign n1304 = ~n1300 & n1303 ;
  assign n1305 = ~n1146 & ~n1148 ;
  assign n1306 = ~x75 & ~x76 ;
  assign n1307 = x75 & x76 ;
  assign n1308 = ~n1306 & ~n1307 ;
  assign n1309 = ~n1305 & n1308 ;
  assign n1310 = n1305 & ~n1308 ;
  assign n1311 = ~n1309 & ~n1310 ;
  assign n1312 = n149 & n1311 ;
  assign n1313 = n1304 & ~n1312 ;
  assign n1314 = x2 & ~n1313 ;
  assign n1315 = x2 & ~n1314 ;
  assign n1316 = ~n1313 & ~n1314 ;
  assign n1317 = ~n1315 & ~n1316 ;
  assign n1318 = n1299 & ~n1317 ;
  assign n1319 = n1299 & ~n1318 ;
  assign n1320 = ~n1317 & ~n1318 ;
  assign n1321 = ~n1319 & ~n1320 ;
  assign n1322 = ~n1138 & ~n1156 ;
  assign n1323 = ~n1160 & ~n1322 ;
  assign n1324 = ~n1321 & ~n1323 ;
  assign n1325 = n1321 & n1323 ;
  assign n1326 = ~n1324 & ~n1325 ;
  assign n1407 = n1326 & x140 ;
  assign n1327 = ~x64 & ~n1244 ;
  assign n1328 = ~n1189 & n1327 ;
  assign n1329 = n1189 & ~n1327 ;
  assign n1330 = ~n1328 & ~n1329 ;
  assign n1331 = ~x67 & n945 ;
  assign n1332 = ~x65 & n1099 ;
  assign n1333 = ~x66 & n940 ;
  assign n1334 = ~n1332 & ~n1333 ;
  assign n1335 = ~n1331 & n1334 ;
  assign n1336 = n266 & n948 ;
  assign n1337 = n1335 & ~n1336 ;
  assign n1338 = ~x11 & ~n1337 ;
  assign n1339 = ~x11 & ~n1338 ;
  assign n1340 = ~n1337 & ~n1338 ;
  assign n1341 = ~n1339 & ~n1340 ;
  assign n1342 = ~n1330 & ~n1341 ;
  assign n1343 = n1330 & n1341 ;
  assign n1344 = ~n1342 & ~n1343 ;
  assign n1345 = ~x70 & n574 ;
  assign n1346 = ~x68 & n673 ;
  assign n1347 = ~x69 & n569 ;
  assign n1348 = ~n1346 & ~n1347 ;
  assign n1349 = ~n1345 & n1348 ;
  assign n1350 = n529 & n577 ;
  assign n1351 = n1349 & ~n1350 ;
  assign n1352 = ~x8 & ~n1351 ;
  assign n1353 = ~x8 & ~n1352 ;
  assign n1354 = ~n1351 & ~n1352 ;
  assign n1355 = ~n1353 & ~n1354 ;
  assign n1356 = n1344 & ~n1355 ;
  assign n1357 = n1344 & ~n1356 ;
  assign n1358 = ~n1355 & ~n1356 ;
  assign n1359 = ~n1357 & ~n1358 ;
  assign n1360 = ~n1202 & ~n1206 ;
  assign n1361 = n1359 & n1360 ;
  assign n1362 = ~n1359 & ~n1360 ;
  assign n1363 = ~n1361 & ~n1362 ;
  assign n1364 = ~x73 & n293 ;
  assign n1365 = ~x71 & n373 ;
  assign n1366 = ~x72 & n288 ;
  assign n1367 = ~n1365 & ~n1366 ;
  assign n1368 = ~n1364 & n1367 ;
  assign n1369 = n296 & n903 ;
  assign n1370 = n1368 & ~n1369 ;
  assign n1371 = ~x5 & ~n1370 ;
  assign n1372 = ~x5 & ~n1371 ;
  assign n1373 = ~n1370 & ~n1371 ;
  assign n1374 = ~n1372 & ~n1373 ;
  assign n1375 = ~n1363 & n1374 ;
  assign n1376 = n1363 & ~n1374 ;
  assign n1377 = ~n1375 & ~n1376 ;
  assign n1378 = ~n1209 & ~n1213 ;
  assign n1379 = n1377 & ~n1378 ;
  assign n1380 = ~n1377 & n1378 ;
  assign n1381 = ~n1379 & ~n1380 ;
  assign n1382 = ~x76 & n164 ;
  assign n1383 = ~x74 & n205 ;
  assign n1384 = ~x75 & n162 ;
  assign n1385 = ~n1383 & ~n1384 ;
  assign n1386 = ~n1382 & n1385 ;
  assign n1387 = ~n1145 & ~n1223 ;
  assign n1388 = n1308 & ~n1387 ;
  assign n1389 = ~n1308 & n1387 ;
  assign n1390 = ~n1388 & ~n1389 ;
  assign n1391 = n167 & n1390 ;
  assign n1392 = n1386 & ~n1391 ;
  assign n1393 = ~x2 & ~n1392 ;
  assign n1394 = ~x2 & ~n1393 ;
  assign n1395 = ~n1392 & ~n1393 ;
  assign n1396 = ~n1394 & ~n1395 ;
  assign n1397 = n1381 & ~n1396 ;
  assign n1398 = n1381 & ~n1397 ;
  assign n1399 = ~n1396 & ~n1397 ;
  assign n1400 = ~n1398 & ~n1399 ;
  assign n1401 = ~n1216 & ~n1231 ;
  assign n1402 = ~n1235 & ~n1401 ;
  assign n1403 = ~n1400 & ~n1402 ;
  assign n1404 = n1400 & n1402 ;
  assign n1405 = ~n1403 & ~n1404 ;
  assign n1408 = ~n1405 & ~x140 ;
  assign n1409 = ~n1407 & ~n1408 ;
  assign n1410 = ~n1318 & ~n1324 ;
  assign n1411 = ~n1294 & ~n1297 ;
  assign n1412 = n1111 & n1245 ;
  assign n1413 = ~n1260 & ~n1412 ;
  assign n1414 = x68 & n945 ;
  assign n1415 = x66 & n1099 ;
  assign n1416 = x67 & n940 ;
  assign n1417 = ~n1415 & ~n1416 ;
  assign n1418 = ~n1414 & n1417 ;
  assign n1419 = n317 & n948 ;
  assign n1420 = n1418 & ~n1419 ;
  assign n1421 = x11 & ~n1420 ;
  assign n1422 = x11 & ~n1421 ;
  assign n1423 = ~n1420 & ~n1421 ;
  assign n1424 = ~n1422 & ~n1423 ;
  assign n1425 = x14 & ~n1245 ;
  assign n1426 = ~x12 & x13 ;
  assign n1427 = x12 & ~x13 ;
  assign n1428 = ~n1426 & ~n1427 ;
  assign n1429 = n1244 & ~n1428 ;
  assign n1430 = x64 & n1429 ;
  assign n1431 = ~x13 & x14 ;
  assign n1432 = x13 & ~x14 ;
  assign n1433 = ~n1431 & ~n1432 ;
  assign n1434 = ~n1244 & n1433 ;
  assign n1435 = x65 & n1434 ;
  assign n1436 = ~n1430 & ~n1435 ;
  assign n1437 = ~n1244 & ~n1433 ;
  assign n1438 = ~n152 & n1437 ;
  assign n1439 = n1436 & ~n1438 ;
  assign n1440 = x14 & ~n1439 ;
  assign n1441 = x14 & ~n1440 ;
  assign n1442 = ~n1439 & ~n1440 ;
  assign n1443 = ~n1441 & ~n1442 ;
  assign n1444 = n1425 & ~n1443 ;
  assign n1445 = ~n1425 & n1443 ;
  assign n1446 = ~n1444 & ~n1445 ;
  assign n1447 = n1424 & ~n1446 ;
  assign n1448 = ~n1424 & n1446 ;
  assign n1449 = ~n1447 & ~n1448 ;
  assign n1450 = ~n1413 & n1449 ;
  assign n1451 = n1413 & ~n1449 ;
  assign n1452 = ~n1450 & ~n1451 ;
  assign n1453 = x71 & n574 ;
  assign n1454 = x69 & n673 ;
  assign n1455 = x70 & n569 ;
  assign n1456 = ~n1454 & ~n1455 ;
  assign n1457 = ~n1453 & n1456 ;
  assign n1458 = n558 & n577 ;
  assign n1459 = n1457 & ~n1458 ;
  assign n1460 = x8 & ~n1459 ;
  assign n1461 = x8 & ~n1460 ;
  assign n1462 = ~n1459 & ~n1460 ;
  assign n1463 = ~n1461 & ~n1462 ;
  assign n1464 = n1452 & ~n1463 ;
  assign n1465 = n1452 & ~n1464 ;
  assign n1466 = ~n1463 & ~n1464 ;
  assign n1467 = ~n1465 & ~n1466 ;
  assign n1468 = ~n1274 & ~n1280 ;
  assign n1469 = n1467 & n1468 ;
  assign n1470 = ~n1467 & ~n1468 ;
  assign n1471 = ~n1469 & ~n1470 ;
  assign n1472 = x74 & n293 ;
  assign n1473 = x72 & n373 ;
  assign n1474 = x73 & n288 ;
  assign n1475 = ~n1473 & ~n1474 ;
  assign n1476 = ~n1472 & n1475 ;
  assign n1477 = n296 & n994 ;
  assign n1478 = n1476 & ~n1477 ;
  assign n1479 = x5 & ~n1478 ;
  assign n1480 = x5 & ~n1479 ;
  assign n1481 = ~n1478 & ~n1479 ;
  assign n1482 = ~n1480 & ~n1481 ;
  assign n1483 = n1471 & ~n1482 ;
  assign n1484 = ~n1471 & n1482 ;
  assign n1485 = ~n1411 & ~n1484 ;
  assign n1486 = ~n1483 & n1485 ;
  assign n1487 = ~n1411 & ~n1486 ;
  assign n1488 = ~n1483 & ~n1486 ;
  assign n1489 = ~n1484 & n1488 ;
  assign n1490 = ~n1487 & ~n1489 ;
  assign n1491 = x77 & n146 ;
  assign n1492 = x75 & n182 ;
  assign n1493 = x76 & n141 ;
  assign n1494 = ~n1492 & ~n1493 ;
  assign n1495 = ~n1491 & n1494 ;
  assign n1496 = ~n1307 & ~n1309 ;
  assign n1497 = ~x76 & ~x77 ;
  assign n1498 = x76 & x77 ;
  assign n1499 = ~n1497 & ~n1498 ;
  assign n1500 = ~n1496 & n1499 ;
  assign n1501 = n1496 & ~n1499 ;
  assign n1502 = ~n1500 & ~n1501 ;
  assign n1503 = n149 & n1502 ;
  assign n1504 = n1495 & ~n1503 ;
  assign n1505 = x2 & ~n1504 ;
  assign n1506 = x2 & ~n1505 ;
  assign n1507 = ~n1504 & ~n1505 ;
  assign n1508 = ~n1506 & ~n1507 ;
  assign n1509 = ~n1490 & n1508 ;
  assign n1510 = n1490 & ~n1508 ;
  assign n1511 = ~n1509 & ~n1510 ;
  assign n1512 = ~n1410 & ~n1511 ;
  assign n1513 = n1410 & n1511 ;
  assign n1514 = ~n1512 & ~n1513 ;
  assign n1608 = n1514 & x141 ;
  assign n1515 = ~n1397 & ~n1403 ;
  assign n1516 = ~n1376 & ~n1379 ;
  assign n1517 = n1189 & n1327 ;
  assign n1518 = ~n1342 & ~n1517 ;
  assign n1519 = ~x68 & n945 ;
  assign n1520 = ~x66 & n1099 ;
  assign n1521 = ~x67 & n940 ;
  assign n1522 = ~n1520 & ~n1521 ;
  assign n1523 = ~n1519 & n1522 ;
  assign n1524 = n352 & n948 ;
  assign n1525 = n1523 & ~n1524 ;
  assign n1526 = ~x11 & ~n1525 ;
  assign n1527 = ~x11 & ~n1526 ;
  assign n1528 = ~n1525 & ~n1526 ;
  assign n1529 = ~n1527 & ~n1528 ;
  assign n1530 = ~x14 & ~n1327 ;
  assign n1531 = ~x64 & n1429 ;
  assign n1532 = ~x65 & n1434 ;
  assign n1533 = ~n1531 & ~n1532 ;
  assign n1534 = ~n1438 & n1533 ;
  assign n1535 = ~x14 & ~n1534 ;
  assign n1536 = ~x14 & ~n1535 ;
  assign n1537 = ~n1534 & ~n1535 ;
  assign n1538 = ~n1536 & ~n1537 ;
  assign n1539 = n1530 & ~n1538 ;
  assign n1540 = ~n1530 & n1538 ;
  assign n1541 = ~n1539 & ~n1540 ;
  assign n1542 = n1529 & ~n1541 ;
  assign n1543 = ~n1529 & n1541 ;
  assign n1544 = ~n1542 & ~n1543 ;
  assign n1545 = ~n1518 & n1544 ;
  assign n1546 = n1518 & ~n1544 ;
  assign n1547 = ~n1545 & ~n1546 ;
  assign n1548 = ~x71 & n574 ;
  assign n1549 = ~x69 & n673 ;
  assign n1550 = ~x70 & n569 ;
  assign n1551 = ~n1549 & ~n1550 ;
  assign n1552 = ~n1548 & n1551 ;
  assign n1553 = n577 & n622 ;
  assign n1554 = n1552 & ~n1553 ;
  assign n1555 = ~x8 & ~n1554 ;
  assign n1556 = ~x8 & ~n1555 ;
  assign n1557 = ~n1554 & ~n1555 ;
  assign n1558 = ~n1556 & ~n1557 ;
  assign n1559 = n1547 & ~n1558 ;
  assign n1560 = n1547 & ~n1559 ;
  assign n1561 = ~n1558 & ~n1559 ;
  assign n1562 = ~n1560 & ~n1561 ;
  assign n1563 = ~n1356 & ~n1362 ;
  assign n1564 = n1562 & n1563 ;
  assign n1565 = ~n1562 & ~n1563 ;
  assign n1566 = ~n1564 & ~n1565 ;
  assign n1567 = ~x74 & n293 ;
  assign n1568 = ~x72 & n373 ;
  assign n1569 = ~x73 & n288 ;
  assign n1570 = ~n1568 & ~n1569 ;
  assign n1571 = ~n1567 & n1570 ;
  assign n1572 = n296 & n1066 ;
  assign n1573 = n1571 & ~n1572 ;
  assign n1574 = ~x5 & ~n1573 ;
  assign n1575 = ~x5 & ~n1574 ;
  assign n1576 = ~n1573 & ~n1574 ;
  assign n1577 = ~n1575 & ~n1576 ;
  assign n1578 = n1566 & ~n1577 ;
  assign n1579 = ~n1566 & n1577 ;
  assign n1580 = ~n1516 & ~n1579 ;
  assign n1581 = ~n1578 & n1580 ;
  assign n1582 = ~n1516 & ~n1581 ;
  assign n1583 = ~n1578 & ~n1581 ;
  assign n1584 = ~n1579 & n1583 ;
  assign n1585 = ~n1582 & ~n1584 ;
  assign n1586 = ~x77 & n164 ;
  assign n1587 = ~x75 & n205 ;
  assign n1588 = ~x76 & n162 ;
  assign n1589 = ~n1587 & ~n1588 ;
  assign n1590 = ~n1586 & n1589 ;
  assign n1591 = ~n1306 & ~n1388 ;
  assign n1592 = n1499 & ~n1591 ;
  assign n1593 = ~n1499 & n1591 ;
  assign n1594 = ~n1592 & ~n1593 ;
  assign n1595 = n167 & n1594 ;
  assign n1596 = n1590 & ~n1595 ;
  assign n1597 = ~x2 & ~n1596 ;
  assign n1598 = ~x2 & ~n1597 ;
  assign n1599 = ~n1596 & ~n1597 ;
  assign n1600 = ~n1598 & ~n1599 ;
  assign n1601 = ~n1585 & n1600 ;
  assign n1602 = n1585 & ~n1600 ;
  assign n1603 = ~n1601 & ~n1602 ;
  assign n1604 = ~n1515 & ~n1603 ;
  assign n1605 = n1515 & n1603 ;
  assign n1606 = ~n1604 & ~n1605 ;
  assign n1609 = ~n1606 & ~x141 ;
  assign n1610 = ~n1608 & ~n1609 ;
  assign n1611 = ~n1490 & ~n1508 ;
  assign n1612 = ~n1512 & ~n1611 ;
  assign n1613 = x78 & n146 ;
  assign n1614 = x76 & n182 ;
  assign n1615 = x77 & n141 ;
  assign n1616 = ~n1614 & ~n1615 ;
  assign n1617 = ~n1613 & n1616 ;
  assign n1618 = ~n1498 & ~n1500 ;
  assign n1619 = ~x77 & ~x78 ;
  assign n1620 = x77 & x78 ;
  assign n1621 = ~n1619 & ~n1620 ;
  assign n1622 = ~n1618 & n1621 ;
  assign n1623 = n1618 & ~n1621 ;
  assign n1624 = ~n1622 & ~n1623 ;
  assign n1625 = n149 & n1624 ;
  assign n1626 = n1617 & ~n1625 ;
  assign n1627 = x2 & ~n1626 ;
  assign n1628 = x2 & ~n1627 ;
  assign n1629 = ~n1626 & ~n1627 ;
  assign n1630 = ~n1628 & ~n1629 ;
  assign n1631 = x75 & n293 ;
  assign n1632 = x73 & n373 ;
  assign n1633 = x74 & n288 ;
  assign n1634 = ~n1632 & ~n1633 ;
  assign n1635 = ~n1631 & n1634 ;
  assign n1636 = n296 & n1150 ;
  assign n1637 = n1635 & ~n1636 ;
  assign n1638 = x5 & ~n1637 ;
  assign n1639 = x5 & ~n1638 ;
  assign n1640 = ~n1637 & ~n1638 ;
  assign n1641 = ~n1639 & ~n1640 ;
  assign n1642 = ~n1464 & ~n1470 ;
  assign n1643 = ~n1448 & ~n1450 ;
  assign n1644 = x66 & n1434 ;
  assign n1645 = n1244 & ~n1433 ;
  assign n1646 = n1428 & n1645 ;
  assign n1647 = x64 & n1646 ;
  assign n1648 = x65 & n1429 ;
  assign n1649 = ~n1647 & ~n1648 ;
  assign n1650 = ~n1644 & n1649 ;
  assign n1651 = n194 & n1437 ;
  assign n1652 = n1650 & ~n1651 ;
  assign n1653 = x14 & ~n1652 ;
  assign n1654 = x14 & ~n1653 ;
  assign n1655 = ~n1652 & ~n1653 ;
  assign n1656 = ~n1654 & ~n1655 ;
  assign n1657 = ~n1444 & n1656 ;
  assign n1658 = n1444 & ~n1656 ;
  assign n1659 = ~n1657 & ~n1658 ;
  assign n1660 = x69 & n945 ;
  assign n1661 = x67 & n1099 ;
  assign n1662 = x68 & n940 ;
  assign n1663 = ~n1661 & ~n1662 ;
  assign n1664 = ~n1660 & n1663 ;
  assign n1665 = n398 & n948 ;
  assign n1666 = n1664 & ~n1665 ;
  assign n1667 = x11 & ~n1666 ;
  assign n1668 = x11 & ~n1667 ;
  assign n1669 = ~n1666 & ~n1667 ;
  assign n1670 = ~n1668 & ~n1669 ;
  assign n1671 = n1659 & ~n1670 ;
  assign n1672 = ~n1659 & n1670 ;
  assign n1673 = ~n1643 & ~n1672 ;
  assign n1674 = ~n1671 & n1673 ;
  assign n1675 = ~n1643 & ~n1674 ;
  assign n1676 = ~n1671 & ~n1674 ;
  assign n1677 = ~n1672 & n1676 ;
  assign n1678 = ~n1675 & ~n1677 ;
  assign n1679 = x72 & n574 ;
  assign n1680 = x70 & n673 ;
  assign n1681 = x71 & n569 ;
  assign n1682 = ~n1680 & ~n1681 ;
  assign n1683 = ~n1679 & n1682 ;
  assign n1684 = n577 & n717 ;
  assign n1685 = n1683 & ~n1684 ;
  assign n1686 = x8 & ~n1685 ;
  assign n1687 = x8 & ~n1686 ;
  assign n1688 = ~n1685 & ~n1686 ;
  assign n1689 = ~n1687 & ~n1688 ;
  assign n1690 = n1678 & n1689 ;
  assign n1691 = ~n1678 & ~n1689 ;
  assign n1692 = ~n1690 & ~n1691 ;
  assign n1693 = ~n1642 & n1692 ;
  assign n1694 = n1642 & ~n1692 ;
  assign n1695 = ~n1693 & ~n1694 ;
  assign n1696 = n1641 & ~n1695 ;
  assign n1697 = ~n1641 & n1695 ;
  assign n1698 = ~n1696 & ~n1697 ;
  assign n1699 = ~n1488 & n1698 ;
  assign n1700 = n1488 & ~n1698 ;
  assign n1701 = ~n1699 & ~n1700 ;
  assign n1702 = n1630 & n1701 ;
  assign n1703 = ~n1630 & ~n1701 ;
  assign n1704 = ~n1702 & ~n1703 ;
  assign n1705 = ~n1612 & ~n1704 ;
  assign n1706 = n1612 & n1704 ;
  assign n1707 = ~n1705 & ~n1706 ;
  assign n1801 = n1707 & x142 ;
  assign n1708 = ~n1585 & ~n1600 ;
  assign n1709 = ~n1604 & ~n1708 ;
  assign n1710 = ~x78 & n164 ;
  assign n1711 = ~x76 & n205 ;
  assign n1712 = ~x77 & n162 ;
  assign n1713 = ~n1711 & ~n1712 ;
  assign n1714 = ~n1710 & n1713 ;
  assign n1715 = ~n1497 & ~n1592 ;
  assign n1716 = n1621 & ~n1715 ;
  assign n1717 = ~n1621 & n1715 ;
  assign n1718 = ~n1716 & ~n1717 ;
  assign n1719 = n167 & n1718 ;
  assign n1720 = n1714 & ~n1719 ;
  assign n1721 = ~x2 & ~n1720 ;
  assign n1722 = ~x2 & ~n1721 ;
  assign n1723 = ~n1720 & ~n1721 ;
  assign n1724 = ~n1722 & ~n1723 ;
  assign n1725 = ~x75 & n293 ;
  assign n1726 = ~x73 & n373 ;
  assign n1727 = ~x74 & n288 ;
  assign n1728 = ~n1726 & ~n1727 ;
  assign n1729 = ~n1725 & n1728 ;
  assign n1730 = n296 & n1225 ;
  assign n1731 = n1729 & ~n1730 ;
  assign n1732 = ~x5 & ~n1731 ;
  assign n1733 = ~x5 & ~n1732 ;
  assign n1734 = ~n1731 & ~n1732 ;
  assign n1735 = ~n1733 & ~n1734 ;
  assign n1736 = ~n1559 & ~n1565 ;
  assign n1737 = ~n1543 & ~n1545 ;
  assign n1738 = ~x66 & n1434 ;
  assign n1739 = ~x64 & n1646 ;
  assign n1740 = ~x65 & n1429 ;
  assign n1741 = ~n1739 & ~n1740 ;
  assign n1742 = ~n1738 & n1741 ;
  assign n1743 = n214 & n1437 ;
  assign n1744 = n1742 & ~n1743 ;
  assign n1745 = ~x14 & ~n1744 ;
  assign n1746 = ~x14 & ~n1745 ;
  assign n1747 = ~n1744 & ~n1745 ;
  assign n1748 = ~n1746 & ~n1747 ;
  assign n1749 = ~n1539 & n1748 ;
  assign n1750 = n1539 & ~n1748 ;
  assign n1751 = ~n1749 & ~n1750 ;
  assign n1752 = ~x69 & n945 ;
  assign n1753 = ~x67 & n1099 ;
  assign n1754 = ~x68 & n940 ;
  assign n1755 = ~n1753 & ~n1754 ;
  assign n1756 = ~n1752 & n1755 ;
  assign n1757 = n435 & n948 ;
  assign n1758 = n1756 & ~n1757 ;
  assign n1759 = ~x11 & ~n1758 ;
  assign n1760 = ~x11 & ~n1759 ;
  assign n1761 = ~n1758 & ~n1759 ;
  assign n1762 = ~n1760 & ~n1761 ;
  assign n1763 = n1751 & ~n1762 ;
  assign n1764 = ~n1751 & n1762 ;
  assign n1765 = ~n1737 & ~n1764 ;
  assign n1766 = ~n1763 & n1765 ;
  assign n1767 = ~n1737 & ~n1766 ;
  assign n1768 = ~n1763 & ~n1766 ;
  assign n1769 = ~n1764 & n1768 ;
  assign n1770 = ~n1767 & ~n1769 ;
  assign n1771 = ~x72 & n574 ;
  assign n1772 = ~x70 & n673 ;
  assign n1773 = ~x71 & n569 ;
  assign n1774 = ~n1772 & ~n1773 ;
  assign n1775 = ~n1771 & n1774 ;
  assign n1776 = n577 & n773 ;
  assign n1777 = n1775 & ~n1776 ;
  assign n1778 = ~x8 & ~n1777 ;
  assign n1779 = ~x8 & ~n1778 ;
  assign n1780 = ~n1777 & ~n1778 ;
  assign n1781 = ~n1779 & ~n1780 ;
  assign n1782 = n1770 & n1781 ;
  assign n1783 = ~n1770 & ~n1781 ;
  assign n1784 = ~n1782 & ~n1783 ;
  assign n1785 = ~n1736 & n1784 ;
  assign n1786 = n1736 & ~n1784 ;
  assign n1787 = ~n1785 & ~n1786 ;
  assign n1788 = n1735 & ~n1787 ;
  assign n1789 = ~n1735 & n1787 ;
  assign n1790 = ~n1788 & ~n1789 ;
  assign n1791 = ~n1583 & n1790 ;
  assign n1792 = n1583 & ~n1790 ;
  assign n1793 = ~n1791 & ~n1792 ;
  assign n1794 = n1724 & n1793 ;
  assign n1795 = ~n1724 & ~n1793 ;
  assign n1796 = ~n1794 & ~n1795 ;
  assign n1797 = ~n1709 & ~n1796 ;
  assign n1798 = n1709 & n1796 ;
  assign n1799 = ~n1797 & ~n1798 ;
  assign n1802 = ~n1799 & ~x142 ;
  assign n1803 = ~n1801 & ~n1802 ;
  assign n1804 = ~n1630 & n1701 ;
  assign n1805 = ~n1705 & ~n1804 ;
  assign n1806 = x79 & n146 ;
  assign n1807 = x77 & n182 ;
  assign n1808 = x78 & n141 ;
  assign n1809 = ~n1807 & ~n1808 ;
  assign n1810 = ~n1806 & n1809 ;
  assign n1811 = ~n1620 & ~n1622 ;
  assign n1812 = ~x78 & ~x79 ;
  assign n1813 = x78 & x79 ;
  assign n1814 = ~n1812 & ~n1813 ;
  assign n1815 = ~n1811 & n1814 ;
  assign n1816 = n1811 & ~n1814 ;
  assign n1817 = ~n1815 & ~n1816 ;
  assign n1818 = n149 & n1817 ;
  assign n1819 = n1810 & ~n1818 ;
  assign n1820 = x2 & ~n1819 ;
  assign n1821 = x2 & ~n1820 ;
  assign n1822 = ~n1819 & ~n1820 ;
  assign n1823 = ~n1821 & ~n1822 ;
  assign n1824 = ~n1697 & ~n1699 ;
  assign n1825 = x76 & n293 ;
  assign n1826 = x74 & n373 ;
  assign n1827 = x75 & n288 ;
  assign n1828 = ~n1826 & ~n1827 ;
  assign n1829 = ~n1825 & n1828 ;
  assign n1830 = n296 & n1311 ;
  assign n1831 = n1829 & ~n1830 ;
  assign n1832 = x5 & ~n1831 ;
  assign n1833 = x5 & ~n1832 ;
  assign n1834 = ~n1831 & ~n1832 ;
  assign n1835 = ~n1833 & ~n1834 ;
  assign n1836 = ~n1691 & ~n1693 ;
  assign n1837 = x73 & n574 ;
  assign n1838 = x71 & n673 ;
  assign n1839 = x72 & n569 ;
  assign n1840 = ~n1838 & ~n1839 ;
  assign n1841 = ~n1837 & n1840 ;
  assign n1842 = n577 & n843 ;
  assign n1843 = n1841 & ~n1842 ;
  assign n1844 = x8 & ~n1843 ;
  assign n1845 = x8 & ~n1844 ;
  assign n1846 = ~n1843 & ~n1844 ;
  assign n1847 = ~n1845 & ~n1846 ;
  assign n1848 = x14 & ~x15 ;
  assign n1849 = ~x14 & x15 ;
  assign n1850 = ~n1848 & ~n1849 ;
  assign n1851 = x64 & ~n1850 ;
  assign n1852 = ~n1658 & n1851 ;
  assign n1853 = n1658 & ~n1851 ;
  assign n1854 = ~n1852 & ~n1853 ;
  assign n1855 = x67 & n1434 ;
  assign n1856 = x65 & n1646 ;
  assign n1857 = x66 & n1429 ;
  assign n1858 = ~n1856 & ~n1857 ;
  assign n1859 = ~n1855 & n1858 ;
  assign n1860 = n240 & n1437 ;
  assign n1861 = n1859 & ~n1860 ;
  assign n1862 = x14 & ~n1861 ;
  assign n1863 = x14 & ~n1862 ;
  assign n1864 = ~n1861 & ~n1862 ;
  assign n1865 = ~n1863 & ~n1864 ;
  assign n1866 = ~n1854 & ~n1865 ;
  assign n1867 = n1854 & n1865 ;
  assign n1868 = ~n1866 & ~n1867 ;
  assign n1869 = x70 & n945 ;
  assign n1870 = x68 & n1099 ;
  assign n1871 = x69 & n940 ;
  assign n1872 = ~n1870 & ~n1871 ;
  assign n1873 = ~n1869 & n1872 ;
  assign n1874 = n488 & n948 ;
  assign n1875 = n1873 & ~n1874 ;
  assign n1876 = x11 & ~n1875 ;
  assign n1877 = x11 & ~n1876 ;
  assign n1878 = ~n1875 & ~n1876 ;
  assign n1879 = ~n1877 & ~n1878 ;
  assign n1880 = n1868 & ~n1879 ;
  assign n1881 = n1868 & ~n1880 ;
  assign n1882 = ~n1879 & ~n1880 ;
  assign n1883 = ~n1881 & ~n1882 ;
  assign n1884 = ~n1676 & ~n1883 ;
  assign n1885 = n1676 & n1883 ;
  assign n1886 = ~n1884 & ~n1885 ;
  assign n1887 = ~n1847 & n1886 ;
  assign n1888 = ~n1847 & ~n1887 ;
  assign n1889 = n1886 & ~n1887 ;
  assign n1890 = ~n1888 & ~n1889 ;
  assign n1891 = ~n1836 & ~n1890 ;
  assign n1892 = n1836 & ~n1889 ;
  assign n1893 = ~n1888 & n1892 ;
  assign n1894 = ~n1891 & ~n1893 ;
  assign n1895 = ~n1835 & n1894 ;
  assign n1896 = ~n1835 & ~n1895 ;
  assign n1897 = n1894 & ~n1895 ;
  assign n1898 = ~n1896 & ~n1897 ;
  assign n1899 = ~n1824 & ~n1898 ;
  assign n1900 = n1824 & ~n1897 ;
  assign n1901 = ~n1896 & n1900 ;
  assign n1902 = ~n1899 & ~n1901 ;
  assign n1903 = ~n1823 & n1902 ;
  assign n1904 = ~n1823 & ~n1903 ;
  assign n1905 = n1902 & ~n1903 ;
  assign n1906 = ~n1904 & ~n1905 ;
  assign n1907 = ~n1805 & ~n1906 ;
  assign n1908 = n1805 & ~n1905 ;
  assign n1909 = ~n1904 & n1908 ;
  assign n1910 = ~n1907 & ~n1909 ;
  assign n2013 = n1910 & x143 ;
  assign n1911 = ~n1724 & n1793 ;
  assign n1912 = ~n1797 & ~n1911 ;
  assign n1913 = ~x79 & n164 ;
  assign n1914 = ~x77 & n205 ;
  assign n1915 = ~x78 & n162 ;
  assign n1916 = ~n1914 & ~n1915 ;
  assign n1917 = ~n1913 & n1916 ;
  assign n1918 = ~n1619 & ~n1716 ;
  assign n1919 = n1814 & ~n1918 ;
  assign n1920 = ~n1814 & n1918 ;
  assign n1921 = ~n1919 & ~n1920 ;
  assign n1922 = n167 & n1921 ;
  assign n1923 = n1917 & ~n1922 ;
  assign n1924 = ~x2 & ~n1923 ;
  assign n1925 = ~x2 & ~n1924 ;
  assign n1926 = ~n1923 & ~n1924 ;
  assign n1927 = ~n1925 & ~n1926 ;
  assign n1928 = ~n1789 & ~n1791 ;
  assign n1929 = ~x76 & n293 ;
  assign n1930 = ~x74 & n373 ;
  assign n1931 = ~x75 & n288 ;
  assign n1932 = ~n1930 & ~n1931 ;
  assign n1933 = ~n1929 & n1932 ;
  assign n1934 = n296 & n1390 ;
  assign n1935 = n1933 & ~n1934 ;
  assign n1936 = ~x5 & ~n1935 ;
  assign n1937 = ~x5 & ~n1936 ;
  assign n1938 = ~n1935 & ~n1936 ;
  assign n1939 = ~n1937 & ~n1938 ;
  assign n1940 = ~n1783 & ~n1785 ;
  assign n1941 = ~x73 & n574 ;
  assign n1942 = ~x71 & n673 ;
  assign n1943 = ~x72 & n569 ;
  assign n1944 = ~n1942 & ~n1943 ;
  assign n1945 = ~n1941 & n1944 ;
  assign n1946 = n577 & n903 ;
  assign n1947 = n1945 & ~n1946 ;
  assign n1948 = ~x8 & ~n1947 ;
  assign n1949 = ~x8 & ~n1948 ;
  assign n1950 = ~n1947 & ~n1948 ;
  assign n1951 = ~n1949 & ~n1950 ;
  assign n1952 = ~x64 & ~n1850 ;
  assign n1953 = ~n1750 & n1952 ;
  assign n1954 = n1750 & ~n1952 ;
  assign n1955 = ~n1953 & ~n1954 ;
  assign n1956 = ~x67 & n1434 ;
  assign n1957 = ~x65 & n1646 ;
  assign n1958 = ~x66 & n1429 ;
  assign n1959 = ~n1957 & ~n1958 ;
  assign n1960 = ~n1956 & n1959 ;
  assign n1961 = n266 & n1437 ;
  assign n1962 = n1960 & ~n1961 ;
  assign n1963 = ~x14 & ~n1962 ;
  assign n1964 = ~x14 & ~n1963 ;
  assign n1965 = ~n1962 & ~n1963 ;
  assign n1966 = ~n1964 & ~n1965 ;
  assign n1967 = ~n1955 & ~n1966 ;
  assign n1968 = n1955 & n1966 ;
  assign n1969 = ~n1967 & ~n1968 ;
  assign n1970 = ~x70 & n945 ;
  assign n1971 = ~x68 & n1099 ;
  assign n1972 = ~x69 & n940 ;
  assign n1973 = ~n1971 & ~n1972 ;
  assign n1974 = ~n1970 & n1973 ;
  assign n1975 = n529 & n948 ;
  assign n1976 = n1974 & ~n1975 ;
  assign n1977 = ~x11 & ~n1976 ;
  assign n1978 = ~x11 & ~n1977 ;
  assign n1979 = ~n1976 & ~n1977 ;
  assign n1980 = ~n1978 & ~n1979 ;
  assign n1981 = n1969 & ~n1980 ;
  assign n1982 = n1969 & ~n1981 ;
  assign n1983 = ~n1980 & ~n1981 ;
  assign n1984 = ~n1982 & ~n1983 ;
  assign n1985 = ~n1768 & ~n1984 ;
  assign n1986 = n1768 & n1984 ;
  assign n1987 = ~n1985 & ~n1986 ;
  assign n1988 = ~n1951 & n1987 ;
  assign n1989 = ~n1951 & ~n1988 ;
  assign n1990 = n1987 & ~n1988 ;
  assign n1991 = ~n1989 & ~n1990 ;
  assign n1992 = ~n1940 & ~n1991 ;
  assign n1993 = n1940 & ~n1990 ;
  assign n1994 = ~n1989 & n1993 ;
  assign n1995 = ~n1992 & ~n1994 ;
  assign n1996 = ~n1939 & n1995 ;
  assign n1997 = ~n1939 & ~n1996 ;
  assign n1998 = n1995 & ~n1996 ;
  assign n1999 = ~n1997 & ~n1998 ;
  assign n2000 = ~n1928 & ~n1999 ;
  assign n2001 = n1928 & ~n1998 ;
  assign n2002 = ~n1997 & n2001 ;
  assign n2003 = ~n2000 & ~n2002 ;
  assign n2004 = ~n1927 & n2003 ;
  assign n2005 = ~n1927 & ~n2004 ;
  assign n2006 = n2003 & ~n2004 ;
  assign n2007 = ~n2005 & ~n2006 ;
  assign n2008 = ~n1912 & ~n2007 ;
  assign n2009 = n1912 & ~n2006 ;
  assign n2010 = ~n2005 & n2009 ;
  assign n2011 = ~n2008 & ~n2010 ;
  assign n2014 = ~n2011 & ~x143 ;
  assign n2015 = ~n2013 & ~n2014 ;
  assign n2016 = ~n1903 & ~n1907 ;
  assign n2017 = x80 & n146 ;
  assign n2018 = x78 & n182 ;
  assign n2019 = x79 & n141 ;
  assign n2020 = ~n2018 & ~n2019 ;
  assign n2021 = ~n2017 & n2020 ;
  assign n2022 = ~n1813 & ~n1815 ;
  assign n2023 = ~x79 & ~x80 ;
  assign n2024 = x79 & x80 ;
  assign n2025 = ~n2023 & ~n2024 ;
  assign n2026 = ~n2022 & n2025 ;
  assign n2027 = n2022 & ~n2025 ;
  assign n2028 = ~n2026 & ~n2027 ;
  assign n2029 = n149 & n2028 ;
  assign n2030 = n2021 & ~n2029 ;
  assign n2031 = x2 & ~n2030 ;
  assign n2032 = x2 & ~n2031 ;
  assign n2033 = ~n2030 & ~n2031 ;
  assign n2034 = ~n2032 & ~n2033 ;
  assign n2035 = ~n1895 & ~n1899 ;
  assign n2036 = x77 & n293 ;
  assign n2037 = x75 & n373 ;
  assign n2038 = x76 & n288 ;
  assign n2039 = ~n2037 & ~n2038 ;
  assign n2040 = ~n2036 & n2039 ;
  assign n2041 = n296 & n1502 ;
  assign n2042 = n2040 & ~n2041 ;
  assign n2043 = x5 & ~n2042 ;
  assign n2044 = x5 & ~n2043 ;
  assign n2045 = ~n2042 & ~n2043 ;
  assign n2046 = ~n2044 & ~n2045 ;
  assign n2047 = ~n1887 & ~n1891 ;
  assign n2048 = x74 & n574 ;
  assign n2049 = x72 & n673 ;
  assign n2050 = x73 & n569 ;
  assign n2051 = ~n2049 & ~n2050 ;
  assign n2052 = ~n2048 & n2051 ;
  assign n2053 = n577 & n994 ;
  assign n2054 = n2052 & ~n2053 ;
  assign n2055 = x8 & ~n2054 ;
  assign n2056 = x8 & ~n2055 ;
  assign n2057 = ~n2054 & ~n2055 ;
  assign n2058 = ~n2056 & ~n2057 ;
  assign n2059 = ~n1880 & ~n1884 ;
  assign n2060 = x71 & n945 ;
  assign n2061 = x69 & n1099 ;
  assign n2062 = x70 & n940 ;
  assign n2063 = ~n2061 & ~n2062 ;
  assign n2064 = ~n2060 & n2063 ;
  assign n2065 = n558 & n948 ;
  assign n2066 = n2064 & ~n2065 ;
  assign n2067 = x11 & ~n2066 ;
  assign n2068 = x11 & ~n2067 ;
  assign n2069 = ~n2066 & ~n2067 ;
  assign n2070 = ~n2068 & ~n2069 ;
  assign n2071 = n1658 & n1851 ;
  assign n2072 = ~n1866 & ~n2071 ;
  assign n2073 = x68 & n1434 ;
  assign n2074 = x66 & n1646 ;
  assign n2075 = x67 & n1429 ;
  assign n2076 = ~n2074 & ~n2075 ;
  assign n2077 = ~n2073 & n2076 ;
  assign n2078 = n317 & n1437 ;
  assign n2079 = n2077 & ~n2078 ;
  assign n2080 = x14 & ~n2079 ;
  assign n2081 = x14 & ~n2080 ;
  assign n2082 = ~n2079 & ~n2080 ;
  assign n2083 = ~n2081 & ~n2082 ;
  assign n2084 = x17 & ~n1851 ;
  assign n2085 = ~x15 & x16 ;
  assign n2086 = x15 & ~x16 ;
  assign n2087 = ~n2085 & ~n2086 ;
  assign n2088 = n1850 & ~n2087 ;
  assign n2089 = x64 & n2088 ;
  assign n2090 = ~x16 & x17 ;
  assign n2091 = x16 & ~x17 ;
  assign n2092 = ~n2090 & ~n2091 ;
  assign n2093 = ~n1850 & n2092 ;
  assign n2094 = x65 & n2093 ;
  assign n2095 = ~n2089 & ~n2094 ;
  assign n2096 = ~n1850 & ~n2092 ;
  assign n2097 = ~n152 & n2096 ;
  assign n2098 = n2095 & ~n2097 ;
  assign n2099 = x17 & ~n2098 ;
  assign n2100 = x17 & ~n2099 ;
  assign n2101 = ~n2098 & ~n2099 ;
  assign n2102 = ~n2100 & ~n2101 ;
  assign n2103 = n2084 & ~n2102 ;
  assign n2104 = ~n2084 & n2102 ;
  assign n2105 = ~n2103 & ~n2104 ;
  assign n2106 = n2083 & ~n2105 ;
  assign n2107 = ~n2083 & n2105 ;
  assign n2108 = ~n2106 & ~n2107 ;
  assign n2109 = ~n2072 & n2108 ;
  assign n2110 = n2072 & ~n2108 ;
  assign n2111 = ~n2109 & ~n2110 ;
  assign n2112 = n2070 & ~n2111 ;
  assign n2113 = ~n2070 & n2111 ;
  assign n2114 = ~n2112 & ~n2113 ;
  assign n2115 = ~n2059 & n2114 ;
  assign n2116 = n2059 & ~n2114 ;
  assign n2117 = ~n2115 & ~n2116 ;
  assign n2118 = n2058 & ~n2117 ;
  assign n2119 = ~n2058 & n2117 ;
  assign n2120 = ~n2118 & ~n2119 ;
  assign n2121 = ~n2047 & n2120 ;
  assign n2122 = n2047 & ~n2120 ;
  assign n2123 = ~n2121 & ~n2122 ;
  assign n2124 = n2046 & ~n2123 ;
  assign n2125 = ~n2046 & n2123 ;
  assign n2126 = ~n2124 & ~n2125 ;
  assign n2127 = ~n2035 & n2126 ;
  assign n2128 = n2035 & ~n2126 ;
  assign n2129 = ~n2127 & ~n2128 ;
  assign n2130 = n2034 & n2129 ;
  assign n2131 = ~n2034 & ~n2129 ;
  assign n2132 = ~n2130 & ~n2131 ;
  assign n2133 = ~n2016 & ~n2132 ;
  assign n2134 = n2016 & n2132 ;
  assign n2135 = ~n2133 & ~n2134 ;
  assign n2244 = n2135 & x144 ;
  assign n2136 = ~n2004 & ~n2008 ;
  assign n2137 = ~x80 & n164 ;
  assign n2138 = ~x78 & n205 ;
  assign n2139 = ~x79 & n162 ;
  assign n2140 = ~n2138 & ~n2139 ;
  assign n2141 = ~n2137 & n2140 ;
  assign n2142 = ~n1812 & ~n1919 ;
  assign n2143 = n2025 & ~n2142 ;
  assign n2144 = ~n2025 & n2142 ;
  assign n2145 = ~n2143 & ~n2144 ;
  assign n2146 = n167 & n2145 ;
  assign n2147 = n2141 & ~n2146 ;
  assign n2148 = ~x2 & ~n2147 ;
  assign n2149 = ~x2 & ~n2148 ;
  assign n2150 = ~n2147 & ~n2148 ;
  assign n2151 = ~n2149 & ~n2150 ;
  assign n2152 = ~n1996 & ~n2000 ;
  assign n2153 = ~x77 & n293 ;
  assign n2154 = ~x75 & n373 ;
  assign n2155 = ~x76 & n288 ;
  assign n2156 = ~n2154 & ~n2155 ;
  assign n2157 = ~n2153 & n2156 ;
  assign n2158 = n296 & n1594 ;
  assign n2159 = n2157 & ~n2158 ;
  assign n2160 = ~x5 & ~n2159 ;
  assign n2161 = ~x5 & ~n2160 ;
  assign n2162 = ~n2159 & ~n2160 ;
  assign n2163 = ~n2161 & ~n2162 ;
  assign n2164 = ~n1988 & ~n1992 ;
  assign n2165 = ~x74 & n574 ;
  assign n2166 = ~x72 & n673 ;
  assign n2167 = ~x73 & n569 ;
  assign n2168 = ~n2166 & ~n2167 ;
  assign n2169 = ~n2165 & n2168 ;
  assign n2170 = n577 & n1066 ;
  assign n2171 = n2169 & ~n2170 ;
  assign n2172 = ~x8 & ~n2171 ;
  assign n2173 = ~x8 & ~n2172 ;
  assign n2174 = ~n2171 & ~n2172 ;
  assign n2175 = ~n2173 & ~n2174 ;
  assign n2176 = ~n1981 & ~n1985 ;
  assign n2177 = ~x71 & n945 ;
  assign n2178 = ~x69 & n1099 ;
  assign n2179 = ~x70 & n940 ;
  assign n2180 = ~n2178 & ~n2179 ;
  assign n2181 = ~n2177 & n2180 ;
  assign n2182 = n622 & n948 ;
  assign n2183 = n2181 & ~n2182 ;
  assign n2184 = ~x11 & ~n2183 ;
  assign n2185 = ~x11 & ~n2184 ;
  assign n2186 = ~n2183 & ~n2184 ;
  assign n2187 = ~n2185 & ~n2186 ;
  assign n2188 = n1750 & n1952 ;
  assign n2189 = ~n1967 & ~n2188 ;
  assign n2190 = ~x68 & n1434 ;
  assign n2191 = ~x66 & n1646 ;
  assign n2192 = ~x67 & n1429 ;
  assign n2193 = ~n2191 & ~n2192 ;
  assign n2194 = ~n2190 & n2193 ;
  assign n2195 = n352 & n1437 ;
  assign n2196 = n2194 & ~n2195 ;
  assign n2197 = ~x14 & ~n2196 ;
  assign n2198 = ~x14 & ~n2197 ;
  assign n2199 = ~n2196 & ~n2197 ;
  assign n2200 = ~n2198 & ~n2199 ;
  assign n2201 = ~x17 & ~n1952 ;
  assign n2202 = ~x64 & n2088 ;
  assign n2203 = ~x65 & n2093 ;
  assign n2204 = ~n2202 & ~n2203 ;
  assign n2205 = ~n2097 & n2204 ;
  assign n2206 = ~x17 & ~n2205 ;
  assign n2207 = ~x17 & ~n2206 ;
  assign n2208 = ~n2205 & ~n2206 ;
  assign n2209 = ~n2207 & ~n2208 ;
  assign n2210 = n2201 & ~n2209 ;
  assign n2211 = ~n2201 & n2209 ;
  assign n2212 = ~n2210 & ~n2211 ;
  assign n2213 = n2200 & ~n2212 ;
  assign n2214 = ~n2200 & n2212 ;
  assign n2215 = ~n2213 & ~n2214 ;
  assign n2216 = ~n2189 & n2215 ;
  assign n2217 = n2189 & ~n2215 ;
  assign n2218 = ~n2216 & ~n2217 ;
  assign n2219 = n2187 & ~n2218 ;
  assign n2220 = ~n2187 & n2218 ;
  assign n2221 = ~n2219 & ~n2220 ;
  assign n2222 = ~n2176 & n2221 ;
  assign n2223 = n2176 & ~n2221 ;
  assign n2224 = ~n2222 & ~n2223 ;
  assign n2225 = n2175 & ~n2224 ;
  assign n2226 = ~n2175 & n2224 ;
  assign n2227 = ~n2225 & ~n2226 ;
  assign n2228 = ~n2164 & n2227 ;
  assign n2229 = n2164 & ~n2227 ;
  assign n2230 = ~n2228 & ~n2229 ;
  assign n2231 = n2163 & ~n2230 ;
  assign n2232 = ~n2163 & n2230 ;
  assign n2233 = ~n2231 & ~n2232 ;
  assign n2234 = ~n2152 & n2233 ;
  assign n2235 = n2152 & ~n2233 ;
  assign n2236 = ~n2234 & ~n2235 ;
  assign n2237 = n2151 & n2236 ;
  assign n2238 = ~n2151 & ~n2236 ;
  assign n2239 = ~n2237 & ~n2238 ;
  assign n2240 = ~n2136 & ~n2239 ;
  assign n2241 = n2136 & n2239 ;
  assign n2242 = ~n2240 & ~n2241 ;
  assign n2245 = ~n2242 & ~x144 ;
  assign n2246 = ~n2244 & ~n2245 ;
  assign n2247 = ~n2125 & ~n2127 ;
  assign n2248 = x78 & n293 ;
  assign n2249 = x76 & n373 ;
  assign n2250 = x77 & n288 ;
  assign n2251 = ~n2249 & ~n2250 ;
  assign n2252 = ~n2248 & n2251 ;
  assign n2253 = n296 & n1624 ;
  assign n2254 = n2252 & ~n2253 ;
  assign n2255 = x5 & ~n2254 ;
  assign n2256 = x5 & ~n2255 ;
  assign n2257 = ~n2254 & ~n2255 ;
  assign n2258 = ~n2256 & ~n2257 ;
  assign n2259 = ~n2119 & ~n2121 ;
  assign n2260 = x75 & n574 ;
  assign n2261 = x73 & n673 ;
  assign n2262 = x74 & n569 ;
  assign n2263 = ~n2261 & ~n2262 ;
  assign n2264 = ~n2260 & n2263 ;
  assign n2265 = n577 & n1150 ;
  assign n2266 = n2264 & ~n2265 ;
  assign n2267 = x8 & ~n2266 ;
  assign n2268 = x8 & ~n2267 ;
  assign n2269 = ~n2266 & ~n2267 ;
  assign n2270 = ~n2268 & ~n2269 ;
  assign n2271 = ~n2113 & ~n2115 ;
  assign n2272 = ~n2107 & ~n2109 ;
  assign n2273 = x66 & n2093 ;
  assign n2274 = n1850 & ~n2092 ;
  assign n2275 = n2087 & n2274 ;
  assign n2276 = x64 & n2275 ;
  assign n2277 = x65 & n2088 ;
  assign n2278 = ~n2276 & ~n2277 ;
  assign n2279 = ~n2273 & n2278 ;
  assign n2280 = n194 & n2096 ;
  assign n2281 = n2279 & ~n2280 ;
  assign n2282 = x17 & ~n2281 ;
  assign n2283 = x17 & ~n2282 ;
  assign n2284 = ~n2281 & ~n2282 ;
  assign n2285 = ~n2283 & ~n2284 ;
  assign n2286 = ~n2103 & n2285 ;
  assign n2287 = n2103 & ~n2285 ;
  assign n2288 = ~n2286 & ~n2287 ;
  assign n2289 = x69 & n1434 ;
  assign n2290 = x67 & n1646 ;
  assign n2291 = x68 & n1429 ;
  assign n2292 = ~n2290 & ~n2291 ;
  assign n2293 = ~n2289 & n2292 ;
  assign n2294 = n398 & n1437 ;
  assign n2295 = n2293 & ~n2294 ;
  assign n2296 = x14 & ~n2295 ;
  assign n2297 = x14 & ~n2296 ;
  assign n2298 = ~n2295 & ~n2296 ;
  assign n2299 = ~n2297 & ~n2298 ;
  assign n2300 = n2288 & ~n2299 ;
  assign n2301 = ~n2288 & n2299 ;
  assign n2302 = ~n2272 & ~n2301 ;
  assign n2303 = ~n2300 & n2302 ;
  assign n2304 = ~n2272 & ~n2303 ;
  assign n2305 = ~n2300 & ~n2303 ;
  assign n2306 = ~n2301 & n2305 ;
  assign n2307 = ~n2304 & ~n2306 ;
  assign n2308 = x72 & n945 ;
  assign n2309 = x70 & n1099 ;
  assign n2310 = x71 & n940 ;
  assign n2311 = ~n2309 & ~n2310 ;
  assign n2312 = ~n2308 & n2311 ;
  assign n2313 = n717 & n948 ;
  assign n2314 = n2312 & ~n2313 ;
  assign n2315 = x11 & ~n2314 ;
  assign n2316 = x11 & ~n2315 ;
  assign n2317 = ~n2314 & ~n2315 ;
  assign n2318 = ~n2316 & ~n2317 ;
  assign n2319 = n2307 & n2318 ;
  assign n2320 = ~n2307 & ~n2318 ;
  assign n2321 = ~n2319 & ~n2320 ;
  assign n2322 = ~n2271 & n2321 ;
  assign n2323 = n2271 & ~n2321 ;
  assign n2324 = ~n2322 & ~n2323 ;
  assign n2325 = n2270 & ~n2324 ;
  assign n2326 = ~n2270 & n2324 ;
  assign n2327 = ~n2325 & ~n2326 ;
  assign n2328 = ~n2259 & n2327 ;
  assign n2329 = n2259 & ~n2327 ;
  assign n2330 = ~n2328 & ~n2329 ;
  assign n2331 = n2258 & ~n2330 ;
  assign n2332 = ~n2258 & n2330 ;
  assign n2333 = ~n2331 & ~n2332 ;
  assign n2334 = ~n2247 & n2333 ;
  assign n2335 = n2247 & ~n2333 ;
  assign n2336 = ~n2334 & ~n2335 ;
  assign n2337 = x81 & n146 ;
  assign n2338 = x79 & n182 ;
  assign n2339 = x80 & n141 ;
  assign n2340 = ~n2338 & ~n2339 ;
  assign n2341 = ~n2337 & n2340 ;
  assign n2342 = ~n2024 & ~n2026 ;
  assign n2343 = ~x80 & ~x81 ;
  assign n2344 = x80 & x81 ;
  assign n2345 = ~n2343 & ~n2344 ;
  assign n2346 = ~n2342 & n2345 ;
  assign n2347 = n2342 & ~n2345 ;
  assign n2348 = ~n2346 & ~n2347 ;
  assign n2349 = n149 & n2348 ;
  assign n2350 = n2341 & ~n2349 ;
  assign n2351 = x2 & ~n2350 ;
  assign n2352 = x2 & ~n2351 ;
  assign n2353 = ~n2350 & ~n2351 ;
  assign n2354 = ~n2352 & ~n2353 ;
  assign n2355 = n2336 & ~n2354 ;
  assign n2356 = n2336 & ~n2355 ;
  assign n2357 = ~n2354 & ~n2355 ;
  assign n2358 = ~n2356 & ~n2357 ;
  assign n2359 = ~n2034 & n2129 ;
  assign n2360 = ~n2133 & ~n2359 ;
  assign n2361 = ~n2358 & ~n2360 ;
  assign n2362 = n2358 & n2360 ;
  assign n2363 = ~n2361 & ~n2362 ;
  assign n2477 = n2363 & x145 ;
  assign n2364 = ~n2232 & ~n2234 ;
  assign n2365 = ~x78 & n293 ;
  assign n2366 = ~x76 & n373 ;
  assign n2367 = ~x77 & n288 ;
  assign n2368 = ~n2366 & ~n2367 ;
  assign n2369 = ~n2365 & n2368 ;
  assign n2370 = n296 & n1718 ;
  assign n2371 = n2369 & ~n2370 ;
  assign n2372 = ~x5 & ~n2371 ;
  assign n2373 = ~x5 & ~n2372 ;
  assign n2374 = ~n2371 & ~n2372 ;
  assign n2375 = ~n2373 & ~n2374 ;
  assign n2376 = ~n2226 & ~n2228 ;
  assign n2377 = ~x75 & n574 ;
  assign n2378 = ~x73 & n673 ;
  assign n2379 = ~x74 & n569 ;
  assign n2380 = ~n2378 & ~n2379 ;
  assign n2381 = ~n2377 & n2380 ;
  assign n2382 = n577 & n1225 ;
  assign n2383 = n2381 & ~n2382 ;
  assign n2384 = ~x8 & ~n2383 ;
  assign n2385 = ~x8 & ~n2384 ;
  assign n2386 = ~n2383 & ~n2384 ;
  assign n2387 = ~n2385 & ~n2386 ;
  assign n2388 = ~n2220 & ~n2222 ;
  assign n2389 = ~n2214 & ~n2216 ;
  assign n2390 = ~x66 & n2093 ;
  assign n2391 = ~x64 & n2275 ;
  assign n2392 = ~x65 & n2088 ;
  assign n2393 = ~n2391 & ~n2392 ;
  assign n2394 = ~n2390 & n2393 ;
  assign n2395 = n214 & n2096 ;
  assign n2396 = n2394 & ~n2395 ;
  assign n2397 = ~x17 & ~n2396 ;
  assign n2398 = ~x17 & ~n2397 ;
  assign n2399 = ~n2396 & ~n2397 ;
  assign n2400 = ~n2398 & ~n2399 ;
  assign n2401 = ~n2210 & n2400 ;
  assign n2402 = n2210 & ~n2400 ;
  assign n2403 = ~n2401 & ~n2402 ;
  assign n2404 = ~x69 & n1434 ;
  assign n2405 = ~x67 & n1646 ;
  assign n2406 = ~x68 & n1429 ;
  assign n2407 = ~n2405 & ~n2406 ;
  assign n2408 = ~n2404 & n2407 ;
  assign n2409 = n435 & n1437 ;
  assign n2410 = n2408 & ~n2409 ;
  assign n2411 = ~x14 & ~n2410 ;
  assign n2412 = ~x14 & ~n2411 ;
  assign n2413 = ~n2410 & ~n2411 ;
  assign n2414 = ~n2412 & ~n2413 ;
  assign n2415 = n2403 & ~n2414 ;
  assign n2416 = ~n2403 & n2414 ;
  assign n2417 = ~n2389 & ~n2416 ;
  assign n2418 = ~n2415 & n2417 ;
  assign n2419 = ~n2389 & ~n2418 ;
  assign n2420 = ~n2415 & ~n2418 ;
  assign n2421 = ~n2416 & n2420 ;
  assign n2422 = ~n2419 & ~n2421 ;
  assign n2423 = ~x72 & n945 ;
  assign n2424 = ~x70 & n1099 ;
  assign n2425 = ~x71 & n940 ;
  assign n2426 = ~n2424 & ~n2425 ;
  assign n2427 = ~n2423 & n2426 ;
  assign n2428 = n773 & n948 ;
  assign n2429 = n2427 & ~n2428 ;
  assign n2430 = ~x11 & ~n2429 ;
  assign n2431 = ~x11 & ~n2430 ;
  assign n2432 = ~n2429 & ~n2430 ;
  assign n2433 = ~n2431 & ~n2432 ;
  assign n2434 = n2422 & n2433 ;
  assign n2435 = ~n2422 & ~n2433 ;
  assign n2436 = ~n2434 & ~n2435 ;
  assign n2437 = ~n2388 & n2436 ;
  assign n2438 = n2388 & ~n2436 ;
  assign n2439 = ~n2437 & ~n2438 ;
  assign n2440 = n2387 & ~n2439 ;
  assign n2441 = ~n2387 & n2439 ;
  assign n2442 = ~n2440 & ~n2441 ;
  assign n2443 = ~n2376 & n2442 ;
  assign n2444 = n2376 & ~n2442 ;
  assign n2445 = ~n2443 & ~n2444 ;
  assign n2446 = n2375 & ~n2445 ;
  assign n2447 = ~n2375 & n2445 ;
  assign n2448 = ~n2446 & ~n2447 ;
  assign n2449 = ~n2364 & n2448 ;
  assign n2450 = n2364 & ~n2448 ;
  assign n2451 = ~n2449 & ~n2450 ;
  assign n2452 = ~x81 & n164 ;
  assign n2453 = ~x79 & n205 ;
  assign n2454 = ~x80 & n162 ;
  assign n2455 = ~n2453 & ~n2454 ;
  assign n2456 = ~n2452 & n2455 ;
  assign n2457 = ~n2023 & ~n2143 ;
  assign n2458 = n2345 & ~n2457 ;
  assign n2459 = ~n2345 & n2457 ;
  assign n2460 = ~n2458 & ~n2459 ;
  assign n2461 = n167 & n2460 ;
  assign n2462 = n2456 & ~n2461 ;
  assign n2463 = ~x2 & ~n2462 ;
  assign n2464 = ~x2 & ~n2463 ;
  assign n2465 = ~n2462 & ~n2463 ;
  assign n2466 = ~n2464 & ~n2465 ;
  assign n2467 = n2451 & ~n2466 ;
  assign n2468 = n2451 & ~n2467 ;
  assign n2469 = ~n2466 & ~n2467 ;
  assign n2470 = ~n2468 & ~n2469 ;
  assign n2471 = ~n2151 & n2236 ;
  assign n2472 = ~n2240 & ~n2471 ;
  assign n2473 = ~n2470 & ~n2472 ;
  assign n2474 = n2470 & n2472 ;
  assign n2475 = ~n2473 & ~n2474 ;
  assign n2478 = ~n2475 & ~x145 ;
  assign n2479 = ~n2477 & ~n2478 ;
  assign n2480 = ~n2332 & ~n2334 ;
  assign n2481 = x79 & n293 ;
  assign n2482 = x77 & n373 ;
  assign n2483 = x78 & n288 ;
  assign n2484 = ~n2482 & ~n2483 ;
  assign n2485 = ~n2481 & n2484 ;
  assign n2486 = n296 & n1817 ;
  assign n2487 = n2485 & ~n2486 ;
  assign n2488 = x5 & ~n2487 ;
  assign n2489 = x5 & ~n2488 ;
  assign n2490 = ~n2487 & ~n2488 ;
  assign n2491 = ~n2489 & ~n2490 ;
  assign n2492 = ~n2326 & ~n2328 ;
  assign n2493 = x76 & n574 ;
  assign n2494 = x74 & n673 ;
  assign n2495 = x75 & n569 ;
  assign n2496 = ~n2494 & ~n2495 ;
  assign n2497 = ~n2493 & n2496 ;
  assign n2498 = n577 & n1311 ;
  assign n2499 = n2497 & ~n2498 ;
  assign n2500 = x8 & ~n2499 ;
  assign n2501 = x8 & ~n2500 ;
  assign n2502 = ~n2499 & ~n2500 ;
  assign n2503 = ~n2501 & ~n2502 ;
  assign n2504 = ~n2320 & ~n2322 ;
  assign n2505 = x17 & ~x18 ;
  assign n2506 = ~x17 & x18 ;
  assign n2507 = ~n2505 & ~n2506 ;
  assign n2508 = x64 & ~n2507 ;
  assign n2509 = ~n2287 & n2508 ;
  assign n2510 = n2287 & ~n2508 ;
  assign n2511 = ~n2509 & ~n2510 ;
  assign n2512 = x67 & n2093 ;
  assign n2513 = x65 & n2275 ;
  assign n2514 = x66 & n2088 ;
  assign n2515 = ~n2513 & ~n2514 ;
  assign n2516 = ~n2512 & n2515 ;
  assign n2517 = n240 & n2096 ;
  assign n2518 = n2516 & ~n2517 ;
  assign n2519 = x17 & ~n2518 ;
  assign n2520 = x17 & ~n2519 ;
  assign n2521 = ~n2518 & ~n2519 ;
  assign n2522 = ~n2520 & ~n2521 ;
  assign n2523 = ~n2511 & ~n2522 ;
  assign n2524 = n2511 & n2522 ;
  assign n2525 = ~n2523 & ~n2524 ;
  assign n2526 = x70 & n1434 ;
  assign n2527 = x68 & n1646 ;
  assign n2528 = x69 & n1429 ;
  assign n2529 = ~n2527 & ~n2528 ;
  assign n2530 = ~n2526 & n2529 ;
  assign n2531 = n488 & n1437 ;
  assign n2532 = n2530 & ~n2531 ;
  assign n2533 = x14 & ~n2532 ;
  assign n2534 = x14 & ~n2533 ;
  assign n2535 = ~n2532 & ~n2533 ;
  assign n2536 = ~n2534 & ~n2535 ;
  assign n2537 = n2525 & ~n2536 ;
  assign n2538 = n2525 & ~n2537 ;
  assign n2539 = ~n2536 & ~n2537 ;
  assign n2540 = ~n2538 & ~n2539 ;
  assign n2541 = ~n2305 & n2540 ;
  assign n2542 = n2305 & ~n2540 ;
  assign n2543 = ~n2541 & ~n2542 ;
  assign n2544 = x73 & n945 ;
  assign n2545 = x71 & n1099 ;
  assign n2546 = x72 & n940 ;
  assign n2547 = ~n2545 & ~n2546 ;
  assign n2548 = ~n2544 & n2547 ;
  assign n2549 = n843 & n948 ;
  assign n2550 = n2548 & ~n2549 ;
  assign n2551 = x11 & ~n2550 ;
  assign n2552 = x11 & ~n2551 ;
  assign n2553 = ~n2550 & ~n2551 ;
  assign n2554 = ~n2552 & ~n2553 ;
  assign n2555 = ~n2543 & ~n2554 ;
  assign n2556 = n2543 & n2554 ;
  assign n2557 = ~n2555 & ~n2556 ;
  assign n2558 = ~n2504 & n2557 ;
  assign n2559 = n2504 & ~n2557 ;
  assign n2560 = ~n2558 & ~n2559 ;
  assign n2561 = n2503 & ~n2560 ;
  assign n2562 = ~n2503 & n2560 ;
  assign n2563 = ~n2561 & ~n2562 ;
  assign n2564 = ~n2492 & n2563 ;
  assign n2565 = n2492 & ~n2563 ;
  assign n2566 = ~n2564 & ~n2565 ;
  assign n2567 = ~n2491 & n2566 ;
  assign n2568 = n2491 & ~n2566 ;
  assign n2569 = ~n2567 & ~n2568 ;
  assign n2570 = ~n2480 & n2569 ;
  assign n2571 = n2480 & ~n2569 ;
  assign n2572 = ~n2570 & ~n2571 ;
  assign n2573 = x82 & n146 ;
  assign n2574 = x80 & n182 ;
  assign n2575 = x81 & n141 ;
  assign n2576 = ~n2574 & ~n2575 ;
  assign n2577 = ~n2573 & n2576 ;
  assign n2578 = ~n2344 & ~n2346 ;
  assign n2579 = ~x81 & ~x82 ;
  assign n2580 = x81 & x82 ;
  assign n2581 = ~n2579 & ~n2580 ;
  assign n2582 = ~n2578 & n2581 ;
  assign n2583 = n2578 & ~n2581 ;
  assign n2584 = ~n2582 & ~n2583 ;
  assign n2585 = n149 & n2584 ;
  assign n2586 = n2577 & ~n2585 ;
  assign n2587 = x2 & ~n2586 ;
  assign n2588 = x2 & ~n2587 ;
  assign n2589 = ~n2586 & ~n2587 ;
  assign n2590 = ~n2588 & ~n2589 ;
  assign n2591 = n2572 & ~n2590 ;
  assign n2592 = n2572 & ~n2591 ;
  assign n2593 = ~n2590 & ~n2591 ;
  assign n2594 = ~n2592 & ~n2593 ;
  assign n2595 = ~n2355 & ~n2361 ;
  assign n2596 = ~n2594 & ~n2595 ;
  assign n2597 = n2594 & n2595 ;
  assign n2598 = ~n2596 & ~n2597 ;
  assign n2713 = n2598 & x146 ;
  assign n2599 = ~n2447 & ~n2449 ;
  assign n2600 = ~x79 & n293 ;
  assign n2601 = ~x77 & n373 ;
  assign n2602 = ~x78 & n288 ;
  assign n2603 = ~n2601 & ~n2602 ;
  assign n2604 = ~n2600 & n2603 ;
  assign n2605 = n296 & n1921 ;
  assign n2606 = n2604 & ~n2605 ;
  assign n2607 = ~x5 & ~n2606 ;
  assign n2608 = ~x5 & ~n2607 ;
  assign n2609 = ~n2606 & ~n2607 ;
  assign n2610 = ~n2608 & ~n2609 ;
  assign n2611 = ~n2441 & ~n2443 ;
  assign n2612 = ~x76 & n574 ;
  assign n2613 = ~x74 & n673 ;
  assign n2614 = ~x75 & n569 ;
  assign n2615 = ~n2613 & ~n2614 ;
  assign n2616 = ~n2612 & n2615 ;
  assign n2617 = n577 & n1390 ;
  assign n2618 = n2616 & ~n2617 ;
  assign n2619 = ~x8 & ~n2618 ;
  assign n2620 = ~x8 & ~n2619 ;
  assign n2621 = ~n2618 & ~n2619 ;
  assign n2622 = ~n2620 & ~n2621 ;
  assign n2623 = ~n2435 & ~n2437 ;
  assign n2624 = ~x64 & ~n2507 ;
  assign n2625 = ~n2402 & n2624 ;
  assign n2626 = n2402 & ~n2624 ;
  assign n2627 = ~n2625 & ~n2626 ;
  assign n2628 = ~x67 & n2093 ;
  assign n2629 = ~x65 & n2275 ;
  assign n2630 = ~x66 & n2088 ;
  assign n2631 = ~n2629 & ~n2630 ;
  assign n2632 = ~n2628 & n2631 ;
  assign n2633 = n266 & n2096 ;
  assign n2634 = n2632 & ~n2633 ;
  assign n2635 = ~x17 & ~n2634 ;
  assign n2636 = ~x17 & ~n2635 ;
  assign n2637 = ~n2634 & ~n2635 ;
  assign n2638 = ~n2636 & ~n2637 ;
  assign n2639 = ~n2627 & ~n2638 ;
  assign n2640 = n2627 & n2638 ;
  assign n2641 = ~n2639 & ~n2640 ;
  assign n2642 = ~x70 & n1434 ;
  assign n2643 = ~x68 & n1646 ;
  assign n2644 = ~x69 & n1429 ;
  assign n2645 = ~n2643 & ~n2644 ;
  assign n2646 = ~n2642 & n2645 ;
  assign n2647 = n529 & n1437 ;
  assign n2648 = n2646 & ~n2647 ;
  assign n2649 = ~x14 & ~n2648 ;
  assign n2650 = ~x14 & ~n2649 ;
  assign n2651 = ~n2648 & ~n2649 ;
  assign n2652 = ~n2650 & ~n2651 ;
  assign n2653 = n2641 & ~n2652 ;
  assign n2654 = n2641 & ~n2653 ;
  assign n2655 = ~n2652 & ~n2653 ;
  assign n2656 = ~n2654 & ~n2655 ;
  assign n2657 = ~n2420 & n2656 ;
  assign n2658 = n2420 & ~n2656 ;
  assign n2659 = ~n2657 & ~n2658 ;
  assign n2660 = ~x73 & n945 ;
  assign n2661 = ~x71 & n1099 ;
  assign n2662 = ~x72 & n940 ;
  assign n2663 = ~n2661 & ~n2662 ;
  assign n2664 = ~n2660 & n2663 ;
  assign n2665 = n903 & n948 ;
  assign n2666 = n2664 & ~n2665 ;
  assign n2667 = ~x11 & ~n2666 ;
  assign n2668 = ~x11 & ~n2667 ;
  assign n2669 = ~n2666 & ~n2667 ;
  assign n2670 = ~n2668 & ~n2669 ;
  assign n2671 = ~n2659 & ~n2670 ;
  assign n2672 = n2659 & n2670 ;
  assign n2673 = ~n2671 & ~n2672 ;
  assign n2674 = ~n2623 & n2673 ;
  assign n2675 = n2623 & ~n2673 ;
  assign n2676 = ~n2674 & ~n2675 ;
  assign n2677 = n2622 & ~n2676 ;
  assign n2678 = ~n2622 & n2676 ;
  assign n2679 = ~n2677 & ~n2678 ;
  assign n2680 = ~n2611 & n2679 ;
  assign n2681 = n2611 & ~n2679 ;
  assign n2682 = ~n2680 & ~n2681 ;
  assign n2683 = ~n2610 & n2682 ;
  assign n2684 = n2610 & ~n2682 ;
  assign n2685 = ~n2683 & ~n2684 ;
  assign n2686 = ~n2599 & n2685 ;
  assign n2687 = n2599 & ~n2685 ;
  assign n2688 = ~n2686 & ~n2687 ;
  assign n2689 = ~x82 & n164 ;
  assign n2690 = ~x80 & n205 ;
  assign n2691 = ~x81 & n162 ;
  assign n2692 = ~n2690 & ~n2691 ;
  assign n2693 = ~n2689 & n2692 ;
  assign n2694 = ~n2343 & ~n2458 ;
  assign n2695 = n2581 & ~n2694 ;
  assign n2696 = ~n2581 & n2694 ;
  assign n2697 = ~n2695 & ~n2696 ;
  assign n2698 = n167 & n2697 ;
  assign n2699 = n2693 & ~n2698 ;
  assign n2700 = ~x2 & ~n2699 ;
  assign n2701 = ~x2 & ~n2700 ;
  assign n2702 = ~n2699 & ~n2700 ;
  assign n2703 = ~n2701 & ~n2702 ;
  assign n2704 = n2688 & ~n2703 ;
  assign n2705 = n2688 & ~n2704 ;
  assign n2706 = ~n2703 & ~n2704 ;
  assign n2707 = ~n2705 & ~n2706 ;
  assign n2708 = ~n2467 & ~n2473 ;
  assign n2709 = ~n2707 & ~n2708 ;
  assign n2710 = n2707 & n2708 ;
  assign n2711 = ~n2709 & ~n2710 ;
  assign n2714 = ~n2711 & ~x146 ;
  assign n2715 = ~n2713 & ~n2714 ;
  assign n2716 = ~n2305 & ~n2540 ;
  assign n2717 = ~n2537 & ~n2716 ;
  assign n2718 = x71 & n1434 ;
  assign n2719 = x69 & n1646 ;
  assign n2720 = x70 & n1429 ;
  assign n2721 = ~n2719 & ~n2720 ;
  assign n2722 = ~n2718 & n2721 ;
  assign n2723 = n558 & n1437 ;
  assign n2724 = n2722 & ~n2723 ;
  assign n2725 = x14 & ~n2724 ;
  assign n2726 = x14 & ~n2725 ;
  assign n2727 = ~n2724 & ~n2725 ;
  assign n2728 = ~n2726 & ~n2727 ;
  assign n2729 = n2287 & n2508 ;
  assign n2730 = ~n2523 & ~n2729 ;
  assign n2731 = x68 & n2093 ;
  assign n2732 = x66 & n2275 ;
  assign n2733 = x67 & n2088 ;
  assign n2734 = ~n2732 & ~n2733 ;
  assign n2735 = ~n2731 & n2734 ;
  assign n2736 = n317 & n2096 ;
  assign n2737 = n2735 & ~n2736 ;
  assign n2738 = x17 & ~n2737 ;
  assign n2739 = x17 & ~n2738 ;
  assign n2740 = ~n2737 & ~n2738 ;
  assign n2741 = ~n2739 & ~n2740 ;
  assign n2742 = x20 & ~n2508 ;
  assign n2743 = ~x18 & x19 ;
  assign n2744 = x18 & ~x19 ;
  assign n2745 = ~n2743 & ~n2744 ;
  assign n2746 = n2507 & ~n2745 ;
  assign n2747 = x64 & n2746 ;
  assign n2748 = ~x19 & x20 ;
  assign n2749 = x19 & ~x20 ;
  assign n2750 = ~n2748 & ~n2749 ;
  assign n2751 = ~n2507 & n2750 ;
  assign n2752 = x65 & n2751 ;
  assign n2753 = ~n2747 & ~n2752 ;
  assign n2754 = ~n2507 & ~n2750 ;
  assign n2755 = ~n152 & n2754 ;
  assign n2756 = n2753 & ~n2755 ;
  assign n2757 = x20 & ~n2756 ;
  assign n2758 = x20 & ~n2757 ;
  assign n2759 = ~n2756 & ~n2757 ;
  assign n2760 = ~n2758 & ~n2759 ;
  assign n2761 = n2742 & ~n2760 ;
  assign n2762 = ~n2742 & n2760 ;
  assign n2763 = ~n2761 & ~n2762 ;
  assign n2764 = n2741 & n2763 ;
  assign n2765 = ~n2741 & ~n2763 ;
  assign n2766 = ~n2764 & ~n2765 ;
  assign n2767 = ~n2730 & ~n2766 ;
  assign n2768 = n2730 & n2766 ;
  assign n2769 = ~n2767 & ~n2768 ;
  assign n2770 = ~n2728 & n2769 ;
  assign n2771 = n2728 & ~n2769 ;
  assign n2772 = ~n2770 & ~n2771 ;
  assign n2773 = ~n2717 & n2772 ;
  assign n2774 = n2717 & ~n2772 ;
  assign n2775 = ~n2773 & ~n2774 ;
  assign n2776 = x74 & n945 ;
  assign n2777 = x72 & n1099 ;
  assign n2778 = x73 & n940 ;
  assign n2779 = ~n2777 & ~n2778 ;
  assign n2780 = ~n2776 & n2779 ;
  assign n2781 = n948 & n994 ;
  assign n2782 = n2780 & ~n2781 ;
  assign n2783 = x11 & ~n2782 ;
  assign n2784 = x11 & ~n2783 ;
  assign n2785 = ~n2782 & ~n2783 ;
  assign n2786 = ~n2784 & ~n2785 ;
  assign n2787 = n2775 & ~n2786 ;
  assign n2788 = n2775 & ~n2787 ;
  assign n2789 = ~n2786 & ~n2787 ;
  assign n2790 = ~n2788 & ~n2789 ;
  assign n2791 = ~n2555 & ~n2558 ;
  assign n2792 = n2790 & n2791 ;
  assign n2793 = ~n2790 & ~n2791 ;
  assign n2794 = ~n2792 & ~n2793 ;
  assign n2795 = x77 & n574 ;
  assign n2796 = x75 & n673 ;
  assign n2797 = x76 & n569 ;
  assign n2798 = ~n2796 & ~n2797 ;
  assign n2799 = ~n2795 & n2798 ;
  assign n2800 = n577 & n1502 ;
  assign n2801 = n2799 & ~n2800 ;
  assign n2802 = x8 & ~n2801 ;
  assign n2803 = x8 & ~n2802 ;
  assign n2804 = ~n2801 & ~n2802 ;
  assign n2805 = ~n2803 & ~n2804 ;
  assign n2806 = ~n2794 & n2805 ;
  assign n2807 = n2794 & ~n2805 ;
  assign n2808 = ~n2806 & ~n2807 ;
  assign n2809 = ~n2562 & ~n2564 ;
  assign n2810 = n2808 & ~n2809 ;
  assign n2811 = ~n2808 & n2809 ;
  assign n2812 = ~n2810 & ~n2811 ;
  assign n2813 = x80 & n293 ;
  assign n2814 = x78 & n373 ;
  assign n2815 = x79 & n288 ;
  assign n2816 = ~n2814 & ~n2815 ;
  assign n2817 = ~n2813 & n2816 ;
  assign n2818 = n296 & n2028 ;
  assign n2819 = n2817 & ~n2818 ;
  assign n2820 = x5 & ~n2819 ;
  assign n2821 = x5 & ~n2820 ;
  assign n2822 = ~n2819 & ~n2820 ;
  assign n2823 = ~n2821 & ~n2822 ;
  assign n2824 = n2812 & ~n2823 ;
  assign n2825 = n2812 & ~n2824 ;
  assign n2826 = ~n2823 & ~n2824 ;
  assign n2827 = ~n2825 & ~n2826 ;
  assign n2828 = ~n2567 & ~n2570 ;
  assign n2829 = n2827 & n2828 ;
  assign n2830 = ~n2827 & ~n2828 ;
  assign n2831 = ~n2829 & ~n2830 ;
  assign n2832 = x83 & n146 ;
  assign n2833 = x81 & n182 ;
  assign n2834 = x82 & n141 ;
  assign n2835 = ~n2833 & ~n2834 ;
  assign n2836 = ~n2832 & n2835 ;
  assign n2837 = ~n2580 & ~n2582 ;
  assign n2838 = ~x82 & ~x83 ;
  assign n2839 = x82 & x83 ;
  assign n2840 = ~n2838 & ~n2839 ;
  assign n2841 = ~n2837 & n2840 ;
  assign n2842 = n2837 & ~n2840 ;
  assign n2843 = ~n2841 & ~n2842 ;
  assign n2844 = n149 & n2843 ;
  assign n2845 = n2836 & ~n2844 ;
  assign n2846 = x2 & ~n2845 ;
  assign n2847 = x2 & ~n2846 ;
  assign n2848 = ~n2845 & ~n2846 ;
  assign n2849 = ~n2847 & ~n2848 ;
  assign n2850 = n2831 & ~n2849 ;
  assign n2851 = n2831 & ~n2850 ;
  assign n2852 = ~n2849 & ~n2850 ;
  assign n2853 = ~n2851 & ~n2852 ;
  assign n2854 = ~n2591 & ~n2596 ;
  assign n2855 = ~n2853 & ~n2854 ;
  assign n2856 = n2853 & n2854 ;
  assign n2857 = ~n2855 & ~n2856 ;
  assign n2988 = n2857 & x147 ;
  assign n2858 = ~n2420 & ~n2656 ;
  assign n2859 = ~n2653 & ~n2858 ;
  assign n2860 = ~x71 & n1434 ;
  assign n2861 = ~x69 & n1646 ;
  assign n2862 = ~x70 & n1429 ;
  assign n2863 = ~n2861 & ~n2862 ;
  assign n2864 = ~n2860 & n2863 ;
  assign n2865 = n622 & n1437 ;
  assign n2866 = n2864 & ~n2865 ;
  assign n2867 = ~x14 & ~n2866 ;
  assign n2868 = ~x14 & ~n2867 ;
  assign n2869 = ~n2866 & ~n2867 ;
  assign n2870 = ~n2868 & ~n2869 ;
  assign n2871 = n2402 & n2624 ;
  assign n2872 = ~n2639 & ~n2871 ;
  assign n2873 = ~x68 & n2093 ;
  assign n2874 = ~x66 & n2275 ;
  assign n2875 = ~x67 & n2088 ;
  assign n2876 = ~n2874 & ~n2875 ;
  assign n2877 = ~n2873 & n2876 ;
  assign n2878 = n352 & n2096 ;
  assign n2879 = n2877 & ~n2878 ;
  assign n2880 = ~x17 & ~n2879 ;
  assign n2881 = ~x17 & ~n2880 ;
  assign n2882 = ~n2879 & ~n2880 ;
  assign n2883 = ~n2881 & ~n2882 ;
  assign n2884 = ~x20 & ~n2624 ;
  assign n2885 = ~x64 & n2746 ;
  assign n2886 = ~x65 & n2751 ;
  assign n2887 = ~n2885 & ~n2886 ;
  assign n2888 = ~n2755 & n2887 ;
  assign n2889 = ~x20 & ~n2888 ;
  assign n2890 = ~x20 & ~n2889 ;
  assign n2891 = ~n2888 & ~n2889 ;
  assign n2892 = ~n2890 & ~n2891 ;
  assign n2893 = n2884 & ~n2892 ;
  assign n2894 = ~n2884 & n2892 ;
  assign n2895 = ~n2893 & ~n2894 ;
  assign n2896 = n2883 & n2895 ;
  assign n2897 = ~n2883 & ~n2895 ;
  assign n2898 = ~n2896 & ~n2897 ;
  assign n2899 = ~n2872 & ~n2898 ;
  assign n2900 = n2872 & n2898 ;
  assign n2901 = ~n2899 & ~n2900 ;
  assign n2902 = ~n2870 & n2901 ;
  assign n2903 = n2870 & ~n2901 ;
  assign n2904 = ~n2902 & ~n2903 ;
  assign n2905 = ~n2859 & n2904 ;
  assign n2906 = n2859 & ~n2904 ;
  assign n2907 = ~n2905 & ~n2906 ;
  assign n2908 = ~x74 & n945 ;
  assign n2909 = ~x72 & n1099 ;
  assign n2910 = ~x73 & n940 ;
  assign n2911 = ~n2909 & ~n2910 ;
  assign n2912 = ~n2908 & n2911 ;
  assign n2913 = n948 & n1066 ;
  assign n2914 = n2912 & ~n2913 ;
  assign n2915 = ~x11 & ~n2914 ;
  assign n2916 = ~x11 & ~n2915 ;
  assign n2917 = ~n2914 & ~n2915 ;
  assign n2918 = ~n2916 & ~n2917 ;
  assign n2919 = n2907 & ~n2918 ;
  assign n2920 = n2907 & ~n2919 ;
  assign n2921 = ~n2918 & ~n2919 ;
  assign n2922 = ~n2920 & ~n2921 ;
  assign n2923 = ~n2671 & ~n2674 ;
  assign n2924 = n2922 & n2923 ;
  assign n2925 = ~n2922 & ~n2923 ;
  assign n2926 = ~n2924 & ~n2925 ;
  assign n2927 = ~x77 & n574 ;
  assign n2928 = ~x75 & n673 ;
  assign n2929 = ~x76 & n569 ;
  assign n2930 = ~n2928 & ~n2929 ;
  assign n2931 = ~n2927 & n2930 ;
  assign n2932 = n577 & n1594 ;
  assign n2933 = n2931 & ~n2932 ;
  assign n2934 = ~x8 & ~n2933 ;
  assign n2935 = ~x8 & ~n2934 ;
  assign n2936 = ~n2933 & ~n2934 ;
  assign n2937 = ~n2935 & ~n2936 ;
  assign n2938 = ~n2926 & n2937 ;
  assign n2939 = n2926 & ~n2937 ;
  assign n2940 = ~n2938 & ~n2939 ;
  assign n2941 = ~n2678 & ~n2680 ;
  assign n2942 = n2940 & ~n2941 ;
  assign n2943 = ~n2940 & n2941 ;
  assign n2944 = ~n2942 & ~n2943 ;
  assign n2945 = ~x80 & n293 ;
  assign n2946 = ~x78 & n373 ;
  assign n2947 = ~x79 & n288 ;
  assign n2948 = ~n2946 & ~n2947 ;
  assign n2949 = ~n2945 & n2948 ;
  assign n2950 = n296 & n2145 ;
  assign n2951 = n2949 & ~n2950 ;
  assign n2952 = ~x5 & ~n2951 ;
  assign n2953 = ~x5 & ~n2952 ;
  assign n2954 = ~n2951 & ~n2952 ;
  assign n2955 = ~n2953 & ~n2954 ;
  assign n2956 = n2944 & ~n2955 ;
  assign n2957 = n2944 & ~n2956 ;
  assign n2958 = ~n2955 & ~n2956 ;
  assign n2959 = ~n2957 & ~n2958 ;
  assign n2960 = ~n2683 & ~n2686 ;
  assign n2961 = n2959 & n2960 ;
  assign n2962 = ~n2959 & ~n2960 ;
  assign n2963 = ~n2961 & ~n2962 ;
  assign n2964 = ~x83 & n164 ;
  assign n2965 = ~x81 & n205 ;
  assign n2966 = ~x82 & n162 ;
  assign n2967 = ~n2965 & ~n2966 ;
  assign n2968 = ~n2964 & n2967 ;
  assign n2969 = ~n2579 & ~n2695 ;
  assign n2970 = n2840 & ~n2969 ;
  assign n2971 = ~n2840 & n2969 ;
  assign n2972 = ~n2970 & ~n2971 ;
  assign n2973 = n167 & n2972 ;
  assign n2974 = n2968 & ~n2973 ;
  assign n2975 = ~x2 & ~n2974 ;
  assign n2976 = ~x2 & ~n2975 ;
  assign n2977 = ~n2974 & ~n2975 ;
  assign n2978 = ~n2976 & ~n2977 ;
  assign n2979 = n2963 & ~n2978 ;
  assign n2980 = n2963 & ~n2979 ;
  assign n2981 = ~n2978 & ~n2979 ;
  assign n2982 = ~n2980 & ~n2981 ;
  assign n2983 = ~n2704 & ~n2709 ;
  assign n2984 = ~n2982 & ~n2983 ;
  assign n2985 = n2982 & n2983 ;
  assign n2986 = ~n2984 & ~n2985 ;
  assign n2989 = ~n2986 & ~x147 ;
  assign n2990 = ~n2988 & ~n2989 ;
  assign n2991 = ~n2824 & ~n2830 ;
  assign n2992 = x81 & n293 ;
  assign n2993 = x79 & n373 ;
  assign n2994 = x80 & n288 ;
  assign n2995 = ~n2993 & ~n2994 ;
  assign n2996 = ~n2992 & n2995 ;
  assign n2997 = n296 & n2348 ;
  assign n2998 = n2996 & ~n2997 ;
  assign n2999 = x5 & ~n2998 ;
  assign n3000 = x5 & ~n2999 ;
  assign n3001 = ~n2998 & ~n2999 ;
  assign n3002 = ~n3000 & ~n3001 ;
  assign n3003 = ~n2787 & ~n2793 ;
  assign n3004 = x75 & n945 ;
  assign n3005 = x73 & n1099 ;
  assign n3006 = x74 & n940 ;
  assign n3007 = ~n3005 & ~n3006 ;
  assign n3008 = ~n3004 & n3007 ;
  assign n3009 = n948 & n1150 ;
  assign n3010 = n3008 & ~n3009 ;
  assign n3011 = x11 & ~n3010 ;
  assign n3012 = x11 & ~n3011 ;
  assign n3013 = ~n3010 & ~n3011 ;
  assign n3014 = ~n3012 & ~n3013 ;
  assign n3015 = ~n2770 & ~n2773 ;
  assign n3016 = ~n2741 & n2763 ;
  assign n3017 = ~n2767 & ~n3016 ;
  assign n3018 = x66 & n2751 ;
  assign n3019 = n2507 & ~n2750 ;
  assign n3020 = n2745 & n3019 ;
  assign n3021 = x64 & n3020 ;
  assign n3022 = x65 & n2746 ;
  assign n3023 = ~n3021 & ~n3022 ;
  assign n3024 = ~n3018 & n3023 ;
  assign n3025 = n194 & n2754 ;
  assign n3026 = n3024 & ~n3025 ;
  assign n3027 = x20 & ~n3026 ;
  assign n3028 = x20 & ~n3027 ;
  assign n3029 = ~n3026 & ~n3027 ;
  assign n3030 = ~n3028 & ~n3029 ;
  assign n3031 = ~n2761 & n3030 ;
  assign n3032 = n2761 & ~n3030 ;
  assign n3033 = ~n3031 & ~n3032 ;
  assign n3034 = x69 & n2093 ;
  assign n3035 = x67 & n2275 ;
  assign n3036 = x68 & n2088 ;
  assign n3037 = ~n3035 & ~n3036 ;
  assign n3038 = ~n3034 & n3037 ;
  assign n3039 = n398 & n2096 ;
  assign n3040 = n3038 & ~n3039 ;
  assign n3041 = x17 & ~n3040 ;
  assign n3042 = x17 & ~n3041 ;
  assign n3043 = ~n3040 & ~n3041 ;
  assign n3044 = ~n3042 & ~n3043 ;
  assign n3045 = n3033 & ~n3044 ;
  assign n3046 = ~n3033 & n3044 ;
  assign n3047 = ~n3017 & ~n3046 ;
  assign n3048 = ~n3045 & n3047 ;
  assign n3049 = ~n3017 & ~n3048 ;
  assign n3050 = ~n3045 & ~n3048 ;
  assign n3051 = ~n3046 & n3050 ;
  assign n3052 = ~n3049 & ~n3051 ;
  assign n3053 = x72 & n1434 ;
  assign n3054 = x70 & n1646 ;
  assign n3055 = x71 & n1429 ;
  assign n3056 = ~n3054 & ~n3055 ;
  assign n3057 = ~n3053 & n3056 ;
  assign n3058 = n717 & n1437 ;
  assign n3059 = n3057 & ~n3058 ;
  assign n3060 = x14 & ~n3059 ;
  assign n3061 = x14 & ~n3060 ;
  assign n3062 = ~n3059 & ~n3060 ;
  assign n3063 = ~n3061 & ~n3062 ;
  assign n3064 = n3052 & n3063 ;
  assign n3065 = ~n3052 & ~n3063 ;
  assign n3066 = ~n3064 & ~n3065 ;
  assign n3067 = ~n3015 & n3066 ;
  assign n3068 = n3015 & ~n3066 ;
  assign n3069 = ~n3067 & ~n3068 ;
  assign n3070 = n3014 & ~n3069 ;
  assign n3071 = ~n3014 & n3069 ;
  assign n3072 = ~n3070 & ~n3071 ;
  assign n3073 = ~n3003 & n3072 ;
  assign n3074 = n3003 & ~n3072 ;
  assign n3075 = ~n3073 & ~n3074 ;
  assign n3076 = x78 & n574 ;
  assign n3077 = x76 & n673 ;
  assign n3078 = x77 & n569 ;
  assign n3079 = ~n3077 & ~n3078 ;
  assign n3080 = ~n3076 & n3079 ;
  assign n3081 = n577 & n1624 ;
  assign n3082 = n3080 & ~n3081 ;
  assign n3083 = x8 & ~n3082 ;
  assign n3084 = x8 & ~n3083 ;
  assign n3085 = ~n3082 & ~n3083 ;
  assign n3086 = ~n3084 & ~n3085 ;
  assign n3087 = n3075 & ~n3086 ;
  assign n3088 = n3075 & ~n3087 ;
  assign n3089 = ~n3086 & ~n3087 ;
  assign n3090 = ~n3088 & ~n3089 ;
  assign n3091 = ~n2807 & ~n2810 ;
  assign n3092 = ~n3090 & ~n3091 ;
  assign n3093 = n3090 & n3091 ;
  assign n3094 = ~n3092 & ~n3093 ;
  assign n3095 = ~n3002 & n3094 ;
  assign n3096 = ~n3002 & ~n3095 ;
  assign n3097 = n3094 & ~n3095 ;
  assign n3098 = ~n3096 & ~n3097 ;
  assign n3099 = ~n2991 & ~n3098 ;
  assign n3100 = ~n2991 & ~n3099 ;
  assign n3101 = ~n3098 & ~n3099 ;
  assign n3102 = ~n3100 & ~n3101 ;
  assign n3103 = x84 & n146 ;
  assign n3104 = x82 & n182 ;
  assign n3105 = x83 & n141 ;
  assign n3106 = ~n3104 & ~n3105 ;
  assign n3107 = ~n3103 & n3106 ;
  assign n3108 = ~n2839 & ~n2841 ;
  assign n3109 = ~x83 & ~x84 ;
  assign n3110 = x83 & x84 ;
  assign n3111 = ~n3109 & ~n3110 ;
  assign n3112 = ~n3108 & n3111 ;
  assign n3113 = n3108 & ~n3111 ;
  assign n3114 = ~n3112 & ~n3113 ;
  assign n3115 = n149 & n3114 ;
  assign n3116 = n3107 & ~n3115 ;
  assign n3117 = x2 & ~n3116 ;
  assign n3118 = x2 & ~n3117 ;
  assign n3119 = ~n3116 & ~n3117 ;
  assign n3120 = ~n3118 & ~n3119 ;
  assign n3121 = ~n3102 & ~n3120 ;
  assign n3122 = ~n3102 & ~n3121 ;
  assign n3123 = ~n3120 & ~n3121 ;
  assign n3124 = ~n3122 & ~n3123 ;
  assign n3125 = ~n2850 & ~n2855 ;
  assign n3126 = ~n3124 & ~n3125 ;
  assign n3127 = n3124 & n3125 ;
  assign n3128 = ~n3126 & ~n3127 ;
  assign n3263 = n3128 & x148 ;
  assign n3129 = ~n2956 & ~n2962 ;
  assign n3130 = ~x81 & n293 ;
  assign n3131 = ~x79 & n373 ;
  assign n3132 = ~x80 & n288 ;
  assign n3133 = ~n3131 & ~n3132 ;
  assign n3134 = ~n3130 & n3133 ;
  assign n3135 = n296 & n2460 ;
  assign n3136 = n3134 & ~n3135 ;
  assign n3137 = ~x5 & ~n3136 ;
  assign n3138 = ~x5 & ~n3137 ;
  assign n3139 = ~n3136 & ~n3137 ;
  assign n3140 = ~n3138 & ~n3139 ;
  assign n3141 = ~n2919 & ~n2925 ;
  assign n3142 = ~x75 & n945 ;
  assign n3143 = ~x73 & n1099 ;
  assign n3144 = ~x74 & n940 ;
  assign n3145 = ~n3143 & ~n3144 ;
  assign n3146 = ~n3142 & n3145 ;
  assign n3147 = n948 & n1225 ;
  assign n3148 = n3146 & ~n3147 ;
  assign n3149 = ~x11 & ~n3148 ;
  assign n3150 = ~x11 & ~n3149 ;
  assign n3151 = ~n3148 & ~n3149 ;
  assign n3152 = ~n3150 & ~n3151 ;
  assign n3153 = ~n2902 & ~n2905 ;
  assign n3154 = ~n2883 & n2895 ;
  assign n3155 = ~n2899 & ~n3154 ;
  assign n3156 = ~x66 & n2751 ;
  assign n3157 = ~x64 & n3020 ;
  assign n3158 = ~x65 & n2746 ;
  assign n3159 = ~n3157 & ~n3158 ;
  assign n3160 = ~n3156 & n3159 ;
  assign n3161 = n214 & n2754 ;
  assign n3162 = n3160 & ~n3161 ;
  assign n3163 = ~x20 & ~n3162 ;
  assign n3164 = ~x20 & ~n3163 ;
  assign n3165 = ~n3162 & ~n3163 ;
  assign n3166 = ~n3164 & ~n3165 ;
  assign n3167 = ~n2893 & n3166 ;
  assign n3168 = n2893 & ~n3166 ;
  assign n3169 = ~n3167 & ~n3168 ;
  assign n3170 = ~x69 & n2093 ;
  assign n3171 = ~x67 & n2275 ;
  assign n3172 = ~x68 & n2088 ;
  assign n3173 = ~n3171 & ~n3172 ;
  assign n3174 = ~n3170 & n3173 ;
  assign n3175 = n435 & n2096 ;
  assign n3176 = n3174 & ~n3175 ;
  assign n3177 = ~x17 & ~n3176 ;
  assign n3178 = ~x17 & ~n3177 ;
  assign n3179 = ~n3176 & ~n3177 ;
  assign n3180 = ~n3178 & ~n3179 ;
  assign n3181 = n3169 & ~n3180 ;
  assign n3182 = ~n3169 & n3180 ;
  assign n3183 = ~n3155 & ~n3182 ;
  assign n3184 = ~n3181 & n3183 ;
  assign n3185 = ~n3155 & ~n3184 ;
  assign n3186 = ~n3181 & ~n3184 ;
  assign n3187 = ~n3182 & n3186 ;
  assign n3188 = ~n3185 & ~n3187 ;
  assign n3189 = ~x72 & n1434 ;
  assign n3190 = ~x70 & n1646 ;
  assign n3191 = ~x71 & n1429 ;
  assign n3192 = ~n3190 & ~n3191 ;
  assign n3193 = ~n3189 & n3192 ;
  assign n3194 = n773 & n1437 ;
  assign n3195 = n3193 & ~n3194 ;
  assign n3196 = ~x14 & ~n3195 ;
  assign n3197 = ~x14 & ~n3196 ;
  assign n3198 = ~n3195 & ~n3196 ;
  assign n3199 = ~n3197 & ~n3198 ;
  assign n3200 = n3188 & n3199 ;
  assign n3201 = ~n3188 & ~n3199 ;
  assign n3202 = ~n3200 & ~n3201 ;
  assign n3203 = ~n3153 & n3202 ;
  assign n3204 = n3153 & ~n3202 ;
  assign n3205 = ~n3203 & ~n3204 ;
  assign n3206 = n3152 & ~n3205 ;
  assign n3207 = ~n3152 & n3205 ;
  assign n3208 = ~n3206 & ~n3207 ;
  assign n3209 = ~n3141 & n3208 ;
  assign n3210 = n3141 & ~n3208 ;
  assign n3211 = ~n3209 & ~n3210 ;
  assign n3212 = ~x78 & n574 ;
  assign n3213 = ~x76 & n673 ;
  assign n3214 = ~x77 & n569 ;
  assign n3215 = ~n3213 & ~n3214 ;
  assign n3216 = ~n3212 & n3215 ;
  assign n3217 = n577 & n1718 ;
  assign n3218 = n3216 & ~n3217 ;
  assign n3219 = ~x8 & ~n3218 ;
  assign n3220 = ~x8 & ~n3219 ;
  assign n3221 = ~n3218 & ~n3219 ;
  assign n3222 = ~n3220 & ~n3221 ;
  assign n3223 = n3211 & ~n3222 ;
  assign n3224 = n3211 & ~n3223 ;
  assign n3225 = ~n3222 & ~n3223 ;
  assign n3226 = ~n3224 & ~n3225 ;
  assign n3227 = ~n2939 & ~n2942 ;
  assign n3228 = ~n3226 & ~n3227 ;
  assign n3229 = n3226 & n3227 ;
  assign n3230 = ~n3228 & ~n3229 ;
  assign n3231 = ~n3140 & n3230 ;
  assign n3232 = ~n3140 & ~n3231 ;
  assign n3233 = n3230 & ~n3231 ;
  assign n3234 = ~n3232 & ~n3233 ;
  assign n3235 = ~n3129 & ~n3234 ;
  assign n3236 = ~n3129 & ~n3235 ;
  assign n3237 = ~n3234 & ~n3235 ;
  assign n3238 = ~n3236 & ~n3237 ;
  assign n3239 = ~x84 & n164 ;
  assign n3240 = ~x82 & n205 ;
  assign n3241 = ~x83 & n162 ;
  assign n3242 = ~n3240 & ~n3241 ;
  assign n3243 = ~n3239 & n3242 ;
  assign n3244 = ~n2838 & ~n2970 ;
  assign n3245 = n3111 & ~n3244 ;
  assign n3246 = ~n3111 & n3244 ;
  assign n3247 = ~n3245 & ~n3246 ;
  assign n3248 = n167 & n3247 ;
  assign n3249 = n3243 & ~n3248 ;
  assign n3250 = ~x2 & ~n3249 ;
  assign n3251 = ~x2 & ~n3250 ;
  assign n3252 = ~n3249 & ~n3250 ;
  assign n3253 = ~n3251 & ~n3252 ;
  assign n3254 = ~n3238 & ~n3253 ;
  assign n3255 = ~n3238 & ~n3254 ;
  assign n3256 = ~n3253 & ~n3254 ;
  assign n3257 = ~n3255 & ~n3256 ;
  assign n3258 = ~n2979 & ~n2984 ;
  assign n3259 = ~n3257 & ~n3258 ;
  assign n3260 = n3257 & n3258 ;
  assign n3261 = ~n3259 & ~n3260 ;
  assign n3264 = ~n3261 & ~x148 ;
  assign n3265 = ~n3263 & ~n3264 ;
  assign n3266 = ~n3087 & ~n3092 ;
  assign n3267 = x79 & n574 ;
  assign n3268 = x77 & n673 ;
  assign n3269 = x78 & n569 ;
  assign n3270 = ~n3268 & ~n3269 ;
  assign n3271 = ~n3267 & n3270 ;
  assign n3272 = n577 & n1817 ;
  assign n3273 = n3271 & ~n3272 ;
  assign n3274 = x8 & ~n3273 ;
  assign n3275 = x8 & ~n3274 ;
  assign n3276 = ~n3273 & ~n3274 ;
  assign n3277 = ~n3275 & ~n3276 ;
  assign n3278 = ~n3071 & ~n3073 ;
  assign n3279 = x76 & n945 ;
  assign n3280 = x74 & n1099 ;
  assign n3281 = x75 & n940 ;
  assign n3282 = ~n3280 & ~n3281 ;
  assign n3283 = ~n3279 & n3282 ;
  assign n3284 = n948 & n1311 ;
  assign n3285 = n3283 & ~n3284 ;
  assign n3286 = x11 & ~n3285 ;
  assign n3287 = x11 & ~n3286 ;
  assign n3288 = ~n3285 & ~n3286 ;
  assign n3289 = ~n3287 & ~n3288 ;
  assign n3290 = ~n3065 & ~n3067 ;
  assign n3291 = x20 & ~x21 ;
  assign n3292 = ~x20 & x21 ;
  assign n3293 = ~n3291 & ~n3292 ;
  assign n3294 = x64 & ~n3293 ;
  assign n3295 = ~n3032 & n3294 ;
  assign n3296 = n3032 & ~n3294 ;
  assign n3297 = ~n3295 & ~n3296 ;
  assign n3298 = x67 & n2751 ;
  assign n3299 = x65 & n3020 ;
  assign n3300 = x66 & n2746 ;
  assign n3301 = ~n3299 & ~n3300 ;
  assign n3302 = ~n3298 & n3301 ;
  assign n3303 = n240 & n2754 ;
  assign n3304 = n3302 & ~n3303 ;
  assign n3305 = x20 & ~n3304 ;
  assign n3306 = x20 & ~n3305 ;
  assign n3307 = ~n3304 & ~n3305 ;
  assign n3308 = ~n3306 & ~n3307 ;
  assign n3309 = ~n3297 & ~n3308 ;
  assign n3310 = n3297 & n3308 ;
  assign n3311 = ~n3309 & ~n3310 ;
  assign n3312 = x70 & n2093 ;
  assign n3313 = x68 & n2275 ;
  assign n3314 = x69 & n2088 ;
  assign n3315 = ~n3313 & ~n3314 ;
  assign n3316 = ~n3312 & n3315 ;
  assign n3317 = n488 & n2096 ;
  assign n3318 = n3316 & ~n3317 ;
  assign n3319 = x17 & ~n3318 ;
  assign n3320 = x17 & ~n3319 ;
  assign n3321 = ~n3318 & ~n3319 ;
  assign n3322 = ~n3320 & ~n3321 ;
  assign n3323 = n3311 & ~n3322 ;
  assign n3324 = n3311 & ~n3323 ;
  assign n3325 = ~n3322 & ~n3323 ;
  assign n3326 = ~n3324 & ~n3325 ;
  assign n3327 = ~n3050 & n3326 ;
  assign n3328 = n3050 & ~n3326 ;
  assign n3329 = ~n3327 & ~n3328 ;
  assign n3330 = x73 & n1434 ;
  assign n3331 = x71 & n1646 ;
  assign n3332 = x72 & n1429 ;
  assign n3333 = ~n3331 & ~n3332 ;
  assign n3334 = ~n3330 & n3333 ;
  assign n3335 = n843 & n1437 ;
  assign n3336 = n3334 & ~n3335 ;
  assign n3337 = x14 & ~n3336 ;
  assign n3338 = x14 & ~n3337 ;
  assign n3339 = ~n3336 & ~n3337 ;
  assign n3340 = ~n3338 & ~n3339 ;
  assign n3341 = ~n3329 & ~n3340 ;
  assign n3342 = n3329 & n3340 ;
  assign n3343 = ~n3341 & ~n3342 ;
  assign n3344 = ~n3290 & n3343 ;
  assign n3345 = n3290 & ~n3343 ;
  assign n3346 = ~n3344 & ~n3345 ;
  assign n3347 = n3289 & ~n3346 ;
  assign n3348 = ~n3289 & n3346 ;
  assign n3349 = ~n3347 & ~n3348 ;
  assign n3350 = ~n3278 & n3349 ;
  assign n3351 = n3278 & ~n3349 ;
  assign n3352 = ~n3350 & ~n3351 ;
  assign n3353 = ~n3277 & n3352 ;
  assign n3354 = n3277 & ~n3352 ;
  assign n3355 = ~n3353 & ~n3354 ;
  assign n3356 = ~n3266 & n3355 ;
  assign n3357 = n3266 & ~n3355 ;
  assign n3358 = ~n3356 & ~n3357 ;
  assign n3359 = x82 & n293 ;
  assign n3360 = x80 & n373 ;
  assign n3361 = x81 & n288 ;
  assign n3362 = ~n3360 & ~n3361 ;
  assign n3363 = ~n3359 & n3362 ;
  assign n3364 = n296 & n2584 ;
  assign n3365 = n3363 & ~n3364 ;
  assign n3366 = x5 & ~n3365 ;
  assign n3367 = x5 & ~n3366 ;
  assign n3368 = ~n3365 & ~n3366 ;
  assign n3369 = ~n3367 & ~n3368 ;
  assign n3370 = n3358 & ~n3369 ;
  assign n3371 = n3358 & ~n3370 ;
  assign n3372 = ~n3369 & ~n3370 ;
  assign n3373 = ~n3371 & ~n3372 ;
  assign n3374 = ~n3095 & ~n3099 ;
  assign n3375 = n3373 & n3374 ;
  assign n3376 = ~n3373 & ~n3374 ;
  assign n3377 = ~n3375 & ~n3376 ;
  assign n3378 = x85 & n146 ;
  assign n3379 = x83 & n182 ;
  assign n3380 = x84 & n141 ;
  assign n3381 = ~n3379 & ~n3380 ;
  assign n3382 = ~n3378 & n3381 ;
  assign n3383 = ~n3110 & ~n3112 ;
  assign n3384 = ~x84 & ~x85 ;
  assign n3385 = x84 & x85 ;
  assign n3386 = ~n3384 & ~n3385 ;
  assign n3387 = ~n3383 & n3386 ;
  assign n3388 = n3383 & ~n3386 ;
  assign n3389 = ~n3387 & ~n3388 ;
  assign n3390 = n149 & n3389 ;
  assign n3391 = n3382 & ~n3390 ;
  assign n3392 = x2 & ~n3391 ;
  assign n3393 = x2 & ~n3392 ;
  assign n3394 = ~n3391 & ~n3392 ;
  assign n3395 = ~n3393 & ~n3394 ;
  assign n3396 = n3377 & ~n3395 ;
  assign n3397 = n3377 & ~n3396 ;
  assign n3398 = ~n3395 & ~n3396 ;
  assign n3399 = ~n3397 & ~n3398 ;
  assign n3400 = ~n3121 & ~n3126 ;
  assign n3401 = ~n3399 & ~n3400 ;
  assign n3402 = n3399 & n3400 ;
  assign n3403 = ~n3401 & ~n3402 ;
  assign n3537 = n3403 & x149 ;
  assign n3404 = ~n3223 & ~n3228 ;
  assign n3405 = ~x79 & n574 ;
  assign n3406 = ~x77 & n673 ;
  assign n3407 = ~x78 & n569 ;
  assign n3408 = ~n3406 & ~n3407 ;
  assign n3409 = ~n3405 & n3408 ;
  assign n3410 = n577 & n1921 ;
  assign n3411 = n3409 & ~n3410 ;
  assign n3412 = ~x8 & ~n3411 ;
  assign n3413 = ~x8 & ~n3412 ;
  assign n3414 = ~n3411 & ~n3412 ;
  assign n3415 = ~n3413 & ~n3414 ;
  assign n3416 = ~n3207 & ~n3209 ;
  assign n3417 = ~x76 & n945 ;
  assign n3418 = ~x74 & n1099 ;
  assign n3419 = ~x75 & n940 ;
  assign n3420 = ~n3418 & ~n3419 ;
  assign n3421 = ~n3417 & n3420 ;
  assign n3422 = n948 & n1390 ;
  assign n3423 = n3421 & ~n3422 ;
  assign n3424 = ~x11 & ~n3423 ;
  assign n3425 = ~x11 & ~n3424 ;
  assign n3426 = ~n3423 & ~n3424 ;
  assign n3427 = ~n3425 & ~n3426 ;
  assign n3428 = ~n3201 & ~n3203 ;
  assign n3429 = ~x64 & ~n3293 ;
  assign n3430 = ~n3168 & n3429 ;
  assign n3431 = n3168 & ~n3429 ;
  assign n3432 = ~n3430 & ~n3431 ;
  assign n3433 = ~x67 & n2751 ;
  assign n3434 = ~x65 & n3020 ;
  assign n3435 = ~x66 & n2746 ;
  assign n3436 = ~n3434 & ~n3435 ;
  assign n3437 = ~n3433 & n3436 ;
  assign n3438 = n266 & n2754 ;
  assign n3439 = n3437 & ~n3438 ;
  assign n3440 = ~x20 & ~n3439 ;
  assign n3441 = ~x20 & ~n3440 ;
  assign n3442 = ~n3439 & ~n3440 ;
  assign n3443 = ~n3441 & ~n3442 ;
  assign n3444 = ~n3432 & ~n3443 ;
  assign n3445 = n3432 & n3443 ;
  assign n3446 = ~n3444 & ~n3445 ;
  assign n3447 = ~x70 & n2093 ;
  assign n3448 = ~x68 & n2275 ;
  assign n3449 = ~x69 & n2088 ;
  assign n3450 = ~n3448 & ~n3449 ;
  assign n3451 = ~n3447 & n3450 ;
  assign n3452 = n529 & n2096 ;
  assign n3453 = n3451 & ~n3452 ;
  assign n3454 = ~x17 & ~n3453 ;
  assign n3455 = ~x17 & ~n3454 ;
  assign n3456 = ~n3453 & ~n3454 ;
  assign n3457 = ~n3455 & ~n3456 ;
  assign n3458 = n3446 & ~n3457 ;
  assign n3459 = n3446 & ~n3458 ;
  assign n3460 = ~n3457 & ~n3458 ;
  assign n3461 = ~n3459 & ~n3460 ;
  assign n3462 = ~n3186 & n3461 ;
  assign n3463 = n3186 & ~n3461 ;
  assign n3464 = ~n3462 & ~n3463 ;
  assign n3465 = ~x73 & n1434 ;
  assign n3466 = ~x71 & n1646 ;
  assign n3467 = ~x72 & n1429 ;
  assign n3468 = ~n3466 & ~n3467 ;
  assign n3469 = ~n3465 & n3468 ;
  assign n3470 = n903 & n1437 ;
  assign n3471 = n3469 & ~n3470 ;
  assign n3472 = ~x14 & ~n3471 ;
  assign n3473 = ~x14 & ~n3472 ;
  assign n3474 = ~n3471 & ~n3472 ;
  assign n3475 = ~n3473 & ~n3474 ;
  assign n3476 = ~n3464 & ~n3475 ;
  assign n3477 = n3464 & n3475 ;
  assign n3478 = ~n3476 & ~n3477 ;
  assign n3479 = ~n3428 & n3478 ;
  assign n3480 = n3428 & ~n3478 ;
  assign n3481 = ~n3479 & ~n3480 ;
  assign n3482 = n3427 & ~n3481 ;
  assign n3483 = ~n3427 & n3481 ;
  assign n3484 = ~n3482 & ~n3483 ;
  assign n3485 = ~n3416 & n3484 ;
  assign n3486 = n3416 & ~n3484 ;
  assign n3487 = ~n3485 & ~n3486 ;
  assign n3488 = ~n3415 & n3487 ;
  assign n3489 = n3415 & ~n3487 ;
  assign n3490 = ~n3488 & ~n3489 ;
  assign n3491 = ~n3404 & n3490 ;
  assign n3492 = n3404 & ~n3490 ;
  assign n3493 = ~n3491 & ~n3492 ;
  assign n3494 = ~x82 & n293 ;
  assign n3495 = ~x80 & n373 ;
  assign n3496 = ~x81 & n288 ;
  assign n3497 = ~n3495 & ~n3496 ;
  assign n3498 = ~n3494 & n3497 ;
  assign n3499 = n296 & n2697 ;
  assign n3500 = n3498 & ~n3499 ;
  assign n3501 = ~x5 & ~n3500 ;
  assign n3502 = ~x5 & ~n3501 ;
  assign n3503 = ~n3500 & ~n3501 ;
  assign n3504 = ~n3502 & ~n3503 ;
  assign n3505 = n3493 & ~n3504 ;
  assign n3506 = n3493 & ~n3505 ;
  assign n3507 = ~n3504 & ~n3505 ;
  assign n3508 = ~n3506 & ~n3507 ;
  assign n3509 = ~n3231 & ~n3235 ;
  assign n3510 = n3508 & n3509 ;
  assign n3511 = ~n3508 & ~n3509 ;
  assign n3512 = ~n3510 & ~n3511 ;
  assign n3513 = ~x85 & n164 ;
  assign n3514 = ~x83 & n205 ;
  assign n3515 = ~x84 & n162 ;
  assign n3516 = ~n3514 & ~n3515 ;
  assign n3517 = ~n3513 & n3516 ;
  assign n3518 = ~n3109 & ~n3245 ;
  assign n3519 = n3386 & ~n3518 ;
  assign n3520 = ~n3386 & n3518 ;
  assign n3521 = ~n3519 & ~n3520 ;
  assign n3522 = n167 & n3521 ;
  assign n3523 = n3517 & ~n3522 ;
  assign n3524 = ~x2 & ~n3523 ;
  assign n3525 = ~x2 & ~n3524 ;
  assign n3526 = ~n3523 & ~n3524 ;
  assign n3527 = ~n3525 & ~n3526 ;
  assign n3528 = n3512 & ~n3527 ;
  assign n3529 = n3512 & ~n3528 ;
  assign n3530 = ~n3527 & ~n3528 ;
  assign n3531 = ~n3529 & ~n3530 ;
  assign n3532 = ~n3254 & ~n3259 ;
  assign n3533 = ~n3531 & ~n3532 ;
  assign n3534 = n3531 & n3532 ;
  assign n3535 = ~n3533 & ~n3534 ;
  assign n3538 = ~n3535 & ~x149 ;
  assign n3539 = ~n3537 & ~n3538 ;
  assign n3540 = ~n3396 & ~n3401 ;
  assign n3541 = ~n3353 & ~n3356 ;
  assign n3542 = x80 & n574 ;
  assign n3543 = x78 & n673 ;
  assign n3544 = x79 & n569 ;
  assign n3545 = ~n3543 & ~n3544 ;
  assign n3546 = ~n3542 & n3545 ;
  assign n3547 = n577 & n2028 ;
  assign n3548 = n3546 & ~n3547 ;
  assign n3549 = x8 & ~n3548 ;
  assign n3550 = x8 & ~n3549 ;
  assign n3551 = ~n3548 & ~n3549 ;
  assign n3552 = ~n3550 & ~n3551 ;
  assign n3553 = ~n3348 & ~n3350 ;
  assign n3554 = ~n3050 & ~n3326 ;
  assign n3555 = ~n3323 & ~n3554 ;
  assign n3556 = x71 & n2093 ;
  assign n3557 = x69 & n2275 ;
  assign n3558 = x70 & n2088 ;
  assign n3559 = ~n3557 & ~n3558 ;
  assign n3560 = ~n3556 & n3559 ;
  assign n3561 = n558 & n2096 ;
  assign n3562 = n3560 & ~n3561 ;
  assign n3563 = x17 & ~n3562 ;
  assign n3564 = x17 & ~n3563 ;
  assign n3565 = ~n3562 & ~n3563 ;
  assign n3566 = ~n3564 & ~n3565 ;
  assign n3567 = n3032 & n3294 ;
  assign n3568 = ~n3309 & ~n3567 ;
  assign n3569 = x68 & n2751 ;
  assign n3570 = x66 & n3020 ;
  assign n3571 = x67 & n2746 ;
  assign n3572 = ~n3570 & ~n3571 ;
  assign n3573 = ~n3569 & n3572 ;
  assign n3574 = n317 & n2754 ;
  assign n3575 = n3573 & ~n3574 ;
  assign n3576 = x20 & ~n3575 ;
  assign n3577 = x20 & ~n3576 ;
  assign n3578 = ~n3575 & ~n3576 ;
  assign n3579 = ~n3577 & ~n3578 ;
  assign n3580 = x23 & ~n3294 ;
  assign n3581 = ~x21 & x22 ;
  assign n3582 = x21 & ~x22 ;
  assign n3583 = ~n3581 & ~n3582 ;
  assign n3584 = n3293 & ~n3583 ;
  assign n3585 = x64 & n3584 ;
  assign n3586 = ~x22 & x23 ;
  assign n3587 = x22 & ~x23 ;
  assign n3588 = ~n3586 & ~n3587 ;
  assign n3589 = ~n3293 & n3588 ;
  assign n3590 = x65 & n3589 ;
  assign n3591 = ~n3585 & ~n3590 ;
  assign n3592 = ~n3293 & ~n3588 ;
  assign n3593 = ~n152 & n3592 ;
  assign n3594 = n3591 & ~n3593 ;
  assign n3595 = x23 & ~n3594 ;
  assign n3596 = x23 & ~n3595 ;
  assign n3597 = ~n3594 & ~n3595 ;
  assign n3598 = ~n3596 & ~n3597 ;
  assign n3599 = n3580 & ~n3598 ;
  assign n3600 = ~n3580 & n3598 ;
  assign n3601 = ~n3599 & ~n3600 ;
  assign n3602 = n3579 & n3601 ;
  assign n3603 = ~n3579 & ~n3601 ;
  assign n3604 = ~n3602 & ~n3603 ;
  assign n3605 = ~n3568 & ~n3604 ;
  assign n3606 = n3568 & n3604 ;
  assign n3607 = ~n3605 & ~n3606 ;
  assign n3608 = ~n3566 & n3607 ;
  assign n3609 = n3566 & ~n3607 ;
  assign n3610 = ~n3608 & ~n3609 ;
  assign n3611 = ~n3555 & n3610 ;
  assign n3612 = n3555 & ~n3610 ;
  assign n3613 = ~n3611 & ~n3612 ;
  assign n3614 = x74 & n1434 ;
  assign n3615 = x72 & n1646 ;
  assign n3616 = x73 & n1429 ;
  assign n3617 = ~n3615 & ~n3616 ;
  assign n3618 = ~n3614 & n3617 ;
  assign n3619 = n994 & n1437 ;
  assign n3620 = n3618 & ~n3619 ;
  assign n3621 = x14 & ~n3620 ;
  assign n3622 = x14 & ~n3621 ;
  assign n3623 = ~n3620 & ~n3621 ;
  assign n3624 = ~n3622 & ~n3623 ;
  assign n3625 = n3613 & ~n3624 ;
  assign n3626 = n3613 & ~n3625 ;
  assign n3627 = ~n3624 & ~n3625 ;
  assign n3628 = ~n3626 & ~n3627 ;
  assign n3629 = ~n3341 & ~n3344 ;
  assign n3630 = n3628 & n3629 ;
  assign n3631 = ~n3628 & ~n3629 ;
  assign n3632 = ~n3630 & ~n3631 ;
  assign n3633 = x77 & n945 ;
  assign n3634 = x75 & n1099 ;
  assign n3635 = x76 & n940 ;
  assign n3636 = ~n3634 & ~n3635 ;
  assign n3637 = ~n3633 & n3636 ;
  assign n3638 = n948 & n1502 ;
  assign n3639 = n3637 & ~n3638 ;
  assign n3640 = x11 & ~n3639 ;
  assign n3641 = x11 & ~n3640 ;
  assign n3642 = ~n3639 & ~n3640 ;
  assign n3643 = ~n3641 & ~n3642 ;
  assign n3644 = ~n3632 & n3643 ;
  assign n3645 = n3632 & ~n3643 ;
  assign n3646 = ~n3644 & ~n3645 ;
  assign n3647 = ~n3553 & n3646 ;
  assign n3648 = n3553 & ~n3646 ;
  assign n3649 = ~n3647 & ~n3648 ;
  assign n3650 = ~n3552 & n3649 ;
  assign n3651 = n3552 & ~n3649 ;
  assign n3652 = ~n3650 & ~n3651 ;
  assign n3653 = ~n3541 & n3652 ;
  assign n3654 = n3541 & ~n3652 ;
  assign n3655 = ~n3653 & ~n3654 ;
  assign n3656 = x83 & n293 ;
  assign n3657 = x81 & n373 ;
  assign n3658 = x82 & n288 ;
  assign n3659 = ~n3657 & ~n3658 ;
  assign n3660 = ~n3656 & n3659 ;
  assign n3661 = n296 & n2843 ;
  assign n3662 = n3660 & ~n3661 ;
  assign n3663 = x5 & ~n3662 ;
  assign n3664 = x5 & ~n3663 ;
  assign n3665 = ~n3662 & ~n3663 ;
  assign n3666 = ~n3664 & ~n3665 ;
  assign n3667 = n3655 & ~n3666 ;
  assign n3668 = n3655 & ~n3667 ;
  assign n3669 = ~n3666 & ~n3667 ;
  assign n3670 = ~n3668 & ~n3669 ;
  assign n3671 = ~n3370 & ~n3376 ;
  assign n3672 = n3670 & n3671 ;
  assign n3673 = ~n3670 & ~n3671 ;
  assign n3674 = ~n3672 & ~n3673 ;
  assign n3675 = x86 & n146 ;
  assign n3676 = x84 & n182 ;
  assign n3677 = x85 & n141 ;
  assign n3678 = ~n3676 & ~n3677 ;
  assign n3679 = ~n3675 & n3678 ;
  assign n3680 = ~n3385 & ~n3387 ;
  assign n3681 = ~x85 & ~x86 ;
  assign n3682 = x85 & x86 ;
  assign n3683 = ~n3681 & ~n3682 ;
  assign n3684 = ~n3680 & n3683 ;
  assign n3685 = n3680 & ~n3683 ;
  assign n3686 = ~n3684 & ~n3685 ;
  assign n3687 = n149 & n3686 ;
  assign n3688 = n3679 & ~n3687 ;
  assign n3689 = x2 & ~n3688 ;
  assign n3690 = x2 & ~n3689 ;
  assign n3691 = ~n3688 & ~n3689 ;
  assign n3692 = ~n3690 & ~n3691 ;
  assign n3693 = ~n3674 & n3692 ;
  assign n3694 = n3674 & ~n3692 ;
  assign n3695 = ~n3693 & ~n3694 ;
  assign n3696 = ~n3540 & n3695 ;
  assign n3697 = n3540 & ~n3695 ;
  assign n3698 = ~n3696 & ~n3697 ;
  assign n3846 = n3698 & x150 ;
  assign n3699 = ~n3528 & ~n3533 ;
  assign n3700 = ~n3488 & ~n3491 ;
  assign n3701 = ~x80 & n574 ;
  assign n3702 = ~x78 & n673 ;
  assign n3703 = ~x79 & n569 ;
  assign n3704 = ~n3702 & ~n3703 ;
  assign n3705 = ~n3701 & n3704 ;
  assign n3706 = n577 & n2145 ;
  assign n3707 = n3705 & ~n3706 ;
  assign n3708 = ~x8 & ~n3707 ;
  assign n3709 = ~x8 & ~n3708 ;
  assign n3710 = ~n3707 & ~n3708 ;
  assign n3711 = ~n3709 & ~n3710 ;
  assign n3712 = ~n3483 & ~n3485 ;
  assign n3713 = ~n3186 & ~n3461 ;
  assign n3714 = ~n3458 & ~n3713 ;
  assign n3715 = ~x71 & n2093 ;
  assign n3716 = ~x69 & n2275 ;
  assign n3717 = ~x70 & n2088 ;
  assign n3718 = ~n3716 & ~n3717 ;
  assign n3719 = ~n3715 & n3718 ;
  assign n3720 = n622 & n2096 ;
  assign n3721 = n3719 & ~n3720 ;
  assign n3722 = ~x17 & ~n3721 ;
  assign n3723 = ~x17 & ~n3722 ;
  assign n3724 = ~n3721 & ~n3722 ;
  assign n3725 = ~n3723 & ~n3724 ;
  assign n3726 = n3168 & n3429 ;
  assign n3727 = ~n3444 & ~n3726 ;
  assign n3728 = ~x68 & n2751 ;
  assign n3729 = ~x66 & n3020 ;
  assign n3730 = ~x67 & n2746 ;
  assign n3731 = ~n3729 & ~n3730 ;
  assign n3732 = ~n3728 & n3731 ;
  assign n3733 = n352 & n2754 ;
  assign n3734 = n3732 & ~n3733 ;
  assign n3735 = ~x20 & ~n3734 ;
  assign n3736 = ~x20 & ~n3735 ;
  assign n3737 = ~n3734 & ~n3735 ;
  assign n3738 = ~n3736 & ~n3737 ;
  assign n3739 = ~x23 & ~n3429 ;
  assign n3740 = ~x64 & n3584 ;
  assign n3741 = ~x65 & n3589 ;
  assign n3742 = ~n3740 & ~n3741 ;
  assign n3743 = ~n3593 & n3742 ;
  assign n3744 = ~x23 & ~n3743 ;
  assign n3745 = ~x23 & ~n3744 ;
  assign n3746 = ~n3743 & ~n3744 ;
  assign n3747 = ~n3745 & ~n3746 ;
  assign n3748 = n3739 & ~n3747 ;
  assign n3749 = ~n3739 & n3747 ;
  assign n3750 = ~n3748 & ~n3749 ;
  assign n3751 = n3738 & n3750 ;
  assign n3752 = ~n3738 & ~n3750 ;
  assign n3753 = ~n3751 & ~n3752 ;
  assign n3754 = ~n3727 & ~n3753 ;
  assign n3755 = n3727 & n3753 ;
  assign n3756 = ~n3754 & ~n3755 ;
  assign n3757 = ~n3725 & n3756 ;
  assign n3758 = n3725 & ~n3756 ;
  assign n3759 = ~n3757 & ~n3758 ;
  assign n3760 = ~n3714 & n3759 ;
  assign n3761 = n3714 & ~n3759 ;
  assign n3762 = ~n3760 & ~n3761 ;
  assign n3763 = ~x74 & n1434 ;
  assign n3764 = ~x72 & n1646 ;
  assign n3765 = ~x73 & n1429 ;
  assign n3766 = ~n3764 & ~n3765 ;
  assign n3767 = ~n3763 & n3766 ;
  assign n3768 = n1066 & n1437 ;
  assign n3769 = n3767 & ~n3768 ;
  assign n3770 = ~x14 & ~n3769 ;
  assign n3771 = ~x14 & ~n3770 ;
  assign n3772 = ~n3769 & ~n3770 ;
  assign n3773 = ~n3771 & ~n3772 ;
  assign n3774 = n3762 & ~n3773 ;
  assign n3775 = n3762 & ~n3774 ;
  assign n3776 = ~n3773 & ~n3774 ;
  assign n3777 = ~n3775 & ~n3776 ;
  assign n3778 = ~n3476 & ~n3479 ;
  assign n3779 = n3777 & n3778 ;
  assign n3780 = ~n3777 & ~n3778 ;
  assign n3781 = ~n3779 & ~n3780 ;
  assign n3782 = ~x77 & n945 ;
  assign n3783 = ~x75 & n1099 ;
  assign n3784 = ~x76 & n940 ;
  assign n3785 = ~n3783 & ~n3784 ;
  assign n3786 = ~n3782 & n3785 ;
  assign n3787 = n948 & n1594 ;
  assign n3788 = n3786 & ~n3787 ;
  assign n3789 = ~x11 & ~n3788 ;
  assign n3790 = ~x11 & ~n3789 ;
  assign n3791 = ~n3788 & ~n3789 ;
  assign n3792 = ~n3790 & ~n3791 ;
  assign n3793 = ~n3781 & n3792 ;
  assign n3794 = n3781 & ~n3792 ;
  assign n3795 = ~n3793 & ~n3794 ;
  assign n3796 = ~n3712 & n3795 ;
  assign n3797 = n3712 & ~n3795 ;
  assign n3798 = ~n3796 & ~n3797 ;
  assign n3799 = ~n3711 & n3798 ;
  assign n3800 = n3711 & ~n3798 ;
  assign n3801 = ~n3799 & ~n3800 ;
  assign n3802 = ~n3700 & n3801 ;
  assign n3803 = n3700 & ~n3801 ;
  assign n3804 = ~n3802 & ~n3803 ;
  assign n3805 = ~x83 & n293 ;
  assign n3806 = ~x81 & n373 ;
  assign n3807 = ~x82 & n288 ;
  assign n3808 = ~n3806 & ~n3807 ;
  assign n3809 = ~n3805 & n3808 ;
  assign n3810 = n296 & n2972 ;
  assign n3811 = n3809 & ~n3810 ;
  assign n3812 = ~x5 & ~n3811 ;
  assign n3813 = ~x5 & ~n3812 ;
  assign n3814 = ~n3811 & ~n3812 ;
  assign n3815 = ~n3813 & ~n3814 ;
  assign n3816 = n3804 & ~n3815 ;
  assign n3817 = n3804 & ~n3816 ;
  assign n3818 = ~n3815 & ~n3816 ;
  assign n3819 = ~n3817 & ~n3818 ;
  assign n3820 = ~n3505 & ~n3511 ;
  assign n3821 = n3819 & n3820 ;
  assign n3822 = ~n3819 & ~n3820 ;
  assign n3823 = ~n3821 & ~n3822 ;
  assign n3824 = ~x86 & n164 ;
  assign n3825 = ~x84 & n205 ;
  assign n3826 = ~x85 & n162 ;
  assign n3827 = ~n3825 & ~n3826 ;
  assign n3828 = ~n3824 & n3827 ;
  assign n3829 = ~n3384 & ~n3519 ;
  assign n3830 = n3683 & ~n3829 ;
  assign n3831 = ~n3683 & n3829 ;
  assign n3832 = ~n3830 & ~n3831 ;
  assign n3833 = n167 & n3832 ;
  assign n3834 = n3828 & ~n3833 ;
  assign n3835 = ~x2 & ~n3834 ;
  assign n3836 = ~x2 & ~n3835 ;
  assign n3837 = ~n3834 & ~n3835 ;
  assign n3838 = ~n3836 & ~n3837 ;
  assign n3839 = ~n3823 & n3838 ;
  assign n3840 = n3823 & ~n3838 ;
  assign n3841 = ~n3839 & ~n3840 ;
  assign n3842 = ~n3699 & n3841 ;
  assign n3843 = n3699 & ~n3841 ;
  assign n3844 = ~n3842 & ~n3843 ;
  assign n3847 = ~n3844 & ~x150 ;
  assign n3848 = ~n3846 & ~n3847 ;
  assign n3849 = ~n3650 & ~n3653 ;
  assign n3850 = x81 & n574 ;
  assign n3851 = x79 & n673 ;
  assign n3852 = x80 & n569 ;
  assign n3853 = ~n3851 & ~n3852 ;
  assign n3854 = ~n3850 & n3853 ;
  assign n3855 = n577 & n2348 ;
  assign n3856 = n3854 & ~n3855 ;
  assign n3857 = x8 & ~n3856 ;
  assign n3858 = x8 & ~n3857 ;
  assign n3859 = ~n3856 & ~n3857 ;
  assign n3860 = ~n3858 & ~n3859 ;
  assign n3861 = ~n3625 & ~n3631 ;
  assign n3862 = x75 & n1434 ;
  assign n3863 = x73 & n1646 ;
  assign n3864 = x74 & n1429 ;
  assign n3865 = ~n3863 & ~n3864 ;
  assign n3866 = ~n3862 & n3865 ;
  assign n3867 = n1150 & n1437 ;
  assign n3868 = n3866 & ~n3867 ;
  assign n3869 = x14 & ~n3868 ;
  assign n3870 = x14 & ~n3869 ;
  assign n3871 = ~n3868 & ~n3869 ;
  assign n3872 = ~n3870 & ~n3871 ;
  assign n3873 = ~n3608 & ~n3611 ;
  assign n3874 = ~n3579 & n3601 ;
  assign n3875 = ~n3605 & ~n3874 ;
  assign n3876 = x66 & n3589 ;
  assign n3877 = n3293 & ~n3588 ;
  assign n3878 = n3583 & n3877 ;
  assign n3879 = x64 & n3878 ;
  assign n3880 = x65 & n3584 ;
  assign n3881 = ~n3879 & ~n3880 ;
  assign n3882 = ~n3876 & n3881 ;
  assign n3883 = n194 & n3592 ;
  assign n3884 = n3882 & ~n3883 ;
  assign n3885 = x23 & ~n3884 ;
  assign n3886 = x23 & ~n3885 ;
  assign n3887 = ~n3884 & ~n3885 ;
  assign n3888 = ~n3886 & ~n3887 ;
  assign n3889 = ~n3599 & n3888 ;
  assign n3890 = n3599 & ~n3888 ;
  assign n3891 = ~n3889 & ~n3890 ;
  assign n3892 = x69 & n2751 ;
  assign n3893 = x67 & n3020 ;
  assign n3894 = x68 & n2746 ;
  assign n3895 = ~n3893 & ~n3894 ;
  assign n3896 = ~n3892 & n3895 ;
  assign n3897 = n398 & n2754 ;
  assign n3898 = n3896 & ~n3897 ;
  assign n3899 = x20 & ~n3898 ;
  assign n3900 = x20 & ~n3899 ;
  assign n3901 = ~n3898 & ~n3899 ;
  assign n3902 = ~n3900 & ~n3901 ;
  assign n3903 = n3891 & ~n3902 ;
  assign n3904 = ~n3891 & n3902 ;
  assign n3905 = ~n3875 & ~n3904 ;
  assign n3906 = ~n3903 & n3905 ;
  assign n3907 = ~n3875 & ~n3906 ;
  assign n3908 = ~n3903 & ~n3906 ;
  assign n3909 = ~n3904 & n3908 ;
  assign n3910 = ~n3907 & ~n3909 ;
  assign n3911 = x72 & n2093 ;
  assign n3912 = x70 & n2275 ;
  assign n3913 = x71 & n2088 ;
  assign n3914 = ~n3912 & ~n3913 ;
  assign n3915 = ~n3911 & n3914 ;
  assign n3916 = n717 & n2096 ;
  assign n3917 = n3915 & ~n3916 ;
  assign n3918 = x17 & ~n3917 ;
  assign n3919 = x17 & ~n3918 ;
  assign n3920 = ~n3917 & ~n3918 ;
  assign n3921 = ~n3919 & ~n3920 ;
  assign n3922 = n3910 & n3921 ;
  assign n3923 = ~n3910 & ~n3921 ;
  assign n3924 = ~n3922 & ~n3923 ;
  assign n3925 = ~n3873 & n3924 ;
  assign n3926 = n3873 & ~n3924 ;
  assign n3927 = ~n3925 & ~n3926 ;
  assign n3928 = n3872 & ~n3927 ;
  assign n3929 = ~n3872 & n3927 ;
  assign n3930 = ~n3928 & ~n3929 ;
  assign n3931 = ~n3861 & n3930 ;
  assign n3932 = n3861 & ~n3930 ;
  assign n3933 = ~n3931 & ~n3932 ;
  assign n3934 = x78 & n945 ;
  assign n3935 = x76 & n1099 ;
  assign n3936 = x77 & n940 ;
  assign n3937 = ~n3935 & ~n3936 ;
  assign n3938 = ~n3934 & n3937 ;
  assign n3939 = n948 & n1624 ;
  assign n3940 = n3938 & ~n3939 ;
  assign n3941 = x11 & ~n3940 ;
  assign n3942 = x11 & ~n3941 ;
  assign n3943 = ~n3940 & ~n3941 ;
  assign n3944 = ~n3942 & ~n3943 ;
  assign n3945 = n3933 & ~n3944 ;
  assign n3946 = n3933 & ~n3945 ;
  assign n3947 = ~n3944 & ~n3945 ;
  assign n3948 = ~n3946 & ~n3947 ;
  assign n3949 = ~n3645 & ~n3647 ;
  assign n3950 = ~n3948 & ~n3949 ;
  assign n3951 = n3948 & n3949 ;
  assign n3952 = ~n3950 & ~n3951 ;
  assign n3953 = ~n3860 & n3952 ;
  assign n3954 = ~n3860 & ~n3953 ;
  assign n3955 = n3952 & ~n3953 ;
  assign n3956 = ~n3954 & ~n3955 ;
  assign n3957 = ~n3849 & ~n3956 ;
  assign n3958 = ~n3849 & ~n3957 ;
  assign n3959 = ~n3956 & ~n3957 ;
  assign n3960 = ~n3958 & ~n3959 ;
  assign n3961 = x84 & n293 ;
  assign n3962 = x82 & n373 ;
  assign n3963 = x83 & n288 ;
  assign n3964 = ~n3962 & ~n3963 ;
  assign n3965 = ~n3961 & n3964 ;
  assign n3966 = n296 & n3114 ;
  assign n3967 = n3965 & ~n3966 ;
  assign n3968 = x5 & ~n3967 ;
  assign n3969 = x5 & ~n3968 ;
  assign n3970 = ~n3967 & ~n3968 ;
  assign n3971 = ~n3969 & ~n3970 ;
  assign n3972 = ~n3960 & ~n3971 ;
  assign n3973 = ~n3960 & ~n3972 ;
  assign n3974 = ~n3971 & ~n3972 ;
  assign n3975 = ~n3973 & ~n3974 ;
  assign n3976 = ~n3667 & ~n3673 ;
  assign n3977 = n3975 & n3976 ;
  assign n3978 = ~n3975 & ~n3976 ;
  assign n3979 = ~n3977 & ~n3978 ;
  assign n3980 = x87 & n146 ;
  assign n3981 = x85 & n182 ;
  assign n3982 = x86 & n141 ;
  assign n3983 = ~n3981 & ~n3982 ;
  assign n3984 = ~n3980 & n3983 ;
  assign n3985 = ~n3682 & ~n3684 ;
  assign n3986 = ~x86 & ~x87 ;
  assign n3987 = x86 & x87 ;
  assign n3988 = ~n3986 & ~n3987 ;
  assign n3989 = ~n3985 & n3988 ;
  assign n3990 = n3985 & ~n3988 ;
  assign n3991 = ~n3989 & ~n3990 ;
  assign n3992 = n149 & n3991 ;
  assign n3993 = n3984 & ~n3992 ;
  assign n3994 = x2 & ~n3993 ;
  assign n3995 = x2 & ~n3994 ;
  assign n3996 = ~n3993 & ~n3994 ;
  assign n3997 = ~n3995 & ~n3996 ;
  assign n3998 = n3979 & ~n3997 ;
  assign n3999 = n3979 & ~n3998 ;
  assign n4000 = ~n3997 & ~n3998 ;
  assign n4001 = ~n3999 & ~n4000 ;
  assign n4002 = ~n3694 & ~n3696 ;
  assign n4003 = ~n4001 & ~n4002 ;
  assign n4004 = n4001 & n4002 ;
  assign n4005 = ~n4003 & ~n4004 ;
  assign n4159 = n4005 & x151 ;
  assign n4006 = ~n3799 & ~n3802 ;
  assign n4007 = ~x81 & n574 ;
  assign n4008 = ~x79 & n673 ;
  assign n4009 = ~x80 & n569 ;
  assign n4010 = ~n4008 & ~n4009 ;
  assign n4011 = ~n4007 & n4010 ;
  assign n4012 = n577 & n2460 ;
  assign n4013 = n4011 & ~n4012 ;
  assign n4014 = ~x8 & ~n4013 ;
  assign n4015 = ~x8 & ~n4014 ;
  assign n4016 = ~n4013 & ~n4014 ;
  assign n4017 = ~n4015 & ~n4016 ;
  assign n4018 = ~n3774 & ~n3780 ;
  assign n4019 = ~x75 & n1434 ;
  assign n4020 = ~x73 & n1646 ;
  assign n4021 = ~x74 & n1429 ;
  assign n4022 = ~n4020 & ~n4021 ;
  assign n4023 = ~n4019 & n4022 ;
  assign n4024 = n1225 & n1437 ;
  assign n4025 = n4023 & ~n4024 ;
  assign n4026 = ~x14 & ~n4025 ;
  assign n4027 = ~x14 & ~n4026 ;
  assign n4028 = ~n4025 & ~n4026 ;
  assign n4029 = ~n4027 & ~n4028 ;
  assign n4030 = ~n3757 & ~n3760 ;
  assign n4031 = ~n3738 & n3750 ;
  assign n4032 = ~n3754 & ~n4031 ;
  assign n4033 = ~x66 & n3589 ;
  assign n4034 = ~x64 & n3878 ;
  assign n4035 = ~x65 & n3584 ;
  assign n4036 = ~n4034 & ~n4035 ;
  assign n4037 = ~n4033 & n4036 ;
  assign n4038 = n214 & n3592 ;
  assign n4039 = n4037 & ~n4038 ;
  assign n4040 = ~x23 & ~n4039 ;
  assign n4041 = ~x23 & ~n4040 ;
  assign n4042 = ~n4039 & ~n4040 ;
  assign n4043 = ~n4041 & ~n4042 ;
  assign n4044 = ~n3748 & n4043 ;
  assign n4045 = n3748 & ~n4043 ;
  assign n4046 = ~n4044 & ~n4045 ;
  assign n4047 = ~x69 & n2751 ;
  assign n4048 = ~x67 & n3020 ;
  assign n4049 = ~x68 & n2746 ;
  assign n4050 = ~n4048 & ~n4049 ;
  assign n4051 = ~n4047 & n4050 ;
  assign n4052 = n435 & n2754 ;
  assign n4053 = n4051 & ~n4052 ;
  assign n4054 = ~x20 & ~n4053 ;
  assign n4055 = ~x20 & ~n4054 ;
  assign n4056 = ~n4053 & ~n4054 ;
  assign n4057 = ~n4055 & ~n4056 ;
  assign n4058 = n4046 & ~n4057 ;
  assign n4059 = ~n4046 & n4057 ;
  assign n4060 = ~n4032 & ~n4059 ;
  assign n4061 = ~n4058 & n4060 ;
  assign n4062 = ~n4032 & ~n4061 ;
  assign n4063 = ~n4058 & ~n4061 ;
  assign n4064 = ~n4059 & n4063 ;
  assign n4065 = ~n4062 & ~n4064 ;
  assign n4066 = ~x72 & n2093 ;
  assign n4067 = ~x70 & n2275 ;
  assign n4068 = ~x71 & n2088 ;
  assign n4069 = ~n4067 & ~n4068 ;
  assign n4070 = ~n4066 & n4069 ;
  assign n4071 = n773 & n2096 ;
  assign n4072 = n4070 & ~n4071 ;
  assign n4073 = ~x17 & ~n4072 ;
  assign n4074 = ~x17 & ~n4073 ;
  assign n4075 = ~n4072 & ~n4073 ;
  assign n4076 = ~n4074 & ~n4075 ;
  assign n4077 = n4065 & n4076 ;
  assign n4078 = ~n4065 & ~n4076 ;
  assign n4079 = ~n4077 & ~n4078 ;
  assign n4080 = ~n4030 & n4079 ;
  assign n4081 = n4030 & ~n4079 ;
  assign n4082 = ~n4080 & ~n4081 ;
  assign n4083 = n4029 & ~n4082 ;
  assign n4084 = ~n4029 & n4082 ;
  assign n4085 = ~n4083 & ~n4084 ;
  assign n4086 = ~n4018 & n4085 ;
  assign n4087 = n4018 & ~n4085 ;
  assign n4088 = ~n4086 & ~n4087 ;
  assign n4089 = ~x78 & n945 ;
  assign n4090 = ~x76 & n1099 ;
  assign n4091 = ~x77 & n940 ;
  assign n4092 = ~n4090 & ~n4091 ;
  assign n4093 = ~n4089 & n4092 ;
  assign n4094 = n948 & n1718 ;
  assign n4095 = n4093 & ~n4094 ;
  assign n4096 = ~x11 & ~n4095 ;
  assign n4097 = ~x11 & ~n4096 ;
  assign n4098 = ~n4095 & ~n4096 ;
  assign n4099 = ~n4097 & ~n4098 ;
  assign n4100 = n4088 & ~n4099 ;
  assign n4101 = n4088 & ~n4100 ;
  assign n4102 = ~n4099 & ~n4100 ;
  assign n4103 = ~n4101 & ~n4102 ;
  assign n4104 = ~n3794 & ~n3796 ;
  assign n4105 = ~n4103 & ~n4104 ;
  assign n4106 = n4103 & n4104 ;
  assign n4107 = ~n4105 & ~n4106 ;
  assign n4108 = ~n4017 & n4107 ;
  assign n4109 = ~n4017 & ~n4108 ;
  assign n4110 = n4107 & ~n4108 ;
  assign n4111 = ~n4109 & ~n4110 ;
  assign n4112 = ~n4006 & ~n4111 ;
  assign n4113 = ~n4006 & ~n4112 ;
  assign n4114 = ~n4111 & ~n4112 ;
  assign n4115 = ~n4113 & ~n4114 ;
  assign n4116 = ~x84 & n293 ;
  assign n4117 = ~x82 & n373 ;
  assign n4118 = ~x83 & n288 ;
  assign n4119 = ~n4117 & ~n4118 ;
  assign n4120 = ~n4116 & n4119 ;
  assign n4121 = n296 & n3247 ;
  assign n4122 = n4120 & ~n4121 ;
  assign n4123 = ~x5 & ~n4122 ;
  assign n4124 = ~x5 & ~n4123 ;
  assign n4125 = ~n4122 & ~n4123 ;
  assign n4126 = ~n4124 & ~n4125 ;
  assign n4127 = ~n4115 & ~n4126 ;
  assign n4128 = ~n4115 & ~n4127 ;
  assign n4129 = ~n4126 & ~n4127 ;
  assign n4130 = ~n4128 & ~n4129 ;
  assign n4131 = ~n3816 & ~n3822 ;
  assign n4132 = n4130 & n4131 ;
  assign n4133 = ~n4130 & ~n4131 ;
  assign n4134 = ~n4132 & ~n4133 ;
  assign n4135 = ~x87 & n164 ;
  assign n4136 = ~x85 & n205 ;
  assign n4137 = ~x86 & n162 ;
  assign n4138 = ~n4136 & ~n4137 ;
  assign n4139 = ~n4135 & n4138 ;
  assign n4140 = ~n3681 & ~n3830 ;
  assign n4141 = n3988 & ~n4140 ;
  assign n4142 = ~n3988 & n4140 ;
  assign n4143 = ~n4141 & ~n4142 ;
  assign n4144 = n167 & n4143 ;
  assign n4145 = n4139 & ~n4144 ;
  assign n4146 = ~x2 & ~n4145 ;
  assign n4147 = ~x2 & ~n4146 ;
  assign n4148 = ~n4145 & ~n4146 ;
  assign n4149 = ~n4147 & ~n4148 ;
  assign n4150 = n4134 & ~n4149 ;
  assign n4151 = n4134 & ~n4150 ;
  assign n4152 = ~n4149 & ~n4150 ;
  assign n4153 = ~n4151 & ~n4152 ;
  assign n4154 = ~n3840 & ~n3842 ;
  assign n4155 = ~n4153 & ~n4154 ;
  assign n4156 = n4153 & n4154 ;
  assign n4157 = ~n4155 & ~n4156 ;
  assign n4160 = ~n4157 & ~x151 ;
  assign n4161 = ~n4159 & ~n4160 ;
  assign n4162 = ~n3972 & ~n3978 ;
  assign n4163 = x85 & n293 ;
  assign n4164 = x83 & n373 ;
  assign n4165 = x84 & n288 ;
  assign n4166 = ~n4164 & ~n4165 ;
  assign n4167 = ~n4163 & n4166 ;
  assign n4168 = n296 & n3389 ;
  assign n4169 = n4167 & ~n4168 ;
  assign n4170 = x5 & ~n4169 ;
  assign n4171 = x5 & ~n4170 ;
  assign n4172 = ~n4169 & ~n4170 ;
  assign n4173 = ~n4171 & ~n4172 ;
  assign n4174 = ~n3953 & ~n3957 ;
  assign n4175 = ~n3929 & ~n3931 ;
  assign n4176 = x76 & n1434 ;
  assign n4177 = x74 & n1646 ;
  assign n4178 = x75 & n1429 ;
  assign n4179 = ~n4177 & ~n4178 ;
  assign n4180 = ~n4176 & n4179 ;
  assign n4181 = n1311 & n1437 ;
  assign n4182 = n4180 & ~n4181 ;
  assign n4183 = x14 & ~n4182 ;
  assign n4184 = x14 & ~n4183 ;
  assign n4185 = ~n4182 & ~n4183 ;
  assign n4186 = ~n4184 & ~n4185 ;
  assign n4187 = ~n3923 & ~n3925 ;
  assign n4188 = x23 & ~x24 ;
  assign n4189 = ~x23 & x24 ;
  assign n4190 = ~n4188 & ~n4189 ;
  assign n4191 = x64 & ~n4190 ;
  assign n4192 = ~n3890 & n4191 ;
  assign n4193 = n3890 & ~n4191 ;
  assign n4194 = ~n4192 & ~n4193 ;
  assign n4195 = x67 & n3589 ;
  assign n4196 = x65 & n3878 ;
  assign n4197 = x66 & n3584 ;
  assign n4198 = ~n4196 & ~n4197 ;
  assign n4199 = ~n4195 & n4198 ;
  assign n4200 = n240 & n3592 ;
  assign n4201 = n4199 & ~n4200 ;
  assign n4202 = x23 & ~n4201 ;
  assign n4203 = x23 & ~n4202 ;
  assign n4204 = ~n4201 & ~n4202 ;
  assign n4205 = ~n4203 & ~n4204 ;
  assign n4206 = ~n4194 & ~n4205 ;
  assign n4207 = n4194 & n4205 ;
  assign n4208 = ~n4206 & ~n4207 ;
  assign n4209 = x70 & n2751 ;
  assign n4210 = x68 & n3020 ;
  assign n4211 = x69 & n2746 ;
  assign n4212 = ~n4210 & ~n4211 ;
  assign n4213 = ~n4209 & n4212 ;
  assign n4214 = n488 & n2754 ;
  assign n4215 = n4213 & ~n4214 ;
  assign n4216 = x20 & ~n4215 ;
  assign n4217 = x20 & ~n4216 ;
  assign n4218 = ~n4215 & ~n4216 ;
  assign n4219 = ~n4217 & ~n4218 ;
  assign n4220 = n4208 & ~n4219 ;
  assign n4221 = n4208 & ~n4220 ;
  assign n4222 = ~n4219 & ~n4220 ;
  assign n4223 = ~n4221 & ~n4222 ;
  assign n4224 = ~n3908 & n4223 ;
  assign n4225 = n3908 & ~n4223 ;
  assign n4226 = ~n4224 & ~n4225 ;
  assign n4227 = x73 & n2093 ;
  assign n4228 = x71 & n2275 ;
  assign n4229 = x72 & n2088 ;
  assign n4230 = ~n4228 & ~n4229 ;
  assign n4231 = ~n4227 & n4230 ;
  assign n4232 = n843 & n2096 ;
  assign n4233 = n4231 & ~n4232 ;
  assign n4234 = x17 & ~n4233 ;
  assign n4235 = x17 & ~n4234 ;
  assign n4236 = ~n4233 & ~n4234 ;
  assign n4237 = ~n4235 & ~n4236 ;
  assign n4238 = ~n4226 & ~n4237 ;
  assign n4239 = n4226 & n4237 ;
  assign n4240 = ~n4238 & ~n4239 ;
  assign n4241 = ~n4187 & n4240 ;
  assign n4242 = n4187 & ~n4240 ;
  assign n4243 = ~n4241 & ~n4242 ;
  assign n4244 = n4186 & ~n4243 ;
  assign n4245 = ~n4186 & n4243 ;
  assign n4246 = ~n4244 & ~n4245 ;
  assign n4247 = ~n4175 & n4246 ;
  assign n4248 = n4175 & ~n4246 ;
  assign n4249 = ~n4247 & ~n4248 ;
  assign n4250 = x79 & n945 ;
  assign n4251 = x77 & n1099 ;
  assign n4252 = x78 & n940 ;
  assign n4253 = ~n4251 & ~n4252 ;
  assign n4254 = ~n4250 & n4253 ;
  assign n4255 = n948 & n1817 ;
  assign n4256 = n4254 & ~n4255 ;
  assign n4257 = x11 & ~n4256 ;
  assign n4258 = x11 & ~n4257 ;
  assign n4259 = ~n4256 & ~n4257 ;
  assign n4260 = ~n4258 & ~n4259 ;
  assign n4261 = n4249 & ~n4260 ;
  assign n4262 = n4249 & ~n4261 ;
  assign n4263 = ~n4260 & ~n4261 ;
  assign n4264 = ~n4262 & ~n4263 ;
  assign n4265 = ~n3945 & ~n3950 ;
  assign n4266 = n4264 & n4265 ;
  assign n4267 = ~n4264 & ~n4265 ;
  assign n4268 = ~n4266 & ~n4267 ;
  assign n4269 = x82 & n574 ;
  assign n4270 = x80 & n673 ;
  assign n4271 = x81 & n569 ;
  assign n4272 = ~n4270 & ~n4271 ;
  assign n4273 = ~n4269 & n4272 ;
  assign n4274 = n577 & n2584 ;
  assign n4275 = n4273 & ~n4274 ;
  assign n4276 = x8 & ~n4275 ;
  assign n4277 = x8 & ~n4276 ;
  assign n4278 = ~n4275 & ~n4276 ;
  assign n4279 = ~n4277 & ~n4278 ;
  assign n4280 = ~n4268 & n4279 ;
  assign n4281 = n4268 & ~n4279 ;
  assign n4282 = ~n4280 & ~n4281 ;
  assign n4283 = ~n4174 & n4282 ;
  assign n4284 = n4174 & ~n4282 ;
  assign n4285 = ~n4283 & ~n4284 ;
  assign n4286 = ~n4173 & n4285 ;
  assign n4287 = ~n4173 & ~n4286 ;
  assign n4288 = n4285 & ~n4286 ;
  assign n4289 = ~n4287 & ~n4288 ;
  assign n4290 = ~n4162 & ~n4289 ;
  assign n4291 = ~n4162 & ~n4290 ;
  assign n4292 = ~n4289 & ~n4290 ;
  assign n4293 = ~n4291 & ~n4292 ;
  assign n4294 = x88 & n146 ;
  assign n4295 = x86 & n182 ;
  assign n4296 = x87 & n141 ;
  assign n4297 = ~n4295 & ~n4296 ;
  assign n4298 = ~n4294 & n4297 ;
  assign n4299 = ~n3987 & ~n3989 ;
  assign n4300 = ~x87 & ~x88 ;
  assign n4301 = x87 & x88 ;
  assign n4302 = ~n4300 & ~n4301 ;
  assign n4303 = ~n4299 & n4302 ;
  assign n4304 = n4299 & ~n4302 ;
  assign n4305 = ~n4303 & ~n4304 ;
  assign n4306 = n149 & n4305 ;
  assign n4307 = n4298 & ~n4306 ;
  assign n4308 = x2 & ~n4307 ;
  assign n4309 = x2 & ~n4308 ;
  assign n4310 = ~n4307 & ~n4308 ;
  assign n4311 = ~n4309 & ~n4310 ;
  assign n4312 = ~n4293 & ~n4311 ;
  assign n4313 = ~n4293 & ~n4312 ;
  assign n4314 = ~n4311 & ~n4312 ;
  assign n4315 = ~n4313 & ~n4314 ;
  assign n4316 = ~n3998 & ~n4003 ;
  assign n4317 = ~n4315 & ~n4316 ;
  assign n4318 = n4315 & n4316 ;
  assign n4319 = ~n4317 & ~n4318 ;
  assign n4473 = n4319 & x152 ;
  assign n4320 = ~n4127 & ~n4133 ;
  assign n4321 = ~x85 & n293 ;
  assign n4322 = ~x83 & n373 ;
  assign n4323 = ~x84 & n288 ;
  assign n4324 = ~n4322 & ~n4323 ;
  assign n4325 = ~n4321 & n4324 ;
  assign n4326 = n296 & n3521 ;
  assign n4327 = n4325 & ~n4326 ;
  assign n4328 = ~x5 & ~n4327 ;
  assign n4329 = ~x5 & ~n4328 ;
  assign n4330 = ~n4327 & ~n4328 ;
  assign n4331 = ~n4329 & ~n4330 ;
  assign n4332 = ~n4108 & ~n4112 ;
  assign n4333 = ~n4084 & ~n4086 ;
  assign n4334 = ~x76 & n1434 ;
  assign n4335 = ~x74 & n1646 ;
  assign n4336 = ~x75 & n1429 ;
  assign n4337 = ~n4335 & ~n4336 ;
  assign n4338 = ~n4334 & n4337 ;
  assign n4339 = n1390 & n1437 ;
  assign n4340 = n4338 & ~n4339 ;
  assign n4341 = ~x14 & ~n4340 ;
  assign n4342 = ~x14 & ~n4341 ;
  assign n4343 = ~n4340 & ~n4341 ;
  assign n4344 = ~n4342 & ~n4343 ;
  assign n4345 = ~n4078 & ~n4080 ;
  assign n4346 = ~x64 & ~n4190 ;
  assign n4347 = ~n4045 & n4346 ;
  assign n4348 = n4045 & ~n4346 ;
  assign n4349 = ~n4347 & ~n4348 ;
  assign n4350 = ~x67 & n3589 ;
  assign n4351 = ~x65 & n3878 ;
  assign n4352 = ~x66 & n3584 ;
  assign n4353 = ~n4351 & ~n4352 ;
  assign n4354 = ~n4350 & n4353 ;
  assign n4355 = n266 & n3592 ;
  assign n4356 = n4354 & ~n4355 ;
  assign n4357 = ~x23 & ~n4356 ;
  assign n4358 = ~x23 & ~n4357 ;
  assign n4359 = ~n4356 & ~n4357 ;
  assign n4360 = ~n4358 & ~n4359 ;
  assign n4361 = ~n4349 & ~n4360 ;
  assign n4362 = n4349 & n4360 ;
  assign n4363 = ~n4361 & ~n4362 ;
  assign n4364 = ~x70 & n2751 ;
  assign n4365 = ~x68 & n3020 ;
  assign n4366 = ~x69 & n2746 ;
  assign n4367 = ~n4365 & ~n4366 ;
  assign n4368 = ~n4364 & n4367 ;
  assign n4369 = n529 & n2754 ;
  assign n4370 = n4368 & ~n4369 ;
  assign n4371 = ~x20 & ~n4370 ;
  assign n4372 = ~x20 & ~n4371 ;
  assign n4373 = ~n4370 & ~n4371 ;
  assign n4374 = ~n4372 & ~n4373 ;
  assign n4375 = n4363 & ~n4374 ;
  assign n4376 = n4363 & ~n4375 ;
  assign n4377 = ~n4374 & ~n4375 ;
  assign n4378 = ~n4376 & ~n4377 ;
  assign n4379 = ~n4063 & n4378 ;
  assign n4380 = n4063 & ~n4378 ;
  assign n4381 = ~n4379 & ~n4380 ;
  assign n4382 = ~x73 & n2093 ;
  assign n4383 = ~x71 & n2275 ;
  assign n4384 = ~x72 & n2088 ;
  assign n4385 = ~n4383 & ~n4384 ;
  assign n4386 = ~n4382 & n4385 ;
  assign n4387 = n903 & n2096 ;
  assign n4388 = n4386 & ~n4387 ;
  assign n4389 = ~x17 & ~n4388 ;
  assign n4390 = ~x17 & ~n4389 ;
  assign n4391 = ~n4388 & ~n4389 ;
  assign n4392 = ~n4390 & ~n4391 ;
  assign n4393 = ~n4381 & ~n4392 ;
  assign n4394 = n4381 & n4392 ;
  assign n4395 = ~n4393 & ~n4394 ;
  assign n4396 = ~n4345 & n4395 ;
  assign n4397 = n4345 & ~n4395 ;
  assign n4398 = ~n4396 & ~n4397 ;
  assign n4399 = n4344 & ~n4398 ;
  assign n4400 = ~n4344 & n4398 ;
  assign n4401 = ~n4399 & ~n4400 ;
  assign n4402 = ~n4333 & n4401 ;
  assign n4403 = n4333 & ~n4401 ;
  assign n4404 = ~n4402 & ~n4403 ;
  assign n4405 = ~x79 & n945 ;
  assign n4406 = ~x77 & n1099 ;
  assign n4407 = ~x78 & n940 ;
  assign n4408 = ~n4406 & ~n4407 ;
  assign n4409 = ~n4405 & n4408 ;
  assign n4410 = n948 & n1921 ;
  assign n4411 = n4409 & ~n4410 ;
  assign n4412 = ~x11 & ~n4411 ;
  assign n4413 = ~x11 & ~n4412 ;
  assign n4414 = ~n4411 & ~n4412 ;
  assign n4415 = ~n4413 & ~n4414 ;
  assign n4416 = n4404 & ~n4415 ;
  assign n4417 = n4404 & ~n4416 ;
  assign n4418 = ~n4415 & ~n4416 ;
  assign n4419 = ~n4417 & ~n4418 ;
  assign n4420 = ~n4100 & ~n4105 ;
  assign n4421 = n4419 & n4420 ;
  assign n4422 = ~n4419 & ~n4420 ;
  assign n4423 = ~n4421 & ~n4422 ;
  assign n4424 = ~x82 & n574 ;
  assign n4425 = ~x80 & n673 ;
  assign n4426 = ~x81 & n569 ;
  assign n4427 = ~n4425 & ~n4426 ;
  assign n4428 = ~n4424 & n4427 ;
  assign n4429 = n577 & n2697 ;
  assign n4430 = n4428 & ~n4429 ;
  assign n4431 = ~x8 & ~n4430 ;
  assign n4432 = ~x8 & ~n4431 ;
  assign n4433 = ~n4430 & ~n4431 ;
  assign n4434 = ~n4432 & ~n4433 ;
  assign n4435 = ~n4423 & n4434 ;
  assign n4436 = n4423 & ~n4434 ;
  assign n4437 = ~n4435 & ~n4436 ;
  assign n4438 = ~n4332 & n4437 ;
  assign n4439 = n4332 & ~n4437 ;
  assign n4440 = ~n4438 & ~n4439 ;
  assign n4441 = ~n4331 & n4440 ;
  assign n4442 = ~n4331 & ~n4441 ;
  assign n4443 = n4440 & ~n4441 ;
  assign n4444 = ~n4442 & ~n4443 ;
  assign n4445 = ~n4320 & ~n4444 ;
  assign n4446 = ~n4320 & ~n4445 ;
  assign n4447 = ~n4444 & ~n4445 ;
  assign n4448 = ~n4446 & ~n4447 ;
  assign n4449 = ~x88 & n164 ;
  assign n4450 = ~x86 & n205 ;
  assign n4451 = ~x87 & n162 ;
  assign n4452 = ~n4450 & ~n4451 ;
  assign n4453 = ~n4449 & n4452 ;
  assign n4454 = ~n3986 & ~n4141 ;
  assign n4455 = n4302 & ~n4454 ;
  assign n4456 = ~n4302 & n4454 ;
  assign n4457 = ~n4455 & ~n4456 ;
  assign n4458 = n167 & n4457 ;
  assign n4459 = n4453 & ~n4458 ;
  assign n4460 = ~x2 & ~n4459 ;
  assign n4461 = ~x2 & ~n4460 ;
  assign n4462 = ~n4459 & ~n4460 ;
  assign n4463 = ~n4461 & ~n4462 ;
  assign n4464 = ~n4448 & ~n4463 ;
  assign n4465 = ~n4448 & ~n4464 ;
  assign n4466 = ~n4463 & ~n4464 ;
  assign n4467 = ~n4465 & ~n4466 ;
  assign n4468 = ~n4150 & ~n4155 ;
  assign n4469 = ~n4467 & ~n4468 ;
  assign n4470 = n4467 & n4468 ;
  assign n4471 = ~n4469 & ~n4470 ;
  assign n4474 = ~n4471 & ~x152 ;
  assign n4475 = ~n4473 & ~n4474 ;
  assign n4476 = ~n4312 & ~n4317 ;
  assign n4477 = x89 & n146 ;
  assign n4478 = x87 & n182 ;
  assign n4479 = x88 & n141 ;
  assign n4480 = ~n4478 & ~n4479 ;
  assign n4481 = ~n4477 & n4480 ;
  assign n4482 = ~n4301 & ~n4303 ;
  assign n4483 = ~x88 & ~x89 ;
  assign n4484 = x88 & x89 ;
  assign n4485 = ~n4483 & ~n4484 ;
  assign n4486 = ~n4482 & n4485 ;
  assign n4487 = n4482 & ~n4485 ;
  assign n4488 = ~n4486 & ~n4487 ;
  assign n4489 = n149 & n4488 ;
  assign n4490 = n4481 & ~n4489 ;
  assign n4491 = x2 & ~n4490 ;
  assign n4492 = x2 & ~n4491 ;
  assign n4493 = ~n4490 & ~n4491 ;
  assign n4494 = ~n4492 & ~n4493 ;
  assign n4495 = ~n4286 & ~n4290 ;
  assign n4496 = ~n3908 & ~n4223 ;
  assign n4497 = ~n4220 & ~n4496 ;
  assign n4498 = x71 & n2751 ;
  assign n4499 = x69 & n3020 ;
  assign n4500 = x70 & n2746 ;
  assign n4501 = ~n4499 & ~n4500 ;
  assign n4502 = ~n4498 & n4501 ;
  assign n4503 = n558 & n2754 ;
  assign n4504 = n4502 & ~n4503 ;
  assign n4505 = x20 & ~n4504 ;
  assign n4506 = x20 & ~n4505 ;
  assign n4507 = ~n4504 & ~n4505 ;
  assign n4508 = ~n4506 & ~n4507 ;
  assign n4509 = n3890 & n4191 ;
  assign n4510 = ~n4206 & ~n4509 ;
  assign n4511 = x68 & n3589 ;
  assign n4512 = x66 & n3878 ;
  assign n4513 = x67 & n3584 ;
  assign n4514 = ~n4512 & ~n4513 ;
  assign n4515 = ~n4511 & n4514 ;
  assign n4516 = n317 & n3592 ;
  assign n4517 = n4515 & ~n4516 ;
  assign n4518 = x23 & ~n4517 ;
  assign n4519 = x23 & ~n4518 ;
  assign n4520 = ~n4517 & ~n4518 ;
  assign n4521 = ~n4519 & ~n4520 ;
  assign n4522 = x26 & ~n4191 ;
  assign n4523 = ~x24 & x25 ;
  assign n4524 = x24 & ~x25 ;
  assign n4525 = ~n4523 & ~n4524 ;
  assign n4526 = n4190 & ~n4525 ;
  assign n4527 = x64 & n4526 ;
  assign n4528 = ~x25 & x26 ;
  assign n4529 = x25 & ~x26 ;
  assign n4530 = ~n4528 & ~n4529 ;
  assign n4531 = ~n4190 & n4530 ;
  assign n4532 = x65 & n4531 ;
  assign n4533 = ~n4527 & ~n4532 ;
  assign n4534 = ~n4190 & ~n4530 ;
  assign n4535 = ~n152 & n4534 ;
  assign n4536 = n4533 & ~n4535 ;
  assign n4537 = x26 & ~n4536 ;
  assign n4538 = x26 & ~n4537 ;
  assign n4539 = ~n4536 & ~n4537 ;
  assign n4540 = ~n4538 & ~n4539 ;
  assign n4541 = n4522 & ~n4540 ;
  assign n4542 = ~n4522 & n4540 ;
  assign n4543 = ~n4541 & ~n4542 ;
  assign n4544 = n4521 & n4543 ;
  assign n4545 = ~n4521 & ~n4543 ;
  assign n4546 = ~n4544 & ~n4545 ;
  assign n4547 = ~n4510 & ~n4546 ;
  assign n4548 = n4510 & n4546 ;
  assign n4549 = ~n4547 & ~n4548 ;
  assign n4550 = ~n4508 & n4549 ;
  assign n4551 = n4508 & ~n4549 ;
  assign n4552 = ~n4550 & ~n4551 ;
  assign n4553 = ~n4497 & n4552 ;
  assign n4554 = n4497 & ~n4552 ;
  assign n4555 = ~n4553 & ~n4554 ;
  assign n4556 = x74 & n2093 ;
  assign n4557 = x72 & n2275 ;
  assign n4558 = x73 & n2088 ;
  assign n4559 = ~n4557 & ~n4558 ;
  assign n4560 = ~n4556 & n4559 ;
  assign n4561 = n994 & n2096 ;
  assign n4562 = n4560 & ~n4561 ;
  assign n4563 = x17 & ~n4562 ;
  assign n4564 = x17 & ~n4563 ;
  assign n4565 = ~n4562 & ~n4563 ;
  assign n4566 = ~n4564 & ~n4565 ;
  assign n4567 = n4555 & ~n4566 ;
  assign n4568 = n4555 & ~n4567 ;
  assign n4569 = ~n4566 & ~n4567 ;
  assign n4570 = ~n4568 & ~n4569 ;
  assign n4571 = ~n4238 & ~n4241 ;
  assign n4572 = n4570 & n4571 ;
  assign n4573 = ~n4570 & ~n4571 ;
  assign n4574 = ~n4572 & ~n4573 ;
  assign n4575 = x77 & n1434 ;
  assign n4576 = x75 & n1646 ;
  assign n4577 = x76 & n1429 ;
  assign n4578 = ~n4576 & ~n4577 ;
  assign n4579 = ~n4575 & n4578 ;
  assign n4580 = n1437 & n1502 ;
  assign n4581 = n4579 & ~n4580 ;
  assign n4582 = x14 & ~n4581 ;
  assign n4583 = x14 & ~n4582 ;
  assign n4584 = ~n4581 & ~n4582 ;
  assign n4585 = ~n4583 & ~n4584 ;
  assign n4586 = ~n4574 & n4585 ;
  assign n4587 = n4574 & ~n4585 ;
  assign n4588 = ~n4586 & ~n4587 ;
  assign n4589 = ~n4245 & ~n4247 ;
  assign n4590 = n4588 & ~n4589 ;
  assign n4591 = ~n4588 & n4589 ;
  assign n4592 = ~n4590 & ~n4591 ;
  assign n4593 = x80 & n945 ;
  assign n4594 = x78 & n1099 ;
  assign n4595 = x79 & n940 ;
  assign n4596 = ~n4594 & ~n4595 ;
  assign n4597 = ~n4593 & n4596 ;
  assign n4598 = n948 & n2028 ;
  assign n4599 = n4597 & ~n4598 ;
  assign n4600 = x11 & ~n4599 ;
  assign n4601 = x11 & ~n4600 ;
  assign n4602 = ~n4599 & ~n4600 ;
  assign n4603 = ~n4601 & ~n4602 ;
  assign n4604 = n4592 & ~n4603 ;
  assign n4605 = n4592 & ~n4604 ;
  assign n4606 = ~n4603 & ~n4604 ;
  assign n4607 = ~n4605 & ~n4606 ;
  assign n4608 = ~n4261 & ~n4267 ;
  assign n4609 = n4607 & n4608 ;
  assign n4610 = ~n4607 & ~n4608 ;
  assign n4611 = ~n4609 & ~n4610 ;
  assign n4612 = x83 & n574 ;
  assign n4613 = x81 & n673 ;
  assign n4614 = x82 & n569 ;
  assign n4615 = ~n4613 & ~n4614 ;
  assign n4616 = ~n4612 & n4615 ;
  assign n4617 = n577 & n2843 ;
  assign n4618 = n4616 & ~n4617 ;
  assign n4619 = x8 & ~n4618 ;
  assign n4620 = x8 & ~n4619 ;
  assign n4621 = ~n4618 & ~n4619 ;
  assign n4622 = ~n4620 & ~n4621 ;
  assign n4623 = n4611 & ~n4622 ;
  assign n4624 = n4611 & ~n4623 ;
  assign n4625 = ~n4622 & ~n4623 ;
  assign n4626 = ~n4624 & ~n4625 ;
  assign n4627 = ~n4281 & ~n4283 ;
  assign n4628 = ~n4626 & ~n4627 ;
  assign n4629 = ~n4626 & ~n4628 ;
  assign n4630 = ~n4627 & ~n4628 ;
  assign n4631 = ~n4629 & ~n4630 ;
  assign n4632 = x86 & n293 ;
  assign n4633 = x84 & n373 ;
  assign n4634 = x85 & n288 ;
  assign n4635 = ~n4633 & ~n4634 ;
  assign n4636 = ~n4632 & n4635 ;
  assign n4637 = n296 & n3686 ;
  assign n4638 = n4636 & ~n4637 ;
  assign n4639 = x5 & ~n4638 ;
  assign n4640 = x5 & ~n4639 ;
  assign n4641 = ~n4638 & ~n4639 ;
  assign n4642 = ~n4640 & ~n4641 ;
  assign n4643 = ~n4631 & n4642 ;
  assign n4644 = n4631 & ~n4642 ;
  assign n4645 = ~n4643 & ~n4644 ;
  assign n4646 = ~n4495 & ~n4645 ;
  assign n4647 = n4495 & n4645 ;
  assign n4648 = ~n4646 & ~n4647 ;
  assign n4649 = ~n4494 & n4648 ;
  assign n4650 = n4494 & ~n4648 ;
  assign n4651 = ~n4649 & ~n4650 ;
  assign n4652 = ~n4476 & n4651 ;
  assign n4653 = n4476 & ~n4651 ;
  assign n4654 = ~n4652 & ~n4653 ;
  assign n4822 = n4654 & x153 ;
  assign n4655 = ~n4464 & ~n4469 ;
  assign n4656 = ~x89 & n164 ;
  assign n4657 = ~x87 & n205 ;
  assign n4658 = ~x88 & n162 ;
  assign n4659 = ~n4657 & ~n4658 ;
  assign n4660 = ~n4656 & n4659 ;
  assign n4661 = ~n4300 & ~n4455 ;
  assign n4662 = n4485 & ~n4661 ;
  assign n4663 = ~n4485 & n4661 ;
  assign n4664 = ~n4662 & ~n4663 ;
  assign n4665 = n167 & n4664 ;
  assign n4666 = n4660 & ~n4665 ;
  assign n4667 = ~x2 & ~n4666 ;
  assign n4668 = ~x2 & ~n4667 ;
  assign n4669 = ~n4666 & ~n4667 ;
  assign n4670 = ~n4668 & ~n4669 ;
  assign n4671 = ~n4441 & ~n4445 ;
  assign n4672 = ~n4063 & ~n4378 ;
  assign n4673 = ~n4375 & ~n4672 ;
  assign n4674 = ~x71 & n2751 ;
  assign n4675 = ~x69 & n3020 ;
  assign n4676 = ~x70 & n2746 ;
  assign n4677 = ~n4675 & ~n4676 ;
  assign n4678 = ~n4674 & n4677 ;
  assign n4679 = n622 & n2754 ;
  assign n4680 = n4678 & ~n4679 ;
  assign n4681 = ~x20 & ~n4680 ;
  assign n4682 = ~x20 & ~n4681 ;
  assign n4683 = ~n4680 & ~n4681 ;
  assign n4684 = ~n4682 & ~n4683 ;
  assign n4685 = n4045 & n4346 ;
  assign n4686 = ~n4361 & ~n4685 ;
  assign n4687 = ~x68 & n3589 ;
  assign n4688 = ~x66 & n3878 ;
  assign n4689 = ~x67 & n3584 ;
  assign n4690 = ~n4688 & ~n4689 ;
  assign n4691 = ~n4687 & n4690 ;
  assign n4692 = n352 & n3592 ;
  assign n4693 = n4691 & ~n4692 ;
  assign n4694 = ~x23 & ~n4693 ;
  assign n4695 = ~x23 & ~n4694 ;
  assign n4696 = ~n4693 & ~n4694 ;
  assign n4697 = ~n4695 & ~n4696 ;
  assign n4698 = ~x26 & ~n4346 ;
  assign n4699 = ~x64 & n4526 ;
  assign n4700 = ~x65 & n4531 ;
  assign n4701 = ~n4699 & ~n4700 ;
  assign n4702 = ~n4535 & n4701 ;
  assign n4703 = ~x26 & ~n4702 ;
  assign n4704 = ~x26 & ~n4703 ;
  assign n4705 = ~n4702 & ~n4703 ;
  assign n4706 = ~n4704 & ~n4705 ;
  assign n4707 = n4698 & ~n4706 ;
  assign n4708 = ~n4698 & n4706 ;
  assign n4709 = ~n4707 & ~n4708 ;
  assign n4710 = n4697 & n4709 ;
  assign n4711 = ~n4697 & ~n4709 ;
  assign n4712 = ~n4710 & ~n4711 ;
  assign n4713 = ~n4686 & ~n4712 ;
  assign n4714 = n4686 & n4712 ;
  assign n4715 = ~n4713 & ~n4714 ;
  assign n4716 = ~n4684 & n4715 ;
  assign n4717 = n4684 & ~n4715 ;
  assign n4718 = ~n4716 & ~n4717 ;
  assign n4719 = ~n4673 & n4718 ;
  assign n4720 = n4673 & ~n4718 ;
  assign n4721 = ~n4719 & ~n4720 ;
  assign n4722 = ~x74 & n2093 ;
  assign n4723 = ~x72 & n2275 ;
  assign n4724 = ~x73 & n2088 ;
  assign n4725 = ~n4723 & ~n4724 ;
  assign n4726 = ~n4722 & n4725 ;
  assign n4727 = n1066 & n2096 ;
  assign n4728 = n4726 & ~n4727 ;
  assign n4729 = ~x17 & ~n4728 ;
  assign n4730 = ~x17 & ~n4729 ;
  assign n4731 = ~n4728 & ~n4729 ;
  assign n4732 = ~n4730 & ~n4731 ;
  assign n4733 = n4721 & ~n4732 ;
  assign n4734 = n4721 & ~n4733 ;
  assign n4735 = ~n4732 & ~n4733 ;
  assign n4736 = ~n4734 & ~n4735 ;
  assign n4737 = ~n4393 & ~n4396 ;
  assign n4738 = n4736 & n4737 ;
  assign n4739 = ~n4736 & ~n4737 ;
  assign n4740 = ~n4738 & ~n4739 ;
  assign n4741 = ~x77 & n1434 ;
  assign n4742 = ~x75 & n1646 ;
  assign n4743 = ~x76 & n1429 ;
  assign n4744 = ~n4742 & ~n4743 ;
  assign n4745 = ~n4741 & n4744 ;
  assign n4746 = n1437 & n1594 ;
  assign n4747 = n4745 & ~n4746 ;
  assign n4748 = ~x14 & ~n4747 ;
  assign n4749 = ~x14 & ~n4748 ;
  assign n4750 = ~n4747 & ~n4748 ;
  assign n4751 = ~n4749 & ~n4750 ;
  assign n4752 = ~n4740 & n4751 ;
  assign n4753 = n4740 & ~n4751 ;
  assign n4754 = ~n4752 & ~n4753 ;
  assign n4755 = ~n4400 & ~n4402 ;
  assign n4756 = n4754 & ~n4755 ;
  assign n4757 = ~n4754 & n4755 ;
  assign n4758 = ~n4756 & ~n4757 ;
  assign n4759 = ~x80 & n945 ;
  assign n4760 = ~x78 & n1099 ;
  assign n4761 = ~x79 & n940 ;
  assign n4762 = ~n4760 & ~n4761 ;
  assign n4763 = ~n4759 & n4762 ;
  assign n4764 = n948 & n2145 ;
  assign n4765 = n4763 & ~n4764 ;
  assign n4766 = ~x11 & ~n4765 ;
  assign n4767 = ~x11 & ~n4766 ;
  assign n4768 = ~n4765 & ~n4766 ;
  assign n4769 = ~n4767 & ~n4768 ;
  assign n4770 = n4758 & ~n4769 ;
  assign n4771 = n4758 & ~n4770 ;
  assign n4772 = ~n4769 & ~n4770 ;
  assign n4773 = ~n4771 & ~n4772 ;
  assign n4774 = ~n4416 & ~n4422 ;
  assign n4775 = n4773 & n4774 ;
  assign n4776 = ~n4773 & ~n4774 ;
  assign n4777 = ~n4775 & ~n4776 ;
  assign n4778 = ~x83 & n574 ;
  assign n4779 = ~x81 & n673 ;
  assign n4780 = ~x82 & n569 ;
  assign n4781 = ~n4779 & ~n4780 ;
  assign n4782 = ~n4778 & n4781 ;
  assign n4783 = n577 & n2972 ;
  assign n4784 = n4782 & ~n4783 ;
  assign n4785 = ~x8 & ~n4784 ;
  assign n4786 = ~x8 & ~n4785 ;
  assign n4787 = ~n4784 & ~n4785 ;
  assign n4788 = ~n4786 & ~n4787 ;
  assign n4789 = n4777 & ~n4788 ;
  assign n4790 = n4777 & ~n4789 ;
  assign n4791 = ~n4788 & ~n4789 ;
  assign n4792 = ~n4790 & ~n4791 ;
  assign n4793 = ~n4436 & ~n4438 ;
  assign n4794 = ~n4792 & ~n4793 ;
  assign n4795 = ~n4792 & ~n4794 ;
  assign n4796 = ~n4793 & ~n4794 ;
  assign n4797 = ~n4795 & ~n4796 ;
  assign n4798 = ~x86 & n293 ;
  assign n4799 = ~x84 & n373 ;
  assign n4800 = ~x85 & n288 ;
  assign n4801 = ~n4799 & ~n4800 ;
  assign n4802 = ~n4798 & n4801 ;
  assign n4803 = n296 & n3832 ;
  assign n4804 = n4802 & ~n4803 ;
  assign n4805 = ~x5 & ~n4804 ;
  assign n4806 = ~x5 & ~n4805 ;
  assign n4807 = ~n4804 & ~n4805 ;
  assign n4808 = ~n4806 & ~n4807 ;
  assign n4809 = ~n4797 & n4808 ;
  assign n4810 = n4797 & ~n4808 ;
  assign n4811 = ~n4809 & ~n4810 ;
  assign n4812 = ~n4671 & ~n4811 ;
  assign n4813 = n4671 & n4811 ;
  assign n4814 = ~n4812 & ~n4813 ;
  assign n4815 = ~n4670 & n4814 ;
  assign n4816 = n4670 & ~n4814 ;
  assign n4817 = ~n4815 & ~n4816 ;
  assign n4818 = ~n4655 & n4817 ;
  assign n4819 = n4655 & ~n4817 ;
  assign n4820 = ~n4818 & ~n4819 ;
  assign n4823 = ~n4820 & ~x153 ;
  assign n4824 = ~n4822 & ~n4823 ;
  assign n4825 = ~n4649 & ~n4652 ;
  assign n4826 = ~n4631 & ~n4642 ;
  assign n4827 = ~n4646 & ~n4826 ;
  assign n4828 = ~n4604 & ~n4610 ;
  assign n4829 = ~n4587 & ~n4590 ;
  assign n4830 = ~n4567 & ~n4573 ;
  assign n4831 = x75 & n2093 ;
  assign n4832 = x73 & n2275 ;
  assign n4833 = x74 & n2088 ;
  assign n4834 = ~n4832 & ~n4833 ;
  assign n4835 = ~n4831 & n4834 ;
  assign n4836 = n1150 & n2096 ;
  assign n4837 = n4835 & ~n4836 ;
  assign n4838 = x17 & ~n4837 ;
  assign n4839 = x17 & ~n4838 ;
  assign n4840 = ~n4837 & ~n4838 ;
  assign n4841 = ~n4839 & ~n4840 ;
  assign n4842 = ~n4550 & ~n4553 ;
  assign n4843 = ~n4521 & n4543 ;
  assign n4844 = ~n4547 & ~n4843 ;
  assign n4845 = x66 & n4531 ;
  assign n4846 = n4190 & ~n4530 ;
  assign n4847 = n4525 & n4846 ;
  assign n4848 = x64 & n4847 ;
  assign n4849 = x65 & n4526 ;
  assign n4850 = ~n4848 & ~n4849 ;
  assign n4851 = ~n4845 & n4850 ;
  assign n4852 = n194 & n4534 ;
  assign n4853 = n4851 & ~n4852 ;
  assign n4854 = x26 & ~n4853 ;
  assign n4855 = x26 & ~n4854 ;
  assign n4856 = ~n4853 & ~n4854 ;
  assign n4857 = ~n4855 & ~n4856 ;
  assign n4858 = ~n4541 & n4857 ;
  assign n4859 = n4541 & ~n4857 ;
  assign n4860 = ~n4858 & ~n4859 ;
  assign n4861 = x69 & n3589 ;
  assign n4862 = x67 & n3878 ;
  assign n4863 = x68 & n3584 ;
  assign n4864 = ~n4862 & ~n4863 ;
  assign n4865 = ~n4861 & n4864 ;
  assign n4866 = n398 & n3592 ;
  assign n4867 = n4865 & ~n4866 ;
  assign n4868 = x23 & ~n4867 ;
  assign n4869 = x23 & ~n4868 ;
  assign n4870 = ~n4867 & ~n4868 ;
  assign n4871 = ~n4869 & ~n4870 ;
  assign n4872 = n4860 & ~n4871 ;
  assign n4873 = ~n4860 & n4871 ;
  assign n4874 = ~n4844 & ~n4873 ;
  assign n4875 = ~n4872 & n4874 ;
  assign n4876 = ~n4844 & ~n4875 ;
  assign n4877 = ~n4872 & ~n4875 ;
  assign n4878 = ~n4873 & n4877 ;
  assign n4879 = ~n4876 & ~n4878 ;
  assign n4880 = x72 & n2751 ;
  assign n4881 = x70 & n3020 ;
  assign n4882 = x71 & n2746 ;
  assign n4883 = ~n4881 & ~n4882 ;
  assign n4884 = ~n4880 & n4883 ;
  assign n4885 = n717 & n2754 ;
  assign n4886 = n4884 & ~n4885 ;
  assign n4887 = x20 & ~n4886 ;
  assign n4888 = x20 & ~n4887 ;
  assign n4889 = ~n4886 & ~n4887 ;
  assign n4890 = ~n4888 & ~n4889 ;
  assign n4891 = n4879 & n4890 ;
  assign n4892 = ~n4879 & ~n4890 ;
  assign n4893 = ~n4891 & ~n4892 ;
  assign n4894 = ~n4842 & n4893 ;
  assign n4895 = n4842 & ~n4893 ;
  assign n4896 = ~n4894 & ~n4895 ;
  assign n4897 = n4841 & ~n4896 ;
  assign n4898 = ~n4841 & n4896 ;
  assign n4899 = ~n4897 & ~n4898 ;
  assign n4900 = ~n4830 & n4899 ;
  assign n4901 = n4830 & ~n4899 ;
  assign n4902 = ~n4900 & ~n4901 ;
  assign n4903 = x78 & n1434 ;
  assign n4904 = x76 & n1646 ;
  assign n4905 = x77 & n1429 ;
  assign n4906 = ~n4904 & ~n4905 ;
  assign n4907 = ~n4903 & n4906 ;
  assign n4908 = n1437 & n1624 ;
  assign n4909 = n4907 & ~n4908 ;
  assign n4910 = x14 & ~n4909 ;
  assign n4911 = x14 & ~n4910 ;
  assign n4912 = ~n4909 & ~n4910 ;
  assign n4913 = ~n4911 & ~n4912 ;
  assign n4914 = n4902 & ~n4913 ;
  assign n4915 = n4902 & ~n4914 ;
  assign n4916 = ~n4913 & ~n4914 ;
  assign n4917 = ~n4915 & ~n4916 ;
  assign n4918 = ~n4829 & n4917 ;
  assign n4919 = n4829 & ~n4917 ;
  assign n4920 = ~n4918 & ~n4919 ;
  assign n4921 = x81 & n945 ;
  assign n4922 = x79 & n1099 ;
  assign n4923 = x80 & n940 ;
  assign n4924 = ~n4922 & ~n4923 ;
  assign n4925 = ~n4921 & n4924 ;
  assign n4926 = n948 & n2348 ;
  assign n4927 = n4925 & ~n4926 ;
  assign n4928 = x11 & ~n4927 ;
  assign n4929 = x11 & ~n4928 ;
  assign n4930 = ~n4927 & ~n4928 ;
  assign n4931 = ~n4929 & ~n4930 ;
  assign n4932 = ~n4920 & ~n4931 ;
  assign n4933 = n4920 & n4931 ;
  assign n4934 = ~n4932 & ~n4933 ;
  assign n4935 = n4828 & ~n4934 ;
  assign n4936 = ~n4828 & n4934 ;
  assign n4937 = ~n4935 & ~n4936 ;
  assign n4938 = x84 & n574 ;
  assign n4939 = x82 & n673 ;
  assign n4940 = x83 & n569 ;
  assign n4941 = ~n4939 & ~n4940 ;
  assign n4942 = ~n4938 & n4941 ;
  assign n4943 = n577 & n3114 ;
  assign n4944 = n4942 & ~n4943 ;
  assign n4945 = x8 & ~n4944 ;
  assign n4946 = x8 & ~n4945 ;
  assign n4947 = ~n4944 & ~n4945 ;
  assign n4948 = ~n4946 & ~n4947 ;
  assign n4949 = n4937 & ~n4948 ;
  assign n4950 = n4937 & ~n4949 ;
  assign n4951 = ~n4948 & ~n4949 ;
  assign n4952 = ~n4950 & ~n4951 ;
  assign n4953 = ~n4623 & ~n4628 ;
  assign n4954 = n4952 & n4953 ;
  assign n4955 = ~n4952 & ~n4953 ;
  assign n4956 = ~n4954 & ~n4955 ;
  assign n4957 = x87 & n293 ;
  assign n4958 = x85 & n373 ;
  assign n4959 = x86 & n288 ;
  assign n4960 = ~n4958 & ~n4959 ;
  assign n4961 = ~n4957 & n4960 ;
  assign n4962 = n296 & n3991 ;
  assign n4963 = n4961 & ~n4962 ;
  assign n4964 = x5 & ~n4963 ;
  assign n4965 = x5 & ~n4964 ;
  assign n4966 = ~n4963 & ~n4964 ;
  assign n4967 = ~n4965 & ~n4966 ;
  assign n4968 = n4956 & ~n4967 ;
  assign n4969 = n4956 & ~n4968 ;
  assign n4970 = ~n4967 & ~n4968 ;
  assign n4971 = ~n4969 & ~n4970 ;
  assign n4972 = ~n4827 & n4971 ;
  assign n4973 = n4827 & ~n4971 ;
  assign n4974 = ~n4972 & ~n4973 ;
  assign n4975 = x90 & n146 ;
  assign n4976 = x88 & n182 ;
  assign n4977 = x89 & n141 ;
  assign n4978 = ~n4976 & ~n4977 ;
  assign n4979 = ~n4975 & n4978 ;
  assign n4980 = ~n4484 & ~n4486 ;
  assign n4981 = ~x89 & ~x90 ;
  assign n4982 = x89 & x90 ;
  assign n4983 = ~n4981 & ~n4982 ;
  assign n4984 = ~n4980 & n4983 ;
  assign n4985 = n4980 & ~n4983 ;
  assign n4986 = ~n4984 & ~n4985 ;
  assign n4987 = n149 & n4986 ;
  assign n4988 = n4979 & ~n4987 ;
  assign n4989 = x2 & ~n4988 ;
  assign n4990 = x2 & ~n4989 ;
  assign n4991 = ~n4988 & ~n4989 ;
  assign n4992 = ~n4990 & ~n4991 ;
  assign n4993 = ~n4974 & ~n4992 ;
  assign n4994 = n4974 & n4992 ;
  assign n4995 = ~n4993 & ~n4994 ;
  assign n4996 = ~n4825 & n4995 ;
  assign n4997 = n4825 & ~n4995 ;
  assign n4998 = ~n4996 & ~n4997 ;
  assign n5169 = n4998 & x154 ;
  assign n4999 = ~n4815 & ~n4818 ;
  assign n5000 = ~n4797 & ~n4808 ;
  assign n5001 = ~n4812 & ~n5000 ;
  assign n5002 = ~n4770 & ~n4776 ;
  assign n5003 = ~n4753 & ~n4756 ;
  assign n5004 = ~n4733 & ~n4739 ;
  assign n5005 = ~x75 & n2093 ;
  assign n5006 = ~x73 & n2275 ;
  assign n5007 = ~x74 & n2088 ;
  assign n5008 = ~n5006 & ~n5007 ;
  assign n5009 = ~n5005 & n5008 ;
  assign n5010 = n1225 & n2096 ;
  assign n5011 = n5009 & ~n5010 ;
  assign n5012 = ~x17 & ~n5011 ;
  assign n5013 = ~x17 & ~n5012 ;
  assign n5014 = ~n5011 & ~n5012 ;
  assign n5015 = ~n5013 & ~n5014 ;
  assign n5016 = ~n4716 & ~n4719 ;
  assign n5017 = ~n4697 & n4709 ;
  assign n5018 = ~n4713 & ~n5017 ;
  assign n5019 = ~x66 & n4531 ;
  assign n5020 = ~x64 & n4847 ;
  assign n5021 = ~x65 & n4526 ;
  assign n5022 = ~n5020 & ~n5021 ;
  assign n5023 = ~n5019 & n5022 ;
  assign n5024 = n214 & n4534 ;
  assign n5025 = n5023 & ~n5024 ;
  assign n5026 = ~x26 & ~n5025 ;
  assign n5027 = ~x26 & ~n5026 ;
  assign n5028 = ~n5025 & ~n5026 ;
  assign n5029 = ~n5027 & ~n5028 ;
  assign n5030 = ~n4707 & n5029 ;
  assign n5031 = n4707 & ~n5029 ;
  assign n5032 = ~n5030 & ~n5031 ;
  assign n5033 = ~x69 & n3589 ;
  assign n5034 = ~x67 & n3878 ;
  assign n5035 = ~x68 & n3584 ;
  assign n5036 = ~n5034 & ~n5035 ;
  assign n5037 = ~n5033 & n5036 ;
  assign n5038 = n435 & n3592 ;
  assign n5039 = n5037 & ~n5038 ;
  assign n5040 = ~x23 & ~n5039 ;
  assign n5041 = ~x23 & ~n5040 ;
  assign n5042 = ~n5039 & ~n5040 ;
  assign n5043 = ~n5041 & ~n5042 ;
  assign n5044 = n5032 & ~n5043 ;
  assign n5045 = ~n5032 & n5043 ;
  assign n5046 = ~n5018 & ~n5045 ;
  assign n5047 = ~n5044 & n5046 ;
  assign n5048 = ~n5018 & ~n5047 ;
  assign n5049 = ~n5044 & ~n5047 ;
  assign n5050 = ~n5045 & n5049 ;
  assign n5051 = ~n5048 & ~n5050 ;
  assign n5052 = ~x72 & n2751 ;
  assign n5053 = ~x70 & n3020 ;
  assign n5054 = ~x71 & n2746 ;
  assign n5055 = ~n5053 & ~n5054 ;
  assign n5056 = ~n5052 & n5055 ;
  assign n5057 = n773 & n2754 ;
  assign n5058 = n5056 & ~n5057 ;
  assign n5059 = ~x20 & ~n5058 ;
  assign n5060 = ~x20 & ~n5059 ;
  assign n5061 = ~n5058 & ~n5059 ;
  assign n5062 = ~n5060 & ~n5061 ;
  assign n5063 = n5051 & n5062 ;
  assign n5064 = ~n5051 & ~n5062 ;
  assign n5065 = ~n5063 & ~n5064 ;
  assign n5066 = ~n5016 & n5065 ;
  assign n5067 = n5016 & ~n5065 ;
  assign n5068 = ~n5066 & ~n5067 ;
  assign n5069 = n5015 & ~n5068 ;
  assign n5070 = ~n5015 & n5068 ;
  assign n5071 = ~n5069 & ~n5070 ;
  assign n5072 = ~n5004 & n5071 ;
  assign n5073 = n5004 & ~n5071 ;
  assign n5074 = ~n5072 & ~n5073 ;
  assign n5075 = ~x78 & n1434 ;
  assign n5076 = ~x76 & n1646 ;
  assign n5077 = ~x77 & n1429 ;
  assign n5078 = ~n5076 & ~n5077 ;
  assign n5079 = ~n5075 & n5078 ;
  assign n5080 = n1437 & n1718 ;
  assign n5081 = n5079 & ~n5080 ;
  assign n5082 = ~x14 & ~n5081 ;
  assign n5083 = ~x14 & ~n5082 ;
  assign n5084 = ~n5081 & ~n5082 ;
  assign n5085 = ~n5083 & ~n5084 ;
  assign n5086 = n5074 & ~n5085 ;
  assign n5087 = n5074 & ~n5086 ;
  assign n5088 = ~n5085 & ~n5086 ;
  assign n5089 = ~n5087 & ~n5088 ;
  assign n5090 = ~n5003 & n5089 ;
  assign n5091 = n5003 & ~n5089 ;
  assign n5092 = ~n5090 & ~n5091 ;
  assign n5093 = ~x81 & n945 ;
  assign n5094 = ~x79 & n1099 ;
  assign n5095 = ~x80 & n940 ;
  assign n5096 = ~n5094 & ~n5095 ;
  assign n5097 = ~n5093 & n5096 ;
  assign n5098 = n948 & n2460 ;
  assign n5099 = n5097 & ~n5098 ;
  assign n5100 = ~x11 & ~n5099 ;
  assign n5101 = ~x11 & ~n5100 ;
  assign n5102 = ~n5099 & ~n5100 ;
  assign n5103 = ~n5101 & ~n5102 ;
  assign n5104 = ~n5092 & ~n5103 ;
  assign n5105 = n5092 & n5103 ;
  assign n5106 = ~n5104 & ~n5105 ;
  assign n5107 = n5002 & ~n5106 ;
  assign n5108 = ~n5002 & n5106 ;
  assign n5109 = ~n5107 & ~n5108 ;
  assign n5110 = ~x84 & n574 ;
  assign n5111 = ~x82 & n673 ;
  assign n5112 = ~x83 & n569 ;
  assign n5113 = ~n5111 & ~n5112 ;
  assign n5114 = ~n5110 & n5113 ;
  assign n5115 = n577 & n3247 ;
  assign n5116 = n5114 & ~n5115 ;
  assign n5117 = ~x8 & ~n5116 ;
  assign n5118 = ~x8 & ~n5117 ;
  assign n5119 = ~n5116 & ~n5117 ;
  assign n5120 = ~n5118 & ~n5119 ;
  assign n5121 = n5109 & ~n5120 ;
  assign n5122 = n5109 & ~n5121 ;
  assign n5123 = ~n5120 & ~n5121 ;
  assign n5124 = ~n5122 & ~n5123 ;
  assign n5125 = ~n4789 & ~n4794 ;
  assign n5126 = n5124 & n5125 ;
  assign n5127 = ~n5124 & ~n5125 ;
  assign n5128 = ~n5126 & ~n5127 ;
  assign n5129 = ~x87 & n293 ;
  assign n5130 = ~x85 & n373 ;
  assign n5131 = ~x86 & n288 ;
  assign n5132 = ~n5130 & ~n5131 ;
  assign n5133 = ~n5129 & n5132 ;
  assign n5134 = n296 & n4143 ;
  assign n5135 = n5133 & ~n5134 ;
  assign n5136 = ~x5 & ~n5135 ;
  assign n5137 = ~x5 & ~n5136 ;
  assign n5138 = ~n5135 & ~n5136 ;
  assign n5139 = ~n5137 & ~n5138 ;
  assign n5140 = n5128 & ~n5139 ;
  assign n5141 = n5128 & ~n5140 ;
  assign n5142 = ~n5139 & ~n5140 ;
  assign n5143 = ~n5141 & ~n5142 ;
  assign n5144 = ~n5001 & n5143 ;
  assign n5145 = n5001 & ~n5143 ;
  assign n5146 = ~n5144 & ~n5145 ;
  assign n5147 = ~x90 & n164 ;
  assign n5148 = ~x88 & n205 ;
  assign n5149 = ~x89 & n162 ;
  assign n5150 = ~n5148 & ~n5149 ;
  assign n5151 = ~n5147 & n5150 ;
  assign n5152 = ~n4483 & ~n4662 ;
  assign n5153 = n4983 & ~n5152 ;
  assign n5154 = ~n4983 & n5152 ;
  assign n5155 = ~n5153 & ~n5154 ;
  assign n5156 = n167 & n5155 ;
  assign n5157 = n5151 & ~n5156 ;
  assign n5158 = ~x2 & ~n5157 ;
  assign n5159 = ~x2 & ~n5158 ;
  assign n5160 = ~n5157 & ~n5158 ;
  assign n5161 = ~n5159 & ~n5160 ;
  assign n5162 = ~n5146 & ~n5161 ;
  assign n5163 = n5146 & n5161 ;
  assign n5164 = ~n5162 & ~n5163 ;
  assign n5165 = ~n4999 & n5164 ;
  assign n5166 = n4999 & ~n5164 ;
  assign n5167 = ~n5165 & ~n5166 ;
  assign n5170 = ~n5167 & ~x154 ;
  assign n5171 = ~n5169 & ~n5170 ;
  assign n5172 = ~n4993 & ~n4996 ;
  assign n5173 = ~n4898 & ~n4900 ;
  assign n5174 = x76 & n2093 ;
  assign n5175 = x74 & n2275 ;
  assign n5176 = x75 & n2088 ;
  assign n5177 = ~n5175 & ~n5176 ;
  assign n5178 = ~n5174 & n5177 ;
  assign n5179 = n1311 & n2096 ;
  assign n5180 = n5178 & ~n5179 ;
  assign n5181 = x17 & ~n5180 ;
  assign n5182 = x17 & ~n5181 ;
  assign n5183 = ~n5180 & ~n5181 ;
  assign n5184 = ~n5182 & ~n5183 ;
  assign n5185 = ~n4892 & ~n4894 ;
  assign n5186 = x26 & ~x27 ;
  assign n5187 = ~x26 & x27 ;
  assign n5188 = ~n5186 & ~n5187 ;
  assign n5189 = x64 & ~n5188 ;
  assign n5190 = ~n4859 & n5189 ;
  assign n5191 = n4859 & ~n5189 ;
  assign n5192 = ~n5190 & ~n5191 ;
  assign n5193 = x67 & n4531 ;
  assign n5194 = x65 & n4847 ;
  assign n5195 = x66 & n4526 ;
  assign n5196 = ~n5194 & ~n5195 ;
  assign n5197 = ~n5193 & n5196 ;
  assign n5198 = n240 & n4534 ;
  assign n5199 = n5197 & ~n5198 ;
  assign n5200 = x26 & ~n5199 ;
  assign n5201 = x26 & ~n5200 ;
  assign n5202 = ~n5199 & ~n5200 ;
  assign n5203 = ~n5201 & ~n5202 ;
  assign n5204 = ~n5192 & ~n5203 ;
  assign n5205 = n5192 & n5203 ;
  assign n5206 = ~n5204 & ~n5205 ;
  assign n5207 = x70 & n3589 ;
  assign n5208 = x68 & n3878 ;
  assign n5209 = x69 & n3584 ;
  assign n5210 = ~n5208 & ~n5209 ;
  assign n5211 = ~n5207 & n5210 ;
  assign n5212 = n488 & n3592 ;
  assign n5213 = n5211 & ~n5212 ;
  assign n5214 = x23 & ~n5213 ;
  assign n5215 = x23 & ~n5214 ;
  assign n5216 = ~n5213 & ~n5214 ;
  assign n5217 = ~n5215 & ~n5216 ;
  assign n5218 = n5206 & ~n5217 ;
  assign n5219 = n5206 & ~n5218 ;
  assign n5220 = ~n5217 & ~n5218 ;
  assign n5221 = ~n5219 & ~n5220 ;
  assign n5222 = ~n4877 & n5221 ;
  assign n5223 = n4877 & ~n5221 ;
  assign n5224 = ~n5222 & ~n5223 ;
  assign n5225 = x73 & n2751 ;
  assign n5226 = x71 & n3020 ;
  assign n5227 = x72 & n2746 ;
  assign n5228 = ~n5226 & ~n5227 ;
  assign n5229 = ~n5225 & n5228 ;
  assign n5230 = n843 & n2754 ;
  assign n5231 = n5229 & ~n5230 ;
  assign n5232 = x20 & ~n5231 ;
  assign n5233 = x20 & ~n5232 ;
  assign n5234 = ~n5231 & ~n5232 ;
  assign n5235 = ~n5233 & ~n5234 ;
  assign n5236 = ~n5224 & ~n5235 ;
  assign n5237 = n5224 & n5235 ;
  assign n5238 = ~n5236 & ~n5237 ;
  assign n5239 = ~n5185 & n5238 ;
  assign n5240 = n5185 & ~n5238 ;
  assign n5241 = ~n5239 & ~n5240 ;
  assign n5242 = n5184 & ~n5241 ;
  assign n5243 = ~n5184 & n5241 ;
  assign n5244 = ~n5242 & ~n5243 ;
  assign n5245 = ~n5173 & n5244 ;
  assign n5246 = n5173 & ~n5244 ;
  assign n5247 = ~n5245 & ~n5246 ;
  assign n5248 = x79 & n1434 ;
  assign n5249 = x77 & n1646 ;
  assign n5250 = x78 & n1429 ;
  assign n5251 = ~n5249 & ~n5250 ;
  assign n5252 = ~n5248 & n5251 ;
  assign n5253 = n1437 & n1817 ;
  assign n5254 = n5252 & ~n5253 ;
  assign n5255 = x14 & ~n5254 ;
  assign n5256 = x14 & ~n5255 ;
  assign n5257 = ~n5254 & ~n5255 ;
  assign n5258 = ~n5256 & ~n5257 ;
  assign n5259 = n5247 & ~n5258 ;
  assign n5260 = n5247 & ~n5259 ;
  assign n5261 = ~n5258 & ~n5259 ;
  assign n5262 = ~n5260 & ~n5261 ;
  assign n5263 = ~n4829 & ~n4917 ;
  assign n5264 = ~n4914 & ~n5263 ;
  assign n5265 = n5262 & n5264 ;
  assign n5266 = ~n5262 & ~n5264 ;
  assign n5267 = ~n5265 & ~n5266 ;
  assign n5268 = x82 & n945 ;
  assign n5269 = x80 & n1099 ;
  assign n5270 = x81 & n940 ;
  assign n5271 = ~n5269 & ~n5270 ;
  assign n5272 = ~n5268 & n5271 ;
  assign n5273 = n948 & n2584 ;
  assign n5274 = n5272 & ~n5273 ;
  assign n5275 = x11 & ~n5274 ;
  assign n5276 = x11 & ~n5275 ;
  assign n5277 = ~n5274 & ~n5275 ;
  assign n5278 = ~n5276 & ~n5277 ;
  assign n5279 = n5267 & ~n5278 ;
  assign n5280 = n5267 & ~n5279 ;
  assign n5281 = ~n5278 & ~n5279 ;
  assign n5282 = ~n5280 & ~n5281 ;
  assign n5283 = ~n4932 & ~n4936 ;
  assign n5284 = n5282 & n5283 ;
  assign n5285 = ~n5282 & ~n5283 ;
  assign n5286 = ~n5284 & ~n5285 ;
  assign n5287 = x85 & n574 ;
  assign n5288 = x83 & n673 ;
  assign n5289 = x84 & n569 ;
  assign n5290 = ~n5288 & ~n5289 ;
  assign n5291 = ~n5287 & n5290 ;
  assign n5292 = n577 & n3389 ;
  assign n5293 = n5291 & ~n5292 ;
  assign n5294 = x8 & ~n5293 ;
  assign n5295 = x8 & ~n5294 ;
  assign n5296 = ~n5293 & ~n5294 ;
  assign n5297 = ~n5295 & ~n5296 ;
  assign n5298 = ~n5286 & n5297 ;
  assign n5299 = n5286 & ~n5297 ;
  assign n5300 = ~n5298 & ~n5299 ;
  assign n5301 = ~n4949 & ~n4955 ;
  assign n5302 = n5300 & ~n5301 ;
  assign n5303 = ~n5300 & n5301 ;
  assign n5304 = ~n5302 & ~n5303 ;
  assign n5305 = x88 & n293 ;
  assign n5306 = x86 & n373 ;
  assign n5307 = x87 & n288 ;
  assign n5308 = ~n5306 & ~n5307 ;
  assign n5309 = ~n5305 & n5308 ;
  assign n5310 = n296 & n4305 ;
  assign n5311 = n5309 & ~n5310 ;
  assign n5312 = x5 & ~n5311 ;
  assign n5313 = x5 & ~n5312 ;
  assign n5314 = ~n5311 & ~n5312 ;
  assign n5315 = ~n5313 & ~n5314 ;
  assign n5316 = n5304 & ~n5315 ;
  assign n5317 = n5304 & ~n5316 ;
  assign n5318 = ~n5315 & ~n5316 ;
  assign n5319 = ~n5317 & ~n5318 ;
  assign n5320 = ~n4827 & ~n4971 ;
  assign n5321 = ~n4968 & ~n5320 ;
  assign n5322 = n5319 & n5321 ;
  assign n5323 = ~n5319 & ~n5321 ;
  assign n5324 = ~n5322 & ~n5323 ;
  assign n5325 = x91 & n146 ;
  assign n5326 = x89 & n182 ;
  assign n5327 = x90 & n141 ;
  assign n5328 = ~n5326 & ~n5327 ;
  assign n5329 = ~n5325 & n5328 ;
  assign n5330 = ~n4982 & ~n4984 ;
  assign n5331 = ~x90 & ~x91 ;
  assign n5332 = x90 & x91 ;
  assign n5333 = ~n5331 & ~n5332 ;
  assign n5334 = ~n5330 & n5333 ;
  assign n5335 = n5330 & ~n5333 ;
  assign n5336 = ~n5334 & ~n5335 ;
  assign n5337 = n149 & n5336 ;
  assign n5338 = n5329 & ~n5337 ;
  assign n5339 = x2 & ~n5338 ;
  assign n5340 = x2 & ~n5339 ;
  assign n5341 = ~n5338 & ~n5339 ;
  assign n5342 = ~n5340 & ~n5341 ;
  assign n5343 = ~n5324 & n5342 ;
  assign n5344 = n5324 & ~n5342 ;
  assign n5345 = ~n5343 & ~n5344 ;
  assign n5346 = ~n5172 & n5345 ;
  assign n5347 = n5172 & ~n5345 ;
  assign n5348 = ~n5346 & ~n5347 ;
  assign n5521 = n5348 & x155 ;
  assign n5349 = ~n5162 & ~n5165 ;
  assign n5350 = ~n5070 & ~n5072 ;
  assign n5351 = ~x76 & n2093 ;
  assign n5352 = ~x74 & n2275 ;
  assign n5353 = ~x75 & n2088 ;
  assign n5354 = ~n5352 & ~n5353 ;
  assign n5355 = ~n5351 & n5354 ;
  assign n5356 = n1390 & n2096 ;
  assign n5357 = n5355 & ~n5356 ;
  assign n5358 = ~x17 & ~n5357 ;
  assign n5359 = ~x17 & ~n5358 ;
  assign n5360 = ~n5357 & ~n5358 ;
  assign n5361 = ~n5359 & ~n5360 ;
  assign n5362 = ~n5064 & ~n5066 ;
  assign n5363 = ~x64 & ~n5188 ;
  assign n5364 = ~n5031 & n5363 ;
  assign n5365 = n5031 & ~n5363 ;
  assign n5366 = ~n5364 & ~n5365 ;
  assign n5367 = ~x67 & n4531 ;
  assign n5368 = ~x65 & n4847 ;
  assign n5369 = ~x66 & n4526 ;
  assign n5370 = ~n5368 & ~n5369 ;
  assign n5371 = ~n5367 & n5370 ;
  assign n5372 = n266 & n4534 ;
  assign n5373 = n5371 & ~n5372 ;
  assign n5374 = ~x26 & ~n5373 ;
  assign n5375 = ~x26 & ~n5374 ;
  assign n5376 = ~n5373 & ~n5374 ;
  assign n5377 = ~n5375 & ~n5376 ;
  assign n5378 = ~n5366 & ~n5377 ;
  assign n5379 = n5366 & n5377 ;
  assign n5380 = ~n5378 & ~n5379 ;
  assign n5381 = ~x70 & n3589 ;
  assign n5382 = ~x68 & n3878 ;
  assign n5383 = ~x69 & n3584 ;
  assign n5384 = ~n5382 & ~n5383 ;
  assign n5385 = ~n5381 & n5384 ;
  assign n5386 = n529 & n3592 ;
  assign n5387 = n5385 & ~n5386 ;
  assign n5388 = ~x23 & ~n5387 ;
  assign n5389 = ~x23 & ~n5388 ;
  assign n5390 = ~n5387 & ~n5388 ;
  assign n5391 = ~n5389 & ~n5390 ;
  assign n5392 = n5380 & ~n5391 ;
  assign n5393 = n5380 & ~n5392 ;
  assign n5394 = ~n5391 & ~n5392 ;
  assign n5395 = ~n5393 & ~n5394 ;
  assign n5396 = ~n5049 & n5395 ;
  assign n5397 = n5049 & ~n5395 ;
  assign n5398 = ~n5396 & ~n5397 ;
  assign n5399 = ~x73 & n2751 ;
  assign n5400 = ~x71 & n3020 ;
  assign n5401 = ~x72 & n2746 ;
  assign n5402 = ~n5400 & ~n5401 ;
  assign n5403 = ~n5399 & n5402 ;
  assign n5404 = n903 & n2754 ;
  assign n5405 = n5403 & ~n5404 ;
  assign n5406 = ~x20 & ~n5405 ;
  assign n5407 = ~x20 & ~n5406 ;
  assign n5408 = ~n5405 & ~n5406 ;
  assign n5409 = ~n5407 & ~n5408 ;
  assign n5410 = ~n5398 & ~n5409 ;
  assign n5411 = n5398 & n5409 ;
  assign n5412 = ~n5410 & ~n5411 ;
  assign n5413 = ~n5362 & n5412 ;
  assign n5414 = n5362 & ~n5412 ;
  assign n5415 = ~n5413 & ~n5414 ;
  assign n5416 = n5361 & ~n5415 ;
  assign n5417 = ~n5361 & n5415 ;
  assign n5418 = ~n5416 & ~n5417 ;
  assign n5419 = ~n5350 & n5418 ;
  assign n5420 = n5350 & ~n5418 ;
  assign n5421 = ~n5419 & ~n5420 ;
  assign n5422 = ~x79 & n1434 ;
  assign n5423 = ~x77 & n1646 ;
  assign n5424 = ~x78 & n1429 ;
  assign n5425 = ~n5423 & ~n5424 ;
  assign n5426 = ~n5422 & n5425 ;
  assign n5427 = n1437 & n1921 ;
  assign n5428 = n5426 & ~n5427 ;
  assign n5429 = ~x14 & ~n5428 ;
  assign n5430 = ~x14 & ~n5429 ;
  assign n5431 = ~n5428 & ~n5429 ;
  assign n5432 = ~n5430 & ~n5431 ;
  assign n5433 = n5421 & ~n5432 ;
  assign n5434 = n5421 & ~n5433 ;
  assign n5435 = ~n5432 & ~n5433 ;
  assign n5436 = ~n5434 & ~n5435 ;
  assign n5437 = ~n5003 & ~n5089 ;
  assign n5438 = ~n5086 & ~n5437 ;
  assign n5439 = n5436 & n5438 ;
  assign n5440 = ~n5436 & ~n5438 ;
  assign n5441 = ~n5439 & ~n5440 ;
  assign n5442 = ~x82 & n945 ;
  assign n5443 = ~x80 & n1099 ;
  assign n5444 = ~x81 & n940 ;
  assign n5445 = ~n5443 & ~n5444 ;
  assign n5446 = ~n5442 & n5445 ;
  assign n5447 = n948 & n2697 ;
  assign n5448 = n5446 & ~n5447 ;
  assign n5449 = ~x11 & ~n5448 ;
  assign n5450 = ~x11 & ~n5449 ;
  assign n5451 = ~n5448 & ~n5449 ;
  assign n5452 = ~n5450 & ~n5451 ;
  assign n5453 = n5441 & ~n5452 ;
  assign n5454 = n5441 & ~n5453 ;
  assign n5455 = ~n5452 & ~n5453 ;
  assign n5456 = ~n5454 & ~n5455 ;
  assign n5457 = ~n5104 & ~n5108 ;
  assign n5458 = n5456 & n5457 ;
  assign n5459 = ~n5456 & ~n5457 ;
  assign n5460 = ~n5458 & ~n5459 ;
  assign n5461 = ~x85 & n574 ;
  assign n5462 = ~x83 & n673 ;
  assign n5463 = ~x84 & n569 ;
  assign n5464 = ~n5462 & ~n5463 ;
  assign n5465 = ~n5461 & n5464 ;
  assign n5466 = n577 & n3521 ;
  assign n5467 = n5465 & ~n5466 ;
  assign n5468 = ~x8 & ~n5467 ;
  assign n5469 = ~x8 & ~n5468 ;
  assign n5470 = ~n5467 & ~n5468 ;
  assign n5471 = ~n5469 & ~n5470 ;
  assign n5472 = ~n5460 & n5471 ;
  assign n5473 = n5460 & ~n5471 ;
  assign n5474 = ~n5472 & ~n5473 ;
  assign n5475 = ~n5121 & ~n5127 ;
  assign n5476 = n5474 & ~n5475 ;
  assign n5477 = ~n5474 & n5475 ;
  assign n5478 = ~n5476 & ~n5477 ;
  assign n5479 = ~x88 & n293 ;
  assign n5480 = ~x86 & n373 ;
  assign n5481 = ~x87 & n288 ;
  assign n5482 = ~n5480 & ~n5481 ;
  assign n5483 = ~n5479 & n5482 ;
  assign n5484 = n296 & n4457 ;
  assign n5485 = n5483 & ~n5484 ;
  assign n5486 = ~x5 & ~n5485 ;
  assign n5487 = ~x5 & ~n5486 ;
  assign n5488 = ~n5485 & ~n5486 ;
  assign n5489 = ~n5487 & ~n5488 ;
  assign n5490 = n5478 & ~n5489 ;
  assign n5491 = n5478 & ~n5490 ;
  assign n5492 = ~n5489 & ~n5490 ;
  assign n5493 = ~n5491 & ~n5492 ;
  assign n5494 = ~n5001 & ~n5143 ;
  assign n5495 = ~n5140 & ~n5494 ;
  assign n5496 = n5493 & n5495 ;
  assign n5497 = ~n5493 & ~n5495 ;
  assign n5498 = ~n5496 & ~n5497 ;
  assign n5499 = ~x91 & n164 ;
  assign n5500 = ~x89 & n205 ;
  assign n5501 = ~x90 & n162 ;
  assign n5502 = ~n5500 & ~n5501 ;
  assign n5503 = ~n5499 & n5502 ;
  assign n5504 = ~n4981 & ~n5153 ;
  assign n5505 = n5333 & ~n5504 ;
  assign n5506 = ~n5333 & n5504 ;
  assign n5507 = ~n5505 & ~n5506 ;
  assign n5508 = n167 & n5507 ;
  assign n5509 = n5503 & ~n5508 ;
  assign n5510 = ~x2 & ~n5509 ;
  assign n5511 = ~x2 & ~n5510 ;
  assign n5512 = ~n5509 & ~n5510 ;
  assign n5513 = ~n5511 & ~n5512 ;
  assign n5514 = ~n5498 & n5513 ;
  assign n5515 = n5498 & ~n5513 ;
  assign n5516 = ~n5514 & ~n5515 ;
  assign n5517 = ~n5349 & n5516 ;
  assign n5518 = n5349 & ~n5516 ;
  assign n5519 = ~n5517 & ~n5518 ;
  assign n5522 = ~n5519 & ~x155 ;
  assign n5523 = ~n5521 & ~n5522 ;
  assign n5524 = ~n5344 & ~n5346 ;
  assign n5525 = ~n4877 & ~n5221 ;
  assign n5526 = ~n5218 & ~n5525 ;
  assign n5527 = x71 & n3589 ;
  assign n5528 = x69 & n3878 ;
  assign n5529 = x70 & n3584 ;
  assign n5530 = ~n5528 & ~n5529 ;
  assign n5531 = ~n5527 & n5530 ;
  assign n5532 = n558 & n3592 ;
  assign n5533 = n5531 & ~n5532 ;
  assign n5534 = x23 & ~n5533 ;
  assign n5535 = x23 & ~n5534 ;
  assign n5536 = ~n5533 & ~n5534 ;
  assign n5537 = ~n5535 & ~n5536 ;
  assign n5538 = n4859 & n5189 ;
  assign n5539 = ~n5204 & ~n5538 ;
  assign n5540 = x68 & n4531 ;
  assign n5541 = x66 & n4847 ;
  assign n5542 = x67 & n4526 ;
  assign n5543 = ~n5541 & ~n5542 ;
  assign n5544 = ~n5540 & n5543 ;
  assign n5545 = n317 & n4534 ;
  assign n5546 = n5544 & ~n5545 ;
  assign n5547 = x26 & ~n5546 ;
  assign n5548 = x26 & ~n5547 ;
  assign n5549 = ~n5546 & ~n5547 ;
  assign n5550 = ~n5548 & ~n5549 ;
  assign n5551 = x29 & ~n5189 ;
  assign n5552 = ~x27 & x28 ;
  assign n5553 = x27 & ~x28 ;
  assign n5554 = ~n5552 & ~n5553 ;
  assign n5555 = n5188 & ~n5554 ;
  assign n5556 = x64 & n5555 ;
  assign n5557 = ~x28 & x29 ;
  assign n5558 = x28 & ~x29 ;
  assign n5559 = ~n5557 & ~n5558 ;
  assign n5560 = ~n5188 & n5559 ;
  assign n5561 = x65 & n5560 ;
  assign n5562 = ~n5556 & ~n5561 ;
  assign n5563 = ~n5188 & ~n5559 ;
  assign n5564 = ~n152 & n5563 ;
  assign n5565 = n5562 & ~n5564 ;
  assign n5566 = x29 & ~n5565 ;
  assign n5567 = x29 & ~n5566 ;
  assign n5568 = ~n5565 & ~n5566 ;
  assign n5569 = ~n5567 & ~n5568 ;
  assign n5570 = n5551 & ~n5569 ;
  assign n5571 = ~n5551 & n5569 ;
  assign n5572 = ~n5570 & ~n5571 ;
  assign n5573 = n5550 & n5572 ;
  assign n5574 = ~n5550 & ~n5572 ;
  assign n5575 = ~n5573 & ~n5574 ;
  assign n5576 = ~n5539 & ~n5575 ;
  assign n5577 = n5539 & n5575 ;
  assign n5578 = ~n5576 & ~n5577 ;
  assign n5579 = ~n5537 & n5578 ;
  assign n5580 = n5537 & ~n5578 ;
  assign n5581 = ~n5579 & ~n5580 ;
  assign n5582 = ~n5526 & n5581 ;
  assign n5583 = n5526 & ~n5581 ;
  assign n5584 = ~n5582 & ~n5583 ;
  assign n5585 = x74 & n2751 ;
  assign n5586 = x72 & n3020 ;
  assign n5587 = x73 & n2746 ;
  assign n5588 = ~n5586 & ~n5587 ;
  assign n5589 = ~n5585 & n5588 ;
  assign n5590 = n994 & n2754 ;
  assign n5591 = n5589 & ~n5590 ;
  assign n5592 = x20 & ~n5591 ;
  assign n5593 = x20 & ~n5592 ;
  assign n5594 = ~n5591 & ~n5592 ;
  assign n5595 = ~n5593 & ~n5594 ;
  assign n5596 = n5584 & ~n5595 ;
  assign n5597 = n5584 & ~n5596 ;
  assign n5598 = ~n5595 & ~n5596 ;
  assign n5599 = ~n5597 & ~n5598 ;
  assign n5600 = ~n5236 & ~n5239 ;
  assign n5601 = n5599 & n5600 ;
  assign n5602 = ~n5599 & ~n5600 ;
  assign n5603 = ~n5601 & ~n5602 ;
  assign n5604 = x77 & n2093 ;
  assign n5605 = x75 & n2275 ;
  assign n5606 = x76 & n2088 ;
  assign n5607 = ~n5605 & ~n5606 ;
  assign n5608 = ~n5604 & n5607 ;
  assign n5609 = n1502 & n2096 ;
  assign n5610 = n5608 & ~n5609 ;
  assign n5611 = x17 & ~n5610 ;
  assign n5612 = x17 & ~n5611 ;
  assign n5613 = ~n5610 & ~n5611 ;
  assign n5614 = ~n5612 & ~n5613 ;
  assign n5615 = n5603 & ~n5614 ;
  assign n5616 = n5603 & ~n5615 ;
  assign n5617 = ~n5614 & ~n5615 ;
  assign n5618 = ~n5616 & ~n5617 ;
  assign n5619 = ~n5243 & ~n5245 ;
  assign n5620 = ~n5618 & ~n5619 ;
  assign n5621 = ~n5618 & ~n5620 ;
  assign n5622 = ~n5619 & ~n5620 ;
  assign n5623 = ~n5621 & ~n5622 ;
  assign n5624 = x80 & n1434 ;
  assign n5625 = x78 & n1646 ;
  assign n5626 = x79 & n1429 ;
  assign n5627 = ~n5625 & ~n5626 ;
  assign n5628 = ~n5624 & n5627 ;
  assign n5629 = n1437 & n2028 ;
  assign n5630 = n5628 & ~n5629 ;
  assign n5631 = x14 & ~n5630 ;
  assign n5632 = x14 & ~n5631 ;
  assign n5633 = ~n5630 & ~n5631 ;
  assign n5634 = ~n5632 & ~n5633 ;
  assign n5635 = ~n5623 & ~n5634 ;
  assign n5636 = ~n5623 & ~n5635 ;
  assign n5637 = ~n5634 & ~n5635 ;
  assign n5638 = ~n5636 & ~n5637 ;
  assign n5639 = ~n5259 & ~n5266 ;
  assign n5640 = n5638 & n5639 ;
  assign n5641 = ~n5638 & ~n5639 ;
  assign n5642 = ~n5640 & ~n5641 ;
  assign n5643 = x83 & n945 ;
  assign n5644 = x81 & n1099 ;
  assign n5645 = x82 & n940 ;
  assign n5646 = ~n5644 & ~n5645 ;
  assign n5647 = ~n5643 & n5646 ;
  assign n5648 = n948 & n2843 ;
  assign n5649 = n5647 & ~n5648 ;
  assign n5650 = x11 & ~n5649 ;
  assign n5651 = x11 & ~n5650 ;
  assign n5652 = ~n5649 & ~n5650 ;
  assign n5653 = ~n5651 & ~n5652 ;
  assign n5654 = n5642 & ~n5653 ;
  assign n5655 = n5642 & ~n5654 ;
  assign n5656 = ~n5653 & ~n5654 ;
  assign n5657 = ~n5655 & ~n5656 ;
  assign n5658 = ~n5279 & ~n5285 ;
  assign n5659 = n5657 & n5658 ;
  assign n5660 = ~n5657 & ~n5658 ;
  assign n5661 = ~n5659 & ~n5660 ;
  assign n5662 = x86 & n574 ;
  assign n5663 = x84 & n673 ;
  assign n5664 = x85 & n569 ;
  assign n5665 = ~n5663 & ~n5664 ;
  assign n5666 = ~n5662 & n5665 ;
  assign n5667 = n577 & n3686 ;
  assign n5668 = n5666 & ~n5667 ;
  assign n5669 = x8 & ~n5668 ;
  assign n5670 = x8 & ~n5669 ;
  assign n5671 = ~n5668 & ~n5669 ;
  assign n5672 = ~n5670 & ~n5671 ;
  assign n5673 = ~n5661 & n5672 ;
  assign n5674 = n5661 & ~n5672 ;
  assign n5675 = ~n5673 & ~n5674 ;
  assign n5676 = ~n5299 & ~n5302 ;
  assign n5677 = n5675 & ~n5676 ;
  assign n5678 = ~n5675 & n5676 ;
  assign n5679 = ~n5677 & ~n5678 ;
  assign n5680 = x89 & n293 ;
  assign n5681 = x87 & n373 ;
  assign n5682 = x88 & n288 ;
  assign n5683 = ~n5681 & ~n5682 ;
  assign n5684 = ~n5680 & n5683 ;
  assign n5685 = n296 & n4488 ;
  assign n5686 = n5684 & ~n5685 ;
  assign n5687 = x5 & ~n5686 ;
  assign n5688 = x5 & ~n5687 ;
  assign n5689 = ~n5686 & ~n5687 ;
  assign n5690 = ~n5688 & ~n5689 ;
  assign n5691 = n5679 & ~n5690 ;
  assign n5692 = n5679 & ~n5691 ;
  assign n5693 = ~n5690 & ~n5691 ;
  assign n5694 = ~n5692 & ~n5693 ;
  assign n5695 = ~n5316 & ~n5323 ;
  assign n5696 = n5694 & n5695 ;
  assign n5697 = ~n5694 & ~n5695 ;
  assign n5698 = ~n5696 & ~n5697 ;
  assign n5699 = x92 & n146 ;
  assign n5700 = x90 & n182 ;
  assign n5701 = x91 & n141 ;
  assign n5702 = ~n5700 & ~n5701 ;
  assign n5703 = ~n5699 & n5702 ;
  assign n5704 = ~n5332 & ~n5334 ;
  assign n5705 = ~x91 & ~x92 ;
  assign n5706 = x91 & x92 ;
  assign n5707 = ~n5705 & ~n5706 ;
  assign n5708 = ~n5704 & n5707 ;
  assign n5709 = n5704 & ~n5707 ;
  assign n5710 = ~n5708 & ~n5709 ;
  assign n5711 = n149 & n5710 ;
  assign n5712 = n5703 & ~n5711 ;
  assign n5713 = x2 & ~n5712 ;
  assign n5714 = x2 & ~n5713 ;
  assign n5715 = ~n5712 & ~n5713 ;
  assign n5716 = ~n5714 & ~n5715 ;
  assign n5717 = ~n5698 & n5716 ;
  assign n5718 = n5698 & ~n5716 ;
  assign n5719 = ~n5717 & ~n5718 ;
  assign n5720 = ~n5524 & n5719 ;
  assign n5721 = n5524 & ~n5719 ;
  assign n5722 = ~n5720 & ~n5721 ;
  assign n5910 = n5722 & x156 ;
  assign n5723 = ~n5515 & ~n5517 ;
  assign n5724 = ~n5049 & ~n5395 ;
  assign n5725 = ~n5392 & ~n5724 ;
  assign n5726 = ~x71 & n3589 ;
  assign n5727 = ~x69 & n3878 ;
  assign n5728 = ~x70 & n3584 ;
  assign n5729 = ~n5727 & ~n5728 ;
  assign n5730 = ~n5726 & n5729 ;
  assign n5731 = n622 & n3592 ;
  assign n5732 = n5730 & ~n5731 ;
  assign n5733 = ~x23 & ~n5732 ;
  assign n5734 = ~x23 & ~n5733 ;
  assign n5735 = ~n5732 & ~n5733 ;
  assign n5736 = ~n5734 & ~n5735 ;
  assign n5737 = n5031 & n5363 ;
  assign n5738 = ~n5378 & ~n5737 ;
  assign n5739 = ~x68 & n4531 ;
  assign n5740 = ~x66 & n4847 ;
  assign n5741 = ~x67 & n4526 ;
  assign n5742 = ~n5740 & ~n5741 ;
  assign n5743 = ~n5739 & n5742 ;
  assign n5744 = n352 & n4534 ;
  assign n5745 = n5743 & ~n5744 ;
  assign n5746 = ~x26 & ~n5745 ;
  assign n5747 = ~x26 & ~n5746 ;
  assign n5748 = ~n5745 & ~n5746 ;
  assign n5749 = ~n5747 & ~n5748 ;
  assign n5750 = ~x29 & ~n5363 ;
  assign n5751 = ~x64 & n5555 ;
  assign n5752 = ~x65 & n5560 ;
  assign n5753 = ~n5751 & ~n5752 ;
  assign n5754 = ~n5564 & n5753 ;
  assign n5755 = ~x29 & ~n5754 ;
  assign n5756 = ~x29 & ~n5755 ;
  assign n5757 = ~n5754 & ~n5755 ;
  assign n5758 = ~n5756 & ~n5757 ;
  assign n5759 = n5750 & ~n5758 ;
  assign n5760 = ~n5750 & n5758 ;
  assign n5761 = ~n5759 & ~n5760 ;
  assign n5762 = n5749 & n5761 ;
  assign n5763 = ~n5749 & ~n5761 ;
  assign n5764 = ~n5762 & ~n5763 ;
  assign n5765 = ~n5738 & ~n5764 ;
  assign n5766 = n5738 & n5764 ;
  assign n5767 = ~n5765 & ~n5766 ;
  assign n5768 = ~n5736 & n5767 ;
  assign n5769 = n5736 & ~n5767 ;
  assign n5770 = ~n5768 & ~n5769 ;
  assign n5771 = ~n5725 & n5770 ;
  assign n5772 = n5725 & ~n5770 ;
  assign n5773 = ~n5771 & ~n5772 ;
  assign n5774 = ~x74 & n2751 ;
  assign n5775 = ~x72 & n3020 ;
  assign n5776 = ~x73 & n2746 ;
  assign n5777 = ~n5775 & ~n5776 ;
  assign n5778 = ~n5774 & n5777 ;
  assign n5779 = n1066 & n2754 ;
  assign n5780 = n5778 & ~n5779 ;
  assign n5781 = ~x20 & ~n5780 ;
  assign n5782 = ~x20 & ~n5781 ;
  assign n5783 = ~n5780 & ~n5781 ;
  assign n5784 = ~n5782 & ~n5783 ;
  assign n5785 = n5773 & ~n5784 ;
  assign n5786 = n5773 & ~n5785 ;
  assign n5787 = ~n5784 & ~n5785 ;
  assign n5788 = ~n5786 & ~n5787 ;
  assign n5789 = ~n5410 & ~n5413 ;
  assign n5790 = n5788 & n5789 ;
  assign n5791 = ~n5788 & ~n5789 ;
  assign n5792 = ~n5790 & ~n5791 ;
  assign n5793 = ~x77 & n2093 ;
  assign n5794 = ~x75 & n2275 ;
  assign n5795 = ~x76 & n2088 ;
  assign n5796 = ~n5794 & ~n5795 ;
  assign n5797 = ~n5793 & n5796 ;
  assign n5798 = n1594 & n2096 ;
  assign n5799 = n5797 & ~n5798 ;
  assign n5800 = ~x17 & ~n5799 ;
  assign n5801 = ~x17 & ~n5800 ;
  assign n5802 = ~n5799 & ~n5800 ;
  assign n5803 = ~n5801 & ~n5802 ;
  assign n5804 = n5792 & ~n5803 ;
  assign n5805 = n5792 & ~n5804 ;
  assign n5806 = ~n5803 & ~n5804 ;
  assign n5807 = ~n5805 & ~n5806 ;
  assign n5808 = ~n5417 & ~n5419 ;
  assign n5809 = ~n5807 & ~n5808 ;
  assign n5810 = ~n5807 & ~n5809 ;
  assign n5811 = ~n5808 & ~n5809 ;
  assign n5812 = ~n5810 & ~n5811 ;
  assign n5813 = ~x80 & n1434 ;
  assign n5814 = ~x78 & n1646 ;
  assign n5815 = ~x79 & n1429 ;
  assign n5816 = ~n5814 & ~n5815 ;
  assign n5817 = ~n5813 & n5816 ;
  assign n5818 = n1437 & n2145 ;
  assign n5819 = n5817 & ~n5818 ;
  assign n5820 = ~x14 & ~n5819 ;
  assign n5821 = ~x14 & ~n5820 ;
  assign n5822 = ~n5819 & ~n5820 ;
  assign n5823 = ~n5821 & ~n5822 ;
  assign n5824 = ~n5812 & ~n5823 ;
  assign n5825 = ~n5812 & ~n5824 ;
  assign n5826 = ~n5823 & ~n5824 ;
  assign n5827 = ~n5825 & ~n5826 ;
  assign n5828 = ~n5433 & ~n5440 ;
  assign n5829 = n5827 & n5828 ;
  assign n5830 = ~n5827 & ~n5828 ;
  assign n5831 = ~n5829 & ~n5830 ;
  assign n5832 = ~x83 & n945 ;
  assign n5833 = ~x81 & n1099 ;
  assign n5834 = ~x82 & n940 ;
  assign n5835 = ~n5833 & ~n5834 ;
  assign n5836 = ~n5832 & n5835 ;
  assign n5837 = n948 & n2972 ;
  assign n5838 = n5836 & ~n5837 ;
  assign n5839 = ~x11 & ~n5838 ;
  assign n5840 = ~x11 & ~n5839 ;
  assign n5841 = ~n5838 & ~n5839 ;
  assign n5842 = ~n5840 & ~n5841 ;
  assign n5843 = n5831 & ~n5842 ;
  assign n5844 = n5831 & ~n5843 ;
  assign n5845 = ~n5842 & ~n5843 ;
  assign n5846 = ~n5844 & ~n5845 ;
  assign n5847 = ~n5453 & ~n5459 ;
  assign n5848 = n5846 & n5847 ;
  assign n5849 = ~n5846 & ~n5847 ;
  assign n5850 = ~n5848 & ~n5849 ;
  assign n5851 = ~x86 & n574 ;
  assign n5852 = ~x84 & n673 ;
  assign n5853 = ~x85 & n569 ;
  assign n5854 = ~n5852 & ~n5853 ;
  assign n5855 = ~n5851 & n5854 ;
  assign n5856 = n577 & n3832 ;
  assign n5857 = n5855 & ~n5856 ;
  assign n5858 = ~x8 & ~n5857 ;
  assign n5859 = ~x8 & ~n5858 ;
  assign n5860 = ~n5857 & ~n5858 ;
  assign n5861 = ~n5859 & ~n5860 ;
  assign n5862 = ~n5850 & n5861 ;
  assign n5863 = n5850 & ~n5861 ;
  assign n5864 = ~n5862 & ~n5863 ;
  assign n5865 = ~n5473 & ~n5476 ;
  assign n5866 = n5864 & ~n5865 ;
  assign n5867 = ~n5864 & n5865 ;
  assign n5868 = ~n5866 & ~n5867 ;
  assign n5869 = ~x89 & n293 ;
  assign n5870 = ~x87 & n373 ;
  assign n5871 = ~x88 & n288 ;
  assign n5872 = ~n5870 & ~n5871 ;
  assign n5873 = ~n5869 & n5872 ;
  assign n5874 = n296 & n4664 ;
  assign n5875 = n5873 & ~n5874 ;
  assign n5876 = ~x5 & ~n5875 ;
  assign n5877 = ~x5 & ~n5876 ;
  assign n5878 = ~n5875 & ~n5876 ;
  assign n5879 = ~n5877 & ~n5878 ;
  assign n5880 = n5868 & ~n5879 ;
  assign n5881 = n5868 & ~n5880 ;
  assign n5882 = ~n5879 & ~n5880 ;
  assign n5883 = ~n5881 & ~n5882 ;
  assign n5884 = ~n5490 & ~n5497 ;
  assign n5885 = n5883 & n5884 ;
  assign n5886 = ~n5883 & ~n5884 ;
  assign n5887 = ~n5885 & ~n5886 ;
  assign n5888 = ~x92 & n164 ;
  assign n5889 = ~x90 & n205 ;
  assign n5890 = ~x91 & n162 ;
  assign n5891 = ~n5889 & ~n5890 ;
  assign n5892 = ~n5888 & n5891 ;
  assign n5893 = ~n5331 & ~n5505 ;
  assign n5894 = n5707 & ~n5893 ;
  assign n5895 = ~n5707 & n5893 ;
  assign n5896 = ~n5894 & ~n5895 ;
  assign n5897 = n167 & n5896 ;
  assign n5898 = n5892 & ~n5897 ;
  assign n5899 = ~x2 & ~n5898 ;
  assign n5900 = ~x2 & ~n5899 ;
  assign n5901 = ~n5898 & ~n5899 ;
  assign n5902 = ~n5900 & ~n5901 ;
  assign n5903 = ~n5887 & n5902 ;
  assign n5904 = n5887 & ~n5902 ;
  assign n5905 = ~n5903 & ~n5904 ;
  assign n5906 = ~n5723 & n5905 ;
  assign n5907 = n5723 & ~n5905 ;
  assign n5908 = ~n5906 & ~n5907 ;
  assign n5911 = ~n5908 & ~x156 ;
  assign n5912 = ~n5910 & ~n5911 ;
  assign n5913 = ~n5691 & ~n5697 ;
  assign n5914 = x90 & n293 ;
  assign n5915 = x88 & n373 ;
  assign n5916 = x89 & n288 ;
  assign n5917 = ~n5915 & ~n5916 ;
  assign n5918 = ~n5914 & n5917 ;
  assign n5919 = n296 & n4986 ;
  assign n5920 = n5918 & ~n5919 ;
  assign n5921 = x5 & ~n5920 ;
  assign n5922 = x5 & ~n5921 ;
  assign n5923 = ~n5920 & ~n5921 ;
  assign n5924 = ~n5922 & ~n5923 ;
  assign n5925 = ~n5654 & ~n5660 ;
  assign n5926 = ~n5596 & ~n5602 ;
  assign n5927 = x75 & n2751 ;
  assign n5928 = x73 & n3020 ;
  assign n5929 = x74 & n2746 ;
  assign n5930 = ~n5928 & ~n5929 ;
  assign n5931 = ~n5927 & n5930 ;
  assign n5932 = n1150 & n2754 ;
  assign n5933 = n5931 & ~n5932 ;
  assign n5934 = x20 & ~n5933 ;
  assign n5935 = x20 & ~n5934 ;
  assign n5936 = ~n5933 & ~n5934 ;
  assign n5937 = ~n5935 & ~n5936 ;
  assign n5938 = ~n5579 & ~n5582 ;
  assign n5939 = ~n5550 & n5572 ;
  assign n5940 = ~n5576 & ~n5939 ;
  assign n5941 = x66 & n5560 ;
  assign n5942 = n5188 & ~n5559 ;
  assign n5943 = n5554 & n5942 ;
  assign n5944 = x64 & n5943 ;
  assign n5945 = x65 & n5555 ;
  assign n5946 = ~n5944 & ~n5945 ;
  assign n5947 = ~n5941 & n5946 ;
  assign n5948 = n194 & n5563 ;
  assign n5949 = n5947 & ~n5948 ;
  assign n5950 = x29 & ~n5949 ;
  assign n5951 = x29 & ~n5950 ;
  assign n5952 = ~n5949 & ~n5950 ;
  assign n5953 = ~n5951 & ~n5952 ;
  assign n5954 = ~n5570 & n5953 ;
  assign n5955 = n5570 & ~n5953 ;
  assign n5956 = ~n5954 & ~n5955 ;
  assign n5957 = x69 & n4531 ;
  assign n5958 = x67 & n4847 ;
  assign n5959 = x68 & n4526 ;
  assign n5960 = ~n5958 & ~n5959 ;
  assign n5961 = ~n5957 & n5960 ;
  assign n5962 = n398 & n4534 ;
  assign n5963 = n5961 & ~n5962 ;
  assign n5964 = x26 & ~n5963 ;
  assign n5965 = x26 & ~n5964 ;
  assign n5966 = ~n5963 & ~n5964 ;
  assign n5967 = ~n5965 & ~n5966 ;
  assign n5968 = n5956 & ~n5967 ;
  assign n5969 = ~n5956 & n5967 ;
  assign n5970 = ~n5940 & ~n5969 ;
  assign n5971 = ~n5968 & n5970 ;
  assign n5972 = ~n5940 & ~n5971 ;
  assign n5973 = ~n5968 & ~n5971 ;
  assign n5974 = ~n5969 & n5973 ;
  assign n5975 = ~n5972 & ~n5974 ;
  assign n5976 = x72 & n3589 ;
  assign n5977 = x70 & n3878 ;
  assign n5978 = x71 & n3584 ;
  assign n5979 = ~n5977 & ~n5978 ;
  assign n5980 = ~n5976 & n5979 ;
  assign n5981 = n717 & n3592 ;
  assign n5982 = n5980 & ~n5981 ;
  assign n5983 = x23 & ~n5982 ;
  assign n5984 = x23 & ~n5983 ;
  assign n5985 = ~n5982 & ~n5983 ;
  assign n5986 = ~n5984 & ~n5985 ;
  assign n5987 = n5975 & n5986 ;
  assign n5988 = ~n5975 & ~n5986 ;
  assign n5989 = ~n5987 & ~n5988 ;
  assign n5990 = ~n5938 & n5989 ;
  assign n5991 = n5938 & ~n5989 ;
  assign n5992 = ~n5990 & ~n5991 ;
  assign n5993 = n5937 & ~n5992 ;
  assign n5994 = ~n5937 & n5992 ;
  assign n5995 = ~n5993 & ~n5994 ;
  assign n5996 = ~n5926 & n5995 ;
  assign n5997 = n5926 & ~n5995 ;
  assign n5998 = ~n5996 & ~n5997 ;
  assign n5999 = x78 & n2093 ;
  assign n6000 = x76 & n2275 ;
  assign n6001 = x77 & n2088 ;
  assign n6002 = ~n6000 & ~n6001 ;
  assign n6003 = ~n5999 & n6002 ;
  assign n6004 = n1624 & n2096 ;
  assign n6005 = n6003 & ~n6004 ;
  assign n6006 = x17 & ~n6005 ;
  assign n6007 = x17 & ~n6006 ;
  assign n6008 = ~n6005 & ~n6006 ;
  assign n6009 = ~n6007 & ~n6008 ;
  assign n6010 = n5998 & ~n6009 ;
  assign n6011 = n5998 & ~n6010 ;
  assign n6012 = ~n6009 & ~n6010 ;
  assign n6013 = ~n6011 & ~n6012 ;
  assign n6014 = ~n5615 & ~n5620 ;
  assign n6015 = n6013 & n6014 ;
  assign n6016 = ~n6013 & ~n6014 ;
  assign n6017 = ~n6015 & ~n6016 ;
  assign n6018 = x81 & n1434 ;
  assign n6019 = x79 & n1646 ;
  assign n6020 = x80 & n1429 ;
  assign n6021 = ~n6019 & ~n6020 ;
  assign n6022 = ~n6018 & n6021 ;
  assign n6023 = n1437 & n2348 ;
  assign n6024 = n6022 & ~n6023 ;
  assign n6025 = x14 & ~n6024 ;
  assign n6026 = x14 & ~n6025 ;
  assign n6027 = ~n6024 & ~n6025 ;
  assign n6028 = ~n6026 & ~n6027 ;
  assign n6029 = n6017 & ~n6028 ;
  assign n6030 = n6017 & ~n6029 ;
  assign n6031 = ~n6028 & ~n6029 ;
  assign n6032 = ~n6030 & ~n6031 ;
  assign n6033 = ~n5635 & ~n5641 ;
  assign n6034 = n6032 & n6033 ;
  assign n6035 = ~n6032 & ~n6033 ;
  assign n6036 = ~n6034 & ~n6035 ;
  assign n6037 = x84 & n945 ;
  assign n6038 = x82 & n1099 ;
  assign n6039 = x83 & n940 ;
  assign n6040 = ~n6038 & ~n6039 ;
  assign n6041 = ~n6037 & n6040 ;
  assign n6042 = n948 & n3114 ;
  assign n6043 = n6041 & ~n6042 ;
  assign n6044 = x11 & ~n6043 ;
  assign n6045 = x11 & ~n6044 ;
  assign n6046 = ~n6043 & ~n6044 ;
  assign n6047 = ~n6045 & ~n6046 ;
  assign n6048 = n6036 & ~n6047 ;
  assign n6049 = ~n6036 & n6047 ;
  assign n6050 = ~n5925 & ~n6049 ;
  assign n6051 = ~n6048 & n6050 ;
  assign n6052 = ~n5925 & ~n6051 ;
  assign n6053 = ~n6048 & ~n6051 ;
  assign n6054 = ~n6049 & n6053 ;
  assign n6055 = ~n6052 & ~n6054 ;
  assign n6056 = x87 & n574 ;
  assign n6057 = x85 & n673 ;
  assign n6058 = x86 & n569 ;
  assign n6059 = ~n6057 & ~n6058 ;
  assign n6060 = ~n6056 & n6059 ;
  assign n6061 = n577 & n3991 ;
  assign n6062 = n6060 & ~n6061 ;
  assign n6063 = x8 & ~n6062 ;
  assign n6064 = x8 & ~n6063 ;
  assign n6065 = ~n6062 & ~n6063 ;
  assign n6066 = ~n6064 & ~n6065 ;
  assign n6067 = ~n6055 & ~n6066 ;
  assign n6068 = ~n6055 & ~n6067 ;
  assign n6069 = ~n6066 & ~n6067 ;
  assign n6070 = ~n6068 & ~n6069 ;
  assign n6071 = ~n5674 & ~n5677 ;
  assign n6072 = ~n6070 & ~n6071 ;
  assign n6073 = n6070 & n6071 ;
  assign n6074 = ~n6072 & ~n6073 ;
  assign n6075 = ~n5924 & n6074 ;
  assign n6076 = ~n5924 & ~n6075 ;
  assign n6077 = n6074 & ~n6075 ;
  assign n6078 = ~n6076 & ~n6077 ;
  assign n6079 = ~n5913 & ~n6078 ;
  assign n6080 = ~n5913 & ~n6079 ;
  assign n6081 = ~n6078 & ~n6079 ;
  assign n6082 = ~n6080 & ~n6081 ;
  assign n6083 = x93 & n146 ;
  assign n6084 = x91 & n182 ;
  assign n6085 = x92 & n141 ;
  assign n6086 = ~n6084 & ~n6085 ;
  assign n6087 = ~n6083 & n6086 ;
  assign n6088 = ~n5706 & ~n5708 ;
  assign n6089 = ~x92 & ~x93 ;
  assign n6090 = x92 & x93 ;
  assign n6091 = ~n6089 & ~n6090 ;
  assign n6092 = ~n6088 & n6091 ;
  assign n6093 = n6088 & ~n6091 ;
  assign n6094 = ~n6092 & ~n6093 ;
  assign n6095 = n149 & n6094 ;
  assign n6096 = n6087 & ~n6095 ;
  assign n6097 = x2 & ~n6096 ;
  assign n6098 = x2 & ~n6097 ;
  assign n6099 = ~n6096 & ~n6097 ;
  assign n6100 = ~n6098 & ~n6099 ;
  assign n6101 = ~n6082 & ~n6100 ;
  assign n6102 = ~n6082 & ~n6101 ;
  assign n6103 = ~n6100 & ~n6101 ;
  assign n6104 = ~n6102 & ~n6103 ;
  assign n6105 = ~n5718 & ~n5720 ;
  assign n6106 = ~n6104 & ~n6105 ;
  assign n6107 = n6104 & n6105 ;
  assign n6108 = ~n6106 & ~n6107 ;
  assign n6301 = n6108 & x157 ;
  assign n6109 = ~n5880 & ~n5886 ;
  assign n6110 = ~x90 & n293 ;
  assign n6111 = ~x88 & n373 ;
  assign n6112 = ~x89 & n288 ;
  assign n6113 = ~n6111 & ~n6112 ;
  assign n6114 = ~n6110 & n6113 ;
  assign n6115 = n296 & n5155 ;
  assign n6116 = n6114 & ~n6115 ;
  assign n6117 = ~x5 & ~n6116 ;
  assign n6118 = ~x5 & ~n6117 ;
  assign n6119 = ~n6116 & ~n6117 ;
  assign n6120 = ~n6118 & ~n6119 ;
  assign n6121 = ~n5843 & ~n5849 ;
  assign n6122 = ~n5785 & ~n5791 ;
  assign n6123 = ~x75 & n2751 ;
  assign n6124 = ~x73 & n3020 ;
  assign n6125 = ~x74 & n2746 ;
  assign n6126 = ~n6124 & ~n6125 ;
  assign n6127 = ~n6123 & n6126 ;
  assign n6128 = n1225 & n2754 ;
  assign n6129 = n6127 & ~n6128 ;
  assign n6130 = ~x20 & ~n6129 ;
  assign n6131 = ~x20 & ~n6130 ;
  assign n6132 = ~n6129 & ~n6130 ;
  assign n6133 = ~n6131 & ~n6132 ;
  assign n6134 = ~n5768 & ~n5771 ;
  assign n6135 = ~n5749 & n5761 ;
  assign n6136 = ~n5765 & ~n6135 ;
  assign n6137 = ~x66 & n5560 ;
  assign n6138 = ~x64 & n5943 ;
  assign n6139 = ~x65 & n5555 ;
  assign n6140 = ~n6138 & ~n6139 ;
  assign n6141 = ~n6137 & n6140 ;
  assign n6142 = n214 & n5563 ;
  assign n6143 = n6141 & ~n6142 ;
  assign n6144 = ~x29 & ~n6143 ;
  assign n6145 = ~x29 & ~n6144 ;
  assign n6146 = ~n6143 & ~n6144 ;
  assign n6147 = ~n6145 & ~n6146 ;
  assign n6148 = ~n5759 & n6147 ;
  assign n6149 = n5759 & ~n6147 ;
  assign n6150 = ~n6148 & ~n6149 ;
  assign n6151 = ~x69 & n4531 ;
  assign n6152 = ~x67 & n4847 ;
  assign n6153 = ~x68 & n4526 ;
  assign n6154 = ~n6152 & ~n6153 ;
  assign n6155 = ~n6151 & n6154 ;
  assign n6156 = n435 & n4534 ;
  assign n6157 = n6155 & ~n6156 ;
  assign n6158 = ~x26 & ~n6157 ;
  assign n6159 = ~x26 & ~n6158 ;
  assign n6160 = ~n6157 & ~n6158 ;
  assign n6161 = ~n6159 & ~n6160 ;
  assign n6162 = n6150 & ~n6161 ;
  assign n6163 = ~n6150 & n6161 ;
  assign n6164 = ~n6136 & ~n6163 ;
  assign n6165 = ~n6162 & n6164 ;
  assign n6166 = ~n6136 & ~n6165 ;
  assign n6167 = ~n6162 & ~n6165 ;
  assign n6168 = ~n6163 & n6167 ;
  assign n6169 = ~n6166 & ~n6168 ;
  assign n6170 = ~x72 & n3589 ;
  assign n6171 = ~x70 & n3878 ;
  assign n6172 = ~x71 & n3584 ;
  assign n6173 = ~n6171 & ~n6172 ;
  assign n6174 = ~n6170 & n6173 ;
  assign n6175 = n773 & n3592 ;
  assign n6176 = n6174 & ~n6175 ;
  assign n6177 = ~x23 & ~n6176 ;
  assign n6178 = ~x23 & ~n6177 ;
  assign n6179 = ~n6176 & ~n6177 ;
  assign n6180 = ~n6178 & ~n6179 ;
  assign n6181 = n6169 & n6180 ;
  assign n6182 = ~n6169 & ~n6180 ;
  assign n6183 = ~n6181 & ~n6182 ;
  assign n6184 = ~n6134 & n6183 ;
  assign n6185 = n6134 & ~n6183 ;
  assign n6186 = ~n6184 & ~n6185 ;
  assign n6187 = n6133 & ~n6186 ;
  assign n6188 = ~n6133 & n6186 ;
  assign n6189 = ~n6187 & ~n6188 ;
  assign n6190 = ~n6122 & n6189 ;
  assign n6191 = n6122 & ~n6189 ;
  assign n6192 = ~n6190 & ~n6191 ;
  assign n6193 = ~x78 & n2093 ;
  assign n6194 = ~x76 & n2275 ;
  assign n6195 = ~x77 & n2088 ;
  assign n6196 = ~n6194 & ~n6195 ;
  assign n6197 = ~n6193 & n6196 ;
  assign n6198 = n1718 & n2096 ;
  assign n6199 = n6197 & ~n6198 ;
  assign n6200 = ~x17 & ~n6199 ;
  assign n6201 = ~x17 & ~n6200 ;
  assign n6202 = ~n6199 & ~n6200 ;
  assign n6203 = ~n6201 & ~n6202 ;
  assign n6204 = n6192 & ~n6203 ;
  assign n6205 = n6192 & ~n6204 ;
  assign n6206 = ~n6203 & ~n6204 ;
  assign n6207 = ~n6205 & ~n6206 ;
  assign n6208 = ~n5804 & ~n5809 ;
  assign n6209 = n6207 & n6208 ;
  assign n6210 = ~n6207 & ~n6208 ;
  assign n6211 = ~n6209 & ~n6210 ;
  assign n6212 = ~x81 & n1434 ;
  assign n6213 = ~x79 & n1646 ;
  assign n6214 = ~x80 & n1429 ;
  assign n6215 = ~n6213 & ~n6214 ;
  assign n6216 = ~n6212 & n6215 ;
  assign n6217 = n1437 & n2460 ;
  assign n6218 = n6216 & ~n6217 ;
  assign n6219 = ~x14 & ~n6218 ;
  assign n6220 = ~x14 & ~n6219 ;
  assign n6221 = ~n6218 & ~n6219 ;
  assign n6222 = ~n6220 & ~n6221 ;
  assign n6223 = n6211 & ~n6222 ;
  assign n6224 = n6211 & ~n6223 ;
  assign n6225 = ~n6222 & ~n6223 ;
  assign n6226 = ~n6224 & ~n6225 ;
  assign n6227 = ~n5824 & ~n5830 ;
  assign n6228 = n6226 & n6227 ;
  assign n6229 = ~n6226 & ~n6227 ;
  assign n6230 = ~n6228 & ~n6229 ;
  assign n6231 = ~x84 & n945 ;
  assign n6232 = ~x82 & n1099 ;
  assign n6233 = ~x83 & n940 ;
  assign n6234 = ~n6232 & ~n6233 ;
  assign n6235 = ~n6231 & n6234 ;
  assign n6236 = n948 & n3247 ;
  assign n6237 = n6235 & ~n6236 ;
  assign n6238 = ~x11 & ~n6237 ;
  assign n6239 = ~x11 & ~n6238 ;
  assign n6240 = ~n6237 & ~n6238 ;
  assign n6241 = ~n6239 & ~n6240 ;
  assign n6242 = n6230 & ~n6241 ;
  assign n6243 = ~n6230 & n6241 ;
  assign n6244 = ~n6121 & ~n6243 ;
  assign n6245 = ~n6242 & n6244 ;
  assign n6246 = ~n6121 & ~n6245 ;
  assign n6247 = ~n6242 & ~n6245 ;
  assign n6248 = ~n6243 & n6247 ;
  assign n6249 = ~n6246 & ~n6248 ;
  assign n6250 = ~x87 & n574 ;
  assign n6251 = ~x85 & n673 ;
  assign n6252 = ~x86 & n569 ;
  assign n6253 = ~n6251 & ~n6252 ;
  assign n6254 = ~n6250 & n6253 ;
  assign n6255 = n577 & n4143 ;
  assign n6256 = n6254 & ~n6255 ;
  assign n6257 = ~x8 & ~n6256 ;
  assign n6258 = ~x8 & ~n6257 ;
  assign n6259 = ~n6256 & ~n6257 ;
  assign n6260 = ~n6258 & ~n6259 ;
  assign n6261 = ~n6249 & ~n6260 ;
  assign n6262 = ~n6249 & ~n6261 ;
  assign n6263 = ~n6260 & ~n6261 ;
  assign n6264 = ~n6262 & ~n6263 ;
  assign n6265 = ~n5863 & ~n5866 ;
  assign n6266 = ~n6264 & ~n6265 ;
  assign n6267 = n6264 & n6265 ;
  assign n6268 = ~n6266 & ~n6267 ;
  assign n6269 = ~n6120 & n6268 ;
  assign n6270 = ~n6120 & ~n6269 ;
  assign n6271 = n6268 & ~n6269 ;
  assign n6272 = ~n6270 & ~n6271 ;
  assign n6273 = ~n6109 & ~n6272 ;
  assign n6274 = ~n6109 & ~n6273 ;
  assign n6275 = ~n6272 & ~n6273 ;
  assign n6276 = ~n6274 & ~n6275 ;
  assign n6277 = ~x93 & n164 ;
  assign n6278 = ~x91 & n205 ;
  assign n6279 = ~x92 & n162 ;
  assign n6280 = ~n6278 & ~n6279 ;
  assign n6281 = ~n6277 & n6280 ;
  assign n6282 = ~n5705 & ~n5894 ;
  assign n6283 = n6091 & ~n6282 ;
  assign n6284 = ~n6091 & n6282 ;
  assign n6285 = ~n6283 & ~n6284 ;
  assign n6286 = n167 & n6285 ;
  assign n6287 = n6281 & ~n6286 ;
  assign n6288 = ~x2 & ~n6287 ;
  assign n6289 = ~x2 & ~n6288 ;
  assign n6290 = ~n6287 & ~n6288 ;
  assign n6291 = ~n6289 & ~n6290 ;
  assign n6292 = ~n6276 & ~n6291 ;
  assign n6293 = ~n6276 & ~n6292 ;
  assign n6294 = ~n6291 & ~n6292 ;
  assign n6295 = ~n6293 & ~n6294 ;
  assign n6296 = ~n5904 & ~n5906 ;
  assign n6297 = ~n6295 & ~n6296 ;
  assign n6298 = n6295 & n6296 ;
  assign n6299 = ~n6297 & ~n6298 ;
  assign n6302 = ~n6299 & ~x157 ;
  assign n6303 = ~n6301 & ~n6302 ;
  assign n6304 = ~n6067 & ~n6072 ;
  assign n6305 = ~n5994 & ~n5996 ;
  assign n6306 = x76 & n2751 ;
  assign n6307 = x74 & n3020 ;
  assign n6308 = x75 & n2746 ;
  assign n6309 = ~n6307 & ~n6308 ;
  assign n6310 = ~n6306 & n6309 ;
  assign n6311 = n1311 & n2754 ;
  assign n6312 = n6310 & ~n6311 ;
  assign n6313 = x20 & ~n6312 ;
  assign n6314 = x20 & ~n6313 ;
  assign n6315 = ~n6312 & ~n6313 ;
  assign n6316 = ~n6314 & ~n6315 ;
  assign n6317 = ~n5988 & ~n5990 ;
  assign n6318 = x29 & ~x30 ;
  assign n6319 = ~x29 & x30 ;
  assign n6320 = ~n6318 & ~n6319 ;
  assign n6321 = x64 & ~n6320 ;
  assign n6322 = ~n5955 & n6321 ;
  assign n6323 = n5955 & ~n6321 ;
  assign n6324 = ~n6322 & ~n6323 ;
  assign n6325 = x67 & n5560 ;
  assign n6326 = x65 & n5943 ;
  assign n6327 = x66 & n5555 ;
  assign n6328 = ~n6326 & ~n6327 ;
  assign n6329 = ~n6325 & n6328 ;
  assign n6330 = n240 & n5563 ;
  assign n6331 = n6329 & ~n6330 ;
  assign n6332 = x29 & ~n6331 ;
  assign n6333 = x29 & ~n6332 ;
  assign n6334 = ~n6331 & ~n6332 ;
  assign n6335 = ~n6333 & ~n6334 ;
  assign n6336 = ~n6324 & ~n6335 ;
  assign n6337 = n6324 & n6335 ;
  assign n6338 = ~n6336 & ~n6337 ;
  assign n6339 = x70 & n4531 ;
  assign n6340 = x68 & n4847 ;
  assign n6341 = x69 & n4526 ;
  assign n6342 = ~n6340 & ~n6341 ;
  assign n6343 = ~n6339 & n6342 ;
  assign n6344 = n488 & n4534 ;
  assign n6345 = n6343 & ~n6344 ;
  assign n6346 = x26 & ~n6345 ;
  assign n6347 = x26 & ~n6346 ;
  assign n6348 = ~n6345 & ~n6346 ;
  assign n6349 = ~n6347 & ~n6348 ;
  assign n6350 = n6338 & ~n6349 ;
  assign n6351 = n6338 & ~n6350 ;
  assign n6352 = ~n6349 & ~n6350 ;
  assign n6353 = ~n6351 & ~n6352 ;
  assign n6354 = ~n5973 & n6353 ;
  assign n6355 = n5973 & ~n6353 ;
  assign n6356 = ~n6354 & ~n6355 ;
  assign n6357 = x73 & n3589 ;
  assign n6358 = x71 & n3878 ;
  assign n6359 = x72 & n3584 ;
  assign n6360 = ~n6358 & ~n6359 ;
  assign n6361 = ~n6357 & n6360 ;
  assign n6362 = n843 & n3592 ;
  assign n6363 = n6361 & ~n6362 ;
  assign n6364 = x23 & ~n6363 ;
  assign n6365 = x23 & ~n6364 ;
  assign n6366 = ~n6363 & ~n6364 ;
  assign n6367 = ~n6365 & ~n6366 ;
  assign n6368 = ~n6356 & ~n6367 ;
  assign n6369 = n6356 & n6367 ;
  assign n6370 = ~n6368 & ~n6369 ;
  assign n6371 = ~n6317 & n6370 ;
  assign n6372 = n6317 & ~n6370 ;
  assign n6373 = ~n6371 & ~n6372 ;
  assign n6374 = n6316 & ~n6373 ;
  assign n6375 = ~n6316 & n6373 ;
  assign n6376 = ~n6374 & ~n6375 ;
  assign n6377 = ~n6305 & n6376 ;
  assign n6378 = n6305 & ~n6376 ;
  assign n6379 = ~n6377 & ~n6378 ;
  assign n6380 = x79 & n2093 ;
  assign n6381 = x77 & n2275 ;
  assign n6382 = x78 & n2088 ;
  assign n6383 = ~n6381 & ~n6382 ;
  assign n6384 = ~n6380 & n6383 ;
  assign n6385 = n1817 & n2096 ;
  assign n6386 = n6384 & ~n6385 ;
  assign n6387 = x17 & ~n6386 ;
  assign n6388 = x17 & ~n6387 ;
  assign n6389 = ~n6386 & ~n6387 ;
  assign n6390 = ~n6388 & ~n6389 ;
  assign n6391 = n6379 & ~n6390 ;
  assign n6392 = n6379 & ~n6391 ;
  assign n6393 = ~n6390 & ~n6391 ;
  assign n6394 = ~n6392 & ~n6393 ;
  assign n6395 = ~n6010 & ~n6016 ;
  assign n6396 = n6394 & n6395 ;
  assign n6397 = ~n6394 & ~n6395 ;
  assign n6398 = ~n6396 & ~n6397 ;
  assign n6399 = x82 & n1434 ;
  assign n6400 = x80 & n1646 ;
  assign n6401 = x81 & n1429 ;
  assign n6402 = ~n6400 & ~n6401 ;
  assign n6403 = ~n6399 & n6402 ;
  assign n6404 = n1437 & n2584 ;
  assign n6405 = n6403 & ~n6404 ;
  assign n6406 = x14 & ~n6405 ;
  assign n6407 = x14 & ~n6406 ;
  assign n6408 = ~n6405 & ~n6406 ;
  assign n6409 = ~n6407 & ~n6408 ;
  assign n6410 = n6398 & ~n6409 ;
  assign n6411 = n6398 & ~n6410 ;
  assign n6412 = ~n6409 & ~n6410 ;
  assign n6413 = ~n6411 & ~n6412 ;
  assign n6414 = ~n6029 & ~n6035 ;
  assign n6415 = n6413 & n6414 ;
  assign n6416 = ~n6413 & ~n6414 ;
  assign n6417 = ~n6415 & ~n6416 ;
  assign n6418 = x85 & n945 ;
  assign n6419 = x83 & n1099 ;
  assign n6420 = x84 & n940 ;
  assign n6421 = ~n6419 & ~n6420 ;
  assign n6422 = ~n6418 & n6421 ;
  assign n6423 = n948 & n3389 ;
  assign n6424 = n6422 & ~n6423 ;
  assign n6425 = x11 & ~n6424 ;
  assign n6426 = x11 & ~n6425 ;
  assign n6427 = ~n6424 & ~n6425 ;
  assign n6428 = ~n6426 & ~n6427 ;
  assign n6429 = n6417 & ~n6428 ;
  assign n6430 = n6417 & ~n6429 ;
  assign n6431 = ~n6428 & ~n6429 ;
  assign n6432 = ~n6430 & ~n6431 ;
  assign n6433 = ~n6053 & n6432 ;
  assign n6434 = n6053 & ~n6432 ;
  assign n6435 = ~n6433 & ~n6434 ;
  assign n6436 = x88 & n574 ;
  assign n6437 = x86 & n673 ;
  assign n6438 = x87 & n569 ;
  assign n6439 = ~n6437 & ~n6438 ;
  assign n6440 = ~n6436 & n6439 ;
  assign n6441 = n577 & n4305 ;
  assign n6442 = n6440 & ~n6441 ;
  assign n6443 = x8 & ~n6442 ;
  assign n6444 = x8 & ~n6443 ;
  assign n6445 = ~n6442 & ~n6443 ;
  assign n6446 = ~n6444 & ~n6445 ;
  assign n6447 = ~n6435 & ~n6446 ;
  assign n6448 = n6435 & n6446 ;
  assign n6449 = ~n6447 & ~n6448 ;
  assign n6450 = n6304 & ~n6449 ;
  assign n6451 = ~n6304 & n6449 ;
  assign n6452 = ~n6450 & ~n6451 ;
  assign n6453 = x91 & n293 ;
  assign n6454 = x89 & n373 ;
  assign n6455 = x90 & n288 ;
  assign n6456 = ~n6454 & ~n6455 ;
  assign n6457 = ~n6453 & n6456 ;
  assign n6458 = n296 & n5336 ;
  assign n6459 = n6457 & ~n6458 ;
  assign n6460 = x5 & ~n6459 ;
  assign n6461 = x5 & ~n6460 ;
  assign n6462 = ~n6459 & ~n6460 ;
  assign n6463 = ~n6461 & ~n6462 ;
  assign n6464 = n6452 & ~n6463 ;
  assign n6465 = n6452 & ~n6464 ;
  assign n6466 = ~n6463 & ~n6464 ;
  assign n6467 = ~n6465 & ~n6466 ;
  assign n6468 = ~n6075 & ~n6079 ;
  assign n6469 = n6467 & n6468 ;
  assign n6470 = ~n6467 & ~n6468 ;
  assign n6471 = ~n6469 & ~n6470 ;
  assign n6472 = x94 & n146 ;
  assign n6473 = x92 & n182 ;
  assign n6474 = x93 & n141 ;
  assign n6475 = ~n6473 & ~n6474 ;
  assign n6476 = ~n6472 & n6475 ;
  assign n6477 = ~n6090 & ~n6092 ;
  assign n6478 = ~x93 & ~x94 ;
  assign n6479 = x93 & x94 ;
  assign n6480 = ~n6478 & ~n6479 ;
  assign n6481 = ~n6477 & n6480 ;
  assign n6482 = n6477 & ~n6480 ;
  assign n6483 = ~n6481 & ~n6482 ;
  assign n6484 = n149 & n6483 ;
  assign n6485 = n6476 & ~n6484 ;
  assign n6486 = x2 & ~n6485 ;
  assign n6487 = x2 & ~n6486 ;
  assign n6488 = ~n6485 & ~n6486 ;
  assign n6489 = ~n6487 & ~n6488 ;
  assign n6490 = n6471 & ~n6489 ;
  assign n6491 = n6471 & ~n6490 ;
  assign n6492 = ~n6489 & ~n6490 ;
  assign n6493 = ~n6491 & ~n6492 ;
  assign n6494 = ~n6101 & ~n6106 ;
  assign n6495 = ~n6493 & ~n6494 ;
  assign n6496 = n6493 & n6494 ;
  assign n6497 = ~n6495 & ~n6496 ;
  assign n6687 = n6497 & x158 ;
  assign n6498 = ~n6261 & ~n6266 ;
  assign n6499 = ~n6188 & ~n6190 ;
  assign n6500 = ~x76 & n2751 ;
  assign n6501 = ~x74 & n3020 ;
  assign n6502 = ~x75 & n2746 ;
  assign n6503 = ~n6501 & ~n6502 ;
  assign n6504 = ~n6500 & n6503 ;
  assign n6505 = n1390 & n2754 ;
  assign n6506 = n6504 & ~n6505 ;
  assign n6507 = ~x20 & ~n6506 ;
  assign n6508 = ~x20 & ~n6507 ;
  assign n6509 = ~n6506 & ~n6507 ;
  assign n6510 = ~n6508 & ~n6509 ;
  assign n6511 = ~n6182 & ~n6184 ;
  assign n6512 = ~x64 & ~n6320 ;
  assign n6513 = ~n6149 & n6512 ;
  assign n6514 = n6149 & ~n6512 ;
  assign n6515 = ~n6513 & ~n6514 ;
  assign n6516 = ~x67 & n5560 ;
  assign n6517 = ~x65 & n5943 ;
  assign n6518 = ~x66 & n5555 ;
  assign n6519 = ~n6517 & ~n6518 ;
  assign n6520 = ~n6516 & n6519 ;
  assign n6521 = n266 & n5563 ;
  assign n6522 = n6520 & ~n6521 ;
  assign n6523 = ~x29 & ~n6522 ;
  assign n6524 = ~x29 & ~n6523 ;
  assign n6525 = ~n6522 & ~n6523 ;
  assign n6526 = ~n6524 & ~n6525 ;
  assign n6527 = ~n6515 & ~n6526 ;
  assign n6528 = n6515 & n6526 ;
  assign n6529 = ~n6527 & ~n6528 ;
  assign n6530 = ~x70 & n4531 ;
  assign n6531 = ~x68 & n4847 ;
  assign n6532 = ~x69 & n4526 ;
  assign n6533 = ~n6531 & ~n6532 ;
  assign n6534 = ~n6530 & n6533 ;
  assign n6535 = n529 & n4534 ;
  assign n6536 = n6534 & ~n6535 ;
  assign n6537 = ~x26 & ~n6536 ;
  assign n6538 = ~x26 & ~n6537 ;
  assign n6539 = ~n6536 & ~n6537 ;
  assign n6540 = ~n6538 & ~n6539 ;
  assign n6541 = n6529 & ~n6540 ;
  assign n6542 = n6529 & ~n6541 ;
  assign n6543 = ~n6540 & ~n6541 ;
  assign n6544 = ~n6542 & ~n6543 ;
  assign n6545 = ~n6167 & n6544 ;
  assign n6546 = n6167 & ~n6544 ;
  assign n6547 = ~n6545 & ~n6546 ;
  assign n6548 = ~x73 & n3589 ;
  assign n6549 = ~x71 & n3878 ;
  assign n6550 = ~x72 & n3584 ;
  assign n6551 = ~n6549 & ~n6550 ;
  assign n6552 = ~n6548 & n6551 ;
  assign n6553 = n903 & n3592 ;
  assign n6554 = n6552 & ~n6553 ;
  assign n6555 = ~x23 & ~n6554 ;
  assign n6556 = ~x23 & ~n6555 ;
  assign n6557 = ~n6554 & ~n6555 ;
  assign n6558 = ~n6556 & ~n6557 ;
  assign n6559 = ~n6547 & ~n6558 ;
  assign n6560 = n6547 & n6558 ;
  assign n6561 = ~n6559 & ~n6560 ;
  assign n6562 = ~n6511 & n6561 ;
  assign n6563 = n6511 & ~n6561 ;
  assign n6564 = ~n6562 & ~n6563 ;
  assign n6565 = n6510 & ~n6564 ;
  assign n6566 = ~n6510 & n6564 ;
  assign n6567 = ~n6565 & ~n6566 ;
  assign n6568 = ~n6499 & n6567 ;
  assign n6569 = n6499 & ~n6567 ;
  assign n6570 = ~n6568 & ~n6569 ;
  assign n6571 = ~x79 & n2093 ;
  assign n6572 = ~x77 & n2275 ;
  assign n6573 = ~x78 & n2088 ;
  assign n6574 = ~n6572 & ~n6573 ;
  assign n6575 = ~n6571 & n6574 ;
  assign n6576 = n1921 & n2096 ;
  assign n6577 = n6575 & ~n6576 ;
  assign n6578 = ~x17 & ~n6577 ;
  assign n6579 = ~x17 & ~n6578 ;
  assign n6580 = ~n6577 & ~n6578 ;
  assign n6581 = ~n6579 & ~n6580 ;
  assign n6582 = n6570 & ~n6581 ;
  assign n6583 = n6570 & ~n6582 ;
  assign n6584 = ~n6581 & ~n6582 ;
  assign n6585 = ~n6583 & ~n6584 ;
  assign n6586 = ~n6204 & ~n6210 ;
  assign n6587 = n6585 & n6586 ;
  assign n6588 = ~n6585 & ~n6586 ;
  assign n6589 = ~n6587 & ~n6588 ;
  assign n6590 = ~x82 & n1434 ;
  assign n6591 = ~x80 & n1646 ;
  assign n6592 = ~x81 & n1429 ;
  assign n6593 = ~n6591 & ~n6592 ;
  assign n6594 = ~n6590 & n6593 ;
  assign n6595 = n1437 & n2697 ;
  assign n6596 = n6594 & ~n6595 ;
  assign n6597 = ~x14 & ~n6596 ;
  assign n6598 = ~x14 & ~n6597 ;
  assign n6599 = ~n6596 & ~n6597 ;
  assign n6600 = ~n6598 & ~n6599 ;
  assign n6601 = n6589 & ~n6600 ;
  assign n6602 = n6589 & ~n6601 ;
  assign n6603 = ~n6600 & ~n6601 ;
  assign n6604 = ~n6602 & ~n6603 ;
  assign n6605 = ~n6223 & ~n6229 ;
  assign n6606 = n6604 & n6605 ;
  assign n6607 = ~n6604 & ~n6605 ;
  assign n6608 = ~n6606 & ~n6607 ;
  assign n6609 = ~x85 & n945 ;
  assign n6610 = ~x83 & n1099 ;
  assign n6611 = ~x84 & n940 ;
  assign n6612 = ~n6610 & ~n6611 ;
  assign n6613 = ~n6609 & n6612 ;
  assign n6614 = n948 & n3521 ;
  assign n6615 = n6613 & ~n6614 ;
  assign n6616 = ~x11 & ~n6615 ;
  assign n6617 = ~x11 & ~n6616 ;
  assign n6618 = ~n6615 & ~n6616 ;
  assign n6619 = ~n6617 & ~n6618 ;
  assign n6620 = n6608 & ~n6619 ;
  assign n6621 = n6608 & ~n6620 ;
  assign n6622 = ~n6619 & ~n6620 ;
  assign n6623 = ~n6621 & ~n6622 ;
  assign n6624 = ~n6247 & n6623 ;
  assign n6625 = n6247 & ~n6623 ;
  assign n6626 = ~n6624 & ~n6625 ;
  assign n6627 = ~x88 & n574 ;
  assign n6628 = ~x86 & n673 ;
  assign n6629 = ~x87 & n569 ;
  assign n6630 = ~n6628 & ~n6629 ;
  assign n6631 = ~n6627 & n6630 ;
  assign n6632 = n577 & n4457 ;
  assign n6633 = n6631 & ~n6632 ;
  assign n6634 = ~x8 & ~n6633 ;
  assign n6635 = ~x8 & ~n6634 ;
  assign n6636 = ~n6633 & ~n6634 ;
  assign n6637 = ~n6635 & ~n6636 ;
  assign n6638 = ~n6626 & ~n6637 ;
  assign n6639 = n6626 & n6637 ;
  assign n6640 = ~n6638 & ~n6639 ;
  assign n6641 = n6498 & ~n6640 ;
  assign n6642 = ~n6498 & n6640 ;
  assign n6643 = ~n6641 & ~n6642 ;
  assign n6644 = ~x91 & n293 ;
  assign n6645 = ~x89 & n373 ;
  assign n6646 = ~x90 & n288 ;
  assign n6647 = ~n6645 & ~n6646 ;
  assign n6648 = ~n6644 & n6647 ;
  assign n6649 = n296 & n5507 ;
  assign n6650 = n6648 & ~n6649 ;
  assign n6651 = ~x5 & ~n6650 ;
  assign n6652 = ~x5 & ~n6651 ;
  assign n6653 = ~n6650 & ~n6651 ;
  assign n6654 = ~n6652 & ~n6653 ;
  assign n6655 = n6643 & ~n6654 ;
  assign n6656 = n6643 & ~n6655 ;
  assign n6657 = ~n6654 & ~n6655 ;
  assign n6658 = ~n6656 & ~n6657 ;
  assign n6659 = ~n6269 & ~n6273 ;
  assign n6660 = n6658 & n6659 ;
  assign n6661 = ~n6658 & ~n6659 ;
  assign n6662 = ~n6660 & ~n6661 ;
  assign n6663 = ~x94 & n164 ;
  assign n6664 = ~x92 & n205 ;
  assign n6665 = ~x93 & n162 ;
  assign n6666 = ~n6664 & ~n6665 ;
  assign n6667 = ~n6663 & n6666 ;
  assign n6668 = ~n6089 & ~n6283 ;
  assign n6669 = n6480 & ~n6668 ;
  assign n6670 = ~n6480 & n6668 ;
  assign n6671 = ~n6669 & ~n6670 ;
  assign n6672 = n167 & n6671 ;
  assign n6673 = n6667 & ~n6672 ;
  assign n6674 = ~x2 & ~n6673 ;
  assign n6675 = ~x2 & ~n6674 ;
  assign n6676 = ~n6673 & ~n6674 ;
  assign n6677 = ~n6675 & ~n6676 ;
  assign n6678 = n6662 & ~n6677 ;
  assign n6679 = n6662 & ~n6678 ;
  assign n6680 = ~n6677 & ~n6678 ;
  assign n6681 = ~n6679 & ~n6680 ;
  assign n6682 = ~n6292 & ~n6297 ;
  assign n6683 = ~n6681 & ~n6682 ;
  assign n6684 = n6681 & n6682 ;
  assign n6685 = ~n6683 & ~n6684 ;
  assign n6688 = ~n6685 & ~x158 ;
  assign n6689 = ~n6687 & ~n6688 ;
  assign n6690 = ~n5973 & ~n6353 ;
  assign n6691 = ~n6350 & ~n6690 ;
  assign n6692 = x71 & n4531 ;
  assign n6693 = x69 & n4847 ;
  assign n6694 = x70 & n4526 ;
  assign n6695 = ~n6693 & ~n6694 ;
  assign n6696 = ~n6692 & n6695 ;
  assign n6697 = n558 & n4534 ;
  assign n6698 = n6696 & ~n6697 ;
  assign n6699 = x26 & ~n6698 ;
  assign n6700 = x26 & ~n6699 ;
  assign n6701 = ~n6698 & ~n6699 ;
  assign n6702 = ~n6700 & ~n6701 ;
  assign n6703 = n5955 & n6321 ;
  assign n6704 = ~n6336 & ~n6703 ;
  assign n6705 = x68 & n5560 ;
  assign n6706 = x66 & n5943 ;
  assign n6707 = x67 & n5555 ;
  assign n6708 = ~n6706 & ~n6707 ;
  assign n6709 = ~n6705 & n6708 ;
  assign n6710 = n317 & n5563 ;
  assign n6711 = n6709 & ~n6710 ;
  assign n6712 = x29 & ~n6711 ;
  assign n6713 = x29 & ~n6712 ;
  assign n6714 = ~n6711 & ~n6712 ;
  assign n6715 = ~n6713 & ~n6714 ;
  assign n6716 = x32 & ~n6321 ;
  assign n6717 = ~x30 & x31 ;
  assign n6718 = x30 & ~x31 ;
  assign n6719 = ~n6717 & ~n6718 ;
  assign n6720 = n6320 & ~n6719 ;
  assign n6721 = x64 & n6720 ;
  assign n6722 = ~x31 & x32 ;
  assign n6723 = x31 & ~x32 ;
  assign n6724 = ~n6722 & ~n6723 ;
  assign n6725 = ~n6320 & n6724 ;
  assign n6726 = x65 & n6725 ;
  assign n6727 = ~n6721 & ~n6726 ;
  assign n6728 = ~n6320 & ~n6724 ;
  assign n6729 = ~n152 & n6728 ;
  assign n6730 = n6727 & ~n6729 ;
  assign n6731 = x32 & ~n6730 ;
  assign n6732 = x32 & ~n6731 ;
  assign n6733 = ~n6730 & ~n6731 ;
  assign n6734 = ~n6732 & ~n6733 ;
  assign n6735 = n6716 & ~n6734 ;
  assign n6736 = ~n6716 & n6734 ;
  assign n6737 = ~n6735 & ~n6736 ;
  assign n6738 = n6715 & n6737 ;
  assign n6739 = ~n6715 & ~n6737 ;
  assign n6740 = ~n6738 & ~n6739 ;
  assign n6741 = ~n6704 & ~n6740 ;
  assign n6742 = n6704 & n6740 ;
  assign n6743 = ~n6741 & ~n6742 ;
  assign n6744 = ~n6702 & n6743 ;
  assign n6745 = n6702 & ~n6743 ;
  assign n6746 = ~n6744 & ~n6745 ;
  assign n6747 = ~n6691 & n6746 ;
  assign n6748 = n6691 & ~n6746 ;
  assign n6749 = ~n6747 & ~n6748 ;
  assign n6750 = x74 & n3589 ;
  assign n6751 = x72 & n3878 ;
  assign n6752 = x73 & n3584 ;
  assign n6753 = ~n6751 & ~n6752 ;
  assign n6754 = ~n6750 & n6753 ;
  assign n6755 = n994 & n3592 ;
  assign n6756 = n6754 & ~n6755 ;
  assign n6757 = x23 & ~n6756 ;
  assign n6758 = x23 & ~n6757 ;
  assign n6759 = ~n6756 & ~n6757 ;
  assign n6760 = ~n6758 & ~n6759 ;
  assign n6761 = n6749 & ~n6760 ;
  assign n6762 = n6749 & ~n6761 ;
  assign n6763 = ~n6760 & ~n6761 ;
  assign n6764 = ~n6762 & ~n6763 ;
  assign n6765 = ~n6368 & ~n6371 ;
  assign n6766 = n6764 & n6765 ;
  assign n6767 = ~n6764 & ~n6765 ;
  assign n6768 = ~n6766 & ~n6767 ;
  assign n6769 = x77 & n2751 ;
  assign n6770 = x75 & n3020 ;
  assign n6771 = x76 & n2746 ;
  assign n6772 = ~n6770 & ~n6771 ;
  assign n6773 = ~n6769 & n6772 ;
  assign n6774 = n1502 & n2754 ;
  assign n6775 = n6773 & ~n6774 ;
  assign n6776 = x20 & ~n6775 ;
  assign n6777 = x20 & ~n6776 ;
  assign n6778 = ~n6775 & ~n6776 ;
  assign n6779 = ~n6777 & ~n6778 ;
  assign n6780 = ~n6768 & n6779 ;
  assign n6781 = n6768 & ~n6779 ;
  assign n6782 = ~n6780 & ~n6781 ;
  assign n6783 = ~n6375 & ~n6377 ;
  assign n6784 = n6782 & ~n6783 ;
  assign n6785 = ~n6782 & n6783 ;
  assign n6786 = ~n6784 & ~n6785 ;
  assign n6787 = x80 & n2093 ;
  assign n6788 = x78 & n2275 ;
  assign n6789 = x79 & n2088 ;
  assign n6790 = ~n6788 & ~n6789 ;
  assign n6791 = ~n6787 & n6790 ;
  assign n6792 = n2028 & n2096 ;
  assign n6793 = n6791 & ~n6792 ;
  assign n6794 = x17 & ~n6793 ;
  assign n6795 = x17 & ~n6794 ;
  assign n6796 = ~n6793 & ~n6794 ;
  assign n6797 = ~n6795 & ~n6796 ;
  assign n6798 = n6786 & ~n6797 ;
  assign n6799 = n6786 & ~n6798 ;
  assign n6800 = ~n6797 & ~n6798 ;
  assign n6801 = ~n6799 & ~n6800 ;
  assign n6802 = ~n6391 & ~n6397 ;
  assign n6803 = n6801 & n6802 ;
  assign n6804 = ~n6801 & ~n6802 ;
  assign n6805 = ~n6803 & ~n6804 ;
  assign n6806 = x83 & n1434 ;
  assign n6807 = x81 & n1646 ;
  assign n6808 = x82 & n1429 ;
  assign n6809 = ~n6807 & ~n6808 ;
  assign n6810 = ~n6806 & n6809 ;
  assign n6811 = n1437 & n2843 ;
  assign n6812 = n6810 & ~n6811 ;
  assign n6813 = x14 & ~n6812 ;
  assign n6814 = x14 & ~n6813 ;
  assign n6815 = ~n6812 & ~n6813 ;
  assign n6816 = ~n6814 & ~n6815 ;
  assign n6817 = n6805 & ~n6816 ;
  assign n6818 = n6805 & ~n6817 ;
  assign n6819 = ~n6816 & ~n6817 ;
  assign n6820 = ~n6818 & ~n6819 ;
  assign n6821 = ~n6410 & ~n6416 ;
  assign n6822 = n6820 & n6821 ;
  assign n6823 = ~n6820 & ~n6821 ;
  assign n6824 = ~n6822 & ~n6823 ;
  assign n6825 = x86 & n945 ;
  assign n6826 = x84 & n1099 ;
  assign n6827 = x85 & n940 ;
  assign n6828 = ~n6826 & ~n6827 ;
  assign n6829 = ~n6825 & n6828 ;
  assign n6830 = n948 & n3686 ;
  assign n6831 = n6829 & ~n6830 ;
  assign n6832 = x11 & ~n6831 ;
  assign n6833 = x11 & ~n6832 ;
  assign n6834 = ~n6831 & ~n6832 ;
  assign n6835 = ~n6833 & ~n6834 ;
  assign n6836 = n6824 & ~n6835 ;
  assign n6837 = n6824 & ~n6836 ;
  assign n6838 = ~n6835 & ~n6836 ;
  assign n6839 = ~n6837 & ~n6838 ;
  assign n6840 = ~n6053 & ~n6432 ;
  assign n6841 = ~n6429 & ~n6840 ;
  assign n6842 = n6839 & n6841 ;
  assign n6843 = ~n6839 & ~n6841 ;
  assign n6844 = ~n6842 & ~n6843 ;
  assign n6845 = x89 & n574 ;
  assign n6846 = x87 & n673 ;
  assign n6847 = x88 & n569 ;
  assign n6848 = ~n6846 & ~n6847 ;
  assign n6849 = ~n6845 & n6848 ;
  assign n6850 = n577 & n4488 ;
  assign n6851 = n6849 & ~n6850 ;
  assign n6852 = x8 & ~n6851 ;
  assign n6853 = x8 & ~n6852 ;
  assign n6854 = ~n6851 & ~n6852 ;
  assign n6855 = ~n6853 & ~n6854 ;
  assign n6856 = n6844 & ~n6855 ;
  assign n6857 = n6844 & ~n6856 ;
  assign n6858 = ~n6855 & ~n6856 ;
  assign n6859 = ~n6857 & ~n6858 ;
  assign n6860 = ~n6447 & ~n6451 ;
  assign n6861 = n6859 & n6860 ;
  assign n6862 = ~n6859 & ~n6860 ;
  assign n6863 = ~n6861 & ~n6862 ;
  assign n6864 = x92 & n293 ;
  assign n6865 = x90 & n373 ;
  assign n6866 = x91 & n288 ;
  assign n6867 = ~n6865 & ~n6866 ;
  assign n6868 = ~n6864 & n6867 ;
  assign n6869 = n296 & n5710 ;
  assign n6870 = n6868 & ~n6869 ;
  assign n6871 = x5 & ~n6870 ;
  assign n6872 = x5 & ~n6871 ;
  assign n6873 = ~n6870 & ~n6871 ;
  assign n6874 = ~n6872 & ~n6873 ;
  assign n6875 = n6863 & ~n6874 ;
  assign n6876 = n6863 & ~n6875 ;
  assign n6877 = ~n6874 & ~n6875 ;
  assign n6878 = ~n6876 & ~n6877 ;
  assign n6879 = ~n6464 & ~n6470 ;
  assign n6880 = n6878 & n6879 ;
  assign n6881 = ~n6878 & ~n6879 ;
  assign n6882 = ~n6880 & ~n6881 ;
  assign n6883 = x95 & n146 ;
  assign n6884 = x93 & n182 ;
  assign n6885 = x94 & n141 ;
  assign n6886 = ~n6884 & ~n6885 ;
  assign n6887 = ~n6883 & n6886 ;
  assign n6888 = ~n6479 & ~n6481 ;
  assign n6889 = ~x94 & ~x95 ;
  assign n6890 = x94 & x95 ;
  assign n6891 = ~n6889 & ~n6890 ;
  assign n6892 = ~n6888 & n6891 ;
  assign n6893 = n6888 & ~n6891 ;
  assign n6894 = ~n6892 & ~n6893 ;
  assign n6895 = n149 & n6894 ;
  assign n6896 = n6887 & ~n6895 ;
  assign n6897 = x2 & ~n6896 ;
  assign n6898 = x2 & ~n6897 ;
  assign n6899 = ~n6896 & ~n6897 ;
  assign n6900 = ~n6898 & ~n6899 ;
  assign n6901 = n6882 & ~n6900 ;
  assign n6902 = n6882 & ~n6901 ;
  assign n6903 = ~n6900 & ~n6901 ;
  assign n6904 = ~n6902 & ~n6903 ;
  assign n6905 = ~n6490 & ~n6495 ;
  assign n6906 = ~n6904 & ~n6905 ;
  assign n6907 = n6904 & n6905 ;
  assign n6908 = ~n6906 & ~n6907 ;
  assign n7116 = n6908 & x159 ;
  assign n6909 = ~n6167 & ~n6544 ;
  assign n6910 = ~n6541 & ~n6909 ;
  assign n6911 = ~x71 & n4531 ;
  assign n6912 = ~x69 & n4847 ;
  assign n6913 = ~x70 & n4526 ;
  assign n6914 = ~n6912 & ~n6913 ;
  assign n6915 = ~n6911 & n6914 ;
  assign n6916 = n622 & n4534 ;
  assign n6917 = n6915 & ~n6916 ;
  assign n6918 = ~x26 & ~n6917 ;
  assign n6919 = ~x26 & ~n6918 ;
  assign n6920 = ~n6917 & ~n6918 ;
  assign n6921 = ~n6919 & ~n6920 ;
  assign n6922 = n6149 & n6512 ;
  assign n6923 = ~n6527 & ~n6922 ;
  assign n6924 = ~x68 & n5560 ;
  assign n6925 = ~x66 & n5943 ;
  assign n6926 = ~x67 & n5555 ;
  assign n6927 = ~n6925 & ~n6926 ;
  assign n6928 = ~n6924 & n6927 ;
  assign n6929 = n352 & n5563 ;
  assign n6930 = n6928 & ~n6929 ;
  assign n6931 = ~x29 & ~n6930 ;
  assign n6932 = ~x29 & ~n6931 ;
  assign n6933 = ~n6930 & ~n6931 ;
  assign n6934 = ~n6932 & ~n6933 ;
  assign n6935 = ~x32 & ~n6512 ;
  assign n6936 = ~x64 & n6720 ;
  assign n6937 = ~x65 & n6725 ;
  assign n6938 = ~n6936 & ~n6937 ;
  assign n6939 = ~n6729 & n6938 ;
  assign n6940 = ~x32 & ~n6939 ;
  assign n6941 = ~x32 & ~n6940 ;
  assign n6942 = ~n6939 & ~n6940 ;
  assign n6943 = ~n6941 & ~n6942 ;
  assign n6944 = n6935 & ~n6943 ;
  assign n6945 = ~n6935 & n6943 ;
  assign n6946 = ~n6944 & ~n6945 ;
  assign n6947 = n6934 & n6946 ;
  assign n6948 = ~n6934 & ~n6946 ;
  assign n6949 = ~n6947 & ~n6948 ;
  assign n6950 = ~n6923 & ~n6949 ;
  assign n6951 = n6923 & n6949 ;
  assign n6952 = ~n6950 & ~n6951 ;
  assign n6953 = ~n6921 & n6952 ;
  assign n6954 = n6921 & ~n6952 ;
  assign n6955 = ~n6953 & ~n6954 ;
  assign n6956 = ~n6910 & n6955 ;
  assign n6957 = n6910 & ~n6955 ;
  assign n6958 = ~n6956 & ~n6957 ;
  assign n6959 = ~x74 & n3589 ;
  assign n6960 = ~x72 & n3878 ;
  assign n6961 = ~x73 & n3584 ;
  assign n6962 = ~n6960 & ~n6961 ;
  assign n6963 = ~n6959 & n6962 ;
  assign n6964 = n1066 & n3592 ;
  assign n6965 = n6963 & ~n6964 ;
  assign n6966 = ~x23 & ~n6965 ;
  assign n6967 = ~x23 & ~n6966 ;
  assign n6968 = ~n6965 & ~n6966 ;
  assign n6969 = ~n6967 & ~n6968 ;
  assign n6970 = n6958 & ~n6969 ;
  assign n6971 = n6958 & ~n6970 ;
  assign n6972 = ~n6969 & ~n6970 ;
  assign n6973 = ~n6971 & ~n6972 ;
  assign n6974 = ~n6559 & ~n6562 ;
  assign n6975 = n6973 & n6974 ;
  assign n6976 = ~n6973 & ~n6974 ;
  assign n6977 = ~n6975 & ~n6976 ;
  assign n6978 = ~x77 & n2751 ;
  assign n6979 = ~x75 & n3020 ;
  assign n6980 = ~x76 & n2746 ;
  assign n6981 = ~n6979 & ~n6980 ;
  assign n6982 = ~n6978 & n6981 ;
  assign n6983 = n1594 & n2754 ;
  assign n6984 = n6982 & ~n6983 ;
  assign n6985 = ~x20 & ~n6984 ;
  assign n6986 = ~x20 & ~n6985 ;
  assign n6987 = ~n6984 & ~n6985 ;
  assign n6988 = ~n6986 & ~n6987 ;
  assign n6989 = ~n6977 & n6988 ;
  assign n6990 = n6977 & ~n6988 ;
  assign n6991 = ~n6989 & ~n6990 ;
  assign n6992 = ~n6566 & ~n6568 ;
  assign n6993 = n6991 & ~n6992 ;
  assign n6994 = ~n6991 & n6992 ;
  assign n6995 = ~n6993 & ~n6994 ;
  assign n6996 = ~x80 & n2093 ;
  assign n6997 = ~x78 & n2275 ;
  assign n6998 = ~x79 & n2088 ;
  assign n6999 = ~n6997 & ~n6998 ;
  assign n7000 = ~n6996 & n6999 ;
  assign n7001 = n2096 & n2145 ;
  assign n7002 = n7000 & ~n7001 ;
  assign n7003 = ~x17 & ~n7002 ;
  assign n7004 = ~x17 & ~n7003 ;
  assign n7005 = ~n7002 & ~n7003 ;
  assign n7006 = ~n7004 & ~n7005 ;
  assign n7007 = n6995 & ~n7006 ;
  assign n7008 = n6995 & ~n7007 ;
  assign n7009 = ~n7006 & ~n7007 ;
  assign n7010 = ~n7008 & ~n7009 ;
  assign n7011 = ~n6582 & ~n6588 ;
  assign n7012 = n7010 & n7011 ;
  assign n7013 = ~n7010 & ~n7011 ;
  assign n7014 = ~n7012 & ~n7013 ;
  assign n7015 = ~x83 & n1434 ;
  assign n7016 = ~x81 & n1646 ;
  assign n7017 = ~x82 & n1429 ;
  assign n7018 = ~n7016 & ~n7017 ;
  assign n7019 = ~n7015 & n7018 ;
  assign n7020 = n1437 & n2972 ;
  assign n7021 = n7019 & ~n7020 ;
  assign n7022 = ~x14 & ~n7021 ;
  assign n7023 = ~x14 & ~n7022 ;
  assign n7024 = ~n7021 & ~n7022 ;
  assign n7025 = ~n7023 & ~n7024 ;
  assign n7026 = n7014 & ~n7025 ;
  assign n7027 = n7014 & ~n7026 ;
  assign n7028 = ~n7025 & ~n7026 ;
  assign n7029 = ~n7027 & ~n7028 ;
  assign n7030 = ~n6601 & ~n6607 ;
  assign n7031 = n7029 & n7030 ;
  assign n7032 = ~n7029 & ~n7030 ;
  assign n7033 = ~n7031 & ~n7032 ;
  assign n7034 = ~x86 & n945 ;
  assign n7035 = ~x84 & n1099 ;
  assign n7036 = ~x85 & n940 ;
  assign n7037 = ~n7035 & ~n7036 ;
  assign n7038 = ~n7034 & n7037 ;
  assign n7039 = n948 & n3832 ;
  assign n7040 = n7038 & ~n7039 ;
  assign n7041 = ~x11 & ~n7040 ;
  assign n7042 = ~x11 & ~n7041 ;
  assign n7043 = ~n7040 & ~n7041 ;
  assign n7044 = ~n7042 & ~n7043 ;
  assign n7045 = n7033 & ~n7044 ;
  assign n7046 = n7033 & ~n7045 ;
  assign n7047 = ~n7044 & ~n7045 ;
  assign n7048 = ~n7046 & ~n7047 ;
  assign n7049 = ~n6247 & ~n6623 ;
  assign n7050 = ~n6620 & ~n7049 ;
  assign n7051 = n7048 & n7050 ;
  assign n7052 = ~n7048 & ~n7050 ;
  assign n7053 = ~n7051 & ~n7052 ;
  assign n7054 = ~x89 & n574 ;
  assign n7055 = ~x87 & n673 ;
  assign n7056 = ~x88 & n569 ;
  assign n7057 = ~n7055 & ~n7056 ;
  assign n7058 = ~n7054 & n7057 ;
  assign n7059 = n577 & n4664 ;
  assign n7060 = n7058 & ~n7059 ;
  assign n7061 = ~x8 & ~n7060 ;
  assign n7062 = ~x8 & ~n7061 ;
  assign n7063 = ~n7060 & ~n7061 ;
  assign n7064 = ~n7062 & ~n7063 ;
  assign n7065 = n7053 & ~n7064 ;
  assign n7066 = n7053 & ~n7065 ;
  assign n7067 = ~n7064 & ~n7065 ;
  assign n7068 = ~n7066 & ~n7067 ;
  assign n7069 = ~n6638 & ~n6642 ;
  assign n7070 = n7068 & n7069 ;
  assign n7071 = ~n7068 & ~n7069 ;
  assign n7072 = ~n7070 & ~n7071 ;
  assign n7073 = ~x92 & n293 ;
  assign n7074 = ~x90 & n373 ;
  assign n7075 = ~x91 & n288 ;
  assign n7076 = ~n7074 & ~n7075 ;
  assign n7077 = ~n7073 & n7076 ;
  assign n7078 = n296 & n5896 ;
  assign n7079 = n7077 & ~n7078 ;
  assign n7080 = ~x5 & ~n7079 ;
  assign n7081 = ~x5 & ~n7080 ;
  assign n7082 = ~n7079 & ~n7080 ;
  assign n7083 = ~n7081 & ~n7082 ;
  assign n7084 = n7072 & ~n7083 ;
  assign n7085 = n7072 & ~n7084 ;
  assign n7086 = ~n7083 & ~n7084 ;
  assign n7087 = ~n7085 & ~n7086 ;
  assign n7088 = ~n6655 & ~n6661 ;
  assign n7089 = n7087 & n7088 ;
  assign n7090 = ~n7087 & ~n7088 ;
  assign n7091 = ~n7089 & ~n7090 ;
  assign n7092 = ~x95 & n164 ;
  assign n7093 = ~x93 & n205 ;
  assign n7094 = ~x94 & n162 ;
  assign n7095 = ~n7093 & ~n7094 ;
  assign n7096 = ~n7092 & n7095 ;
  assign n7097 = ~n6478 & ~n6669 ;
  assign n7098 = n6891 & ~n7097 ;
  assign n7099 = ~n6891 & n7097 ;
  assign n7100 = ~n7098 & ~n7099 ;
  assign n7101 = n167 & n7100 ;
  assign n7102 = n7096 & ~n7101 ;
  assign n7103 = ~x2 & ~n7102 ;
  assign n7104 = ~x2 & ~n7103 ;
  assign n7105 = ~n7102 & ~n7103 ;
  assign n7106 = ~n7104 & ~n7105 ;
  assign n7107 = n7091 & ~n7106 ;
  assign n7108 = n7091 & ~n7107 ;
  assign n7109 = ~n7106 & ~n7107 ;
  assign n7110 = ~n7108 & ~n7109 ;
  assign n7111 = ~n6678 & ~n6683 ;
  assign n7112 = ~n7110 & ~n7111 ;
  assign n7113 = n7110 & n7111 ;
  assign n7114 = ~n7112 & ~n7113 ;
  assign n7117 = ~n7114 & ~x159 ;
  assign n7118 = ~n7116 & ~n7117 ;
  assign n7119 = ~n6901 & ~n6906 ;
  assign n7120 = ~n6875 & ~n6881 ;
  assign n7121 = ~n6836 & ~n6843 ;
  assign n7122 = ~n6817 & ~n6823 ;
  assign n7123 = ~n6781 & ~n6784 ;
  assign n7124 = ~n6761 & ~n6767 ;
  assign n7125 = ~n6715 & n6737 ;
  assign n7126 = ~n6741 & ~n7125 ;
  assign n7127 = x66 & n6725 ;
  assign n7128 = n6320 & ~n6724 ;
  assign n7129 = n6719 & n7128 ;
  assign n7130 = x64 & n7129 ;
  assign n7131 = x65 & n6720 ;
  assign n7132 = ~n7130 & ~n7131 ;
  assign n7133 = ~n7127 & n7132 ;
  assign n7134 = n194 & n6728 ;
  assign n7135 = n7133 & ~n7134 ;
  assign n7136 = x32 & ~n7135 ;
  assign n7137 = x32 & ~n7136 ;
  assign n7138 = ~n7135 & ~n7136 ;
  assign n7139 = ~n7137 & ~n7138 ;
  assign n7140 = ~n6735 & n7139 ;
  assign n7141 = n6735 & ~n7139 ;
  assign n7142 = ~n7140 & ~n7141 ;
  assign n7143 = x69 & n5560 ;
  assign n7144 = x67 & n5943 ;
  assign n7145 = x68 & n5555 ;
  assign n7146 = ~n7144 & ~n7145 ;
  assign n7147 = ~n7143 & n7146 ;
  assign n7148 = n398 & n5563 ;
  assign n7149 = n7147 & ~n7148 ;
  assign n7150 = x29 & ~n7149 ;
  assign n7151 = x29 & ~n7150 ;
  assign n7152 = ~n7149 & ~n7150 ;
  assign n7153 = ~n7151 & ~n7152 ;
  assign n7154 = n7142 & ~n7153 ;
  assign n7155 = ~n7142 & n7153 ;
  assign n7156 = ~n7126 & ~n7155 ;
  assign n7157 = ~n7154 & n7156 ;
  assign n7158 = ~n7126 & ~n7157 ;
  assign n7159 = ~n7154 & ~n7157 ;
  assign n7160 = ~n7155 & n7159 ;
  assign n7161 = ~n7158 & ~n7160 ;
  assign n7162 = x72 & n4531 ;
  assign n7163 = x70 & n4847 ;
  assign n7164 = x71 & n4526 ;
  assign n7165 = ~n7163 & ~n7164 ;
  assign n7166 = ~n7162 & n7165 ;
  assign n7167 = n717 & n4534 ;
  assign n7168 = n7166 & ~n7167 ;
  assign n7169 = x26 & ~n7168 ;
  assign n7170 = x26 & ~n7169 ;
  assign n7171 = ~n7168 & ~n7169 ;
  assign n7172 = ~n7170 & ~n7171 ;
  assign n7173 = ~n7161 & ~n7172 ;
  assign n7174 = ~n7161 & ~n7173 ;
  assign n7175 = ~n7172 & ~n7173 ;
  assign n7176 = ~n7174 & ~n7175 ;
  assign n7177 = ~n6744 & ~n6747 ;
  assign n7178 = n7176 & n7177 ;
  assign n7179 = ~n7176 & ~n7177 ;
  assign n7180 = ~n7178 & ~n7179 ;
  assign n7181 = x75 & n3589 ;
  assign n7182 = x73 & n3878 ;
  assign n7183 = x74 & n3584 ;
  assign n7184 = ~n7182 & ~n7183 ;
  assign n7185 = ~n7181 & n7184 ;
  assign n7186 = n1150 & n3592 ;
  assign n7187 = n7185 & ~n7186 ;
  assign n7188 = x23 & ~n7187 ;
  assign n7189 = x23 & ~n7188 ;
  assign n7190 = ~n7187 & ~n7188 ;
  assign n7191 = ~n7189 & ~n7190 ;
  assign n7192 = n7180 & ~n7191 ;
  assign n7193 = ~n7180 & n7191 ;
  assign n7194 = ~n7124 & ~n7193 ;
  assign n7195 = ~n7192 & n7194 ;
  assign n7196 = ~n7124 & ~n7195 ;
  assign n7197 = ~n7192 & ~n7195 ;
  assign n7198 = ~n7193 & n7197 ;
  assign n7199 = ~n7196 & ~n7198 ;
  assign n7200 = x78 & n2751 ;
  assign n7201 = x76 & n3020 ;
  assign n7202 = x77 & n2746 ;
  assign n7203 = ~n7201 & ~n7202 ;
  assign n7204 = ~n7200 & n7203 ;
  assign n7205 = n1624 & n2754 ;
  assign n7206 = n7204 & ~n7205 ;
  assign n7207 = x20 & ~n7206 ;
  assign n7208 = x20 & ~n7207 ;
  assign n7209 = ~n7206 & ~n7207 ;
  assign n7210 = ~n7208 & ~n7209 ;
  assign n7211 = n7199 & n7210 ;
  assign n7212 = ~n7199 & ~n7210 ;
  assign n7213 = ~n7211 & ~n7212 ;
  assign n7214 = ~n7123 & n7213 ;
  assign n7215 = n7123 & ~n7213 ;
  assign n7216 = ~n7214 & ~n7215 ;
  assign n7217 = x81 & n2093 ;
  assign n7218 = x79 & n2275 ;
  assign n7219 = x80 & n2088 ;
  assign n7220 = ~n7218 & ~n7219 ;
  assign n7221 = ~n7217 & n7220 ;
  assign n7222 = n2096 & n2348 ;
  assign n7223 = n7221 & ~n7222 ;
  assign n7224 = x17 & ~n7223 ;
  assign n7225 = x17 & ~n7224 ;
  assign n7226 = ~n7223 & ~n7224 ;
  assign n7227 = ~n7225 & ~n7226 ;
  assign n7228 = n7216 & ~n7227 ;
  assign n7229 = n7216 & ~n7228 ;
  assign n7230 = ~n7227 & ~n7228 ;
  assign n7231 = ~n7229 & ~n7230 ;
  assign n7232 = ~n6798 & ~n6804 ;
  assign n7233 = n7231 & n7232 ;
  assign n7234 = ~n7231 & ~n7232 ;
  assign n7235 = ~n7233 & ~n7234 ;
  assign n7236 = x84 & n1434 ;
  assign n7237 = x82 & n1646 ;
  assign n7238 = x83 & n1429 ;
  assign n7239 = ~n7237 & ~n7238 ;
  assign n7240 = ~n7236 & n7239 ;
  assign n7241 = n1437 & n3114 ;
  assign n7242 = n7240 & ~n7241 ;
  assign n7243 = x14 & ~n7242 ;
  assign n7244 = x14 & ~n7243 ;
  assign n7245 = ~n7242 & ~n7243 ;
  assign n7246 = ~n7244 & ~n7245 ;
  assign n7247 = n7235 & ~n7246 ;
  assign n7248 = ~n7235 & n7246 ;
  assign n7249 = ~n7122 & ~n7248 ;
  assign n7250 = ~n7247 & n7249 ;
  assign n7251 = ~n7122 & ~n7250 ;
  assign n7252 = ~n7247 & ~n7250 ;
  assign n7253 = ~n7248 & n7252 ;
  assign n7254 = ~n7251 & ~n7253 ;
  assign n7255 = x87 & n945 ;
  assign n7256 = x85 & n1099 ;
  assign n7257 = x86 & n940 ;
  assign n7258 = ~n7256 & ~n7257 ;
  assign n7259 = ~n7255 & n7258 ;
  assign n7260 = n948 & n3991 ;
  assign n7261 = n7259 & ~n7260 ;
  assign n7262 = x11 & ~n7261 ;
  assign n7263 = x11 & ~n7262 ;
  assign n7264 = ~n7261 & ~n7262 ;
  assign n7265 = ~n7263 & ~n7264 ;
  assign n7266 = n7254 & n7265 ;
  assign n7267 = ~n7254 & ~n7265 ;
  assign n7268 = ~n7266 & ~n7267 ;
  assign n7269 = ~n7121 & n7268 ;
  assign n7270 = n7121 & ~n7268 ;
  assign n7271 = ~n7269 & ~n7270 ;
  assign n7272 = x90 & n574 ;
  assign n7273 = x88 & n673 ;
  assign n7274 = x89 & n569 ;
  assign n7275 = ~n7273 & ~n7274 ;
  assign n7276 = ~n7272 & n7275 ;
  assign n7277 = n577 & n4986 ;
  assign n7278 = n7276 & ~n7277 ;
  assign n7279 = x8 & ~n7278 ;
  assign n7280 = x8 & ~n7279 ;
  assign n7281 = ~n7278 & ~n7279 ;
  assign n7282 = ~n7280 & ~n7281 ;
  assign n7283 = n7271 & ~n7282 ;
  assign n7284 = n7271 & ~n7283 ;
  assign n7285 = ~n7282 & ~n7283 ;
  assign n7286 = ~n7284 & ~n7285 ;
  assign n7287 = ~n6856 & ~n6862 ;
  assign n7288 = n7286 & n7287 ;
  assign n7289 = ~n7286 & ~n7287 ;
  assign n7290 = ~n7288 & ~n7289 ;
  assign n7291 = x93 & n293 ;
  assign n7292 = x91 & n373 ;
  assign n7293 = x92 & n288 ;
  assign n7294 = ~n7292 & ~n7293 ;
  assign n7295 = ~n7291 & n7294 ;
  assign n7296 = n296 & n6094 ;
  assign n7297 = n7295 & ~n7296 ;
  assign n7298 = x5 & ~n7297 ;
  assign n7299 = x5 & ~n7298 ;
  assign n7300 = ~n7297 & ~n7298 ;
  assign n7301 = ~n7299 & ~n7300 ;
  assign n7302 = n7290 & ~n7301 ;
  assign n7303 = ~n7290 & n7301 ;
  assign n7304 = ~n7120 & ~n7303 ;
  assign n7305 = ~n7302 & n7304 ;
  assign n7306 = ~n7120 & ~n7305 ;
  assign n7307 = ~n7302 & ~n7305 ;
  assign n7308 = ~n7303 & n7307 ;
  assign n7309 = ~n7306 & ~n7308 ;
  assign n7310 = x96 & n146 ;
  assign n7311 = x94 & n182 ;
  assign n7312 = x95 & n141 ;
  assign n7313 = ~n7311 & ~n7312 ;
  assign n7314 = ~n7310 & n7313 ;
  assign n7315 = ~n6890 & ~n6892 ;
  assign n7316 = ~x95 & ~x96 ;
  assign n7317 = x95 & x96 ;
  assign n7318 = ~n7316 & ~n7317 ;
  assign n7319 = ~n7315 & n7318 ;
  assign n7320 = n7315 & ~n7318 ;
  assign n7321 = ~n7319 & ~n7320 ;
  assign n7322 = n149 & n7321 ;
  assign n7323 = n7314 & ~n7322 ;
  assign n7324 = x2 & ~n7323 ;
  assign n7325 = x2 & ~n7324 ;
  assign n7326 = ~n7323 & ~n7324 ;
  assign n7327 = ~n7325 & ~n7326 ;
  assign n7328 = ~n7309 & n7327 ;
  assign n7329 = n7309 & ~n7327 ;
  assign n7330 = ~n7328 & ~n7329 ;
  assign n7331 = ~n7119 & ~n7330 ;
  assign n7332 = n7119 & n7330 ;
  assign n7333 = ~n7331 & ~n7332 ;
  assign n7545 = n7333 & x160 ;
  assign n7334 = ~n7107 & ~n7112 ;
  assign n7335 = ~n7084 & ~n7090 ;
  assign n7336 = ~n7045 & ~n7052 ;
  assign n7337 = ~n7026 & ~n7032 ;
  assign n7338 = ~n6990 & ~n6993 ;
  assign n7339 = ~n6970 & ~n6976 ;
  assign n7340 = ~n6934 & n6946 ;
  assign n7341 = ~n6950 & ~n7340 ;
  assign n7342 = ~x66 & n6725 ;
  assign n7343 = ~x64 & n7129 ;
  assign n7344 = ~x65 & n6720 ;
  assign n7345 = ~n7343 & ~n7344 ;
  assign n7346 = ~n7342 & n7345 ;
  assign n7347 = n214 & n6728 ;
  assign n7348 = n7346 & ~n7347 ;
  assign n7349 = ~x32 & ~n7348 ;
  assign n7350 = ~x32 & ~n7349 ;
  assign n7351 = ~n7348 & ~n7349 ;
  assign n7352 = ~n7350 & ~n7351 ;
  assign n7353 = ~n6944 & n7352 ;
  assign n7354 = n6944 & ~n7352 ;
  assign n7355 = ~n7353 & ~n7354 ;
  assign n7356 = ~x69 & n5560 ;
  assign n7357 = ~x67 & n5943 ;
  assign n7358 = ~x68 & n5555 ;
  assign n7359 = ~n7357 & ~n7358 ;
  assign n7360 = ~n7356 & n7359 ;
  assign n7361 = n435 & n5563 ;
  assign n7362 = n7360 & ~n7361 ;
  assign n7363 = ~x29 & ~n7362 ;
  assign n7364 = ~x29 & ~n7363 ;
  assign n7365 = ~n7362 & ~n7363 ;
  assign n7366 = ~n7364 & ~n7365 ;
  assign n7367 = n7355 & ~n7366 ;
  assign n7368 = ~n7355 & n7366 ;
  assign n7369 = ~n7341 & ~n7368 ;
  assign n7370 = ~n7367 & n7369 ;
  assign n7371 = ~n7341 & ~n7370 ;
  assign n7372 = ~n7367 & ~n7370 ;
  assign n7373 = ~n7368 & n7372 ;
  assign n7374 = ~n7371 & ~n7373 ;
  assign n7375 = ~x72 & n4531 ;
  assign n7376 = ~x70 & n4847 ;
  assign n7377 = ~x71 & n4526 ;
  assign n7378 = ~n7376 & ~n7377 ;
  assign n7379 = ~n7375 & n7378 ;
  assign n7380 = n773 & n4534 ;
  assign n7381 = n7379 & ~n7380 ;
  assign n7382 = ~x26 & ~n7381 ;
  assign n7383 = ~x26 & ~n7382 ;
  assign n7384 = ~n7381 & ~n7382 ;
  assign n7385 = ~n7383 & ~n7384 ;
  assign n7386 = ~n7374 & ~n7385 ;
  assign n7387 = ~n7374 & ~n7386 ;
  assign n7388 = ~n7385 & ~n7386 ;
  assign n7389 = ~n7387 & ~n7388 ;
  assign n7390 = ~n6953 & ~n6956 ;
  assign n7391 = n7389 & n7390 ;
  assign n7392 = ~n7389 & ~n7390 ;
  assign n7393 = ~n7391 & ~n7392 ;
  assign n7394 = ~x75 & n3589 ;
  assign n7395 = ~x73 & n3878 ;
  assign n7396 = ~x74 & n3584 ;
  assign n7397 = ~n7395 & ~n7396 ;
  assign n7398 = ~n7394 & n7397 ;
  assign n7399 = n1225 & n3592 ;
  assign n7400 = n7398 & ~n7399 ;
  assign n7401 = ~x23 & ~n7400 ;
  assign n7402 = ~x23 & ~n7401 ;
  assign n7403 = ~n7400 & ~n7401 ;
  assign n7404 = ~n7402 & ~n7403 ;
  assign n7405 = n7393 & ~n7404 ;
  assign n7406 = ~n7393 & n7404 ;
  assign n7407 = ~n7339 & ~n7406 ;
  assign n7408 = ~n7405 & n7407 ;
  assign n7409 = ~n7339 & ~n7408 ;
  assign n7410 = ~n7405 & ~n7408 ;
  assign n7411 = ~n7406 & n7410 ;
  assign n7412 = ~n7409 & ~n7411 ;
  assign n7413 = ~x78 & n2751 ;
  assign n7414 = ~x76 & n3020 ;
  assign n7415 = ~x77 & n2746 ;
  assign n7416 = ~n7414 & ~n7415 ;
  assign n7417 = ~n7413 & n7416 ;
  assign n7418 = n1718 & n2754 ;
  assign n7419 = n7417 & ~n7418 ;
  assign n7420 = ~x20 & ~n7419 ;
  assign n7421 = ~x20 & ~n7420 ;
  assign n7422 = ~n7419 & ~n7420 ;
  assign n7423 = ~n7421 & ~n7422 ;
  assign n7424 = n7412 & n7423 ;
  assign n7425 = ~n7412 & ~n7423 ;
  assign n7426 = ~n7424 & ~n7425 ;
  assign n7427 = ~n7338 & n7426 ;
  assign n7428 = n7338 & ~n7426 ;
  assign n7429 = ~n7427 & ~n7428 ;
  assign n7430 = ~x81 & n2093 ;
  assign n7431 = ~x79 & n2275 ;
  assign n7432 = ~x80 & n2088 ;
  assign n7433 = ~n7431 & ~n7432 ;
  assign n7434 = ~n7430 & n7433 ;
  assign n7435 = n2096 & n2460 ;
  assign n7436 = n7434 & ~n7435 ;
  assign n7437 = ~x17 & ~n7436 ;
  assign n7438 = ~x17 & ~n7437 ;
  assign n7439 = ~n7436 & ~n7437 ;
  assign n7440 = ~n7438 & ~n7439 ;
  assign n7441 = n7429 & ~n7440 ;
  assign n7442 = n7429 & ~n7441 ;
  assign n7443 = ~n7440 & ~n7441 ;
  assign n7444 = ~n7442 & ~n7443 ;
  assign n7445 = ~n7007 & ~n7013 ;
  assign n7446 = n7444 & n7445 ;
  assign n7447 = ~n7444 & ~n7445 ;
  assign n7448 = ~n7446 & ~n7447 ;
  assign n7449 = ~x84 & n1434 ;
  assign n7450 = ~x82 & n1646 ;
  assign n7451 = ~x83 & n1429 ;
  assign n7452 = ~n7450 & ~n7451 ;
  assign n7453 = ~n7449 & n7452 ;
  assign n7454 = n1437 & n3247 ;
  assign n7455 = n7453 & ~n7454 ;
  assign n7456 = ~x14 & ~n7455 ;
  assign n7457 = ~x14 & ~n7456 ;
  assign n7458 = ~n7455 & ~n7456 ;
  assign n7459 = ~n7457 & ~n7458 ;
  assign n7460 = n7448 & ~n7459 ;
  assign n7461 = ~n7448 & n7459 ;
  assign n7462 = ~n7337 & ~n7461 ;
  assign n7463 = ~n7460 & n7462 ;
  assign n7464 = ~n7337 & ~n7463 ;
  assign n7465 = ~n7460 & ~n7463 ;
  assign n7466 = ~n7461 & n7465 ;
  assign n7467 = ~n7464 & ~n7466 ;
  assign n7468 = ~x87 & n945 ;
  assign n7469 = ~x85 & n1099 ;
  assign n7470 = ~x86 & n940 ;
  assign n7471 = ~n7469 & ~n7470 ;
  assign n7472 = ~n7468 & n7471 ;
  assign n7473 = n948 & n4143 ;
  assign n7474 = n7472 & ~n7473 ;
  assign n7475 = ~x11 & ~n7474 ;
  assign n7476 = ~x11 & ~n7475 ;
  assign n7477 = ~n7474 & ~n7475 ;
  assign n7478 = ~n7476 & ~n7477 ;
  assign n7479 = n7467 & n7478 ;
  assign n7480 = ~n7467 & ~n7478 ;
  assign n7481 = ~n7479 & ~n7480 ;
  assign n7482 = ~n7336 & n7481 ;
  assign n7483 = n7336 & ~n7481 ;
  assign n7484 = ~n7482 & ~n7483 ;
  assign n7485 = ~x90 & n574 ;
  assign n7486 = ~x88 & n673 ;
  assign n7487 = ~x89 & n569 ;
  assign n7488 = ~n7486 & ~n7487 ;
  assign n7489 = ~n7485 & n7488 ;
  assign n7490 = n577 & n5155 ;
  assign n7491 = n7489 & ~n7490 ;
  assign n7492 = ~x8 & ~n7491 ;
  assign n7493 = ~x8 & ~n7492 ;
  assign n7494 = ~n7491 & ~n7492 ;
  assign n7495 = ~n7493 & ~n7494 ;
  assign n7496 = n7484 & ~n7495 ;
  assign n7497 = n7484 & ~n7496 ;
  assign n7498 = ~n7495 & ~n7496 ;
  assign n7499 = ~n7497 & ~n7498 ;
  assign n7500 = ~n7065 & ~n7071 ;
  assign n7501 = n7499 & n7500 ;
  assign n7502 = ~n7499 & ~n7500 ;
  assign n7503 = ~n7501 & ~n7502 ;
  assign n7504 = ~x93 & n293 ;
  assign n7505 = ~x91 & n373 ;
  assign n7506 = ~x92 & n288 ;
  assign n7507 = ~n7505 & ~n7506 ;
  assign n7508 = ~n7504 & n7507 ;
  assign n7509 = n296 & n6285 ;
  assign n7510 = n7508 & ~n7509 ;
  assign n7511 = ~x5 & ~n7510 ;
  assign n7512 = ~x5 & ~n7511 ;
  assign n7513 = ~n7510 & ~n7511 ;
  assign n7514 = ~n7512 & ~n7513 ;
  assign n7515 = n7503 & ~n7514 ;
  assign n7516 = ~n7503 & n7514 ;
  assign n7517 = ~n7335 & ~n7516 ;
  assign n7518 = ~n7515 & n7517 ;
  assign n7519 = ~n7335 & ~n7518 ;
  assign n7520 = ~n7515 & ~n7518 ;
  assign n7521 = ~n7516 & n7520 ;
  assign n7522 = ~n7519 & ~n7521 ;
  assign n7523 = ~x96 & n164 ;
  assign n7524 = ~x94 & n205 ;
  assign n7525 = ~x95 & n162 ;
  assign n7526 = ~n7524 & ~n7525 ;
  assign n7527 = ~n7523 & n7526 ;
  assign n7528 = ~n6889 & ~n7098 ;
  assign n7529 = n7318 & ~n7528 ;
  assign n7530 = ~n7318 & n7528 ;
  assign n7531 = ~n7529 & ~n7530 ;
  assign n7532 = n167 & n7531 ;
  assign n7533 = n7527 & ~n7532 ;
  assign n7534 = ~x2 & ~n7533 ;
  assign n7535 = ~x2 & ~n7534 ;
  assign n7536 = ~n7533 & ~n7534 ;
  assign n7537 = ~n7535 & ~n7536 ;
  assign n7538 = ~n7522 & n7537 ;
  assign n7539 = n7522 & ~n7537 ;
  assign n7540 = ~n7538 & ~n7539 ;
  assign n7541 = ~n7334 & ~n7540 ;
  assign n7542 = n7334 & n7540 ;
  assign n7543 = ~n7541 & ~n7542 ;
  assign n7546 = ~n7543 & ~x160 ;
  assign n7547 = ~n7545 & ~n7546 ;
  assign n7548 = ~n7309 & ~n7327 ;
  assign n7549 = ~n7331 & ~n7548 ;
  assign n7550 = ~n7267 & ~n7269 ;
  assign n7551 = ~n7228 & ~n7234 ;
  assign n7552 = ~n7212 & ~n7214 ;
  assign n7553 = ~n7173 & ~n7179 ;
  assign n7554 = x32 & ~x33 ;
  assign n7555 = ~x32 & x33 ;
  assign n7556 = ~n7554 & ~n7555 ;
  assign n7557 = x64 & ~n7556 ;
  assign n7558 = ~n7141 & n7557 ;
  assign n7559 = n7141 & ~n7557 ;
  assign n7560 = ~n7558 & ~n7559 ;
  assign n7561 = x67 & n6725 ;
  assign n7562 = x65 & n7129 ;
  assign n7563 = x66 & n6720 ;
  assign n7564 = ~n7562 & ~n7563 ;
  assign n7565 = ~n7561 & n7564 ;
  assign n7566 = n240 & n6728 ;
  assign n7567 = n7565 & ~n7566 ;
  assign n7568 = x32 & ~n7567 ;
  assign n7569 = x32 & ~n7568 ;
  assign n7570 = ~n7567 & ~n7568 ;
  assign n7571 = ~n7569 & ~n7570 ;
  assign n7572 = ~n7560 & ~n7571 ;
  assign n7573 = n7560 & n7571 ;
  assign n7574 = ~n7572 & ~n7573 ;
  assign n7575 = x70 & n5560 ;
  assign n7576 = x68 & n5943 ;
  assign n7577 = x69 & n5555 ;
  assign n7578 = ~n7576 & ~n7577 ;
  assign n7579 = ~n7575 & n7578 ;
  assign n7580 = n488 & n5563 ;
  assign n7581 = n7579 & ~n7580 ;
  assign n7582 = x29 & ~n7581 ;
  assign n7583 = x29 & ~n7582 ;
  assign n7584 = ~n7581 & ~n7582 ;
  assign n7585 = ~n7583 & ~n7584 ;
  assign n7586 = n7574 & ~n7585 ;
  assign n7587 = n7574 & ~n7586 ;
  assign n7588 = ~n7585 & ~n7586 ;
  assign n7589 = ~n7587 & ~n7588 ;
  assign n7590 = ~n7159 & n7589 ;
  assign n7591 = n7159 & ~n7589 ;
  assign n7592 = ~n7590 & ~n7591 ;
  assign n7593 = x73 & n4531 ;
  assign n7594 = x71 & n4847 ;
  assign n7595 = x72 & n4526 ;
  assign n7596 = ~n7594 & ~n7595 ;
  assign n7597 = ~n7593 & n7596 ;
  assign n7598 = n843 & n4534 ;
  assign n7599 = n7597 & ~n7598 ;
  assign n7600 = x26 & ~n7599 ;
  assign n7601 = x26 & ~n7600 ;
  assign n7602 = ~n7599 & ~n7600 ;
  assign n7603 = ~n7601 & ~n7602 ;
  assign n7604 = ~n7592 & ~n7603 ;
  assign n7605 = n7592 & n7603 ;
  assign n7606 = ~n7604 & ~n7605 ;
  assign n7607 = n7553 & ~n7606 ;
  assign n7608 = ~n7553 & n7606 ;
  assign n7609 = ~n7607 & ~n7608 ;
  assign n7610 = x76 & n3589 ;
  assign n7611 = x74 & n3878 ;
  assign n7612 = x75 & n3584 ;
  assign n7613 = ~n7611 & ~n7612 ;
  assign n7614 = ~n7610 & n7613 ;
  assign n7615 = n1311 & n3592 ;
  assign n7616 = n7614 & ~n7615 ;
  assign n7617 = x23 & ~n7616 ;
  assign n7618 = x23 & ~n7617 ;
  assign n7619 = ~n7616 & ~n7617 ;
  assign n7620 = ~n7618 & ~n7619 ;
  assign n7621 = ~n7609 & n7620 ;
  assign n7622 = n7609 & ~n7620 ;
  assign n7623 = ~n7621 & ~n7622 ;
  assign n7624 = ~n7197 & n7623 ;
  assign n7625 = n7197 & ~n7623 ;
  assign n7626 = ~n7624 & ~n7625 ;
  assign n7627 = x79 & n2751 ;
  assign n7628 = x77 & n3020 ;
  assign n7629 = x78 & n2746 ;
  assign n7630 = ~n7628 & ~n7629 ;
  assign n7631 = ~n7627 & n7630 ;
  assign n7632 = n1817 & n2754 ;
  assign n7633 = n7631 & ~n7632 ;
  assign n7634 = x20 & ~n7633 ;
  assign n7635 = x20 & ~n7634 ;
  assign n7636 = ~n7633 & ~n7634 ;
  assign n7637 = ~n7635 & ~n7636 ;
  assign n7638 = n7626 & ~n7637 ;
  assign n7639 = n7626 & ~n7638 ;
  assign n7640 = ~n7637 & ~n7638 ;
  assign n7641 = ~n7639 & ~n7640 ;
  assign n7642 = ~n7552 & n7641 ;
  assign n7643 = n7552 & ~n7641 ;
  assign n7644 = ~n7642 & ~n7643 ;
  assign n7645 = x82 & n2093 ;
  assign n7646 = x80 & n2275 ;
  assign n7647 = x81 & n2088 ;
  assign n7648 = ~n7646 & ~n7647 ;
  assign n7649 = ~n7645 & n7648 ;
  assign n7650 = n2096 & n2584 ;
  assign n7651 = n7649 & ~n7650 ;
  assign n7652 = x17 & ~n7651 ;
  assign n7653 = x17 & ~n7652 ;
  assign n7654 = ~n7651 & ~n7652 ;
  assign n7655 = ~n7653 & ~n7654 ;
  assign n7656 = ~n7644 & ~n7655 ;
  assign n7657 = n7644 & n7655 ;
  assign n7658 = ~n7656 & ~n7657 ;
  assign n7659 = n7551 & ~n7658 ;
  assign n7660 = ~n7551 & n7658 ;
  assign n7661 = ~n7659 & ~n7660 ;
  assign n7662 = x85 & n1434 ;
  assign n7663 = x83 & n1646 ;
  assign n7664 = x84 & n1429 ;
  assign n7665 = ~n7663 & ~n7664 ;
  assign n7666 = ~n7662 & n7665 ;
  assign n7667 = n1437 & n3389 ;
  assign n7668 = n7666 & ~n7667 ;
  assign n7669 = x14 & ~n7668 ;
  assign n7670 = x14 & ~n7669 ;
  assign n7671 = ~n7668 & ~n7669 ;
  assign n7672 = ~n7670 & ~n7671 ;
  assign n7673 = n7661 & ~n7672 ;
  assign n7674 = n7661 & ~n7673 ;
  assign n7675 = ~n7672 & ~n7673 ;
  assign n7676 = ~n7674 & ~n7675 ;
  assign n7677 = ~n7252 & n7676 ;
  assign n7678 = n7252 & ~n7676 ;
  assign n7679 = ~n7677 & ~n7678 ;
  assign n7680 = x88 & n945 ;
  assign n7681 = x86 & n1099 ;
  assign n7682 = x87 & n940 ;
  assign n7683 = ~n7681 & ~n7682 ;
  assign n7684 = ~n7680 & n7683 ;
  assign n7685 = n948 & n4305 ;
  assign n7686 = n7684 & ~n7685 ;
  assign n7687 = x11 & ~n7686 ;
  assign n7688 = x11 & ~n7687 ;
  assign n7689 = ~n7686 & ~n7687 ;
  assign n7690 = ~n7688 & ~n7689 ;
  assign n7691 = n7679 & n7690 ;
  assign n7692 = ~n7679 & ~n7690 ;
  assign n7693 = ~n7691 & ~n7692 ;
  assign n7694 = ~n7550 & n7693 ;
  assign n7695 = n7550 & ~n7693 ;
  assign n7696 = ~n7694 & ~n7695 ;
  assign n7697 = x91 & n574 ;
  assign n7698 = x89 & n673 ;
  assign n7699 = x90 & n569 ;
  assign n7700 = ~n7698 & ~n7699 ;
  assign n7701 = ~n7697 & n7700 ;
  assign n7702 = n577 & n5336 ;
  assign n7703 = n7701 & ~n7702 ;
  assign n7704 = x8 & ~n7703 ;
  assign n7705 = x8 & ~n7704 ;
  assign n7706 = ~n7703 & ~n7704 ;
  assign n7707 = ~n7705 & ~n7706 ;
  assign n7708 = n7696 & ~n7707 ;
  assign n7709 = n7696 & ~n7708 ;
  assign n7710 = ~n7707 & ~n7708 ;
  assign n7711 = ~n7709 & ~n7710 ;
  assign n7712 = ~n7283 & ~n7289 ;
  assign n7713 = n7711 & n7712 ;
  assign n7714 = ~n7711 & ~n7712 ;
  assign n7715 = ~n7713 & ~n7714 ;
  assign n7716 = x94 & n293 ;
  assign n7717 = x92 & n373 ;
  assign n7718 = x93 & n288 ;
  assign n7719 = ~n7717 & ~n7718 ;
  assign n7720 = ~n7716 & n7719 ;
  assign n7721 = n296 & n6483 ;
  assign n7722 = n7720 & ~n7721 ;
  assign n7723 = x5 & ~n7722 ;
  assign n7724 = x5 & ~n7723 ;
  assign n7725 = ~n7722 & ~n7723 ;
  assign n7726 = ~n7724 & ~n7725 ;
  assign n7727 = n7715 & ~n7726 ;
  assign n7728 = n7715 & ~n7727 ;
  assign n7729 = ~n7726 & ~n7727 ;
  assign n7730 = ~n7728 & ~n7729 ;
  assign n7731 = ~n7307 & n7730 ;
  assign n7732 = n7307 & ~n7730 ;
  assign n7733 = ~n7731 & ~n7732 ;
  assign n7734 = x97 & n146 ;
  assign n7735 = x95 & n182 ;
  assign n7736 = x96 & n141 ;
  assign n7737 = ~n7735 & ~n7736 ;
  assign n7738 = ~n7734 & n7737 ;
  assign n7739 = ~n7317 & ~n7319 ;
  assign n7740 = ~x96 & ~x97 ;
  assign n7741 = x96 & x97 ;
  assign n7742 = ~n7740 & ~n7741 ;
  assign n7743 = ~n7739 & n7742 ;
  assign n7744 = n7739 & ~n7742 ;
  assign n7745 = ~n7743 & ~n7744 ;
  assign n7746 = n149 & n7745 ;
  assign n7747 = n7738 & ~n7746 ;
  assign n7748 = x2 & ~n7747 ;
  assign n7749 = x2 & ~n7748 ;
  assign n7750 = ~n7747 & ~n7748 ;
  assign n7751 = ~n7749 & ~n7750 ;
  assign n7752 = ~n7733 & ~n7751 ;
  assign n7753 = n7733 & n7751 ;
  assign n7754 = ~n7752 & ~n7753 ;
  assign n7755 = ~n7549 & n7754 ;
  assign n7756 = n7549 & ~n7754 ;
  assign n7757 = ~n7755 & ~n7756 ;
  assign n7963 = n7757 & x161 ;
  assign n7758 = ~n7522 & ~n7537 ;
  assign n7759 = ~n7541 & ~n7758 ;
  assign n7760 = ~n7480 & ~n7482 ;
  assign n7761 = ~n7441 & ~n7447 ;
  assign n7762 = ~n7425 & ~n7427 ;
  assign n7763 = ~n7386 & ~n7392 ;
  assign n7764 = ~x64 & ~n7556 ;
  assign n7765 = ~n7354 & n7764 ;
  assign n7766 = n7354 & ~n7764 ;
  assign n7767 = ~n7765 & ~n7766 ;
  assign n7768 = ~x67 & n6725 ;
  assign n7769 = ~x65 & n7129 ;
  assign n7770 = ~x66 & n6720 ;
  assign n7771 = ~n7769 & ~n7770 ;
  assign n7772 = ~n7768 & n7771 ;
  assign n7773 = n266 & n6728 ;
  assign n7774 = n7772 & ~n7773 ;
  assign n7775 = ~x32 & ~n7774 ;
  assign n7776 = ~x32 & ~n7775 ;
  assign n7777 = ~n7774 & ~n7775 ;
  assign n7778 = ~n7776 & ~n7777 ;
  assign n7779 = ~n7767 & ~n7778 ;
  assign n7780 = n7767 & n7778 ;
  assign n7781 = ~n7779 & ~n7780 ;
  assign n7782 = ~x70 & n5560 ;
  assign n7783 = ~x68 & n5943 ;
  assign n7784 = ~x69 & n5555 ;
  assign n7785 = ~n7783 & ~n7784 ;
  assign n7786 = ~n7782 & n7785 ;
  assign n7787 = n529 & n5563 ;
  assign n7788 = n7786 & ~n7787 ;
  assign n7789 = ~x29 & ~n7788 ;
  assign n7790 = ~x29 & ~n7789 ;
  assign n7791 = ~n7788 & ~n7789 ;
  assign n7792 = ~n7790 & ~n7791 ;
  assign n7793 = n7781 & ~n7792 ;
  assign n7794 = n7781 & ~n7793 ;
  assign n7795 = ~n7792 & ~n7793 ;
  assign n7796 = ~n7794 & ~n7795 ;
  assign n7797 = ~n7372 & n7796 ;
  assign n7798 = n7372 & ~n7796 ;
  assign n7799 = ~n7797 & ~n7798 ;
  assign n7800 = ~x73 & n4531 ;
  assign n7801 = ~x71 & n4847 ;
  assign n7802 = ~x72 & n4526 ;
  assign n7803 = ~n7801 & ~n7802 ;
  assign n7804 = ~n7800 & n7803 ;
  assign n7805 = n903 & n4534 ;
  assign n7806 = n7804 & ~n7805 ;
  assign n7807 = ~x26 & ~n7806 ;
  assign n7808 = ~x26 & ~n7807 ;
  assign n7809 = ~n7806 & ~n7807 ;
  assign n7810 = ~n7808 & ~n7809 ;
  assign n7811 = ~n7799 & ~n7810 ;
  assign n7812 = n7799 & n7810 ;
  assign n7813 = ~n7811 & ~n7812 ;
  assign n7814 = n7763 & ~n7813 ;
  assign n7815 = ~n7763 & n7813 ;
  assign n7816 = ~n7814 & ~n7815 ;
  assign n7817 = ~x76 & n3589 ;
  assign n7818 = ~x74 & n3878 ;
  assign n7819 = ~x75 & n3584 ;
  assign n7820 = ~n7818 & ~n7819 ;
  assign n7821 = ~n7817 & n7820 ;
  assign n7822 = n1390 & n3592 ;
  assign n7823 = n7821 & ~n7822 ;
  assign n7824 = ~x23 & ~n7823 ;
  assign n7825 = ~x23 & ~n7824 ;
  assign n7826 = ~n7823 & ~n7824 ;
  assign n7827 = ~n7825 & ~n7826 ;
  assign n7828 = ~n7816 & n7827 ;
  assign n7829 = n7816 & ~n7827 ;
  assign n7830 = ~n7828 & ~n7829 ;
  assign n7831 = ~n7410 & n7830 ;
  assign n7832 = n7410 & ~n7830 ;
  assign n7833 = ~n7831 & ~n7832 ;
  assign n7834 = ~x79 & n2751 ;
  assign n7835 = ~x77 & n3020 ;
  assign n7836 = ~x78 & n2746 ;
  assign n7837 = ~n7835 & ~n7836 ;
  assign n7838 = ~n7834 & n7837 ;
  assign n7839 = n1921 & n2754 ;
  assign n7840 = n7838 & ~n7839 ;
  assign n7841 = ~x20 & ~n7840 ;
  assign n7842 = ~x20 & ~n7841 ;
  assign n7843 = ~n7840 & ~n7841 ;
  assign n7844 = ~n7842 & ~n7843 ;
  assign n7845 = n7833 & ~n7844 ;
  assign n7846 = n7833 & ~n7845 ;
  assign n7847 = ~n7844 & ~n7845 ;
  assign n7848 = ~n7846 & ~n7847 ;
  assign n7849 = ~n7762 & n7848 ;
  assign n7850 = n7762 & ~n7848 ;
  assign n7851 = ~n7849 & ~n7850 ;
  assign n7852 = ~x82 & n2093 ;
  assign n7853 = ~x80 & n2275 ;
  assign n7854 = ~x81 & n2088 ;
  assign n7855 = ~n7853 & ~n7854 ;
  assign n7856 = ~n7852 & n7855 ;
  assign n7857 = n2096 & n2697 ;
  assign n7858 = n7856 & ~n7857 ;
  assign n7859 = ~x17 & ~n7858 ;
  assign n7860 = ~x17 & ~n7859 ;
  assign n7861 = ~n7858 & ~n7859 ;
  assign n7862 = ~n7860 & ~n7861 ;
  assign n7863 = ~n7851 & ~n7862 ;
  assign n7864 = n7851 & n7862 ;
  assign n7865 = ~n7863 & ~n7864 ;
  assign n7866 = n7761 & ~n7865 ;
  assign n7867 = ~n7761 & n7865 ;
  assign n7868 = ~n7866 & ~n7867 ;
  assign n7869 = ~x85 & n1434 ;
  assign n7870 = ~x83 & n1646 ;
  assign n7871 = ~x84 & n1429 ;
  assign n7872 = ~n7870 & ~n7871 ;
  assign n7873 = ~n7869 & n7872 ;
  assign n7874 = n1437 & n3521 ;
  assign n7875 = n7873 & ~n7874 ;
  assign n7876 = ~x14 & ~n7875 ;
  assign n7877 = ~x14 & ~n7876 ;
  assign n7878 = ~n7875 & ~n7876 ;
  assign n7879 = ~n7877 & ~n7878 ;
  assign n7880 = n7868 & ~n7879 ;
  assign n7881 = n7868 & ~n7880 ;
  assign n7882 = ~n7879 & ~n7880 ;
  assign n7883 = ~n7881 & ~n7882 ;
  assign n7884 = ~n7465 & n7883 ;
  assign n7885 = n7465 & ~n7883 ;
  assign n7886 = ~n7884 & ~n7885 ;
  assign n7887 = ~x88 & n945 ;
  assign n7888 = ~x86 & n1099 ;
  assign n7889 = ~x87 & n940 ;
  assign n7890 = ~n7888 & ~n7889 ;
  assign n7891 = ~n7887 & n7890 ;
  assign n7892 = n948 & n4457 ;
  assign n7893 = n7891 & ~n7892 ;
  assign n7894 = ~x11 & ~n7893 ;
  assign n7895 = ~x11 & ~n7894 ;
  assign n7896 = ~n7893 & ~n7894 ;
  assign n7897 = ~n7895 & ~n7896 ;
  assign n7898 = n7886 & n7897 ;
  assign n7899 = ~n7886 & ~n7897 ;
  assign n7900 = ~n7898 & ~n7899 ;
  assign n7901 = ~n7760 & n7900 ;
  assign n7902 = n7760 & ~n7900 ;
  assign n7903 = ~n7901 & ~n7902 ;
  assign n7904 = ~x91 & n574 ;
  assign n7905 = ~x89 & n673 ;
  assign n7906 = ~x90 & n569 ;
  assign n7907 = ~n7905 & ~n7906 ;
  assign n7908 = ~n7904 & n7907 ;
  assign n7909 = n577 & n5507 ;
  assign n7910 = n7908 & ~n7909 ;
  assign n7911 = ~x8 & ~n7910 ;
  assign n7912 = ~x8 & ~n7911 ;
  assign n7913 = ~n7910 & ~n7911 ;
  assign n7914 = ~n7912 & ~n7913 ;
  assign n7915 = n7903 & ~n7914 ;
  assign n7916 = n7903 & ~n7915 ;
  assign n7917 = ~n7914 & ~n7915 ;
  assign n7918 = ~n7916 & ~n7917 ;
  assign n7919 = ~n7496 & ~n7502 ;
  assign n7920 = n7918 & n7919 ;
  assign n7921 = ~n7918 & ~n7919 ;
  assign n7922 = ~n7920 & ~n7921 ;
  assign n7923 = ~x94 & n293 ;
  assign n7924 = ~x92 & n373 ;
  assign n7925 = ~x93 & n288 ;
  assign n7926 = ~n7924 & ~n7925 ;
  assign n7927 = ~n7923 & n7926 ;
  assign n7928 = n296 & n6671 ;
  assign n7929 = n7927 & ~n7928 ;
  assign n7930 = ~x5 & ~n7929 ;
  assign n7931 = ~x5 & ~n7930 ;
  assign n7932 = ~n7929 & ~n7930 ;
  assign n7933 = ~n7931 & ~n7932 ;
  assign n7934 = n7922 & ~n7933 ;
  assign n7935 = n7922 & ~n7934 ;
  assign n7936 = ~n7933 & ~n7934 ;
  assign n7937 = ~n7935 & ~n7936 ;
  assign n7938 = ~n7520 & n7937 ;
  assign n7939 = n7520 & ~n7937 ;
  assign n7940 = ~n7938 & ~n7939 ;
  assign n7941 = ~x97 & n164 ;
  assign n7942 = ~x95 & n205 ;
  assign n7943 = ~x96 & n162 ;
  assign n7944 = ~n7942 & ~n7943 ;
  assign n7945 = ~n7941 & n7944 ;
  assign n7946 = ~n7316 & ~n7529 ;
  assign n7947 = n7742 & ~n7946 ;
  assign n7948 = ~n7742 & n7946 ;
  assign n7949 = ~n7947 & ~n7948 ;
  assign n7950 = n167 & n7949 ;
  assign n7951 = n7945 & ~n7950 ;
  assign n7952 = ~x2 & ~n7951 ;
  assign n7953 = ~x2 & ~n7952 ;
  assign n7954 = ~n7951 & ~n7952 ;
  assign n7955 = ~n7953 & ~n7954 ;
  assign n7956 = ~n7940 & ~n7955 ;
  assign n7957 = n7940 & n7955 ;
  assign n7958 = ~n7956 & ~n7957 ;
  assign n7959 = ~n7759 & n7958 ;
  assign n7960 = n7759 & ~n7958 ;
  assign n7961 = ~n7959 & ~n7960 ;
  assign n7964 = ~n7961 & ~x161 ;
  assign n7965 = ~n7963 & ~n7964 ;
  assign n7966 = ~n7752 & ~n7755 ;
  assign n7967 = ~n7307 & ~n7730 ;
  assign n7968 = ~n7727 & ~n7967 ;
  assign n7969 = ~n7692 & ~n7694 ;
  assign n7970 = ~n7622 & ~n7624 ;
  assign n7971 = ~n7159 & ~n7589 ;
  assign n7972 = ~n7586 & ~n7971 ;
  assign n7973 = x71 & n5560 ;
  assign n7974 = x69 & n5943 ;
  assign n7975 = x70 & n5555 ;
  assign n7976 = ~n7974 & ~n7975 ;
  assign n7977 = ~n7973 & n7976 ;
  assign n7978 = n558 & n5563 ;
  assign n7979 = n7977 & ~n7978 ;
  assign n7980 = x29 & ~n7979 ;
  assign n7981 = x29 & ~n7980 ;
  assign n7982 = ~n7979 & ~n7980 ;
  assign n7983 = ~n7981 & ~n7982 ;
  assign n7984 = n7141 & n7557 ;
  assign n7985 = ~n7572 & ~n7984 ;
  assign n7986 = x68 & n6725 ;
  assign n7987 = x66 & n7129 ;
  assign n7988 = x67 & n6720 ;
  assign n7989 = ~n7987 & ~n7988 ;
  assign n7990 = ~n7986 & n7989 ;
  assign n7991 = n317 & n6728 ;
  assign n7992 = n7990 & ~n7991 ;
  assign n7993 = x32 & ~n7992 ;
  assign n7994 = x32 & ~n7993 ;
  assign n7995 = ~n7992 & ~n7993 ;
  assign n7996 = ~n7994 & ~n7995 ;
  assign n7997 = x35 & ~n7557 ;
  assign n7998 = ~x33 & x34 ;
  assign n7999 = x33 & ~x34 ;
  assign n8000 = ~n7998 & ~n7999 ;
  assign n8001 = n7556 & ~n8000 ;
  assign n8002 = x64 & n8001 ;
  assign n8003 = ~x34 & x35 ;
  assign n8004 = x34 & ~x35 ;
  assign n8005 = ~n8003 & ~n8004 ;
  assign n8006 = ~n7556 & n8005 ;
  assign n8007 = x65 & n8006 ;
  assign n8008 = ~n8002 & ~n8007 ;
  assign n8009 = ~n7556 & ~n8005 ;
  assign n8010 = ~n152 & n8009 ;
  assign n8011 = n8008 & ~n8010 ;
  assign n8012 = x35 & ~n8011 ;
  assign n8013 = x35 & ~n8012 ;
  assign n8014 = ~n8011 & ~n8012 ;
  assign n8015 = ~n8013 & ~n8014 ;
  assign n8016 = n7997 & ~n8015 ;
  assign n8017 = ~n7997 & n8015 ;
  assign n8018 = ~n8016 & ~n8017 ;
  assign n8019 = n7996 & ~n8018 ;
  assign n8020 = ~n7996 & n8018 ;
  assign n8021 = ~n8019 & ~n8020 ;
  assign n8022 = ~n7985 & n8021 ;
  assign n8023 = n7985 & ~n8021 ;
  assign n8024 = ~n8022 & ~n8023 ;
  assign n8025 = n7983 & ~n8024 ;
  assign n8026 = ~n7983 & n8024 ;
  assign n8027 = ~n8025 & ~n8026 ;
  assign n8028 = ~n7972 & n8027 ;
  assign n8029 = n7972 & ~n8027 ;
  assign n8030 = ~n8028 & ~n8029 ;
  assign n8031 = x74 & n4531 ;
  assign n8032 = x72 & n4847 ;
  assign n8033 = x73 & n4526 ;
  assign n8034 = ~n8032 & ~n8033 ;
  assign n8035 = ~n8031 & n8034 ;
  assign n8036 = n994 & n4534 ;
  assign n8037 = n8035 & ~n8036 ;
  assign n8038 = x26 & ~n8037 ;
  assign n8039 = x26 & ~n8038 ;
  assign n8040 = ~n8037 & ~n8038 ;
  assign n8041 = ~n8039 & ~n8040 ;
  assign n8042 = n8030 & ~n8041 ;
  assign n8043 = n8030 & ~n8042 ;
  assign n8044 = ~n8041 & ~n8042 ;
  assign n8045 = ~n8043 & ~n8044 ;
  assign n8046 = ~n7604 & ~n7608 ;
  assign n8047 = n8045 & n8046 ;
  assign n8048 = ~n8045 & ~n8046 ;
  assign n8049 = ~n8047 & ~n8048 ;
  assign n8050 = x77 & n3589 ;
  assign n8051 = x75 & n3878 ;
  assign n8052 = x76 & n3584 ;
  assign n8053 = ~n8051 & ~n8052 ;
  assign n8054 = ~n8050 & n8053 ;
  assign n8055 = n1502 & n3592 ;
  assign n8056 = n8054 & ~n8055 ;
  assign n8057 = x23 & ~n8056 ;
  assign n8058 = x23 & ~n8057 ;
  assign n8059 = ~n8056 & ~n8057 ;
  assign n8060 = ~n8058 & ~n8059 ;
  assign n8061 = n8049 & ~n8060 ;
  assign n8062 = ~n8049 & n8060 ;
  assign n8063 = ~n7970 & ~n8062 ;
  assign n8064 = ~n8061 & n8063 ;
  assign n8065 = ~n7970 & ~n8064 ;
  assign n8066 = ~n8061 & ~n8064 ;
  assign n8067 = ~n8062 & n8066 ;
  assign n8068 = ~n8065 & ~n8067 ;
  assign n8069 = x80 & n2751 ;
  assign n8070 = x78 & n3020 ;
  assign n8071 = x79 & n2746 ;
  assign n8072 = ~n8070 & ~n8071 ;
  assign n8073 = ~n8069 & n8072 ;
  assign n8074 = n2028 & n2754 ;
  assign n8075 = n8073 & ~n8074 ;
  assign n8076 = x20 & ~n8075 ;
  assign n8077 = x20 & ~n8076 ;
  assign n8078 = ~n8075 & ~n8076 ;
  assign n8079 = ~n8077 & ~n8078 ;
  assign n8080 = ~n8068 & ~n8079 ;
  assign n8081 = ~n8068 & ~n8080 ;
  assign n8082 = ~n8079 & ~n8080 ;
  assign n8083 = ~n8081 & ~n8082 ;
  assign n8084 = ~n7552 & ~n7641 ;
  assign n8085 = ~n7638 & ~n8084 ;
  assign n8086 = n8083 & n8085 ;
  assign n8087 = ~n8083 & ~n8085 ;
  assign n8088 = ~n8086 & ~n8087 ;
  assign n8089 = x83 & n2093 ;
  assign n8090 = x81 & n2275 ;
  assign n8091 = x82 & n2088 ;
  assign n8092 = ~n8090 & ~n8091 ;
  assign n8093 = ~n8089 & n8092 ;
  assign n8094 = n2096 & n2843 ;
  assign n8095 = n8093 & ~n8094 ;
  assign n8096 = x17 & ~n8095 ;
  assign n8097 = x17 & ~n8096 ;
  assign n8098 = ~n8095 & ~n8096 ;
  assign n8099 = ~n8097 & ~n8098 ;
  assign n8100 = n8088 & ~n8099 ;
  assign n8101 = n8088 & ~n8100 ;
  assign n8102 = ~n8099 & ~n8100 ;
  assign n8103 = ~n8101 & ~n8102 ;
  assign n8104 = ~n7656 & ~n7660 ;
  assign n8105 = n8103 & n8104 ;
  assign n8106 = ~n8103 & ~n8104 ;
  assign n8107 = ~n8105 & ~n8106 ;
  assign n8108 = x86 & n1434 ;
  assign n8109 = x84 & n1646 ;
  assign n8110 = x85 & n1429 ;
  assign n8111 = ~n8109 & ~n8110 ;
  assign n8112 = ~n8108 & n8111 ;
  assign n8113 = n1437 & n3686 ;
  assign n8114 = n8112 & ~n8113 ;
  assign n8115 = x14 & ~n8114 ;
  assign n8116 = x14 & ~n8115 ;
  assign n8117 = ~n8114 & ~n8115 ;
  assign n8118 = ~n8116 & ~n8117 ;
  assign n8119 = n8107 & ~n8118 ;
  assign n8120 = n8107 & ~n8119 ;
  assign n8121 = ~n8118 & ~n8119 ;
  assign n8122 = ~n8120 & ~n8121 ;
  assign n8123 = ~n7252 & ~n7676 ;
  assign n8124 = ~n7673 & ~n8123 ;
  assign n8125 = n8122 & n8124 ;
  assign n8126 = ~n8122 & ~n8124 ;
  assign n8127 = ~n8125 & ~n8126 ;
  assign n8128 = x89 & n945 ;
  assign n8129 = x87 & n1099 ;
  assign n8130 = x88 & n940 ;
  assign n8131 = ~n8129 & ~n8130 ;
  assign n8132 = ~n8128 & n8131 ;
  assign n8133 = n948 & n4488 ;
  assign n8134 = n8132 & ~n8133 ;
  assign n8135 = x11 & ~n8134 ;
  assign n8136 = x11 & ~n8135 ;
  assign n8137 = ~n8134 & ~n8135 ;
  assign n8138 = ~n8136 & ~n8137 ;
  assign n8139 = n8127 & ~n8138 ;
  assign n8140 = ~n8127 & n8138 ;
  assign n8141 = ~n7969 & ~n8140 ;
  assign n8142 = ~n8139 & n8141 ;
  assign n8143 = ~n7969 & ~n8142 ;
  assign n8144 = ~n8139 & ~n8142 ;
  assign n8145 = ~n8140 & n8144 ;
  assign n8146 = ~n8143 & ~n8145 ;
  assign n8147 = x92 & n574 ;
  assign n8148 = x90 & n673 ;
  assign n8149 = x91 & n569 ;
  assign n8150 = ~n8148 & ~n8149 ;
  assign n8151 = ~n8147 & n8150 ;
  assign n8152 = n577 & n5710 ;
  assign n8153 = n8151 & ~n8152 ;
  assign n8154 = x8 & ~n8153 ;
  assign n8155 = x8 & ~n8154 ;
  assign n8156 = ~n8153 & ~n8154 ;
  assign n8157 = ~n8155 & ~n8156 ;
  assign n8158 = ~n8146 & ~n8157 ;
  assign n8159 = ~n8146 & ~n8158 ;
  assign n8160 = ~n8157 & ~n8158 ;
  assign n8161 = ~n8159 & ~n8160 ;
  assign n8162 = ~n7708 & ~n7714 ;
  assign n8163 = n8161 & n8162 ;
  assign n8164 = ~n8161 & ~n8162 ;
  assign n8165 = ~n8163 & ~n8164 ;
  assign n8166 = x95 & n293 ;
  assign n8167 = x93 & n373 ;
  assign n8168 = x94 & n288 ;
  assign n8169 = ~n8167 & ~n8168 ;
  assign n8170 = ~n8166 & n8169 ;
  assign n8171 = n296 & n6894 ;
  assign n8172 = n8170 & ~n8171 ;
  assign n8173 = x5 & ~n8172 ;
  assign n8174 = x5 & ~n8173 ;
  assign n8175 = ~n8172 & ~n8173 ;
  assign n8176 = ~n8174 & ~n8175 ;
  assign n8177 = n8165 & ~n8176 ;
  assign n8178 = ~n8165 & n8176 ;
  assign n8179 = ~n7968 & ~n8178 ;
  assign n8180 = ~n8177 & n8179 ;
  assign n8181 = ~n7968 & ~n8180 ;
  assign n8182 = ~n8177 & ~n8180 ;
  assign n8183 = ~n8178 & n8182 ;
  assign n8184 = ~n8181 & ~n8183 ;
  assign n8185 = x98 & n146 ;
  assign n8186 = x96 & n182 ;
  assign n8187 = x97 & n141 ;
  assign n8188 = ~n8186 & ~n8187 ;
  assign n8189 = ~n8185 & n8188 ;
  assign n8190 = ~n7741 & ~n7743 ;
  assign n8191 = ~x97 & ~x98 ;
  assign n8192 = x97 & x98 ;
  assign n8193 = ~n8191 & ~n8192 ;
  assign n8194 = ~n8190 & n8193 ;
  assign n8195 = n8190 & ~n8193 ;
  assign n8196 = ~n8194 & ~n8195 ;
  assign n8197 = n149 & n8196 ;
  assign n8198 = n8189 & ~n8197 ;
  assign n8199 = x2 & ~n8198 ;
  assign n8200 = x2 & ~n8199 ;
  assign n8201 = ~n8198 & ~n8199 ;
  assign n8202 = ~n8200 & ~n8201 ;
  assign n8203 = ~n8184 & n8202 ;
  assign n8204 = n8184 & ~n8202 ;
  assign n8205 = ~n8203 & ~n8204 ;
  assign n8206 = ~n7966 & ~n8205 ;
  assign n8207 = n7966 & n8205 ;
  assign n8208 = ~n8206 & ~n8207 ;
  assign n8440 = n8208 & x162 ;
  assign n8209 = ~n7956 & ~n7959 ;
  assign n8210 = ~n7520 & ~n7937 ;
  assign n8211 = ~n7934 & ~n8210 ;
  assign n8212 = ~n7899 & ~n7901 ;
  assign n8213 = ~n7829 & ~n7831 ;
  assign n8214 = ~n7372 & ~n7796 ;
  assign n8215 = ~n7793 & ~n8214 ;
  assign n8216 = ~x71 & n5560 ;
  assign n8217 = ~x69 & n5943 ;
  assign n8218 = ~x70 & n5555 ;
  assign n8219 = ~n8217 & ~n8218 ;
  assign n8220 = ~n8216 & n8219 ;
  assign n8221 = n622 & n5563 ;
  assign n8222 = n8220 & ~n8221 ;
  assign n8223 = ~x29 & ~n8222 ;
  assign n8224 = ~x29 & ~n8223 ;
  assign n8225 = ~n8222 & ~n8223 ;
  assign n8226 = ~n8224 & ~n8225 ;
  assign n8227 = n7354 & n7764 ;
  assign n8228 = ~n7779 & ~n8227 ;
  assign n8229 = ~x68 & n6725 ;
  assign n8230 = ~x66 & n7129 ;
  assign n8231 = ~x67 & n6720 ;
  assign n8232 = ~n8230 & ~n8231 ;
  assign n8233 = ~n8229 & n8232 ;
  assign n8234 = n352 & n6728 ;
  assign n8235 = n8233 & ~n8234 ;
  assign n8236 = ~x32 & ~n8235 ;
  assign n8237 = ~x32 & ~n8236 ;
  assign n8238 = ~n8235 & ~n8236 ;
  assign n8239 = ~n8237 & ~n8238 ;
  assign n8240 = ~x35 & ~n7764 ;
  assign n8241 = ~x64 & n8001 ;
  assign n8242 = ~x65 & n8006 ;
  assign n8243 = ~n8241 & ~n8242 ;
  assign n8244 = ~n8010 & n8243 ;
  assign n8245 = ~x35 & ~n8244 ;
  assign n8246 = ~x35 & ~n8245 ;
  assign n8247 = ~n8244 & ~n8245 ;
  assign n8248 = ~n8246 & ~n8247 ;
  assign n8249 = n8240 & ~n8248 ;
  assign n8250 = ~n8240 & n8248 ;
  assign n8251 = ~n8249 & ~n8250 ;
  assign n8252 = n8239 & ~n8251 ;
  assign n8253 = ~n8239 & n8251 ;
  assign n8254 = ~n8252 & ~n8253 ;
  assign n8255 = ~n8228 & n8254 ;
  assign n8256 = n8228 & ~n8254 ;
  assign n8257 = ~n8255 & ~n8256 ;
  assign n8258 = n8226 & ~n8257 ;
  assign n8259 = ~n8226 & n8257 ;
  assign n8260 = ~n8258 & ~n8259 ;
  assign n8261 = ~n8215 & n8260 ;
  assign n8262 = n8215 & ~n8260 ;
  assign n8263 = ~n8261 & ~n8262 ;
  assign n8264 = ~x74 & n4531 ;
  assign n8265 = ~x72 & n4847 ;
  assign n8266 = ~x73 & n4526 ;
  assign n8267 = ~n8265 & ~n8266 ;
  assign n8268 = ~n8264 & n8267 ;
  assign n8269 = n1066 & n4534 ;
  assign n8270 = n8268 & ~n8269 ;
  assign n8271 = ~x26 & ~n8270 ;
  assign n8272 = ~x26 & ~n8271 ;
  assign n8273 = ~n8270 & ~n8271 ;
  assign n8274 = ~n8272 & ~n8273 ;
  assign n8275 = n8263 & ~n8274 ;
  assign n8276 = n8263 & ~n8275 ;
  assign n8277 = ~n8274 & ~n8275 ;
  assign n8278 = ~n8276 & ~n8277 ;
  assign n8279 = ~n7811 & ~n7815 ;
  assign n8280 = n8278 & n8279 ;
  assign n8281 = ~n8278 & ~n8279 ;
  assign n8282 = ~n8280 & ~n8281 ;
  assign n8283 = ~x77 & n3589 ;
  assign n8284 = ~x75 & n3878 ;
  assign n8285 = ~x76 & n3584 ;
  assign n8286 = ~n8284 & ~n8285 ;
  assign n8287 = ~n8283 & n8286 ;
  assign n8288 = n1594 & n3592 ;
  assign n8289 = n8287 & ~n8288 ;
  assign n8290 = ~x23 & ~n8289 ;
  assign n8291 = ~x23 & ~n8290 ;
  assign n8292 = ~n8289 & ~n8290 ;
  assign n8293 = ~n8291 & ~n8292 ;
  assign n8294 = n8282 & ~n8293 ;
  assign n8295 = ~n8282 & n8293 ;
  assign n8296 = ~n8213 & ~n8295 ;
  assign n8297 = ~n8294 & n8296 ;
  assign n8298 = ~n8213 & ~n8297 ;
  assign n8299 = ~n8294 & ~n8297 ;
  assign n8300 = ~n8295 & n8299 ;
  assign n8301 = ~n8298 & ~n8300 ;
  assign n8302 = ~x80 & n2751 ;
  assign n8303 = ~x78 & n3020 ;
  assign n8304 = ~x79 & n2746 ;
  assign n8305 = ~n8303 & ~n8304 ;
  assign n8306 = ~n8302 & n8305 ;
  assign n8307 = n2145 & n2754 ;
  assign n8308 = n8306 & ~n8307 ;
  assign n8309 = ~x20 & ~n8308 ;
  assign n8310 = ~x20 & ~n8309 ;
  assign n8311 = ~n8308 & ~n8309 ;
  assign n8312 = ~n8310 & ~n8311 ;
  assign n8313 = ~n8301 & ~n8312 ;
  assign n8314 = ~n8301 & ~n8313 ;
  assign n8315 = ~n8312 & ~n8313 ;
  assign n8316 = ~n8314 & ~n8315 ;
  assign n8317 = ~n7762 & ~n7848 ;
  assign n8318 = ~n7845 & ~n8317 ;
  assign n8319 = n8316 & n8318 ;
  assign n8320 = ~n8316 & ~n8318 ;
  assign n8321 = ~n8319 & ~n8320 ;
  assign n8322 = ~x83 & n2093 ;
  assign n8323 = ~x81 & n2275 ;
  assign n8324 = ~x82 & n2088 ;
  assign n8325 = ~n8323 & ~n8324 ;
  assign n8326 = ~n8322 & n8325 ;
  assign n8327 = n2096 & n2972 ;
  assign n8328 = n8326 & ~n8327 ;
  assign n8329 = ~x17 & ~n8328 ;
  assign n8330 = ~x17 & ~n8329 ;
  assign n8331 = ~n8328 & ~n8329 ;
  assign n8332 = ~n8330 & ~n8331 ;
  assign n8333 = n8321 & ~n8332 ;
  assign n8334 = n8321 & ~n8333 ;
  assign n8335 = ~n8332 & ~n8333 ;
  assign n8336 = ~n8334 & ~n8335 ;
  assign n8337 = ~n7863 & ~n7867 ;
  assign n8338 = n8336 & n8337 ;
  assign n8339 = ~n8336 & ~n8337 ;
  assign n8340 = ~n8338 & ~n8339 ;
  assign n8341 = ~x86 & n1434 ;
  assign n8342 = ~x84 & n1646 ;
  assign n8343 = ~x85 & n1429 ;
  assign n8344 = ~n8342 & ~n8343 ;
  assign n8345 = ~n8341 & n8344 ;
  assign n8346 = n1437 & n3832 ;
  assign n8347 = n8345 & ~n8346 ;
  assign n8348 = ~x14 & ~n8347 ;
  assign n8349 = ~x14 & ~n8348 ;
  assign n8350 = ~n8347 & ~n8348 ;
  assign n8351 = ~n8349 & ~n8350 ;
  assign n8352 = n8340 & ~n8351 ;
  assign n8353 = n8340 & ~n8352 ;
  assign n8354 = ~n8351 & ~n8352 ;
  assign n8355 = ~n8353 & ~n8354 ;
  assign n8356 = ~n7465 & ~n7883 ;
  assign n8357 = ~n7880 & ~n8356 ;
  assign n8358 = n8355 & n8357 ;
  assign n8359 = ~n8355 & ~n8357 ;
  assign n8360 = ~n8358 & ~n8359 ;
  assign n8361 = ~x89 & n945 ;
  assign n8362 = ~x87 & n1099 ;
  assign n8363 = ~x88 & n940 ;
  assign n8364 = ~n8362 & ~n8363 ;
  assign n8365 = ~n8361 & n8364 ;
  assign n8366 = n948 & n4664 ;
  assign n8367 = n8365 & ~n8366 ;
  assign n8368 = ~x11 & ~n8367 ;
  assign n8369 = ~x11 & ~n8368 ;
  assign n8370 = ~n8367 & ~n8368 ;
  assign n8371 = ~n8369 & ~n8370 ;
  assign n8372 = n8360 & ~n8371 ;
  assign n8373 = ~n8360 & n8371 ;
  assign n8374 = ~n8212 & ~n8373 ;
  assign n8375 = ~n8372 & n8374 ;
  assign n8376 = ~n8212 & ~n8375 ;
  assign n8377 = ~n8372 & ~n8375 ;
  assign n8378 = ~n8373 & n8377 ;
  assign n8379 = ~n8376 & ~n8378 ;
  assign n8380 = ~x92 & n574 ;
  assign n8381 = ~x90 & n673 ;
  assign n8382 = ~x91 & n569 ;
  assign n8383 = ~n8381 & ~n8382 ;
  assign n8384 = ~n8380 & n8383 ;
  assign n8385 = n577 & n5896 ;
  assign n8386 = n8384 & ~n8385 ;
  assign n8387 = ~x8 & ~n8386 ;
  assign n8388 = ~x8 & ~n8387 ;
  assign n8389 = ~n8386 & ~n8387 ;
  assign n8390 = ~n8388 & ~n8389 ;
  assign n8391 = ~n8379 & ~n8390 ;
  assign n8392 = ~n8379 & ~n8391 ;
  assign n8393 = ~n8390 & ~n8391 ;
  assign n8394 = ~n8392 & ~n8393 ;
  assign n8395 = ~n7915 & ~n7921 ;
  assign n8396 = n8394 & n8395 ;
  assign n8397 = ~n8394 & ~n8395 ;
  assign n8398 = ~n8396 & ~n8397 ;
  assign n8399 = ~x95 & n293 ;
  assign n8400 = ~x93 & n373 ;
  assign n8401 = ~x94 & n288 ;
  assign n8402 = ~n8400 & ~n8401 ;
  assign n8403 = ~n8399 & n8402 ;
  assign n8404 = n296 & n7100 ;
  assign n8405 = n8403 & ~n8404 ;
  assign n8406 = ~x5 & ~n8405 ;
  assign n8407 = ~x5 & ~n8406 ;
  assign n8408 = ~n8405 & ~n8406 ;
  assign n8409 = ~n8407 & ~n8408 ;
  assign n8410 = n8398 & ~n8409 ;
  assign n8411 = ~n8398 & n8409 ;
  assign n8412 = ~n8211 & ~n8411 ;
  assign n8413 = ~n8410 & n8412 ;
  assign n8414 = ~n8211 & ~n8413 ;
  assign n8415 = ~n8410 & ~n8413 ;
  assign n8416 = ~n8411 & n8415 ;
  assign n8417 = ~n8414 & ~n8416 ;
  assign n8418 = ~x98 & n164 ;
  assign n8419 = ~x96 & n205 ;
  assign n8420 = ~x97 & n162 ;
  assign n8421 = ~n8419 & ~n8420 ;
  assign n8422 = ~n8418 & n8421 ;
  assign n8423 = ~n7740 & ~n7947 ;
  assign n8424 = n8193 & ~n8423 ;
  assign n8425 = ~n8193 & n8423 ;
  assign n8426 = ~n8424 & ~n8425 ;
  assign n8427 = n167 & n8426 ;
  assign n8428 = n8422 & ~n8427 ;
  assign n8429 = ~x2 & ~n8428 ;
  assign n8430 = ~x2 & ~n8429 ;
  assign n8431 = ~n8428 & ~n8429 ;
  assign n8432 = ~n8430 & ~n8431 ;
  assign n8433 = ~n8417 & n8432 ;
  assign n8434 = n8417 & ~n8432 ;
  assign n8435 = ~n8433 & ~n8434 ;
  assign n8436 = ~n8209 & ~n8435 ;
  assign n8437 = n8209 & n8435 ;
  assign n8438 = ~n8436 & ~n8437 ;
  assign n8441 = ~n8438 & ~x162 ;
  assign n8442 = ~n8440 & ~n8441 ;
  assign n8443 = ~n8184 & ~n8202 ;
  assign n8444 = ~n8206 & ~n8443 ;
  assign n8445 = x90 & n945 ;
  assign n8446 = x88 & n1099 ;
  assign n8447 = x89 & n940 ;
  assign n8448 = ~n8446 & ~n8447 ;
  assign n8449 = ~n8445 & n8448 ;
  assign n8450 = n948 & n4986 ;
  assign n8451 = n8449 & ~n8450 ;
  assign n8452 = x11 & ~n8451 ;
  assign n8453 = x11 & ~n8452 ;
  assign n8454 = ~n8451 & ~n8452 ;
  assign n8455 = ~n8453 & ~n8454 ;
  assign n8456 = ~n8119 & ~n8126 ;
  assign n8457 = ~n8100 & ~n8106 ;
  assign n8458 = ~n8042 & ~n8048 ;
  assign n8459 = x75 & n4531 ;
  assign n8460 = x73 & n4847 ;
  assign n8461 = x74 & n4526 ;
  assign n8462 = ~n8460 & ~n8461 ;
  assign n8463 = ~n8459 & n8462 ;
  assign n8464 = n1150 & n4534 ;
  assign n8465 = n8463 & ~n8464 ;
  assign n8466 = x26 & ~n8465 ;
  assign n8467 = x26 & ~n8466 ;
  assign n8468 = ~n8465 & ~n8466 ;
  assign n8469 = ~n8467 & ~n8468 ;
  assign n8470 = ~n8026 & ~n8028 ;
  assign n8471 = ~n8020 & ~n8022 ;
  assign n8472 = x66 & n8006 ;
  assign n8473 = n7556 & ~n8005 ;
  assign n8474 = n8000 & n8473 ;
  assign n8475 = x64 & n8474 ;
  assign n8476 = x65 & n8001 ;
  assign n8477 = ~n8475 & ~n8476 ;
  assign n8478 = ~n8472 & n8477 ;
  assign n8479 = n194 & n8009 ;
  assign n8480 = n8478 & ~n8479 ;
  assign n8481 = x35 & ~n8480 ;
  assign n8482 = x35 & ~n8481 ;
  assign n8483 = ~n8480 & ~n8481 ;
  assign n8484 = ~n8482 & ~n8483 ;
  assign n8485 = ~n8016 & n8484 ;
  assign n8486 = n8016 & ~n8484 ;
  assign n8487 = ~n8485 & ~n8486 ;
  assign n8488 = x69 & n6725 ;
  assign n8489 = x67 & n7129 ;
  assign n8490 = x68 & n6720 ;
  assign n8491 = ~n8489 & ~n8490 ;
  assign n8492 = ~n8488 & n8491 ;
  assign n8493 = n398 & n6728 ;
  assign n8494 = n8492 & ~n8493 ;
  assign n8495 = x32 & ~n8494 ;
  assign n8496 = x32 & ~n8495 ;
  assign n8497 = ~n8494 & ~n8495 ;
  assign n8498 = ~n8496 & ~n8497 ;
  assign n8499 = n8487 & ~n8498 ;
  assign n8500 = ~n8487 & n8498 ;
  assign n8501 = ~n8471 & ~n8500 ;
  assign n8502 = ~n8499 & n8501 ;
  assign n8503 = ~n8471 & ~n8502 ;
  assign n8504 = ~n8499 & ~n8502 ;
  assign n8505 = ~n8500 & n8504 ;
  assign n8506 = ~n8503 & ~n8505 ;
  assign n8507 = x72 & n5560 ;
  assign n8508 = x70 & n5943 ;
  assign n8509 = x71 & n5555 ;
  assign n8510 = ~n8508 & ~n8509 ;
  assign n8511 = ~n8507 & n8510 ;
  assign n8512 = n717 & n5563 ;
  assign n8513 = n8511 & ~n8512 ;
  assign n8514 = x29 & ~n8513 ;
  assign n8515 = x29 & ~n8514 ;
  assign n8516 = ~n8513 & ~n8514 ;
  assign n8517 = ~n8515 & ~n8516 ;
  assign n8518 = ~n8506 & ~n8517 ;
  assign n8519 = ~n8506 & ~n8518 ;
  assign n8520 = ~n8517 & ~n8518 ;
  assign n8521 = ~n8519 & ~n8520 ;
  assign n8522 = ~n8470 & ~n8521 ;
  assign n8523 = n8470 & n8521 ;
  assign n8524 = ~n8522 & ~n8523 ;
  assign n8525 = ~n8469 & n8524 ;
  assign n8526 = ~n8469 & ~n8525 ;
  assign n8527 = n8524 & ~n8525 ;
  assign n8528 = ~n8526 & ~n8527 ;
  assign n8529 = ~n8458 & ~n8528 ;
  assign n8530 = ~n8458 & ~n8529 ;
  assign n8531 = ~n8528 & ~n8529 ;
  assign n8532 = ~n8530 & ~n8531 ;
  assign n8533 = x78 & n3589 ;
  assign n8534 = x76 & n3878 ;
  assign n8535 = x77 & n3584 ;
  assign n8536 = ~n8534 & ~n8535 ;
  assign n8537 = ~n8533 & n8536 ;
  assign n8538 = n1624 & n3592 ;
  assign n8539 = n8537 & ~n8538 ;
  assign n8540 = x23 & ~n8539 ;
  assign n8541 = x23 & ~n8540 ;
  assign n8542 = ~n8539 & ~n8540 ;
  assign n8543 = ~n8541 & ~n8542 ;
  assign n8544 = n8532 & n8543 ;
  assign n8545 = ~n8532 & ~n8543 ;
  assign n8546 = ~n8544 & ~n8545 ;
  assign n8547 = ~n8066 & n8546 ;
  assign n8548 = n8066 & ~n8546 ;
  assign n8549 = ~n8547 & ~n8548 ;
  assign n8550 = x81 & n2751 ;
  assign n8551 = x79 & n3020 ;
  assign n8552 = x80 & n2746 ;
  assign n8553 = ~n8551 & ~n8552 ;
  assign n8554 = ~n8550 & n8553 ;
  assign n8555 = n2348 & n2754 ;
  assign n8556 = n8554 & ~n8555 ;
  assign n8557 = x20 & ~n8556 ;
  assign n8558 = x20 & ~n8557 ;
  assign n8559 = ~n8556 & ~n8557 ;
  assign n8560 = ~n8558 & ~n8559 ;
  assign n8561 = n8549 & ~n8560 ;
  assign n8562 = n8549 & ~n8561 ;
  assign n8563 = ~n8560 & ~n8561 ;
  assign n8564 = ~n8562 & ~n8563 ;
  assign n8565 = ~n8080 & ~n8087 ;
  assign n8566 = n8564 & n8565 ;
  assign n8567 = ~n8564 & ~n8565 ;
  assign n8568 = ~n8566 & ~n8567 ;
  assign n8569 = x84 & n2093 ;
  assign n8570 = x82 & n2275 ;
  assign n8571 = x83 & n2088 ;
  assign n8572 = ~n8570 & ~n8571 ;
  assign n8573 = ~n8569 & n8572 ;
  assign n8574 = n2096 & n3114 ;
  assign n8575 = n8573 & ~n8574 ;
  assign n8576 = x17 & ~n8575 ;
  assign n8577 = x17 & ~n8576 ;
  assign n8578 = ~n8575 & ~n8576 ;
  assign n8579 = ~n8577 & ~n8578 ;
  assign n8580 = n8568 & ~n8579 ;
  assign n8581 = ~n8568 & n8579 ;
  assign n8582 = ~n8457 & ~n8581 ;
  assign n8583 = ~n8580 & n8582 ;
  assign n8584 = ~n8457 & ~n8583 ;
  assign n8585 = ~n8580 & ~n8583 ;
  assign n8586 = ~n8581 & n8585 ;
  assign n8587 = ~n8584 & ~n8586 ;
  assign n8588 = x87 & n1434 ;
  assign n8589 = x85 & n1646 ;
  assign n8590 = x86 & n1429 ;
  assign n8591 = ~n8589 & ~n8590 ;
  assign n8592 = ~n8588 & n8591 ;
  assign n8593 = n1437 & n3991 ;
  assign n8594 = n8592 & ~n8593 ;
  assign n8595 = x14 & ~n8594 ;
  assign n8596 = x14 & ~n8595 ;
  assign n8597 = ~n8594 & ~n8595 ;
  assign n8598 = ~n8596 & ~n8597 ;
  assign n8599 = n8587 & n8598 ;
  assign n8600 = ~n8587 & ~n8598 ;
  assign n8601 = ~n8599 & ~n8600 ;
  assign n8602 = ~n8456 & n8601 ;
  assign n8603 = n8456 & ~n8601 ;
  assign n8604 = ~n8602 & ~n8603 ;
  assign n8605 = n8455 & ~n8604 ;
  assign n8606 = ~n8455 & n8604 ;
  assign n8607 = ~n8605 & ~n8606 ;
  assign n8608 = ~n8144 & n8607 ;
  assign n8609 = n8144 & ~n8607 ;
  assign n8610 = ~n8608 & ~n8609 ;
  assign n8611 = x93 & n574 ;
  assign n8612 = x91 & n673 ;
  assign n8613 = x92 & n569 ;
  assign n8614 = ~n8612 & ~n8613 ;
  assign n8615 = ~n8611 & n8614 ;
  assign n8616 = n577 & n6094 ;
  assign n8617 = n8615 & ~n8616 ;
  assign n8618 = x8 & ~n8617 ;
  assign n8619 = x8 & ~n8618 ;
  assign n8620 = ~n8617 & ~n8618 ;
  assign n8621 = ~n8619 & ~n8620 ;
  assign n8622 = n8610 & ~n8621 ;
  assign n8623 = n8610 & ~n8622 ;
  assign n8624 = ~n8621 & ~n8622 ;
  assign n8625 = ~n8623 & ~n8624 ;
  assign n8626 = ~n8158 & ~n8164 ;
  assign n8627 = n8625 & n8626 ;
  assign n8628 = ~n8625 & ~n8626 ;
  assign n8629 = ~n8627 & ~n8628 ;
  assign n8630 = x96 & n293 ;
  assign n8631 = x94 & n373 ;
  assign n8632 = x95 & n288 ;
  assign n8633 = ~n8631 & ~n8632 ;
  assign n8634 = ~n8630 & n8633 ;
  assign n8635 = n296 & n7321 ;
  assign n8636 = n8634 & ~n8635 ;
  assign n8637 = x5 & ~n8636 ;
  assign n8638 = x5 & ~n8637 ;
  assign n8639 = ~n8636 & ~n8637 ;
  assign n8640 = ~n8638 & ~n8639 ;
  assign n8641 = n8629 & ~n8640 ;
  assign n8642 = ~n8629 & n8640 ;
  assign n8643 = ~n8182 & ~n8642 ;
  assign n8644 = ~n8641 & n8643 ;
  assign n8645 = ~n8182 & ~n8644 ;
  assign n8646 = ~n8641 & ~n8644 ;
  assign n8647 = ~n8642 & n8646 ;
  assign n8648 = ~n8645 & ~n8647 ;
  assign n8649 = x99 & n146 ;
  assign n8650 = x97 & n182 ;
  assign n8651 = x98 & n141 ;
  assign n8652 = ~n8650 & ~n8651 ;
  assign n8653 = ~n8649 & n8652 ;
  assign n8654 = ~n8192 & ~n8194 ;
  assign n8655 = ~x98 & ~x99 ;
  assign n8656 = x98 & x99 ;
  assign n8657 = ~n8655 & ~n8656 ;
  assign n8658 = ~n8654 & n8657 ;
  assign n8659 = n8654 & ~n8657 ;
  assign n8660 = ~n8658 & ~n8659 ;
  assign n8661 = n149 & n8660 ;
  assign n8662 = n8653 & ~n8661 ;
  assign n8663 = x2 & ~n8662 ;
  assign n8664 = x2 & ~n8663 ;
  assign n8665 = ~n8662 & ~n8663 ;
  assign n8666 = ~n8664 & ~n8665 ;
  assign n8667 = ~n8648 & n8666 ;
  assign n8668 = n8648 & ~n8666 ;
  assign n8669 = ~n8667 & ~n8668 ;
  assign n8670 = ~n8444 & ~n8669 ;
  assign n8671 = n8444 & n8669 ;
  assign n8672 = ~n8670 & ~n8671 ;
  assign n8899 = n8672 & x163 ;
  assign n8673 = ~n8417 & ~n8432 ;
  assign n8674 = ~n8436 & ~n8673 ;
  assign n8675 = ~x90 & n945 ;
  assign n8676 = ~x88 & n1099 ;
  assign n8677 = ~x89 & n940 ;
  assign n8678 = ~n8676 & ~n8677 ;
  assign n8679 = ~n8675 & n8678 ;
  assign n8680 = n948 & n5155 ;
  assign n8681 = n8679 & ~n8680 ;
  assign n8682 = ~x11 & ~n8681 ;
  assign n8683 = ~x11 & ~n8682 ;
  assign n8684 = ~n8681 & ~n8682 ;
  assign n8685 = ~n8683 & ~n8684 ;
  assign n8686 = ~n8352 & ~n8359 ;
  assign n8687 = ~n8333 & ~n8339 ;
  assign n8688 = ~n8275 & ~n8281 ;
  assign n8689 = ~x75 & n4531 ;
  assign n8690 = ~x73 & n4847 ;
  assign n8691 = ~x74 & n4526 ;
  assign n8692 = ~n8690 & ~n8691 ;
  assign n8693 = ~n8689 & n8692 ;
  assign n8694 = n1225 & n4534 ;
  assign n8695 = n8693 & ~n8694 ;
  assign n8696 = ~x26 & ~n8695 ;
  assign n8697 = ~x26 & ~n8696 ;
  assign n8698 = ~n8695 & ~n8696 ;
  assign n8699 = ~n8697 & ~n8698 ;
  assign n8700 = ~n8259 & ~n8261 ;
  assign n8701 = ~n8253 & ~n8255 ;
  assign n8702 = ~x66 & n8006 ;
  assign n8703 = ~x64 & n8474 ;
  assign n8704 = ~x65 & n8001 ;
  assign n8705 = ~n8703 & ~n8704 ;
  assign n8706 = ~n8702 & n8705 ;
  assign n8707 = n214 & n8009 ;
  assign n8708 = n8706 & ~n8707 ;
  assign n8709 = ~x35 & ~n8708 ;
  assign n8710 = ~x35 & ~n8709 ;
  assign n8711 = ~n8708 & ~n8709 ;
  assign n8712 = ~n8710 & ~n8711 ;
  assign n8713 = ~n8249 & n8712 ;
  assign n8714 = n8249 & ~n8712 ;
  assign n8715 = ~n8713 & ~n8714 ;
  assign n8716 = ~x69 & n6725 ;
  assign n8717 = ~x67 & n7129 ;
  assign n8718 = ~x68 & n6720 ;
  assign n8719 = ~n8717 & ~n8718 ;
  assign n8720 = ~n8716 & n8719 ;
  assign n8721 = n435 & n6728 ;
  assign n8722 = n8720 & ~n8721 ;
  assign n8723 = ~x32 & ~n8722 ;
  assign n8724 = ~x32 & ~n8723 ;
  assign n8725 = ~n8722 & ~n8723 ;
  assign n8726 = ~n8724 & ~n8725 ;
  assign n8727 = n8715 & ~n8726 ;
  assign n8728 = ~n8715 & n8726 ;
  assign n8729 = ~n8701 & ~n8728 ;
  assign n8730 = ~n8727 & n8729 ;
  assign n8731 = ~n8701 & ~n8730 ;
  assign n8732 = ~n8727 & ~n8730 ;
  assign n8733 = ~n8728 & n8732 ;
  assign n8734 = ~n8731 & ~n8733 ;
  assign n8735 = ~x72 & n5560 ;
  assign n8736 = ~x70 & n5943 ;
  assign n8737 = ~x71 & n5555 ;
  assign n8738 = ~n8736 & ~n8737 ;
  assign n8739 = ~n8735 & n8738 ;
  assign n8740 = n773 & n5563 ;
  assign n8741 = n8739 & ~n8740 ;
  assign n8742 = ~x29 & ~n8741 ;
  assign n8743 = ~x29 & ~n8742 ;
  assign n8744 = ~n8741 & ~n8742 ;
  assign n8745 = ~n8743 & ~n8744 ;
  assign n8746 = ~n8734 & ~n8745 ;
  assign n8747 = ~n8734 & ~n8746 ;
  assign n8748 = ~n8745 & ~n8746 ;
  assign n8749 = ~n8747 & ~n8748 ;
  assign n8750 = ~n8700 & ~n8749 ;
  assign n8751 = n8700 & n8749 ;
  assign n8752 = ~n8750 & ~n8751 ;
  assign n8753 = ~n8699 & n8752 ;
  assign n8754 = ~n8699 & ~n8753 ;
  assign n8755 = n8752 & ~n8753 ;
  assign n8756 = ~n8754 & ~n8755 ;
  assign n8757 = ~n8688 & ~n8756 ;
  assign n8758 = ~n8688 & ~n8757 ;
  assign n8759 = ~n8756 & ~n8757 ;
  assign n8760 = ~n8758 & ~n8759 ;
  assign n8761 = ~x78 & n3589 ;
  assign n8762 = ~x76 & n3878 ;
  assign n8763 = ~x77 & n3584 ;
  assign n8764 = ~n8762 & ~n8763 ;
  assign n8765 = ~n8761 & n8764 ;
  assign n8766 = n1718 & n3592 ;
  assign n8767 = n8765 & ~n8766 ;
  assign n8768 = ~x23 & ~n8767 ;
  assign n8769 = ~x23 & ~n8768 ;
  assign n8770 = ~n8767 & ~n8768 ;
  assign n8771 = ~n8769 & ~n8770 ;
  assign n8772 = n8760 & n8771 ;
  assign n8773 = ~n8760 & ~n8771 ;
  assign n8774 = ~n8772 & ~n8773 ;
  assign n8775 = ~n8299 & n8774 ;
  assign n8776 = n8299 & ~n8774 ;
  assign n8777 = ~n8775 & ~n8776 ;
  assign n8778 = ~x81 & n2751 ;
  assign n8779 = ~x79 & n3020 ;
  assign n8780 = ~x80 & n2746 ;
  assign n8781 = ~n8779 & ~n8780 ;
  assign n8782 = ~n8778 & n8781 ;
  assign n8783 = n2460 & n2754 ;
  assign n8784 = n8782 & ~n8783 ;
  assign n8785 = ~x20 & ~n8784 ;
  assign n8786 = ~x20 & ~n8785 ;
  assign n8787 = ~n8784 & ~n8785 ;
  assign n8788 = ~n8786 & ~n8787 ;
  assign n8789 = n8777 & ~n8788 ;
  assign n8790 = n8777 & ~n8789 ;
  assign n8791 = ~n8788 & ~n8789 ;
  assign n8792 = ~n8790 & ~n8791 ;
  assign n8793 = ~n8313 & ~n8320 ;
  assign n8794 = n8792 & n8793 ;
  assign n8795 = ~n8792 & ~n8793 ;
  assign n8796 = ~n8794 & ~n8795 ;
  assign n8797 = ~x84 & n2093 ;
  assign n8798 = ~x82 & n2275 ;
  assign n8799 = ~x83 & n2088 ;
  assign n8800 = ~n8798 & ~n8799 ;
  assign n8801 = ~n8797 & n8800 ;
  assign n8802 = n2096 & n3247 ;
  assign n8803 = n8801 & ~n8802 ;
  assign n8804 = ~x17 & ~n8803 ;
  assign n8805 = ~x17 & ~n8804 ;
  assign n8806 = ~n8803 & ~n8804 ;
  assign n8807 = ~n8805 & ~n8806 ;
  assign n8808 = n8796 & ~n8807 ;
  assign n8809 = ~n8796 & n8807 ;
  assign n8810 = ~n8687 & ~n8809 ;
  assign n8811 = ~n8808 & n8810 ;
  assign n8812 = ~n8687 & ~n8811 ;
  assign n8813 = ~n8808 & ~n8811 ;
  assign n8814 = ~n8809 & n8813 ;
  assign n8815 = ~n8812 & ~n8814 ;
  assign n8816 = ~x87 & n1434 ;
  assign n8817 = ~x85 & n1646 ;
  assign n8818 = ~x86 & n1429 ;
  assign n8819 = ~n8817 & ~n8818 ;
  assign n8820 = ~n8816 & n8819 ;
  assign n8821 = n1437 & n4143 ;
  assign n8822 = n8820 & ~n8821 ;
  assign n8823 = ~x14 & ~n8822 ;
  assign n8824 = ~x14 & ~n8823 ;
  assign n8825 = ~n8822 & ~n8823 ;
  assign n8826 = ~n8824 & ~n8825 ;
  assign n8827 = n8815 & n8826 ;
  assign n8828 = ~n8815 & ~n8826 ;
  assign n8829 = ~n8827 & ~n8828 ;
  assign n8830 = ~n8686 & n8829 ;
  assign n8831 = n8686 & ~n8829 ;
  assign n8832 = ~n8830 & ~n8831 ;
  assign n8833 = n8685 & ~n8832 ;
  assign n8834 = ~n8685 & n8832 ;
  assign n8835 = ~n8833 & ~n8834 ;
  assign n8836 = ~n8377 & n8835 ;
  assign n8837 = n8377 & ~n8835 ;
  assign n8838 = ~n8836 & ~n8837 ;
  assign n8839 = ~x93 & n574 ;
  assign n8840 = ~x91 & n673 ;
  assign n8841 = ~x92 & n569 ;
  assign n8842 = ~n8840 & ~n8841 ;
  assign n8843 = ~n8839 & n8842 ;
  assign n8844 = n577 & n6285 ;
  assign n8845 = n8843 & ~n8844 ;
  assign n8846 = ~x8 & ~n8845 ;
  assign n8847 = ~x8 & ~n8846 ;
  assign n8848 = ~n8845 & ~n8846 ;
  assign n8849 = ~n8847 & ~n8848 ;
  assign n8850 = n8838 & ~n8849 ;
  assign n8851 = n8838 & ~n8850 ;
  assign n8852 = ~n8849 & ~n8850 ;
  assign n8853 = ~n8851 & ~n8852 ;
  assign n8854 = ~n8391 & ~n8397 ;
  assign n8855 = n8853 & n8854 ;
  assign n8856 = ~n8853 & ~n8854 ;
  assign n8857 = ~n8855 & ~n8856 ;
  assign n8858 = ~x96 & n293 ;
  assign n8859 = ~x94 & n373 ;
  assign n8860 = ~x95 & n288 ;
  assign n8861 = ~n8859 & ~n8860 ;
  assign n8862 = ~n8858 & n8861 ;
  assign n8863 = n296 & n7531 ;
  assign n8864 = n8862 & ~n8863 ;
  assign n8865 = ~x5 & ~n8864 ;
  assign n8866 = ~x5 & ~n8865 ;
  assign n8867 = ~n8864 & ~n8865 ;
  assign n8868 = ~n8866 & ~n8867 ;
  assign n8869 = n8857 & ~n8868 ;
  assign n8870 = ~n8857 & n8868 ;
  assign n8871 = ~n8415 & ~n8870 ;
  assign n8872 = ~n8869 & n8871 ;
  assign n8873 = ~n8415 & ~n8872 ;
  assign n8874 = ~n8869 & ~n8872 ;
  assign n8875 = ~n8870 & n8874 ;
  assign n8876 = ~n8873 & ~n8875 ;
  assign n8877 = ~x99 & n164 ;
  assign n8878 = ~x97 & n205 ;
  assign n8879 = ~x98 & n162 ;
  assign n8880 = ~n8878 & ~n8879 ;
  assign n8881 = ~n8877 & n8880 ;
  assign n8882 = ~n8191 & ~n8424 ;
  assign n8883 = n8657 & ~n8882 ;
  assign n8884 = ~n8657 & n8882 ;
  assign n8885 = ~n8883 & ~n8884 ;
  assign n8886 = n167 & n8885 ;
  assign n8887 = n8881 & ~n8886 ;
  assign n8888 = ~x2 & ~n8887 ;
  assign n8889 = ~x2 & ~n8888 ;
  assign n8890 = ~n8887 & ~n8888 ;
  assign n8891 = ~n8889 & ~n8890 ;
  assign n8892 = ~n8876 & n8891 ;
  assign n8893 = n8876 & ~n8891 ;
  assign n8894 = ~n8892 & ~n8893 ;
  assign n8895 = ~n8674 & ~n8894 ;
  assign n8896 = n8674 & n8894 ;
  assign n8897 = ~n8895 & ~n8896 ;
  assign n8900 = ~n8897 & ~x163 ;
  assign n8901 = ~n8899 & ~n8900 ;
  assign n8902 = x97 & n293 ;
  assign n8903 = x95 & n373 ;
  assign n8904 = x96 & n288 ;
  assign n8905 = ~n8903 & ~n8904 ;
  assign n8906 = ~n8902 & n8905 ;
  assign n8907 = n296 & n7745 ;
  assign n8908 = n8906 & ~n8907 ;
  assign n8909 = x5 & ~n8908 ;
  assign n8910 = x5 & ~n8909 ;
  assign n8911 = ~n8908 & ~n8909 ;
  assign n8912 = ~n8910 & ~n8911 ;
  assign n8913 = ~n8622 & ~n8628 ;
  assign n8914 = ~n8606 & ~n8608 ;
  assign n8915 = ~n8600 & ~n8602 ;
  assign n8916 = ~n8561 & ~n8567 ;
  assign n8917 = ~n8545 & ~n8547 ;
  assign n8918 = ~n8518 & ~n8522 ;
  assign n8919 = x35 & ~x36 ;
  assign n8920 = ~x35 & x36 ;
  assign n8921 = ~n8919 & ~n8920 ;
  assign n8922 = x64 & ~n8921 ;
  assign n8923 = ~n8486 & n8922 ;
  assign n8924 = n8486 & ~n8922 ;
  assign n8925 = ~n8923 & ~n8924 ;
  assign n8926 = x67 & n8006 ;
  assign n8927 = x65 & n8474 ;
  assign n8928 = x66 & n8001 ;
  assign n8929 = ~n8927 & ~n8928 ;
  assign n8930 = ~n8926 & n8929 ;
  assign n8931 = n240 & n8009 ;
  assign n8932 = n8930 & ~n8931 ;
  assign n8933 = x35 & ~n8932 ;
  assign n8934 = x35 & ~n8933 ;
  assign n8935 = ~n8932 & ~n8933 ;
  assign n8936 = ~n8934 & ~n8935 ;
  assign n8937 = ~n8925 & ~n8936 ;
  assign n8938 = n8925 & n8936 ;
  assign n8939 = ~n8937 & ~n8938 ;
  assign n8940 = x70 & n6725 ;
  assign n8941 = x68 & n7129 ;
  assign n8942 = x69 & n6720 ;
  assign n8943 = ~n8941 & ~n8942 ;
  assign n8944 = ~n8940 & n8943 ;
  assign n8945 = n488 & n6728 ;
  assign n8946 = n8944 & ~n8945 ;
  assign n8947 = x32 & ~n8946 ;
  assign n8948 = x32 & ~n8947 ;
  assign n8949 = ~n8946 & ~n8947 ;
  assign n8950 = ~n8948 & ~n8949 ;
  assign n8951 = n8939 & ~n8950 ;
  assign n8952 = n8939 & ~n8951 ;
  assign n8953 = ~n8950 & ~n8951 ;
  assign n8954 = ~n8952 & ~n8953 ;
  assign n8955 = ~n8504 & n8954 ;
  assign n8956 = n8504 & ~n8954 ;
  assign n8957 = ~n8955 & ~n8956 ;
  assign n8958 = x73 & n5560 ;
  assign n8959 = x71 & n5943 ;
  assign n8960 = x72 & n5555 ;
  assign n8961 = ~n8959 & ~n8960 ;
  assign n8962 = ~n8958 & n8961 ;
  assign n8963 = n843 & n5563 ;
  assign n8964 = n8962 & ~n8963 ;
  assign n8965 = x29 & ~n8964 ;
  assign n8966 = x29 & ~n8965 ;
  assign n8967 = ~n8964 & ~n8965 ;
  assign n8968 = ~n8966 & ~n8967 ;
  assign n8969 = ~n8957 & ~n8968 ;
  assign n8970 = n8957 & n8968 ;
  assign n8971 = ~n8969 & ~n8970 ;
  assign n8972 = n8918 & ~n8971 ;
  assign n8973 = ~n8918 & n8971 ;
  assign n8974 = ~n8972 & ~n8973 ;
  assign n8975 = x76 & n4531 ;
  assign n8976 = x74 & n4847 ;
  assign n8977 = x75 & n4526 ;
  assign n8978 = ~n8976 & ~n8977 ;
  assign n8979 = ~n8975 & n8978 ;
  assign n8980 = n1311 & n4534 ;
  assign n8981 = n8979 & ~n8980 ;
  assign n8982 = x26 & ~n8981 ;
  assign n8983 = x26 & ~n8982 ;
  assign n8984 = ~n8981 & ~n8982 ;
  assign n8985 = ~n8983 & ~n8984 ;
  assign n8986 = ~n8974 & n8985 ;
  assign n8987 = n8974 & ~n8985 ;
  assign n8988 = ~n8986 & ~n8987 ;
  assign n8989 = ~n8525 & ~n8529 ;
  assign n8990 = n8988 & ~n8989 ;
  assign n8991 = ~n8988 & n8989 ;
  assign n8992 = ~n8990 & ~n8991 ;
  assign n8993 = x79 & n3589 ;
  assign n8994 = x77 & n3878 ;
  assign n8995 = x78 & n3584 ;
  assign n8996 = ~n8994 & ~n8995 ;
  assign n8997 = ~n8993 & n8996 ;
  assign n8998 = n1817 & n3592 ;
  assign n8999 = n8997 & ~n8998 ;
  assign n9000 = x23 & ~n8999 ;
  assign n9001 = x23 & ~n9000 ;
  assign n9002 = ~n8999 & ~n9000 ;
  assign n9003 = ~n9001 & ~n9002 ;
  assign n9004 = n8992 & ~n9003 ;
  assign n9005 = n8992 & ~n9004 ;
  assign n9006 = ~n9003 & ~n9004 ;
  assign n9007 = ~n9005 & ~n9006 ;
  assign n9008 = ~n8917 & n9007 ;
  assign n9009 = n8917 & ~n9007 ;
  assign n9010 = ~n9008 & ~n9009 ;
  assign n9011 = x82 & n2751 ;
  assign n9012 = x80 & n3020 ;
  assign n9013 = x81 & n2746 ;
  assign n9014 = ~n9012 & ~n9013 ;
  assign n9015 = ~n9011 & n9014 ;
  assign n9016 = n2584 & n2754 ;
  assign n9017 = n9015 & ~n9016 ;
  assign n9018 = x20 & ~n9017 ;
  assign n9019 = x20 & ~n9018 ;
  assign n9020 = ~n9017 & ~n9018 ;
  assign n9021 = ~n9019 & ~n9020 ;
  assign n9022 = ~n9010 & ~n9021 ;
  assign n9023 = n9010 & n9021 ;
  assign n9024 = ~n9022 & ~n9023 ;
  assign n9025 = n8916 & ~n9024 ;
  assign n9026 = ~n8916 & n9024 ;
  assign n9027 = ~n9025 & ~n9026 ;
  assign n9028 = x85 & n2093 ;
  assign n9029 = x83 & n2275 ;
  assign n9030 = x84 & n2088 ;
  assign n9031 = ~n9029 & ~n9030 ;
  assign n9032 = ~n9028 & n9031 ;
  assign n9033 = n2096 & n3389 ;
  assign n9034 = n9032 & ~n9033 ;
  assign n9035 = x17 & ~n9034 ;
  assign n9036 = x17 & ~n9035 ;
  assign n9037 = ~n9034 & ~n9035 ;
  assign n9038 = ~n9036 & ~n9037 ;
  assign n9039 = n9027 & ~n9038 ;
  assign n9040 = n9027 & ~n9039 ;
  assign n9041 = ~n9038 & ~n9039 ;
  assign n9042 = ~n9040 & ~n9041 ;
  assign n9043 = ~n8585 & n9042 ;
  assign n9044 = n8585 & ~n9042 ;
  assign n9045 = ~n9043 & ~n9044 ;
  assign n9046 = x88 & n1434 ;
  assign n9047 = x86 & n1646 ;
  assign n9048 = x87 & n1429 ;
  assign n9049 = ~n9047 & ~n9048 ;
  assign n9050 = ~n9046 & n9049 ;
  assign n9051 = n1437 & n4305 ;
  assign n9052 = n9050 & ~n9051 ;
  assign n9053 = x14 & ~n9052 ;
  assign n9054 = x14 & ~n9053 ;
  assign n9055 = ~n9052 & ~n9053 ;
  assign n9056 = ~n9054 & ~n9055 ;
  assign n9057 = n9045 & n9056 ;
  assign n9058 = ~n9045 & ~n9056 ;
  assign n9059 = ~n9057 & ~n9058 ;
  assign n9060 = ~n8915 & n9059 ;
  assign n9061 = n8915 & ~n9059 ;
  assign n9062 = ~n9060 & ~n9061 ;
  assign n9063 = x91 & n945 ;
  assign n9064 = x89 & n1099 ;
  assign n9065 = x90 & n940 ;
  assign n9066 = ~n9064 & ~n9065 ;
  assign n9067 = ~n9063 & n9066 ;
  assign n9068 = n948 & n5336 ;
  assign n9069 = n9067 & ~n9068 ;
  assign n9070 = x11 & ~n9069 ;
  assign n9071 = x11 & ~n9070 ;
  assign n9072 = ~n9069 & ~n9070 ;
  assign n9073 = ~n9071 & ~n9072 ;
  assign n9074 = n9062 & ~n9073 ;
  assign n9075 = n9062 & ~n9074 ;
  assign n9076 = ~n9073 & ~n9074 ;
  assign n9077 = ~n9075 & ~n9076 ;
  assign n9078 = ~n8914 & n9077 ;
  assign n9079 = n8914 & ~n9077 ;
  assign n9080 = ~n9078 & ~n9079 ;
  assign n9081 = x94 & n574 ;
  assign n9082 = x92 & n673 ;
  assign n9083 = x93 & n569 ;
  assign n9084 = ~n9082 & ~n9083 ;
  assign n9085 = ~n9081 & n9084 ;
  assign n9086 = n577 & n6483 ;
  assign n9087 = n9085 & ~n9086 ;
  assign n9088 = x8 & ~n9087 ;
  assign n9089 = x8 & ~n9088 ;
  assign n9090 = ~n9087 & ~n9088 ;
  assign n9091 = ~n9089 & ~n9090 ;
  assign n9092 = n9080 & n9091 ;
  assign n9093 = ~n9080 & ~n9091 ;
  assign n9094 = ~n9092 & ~n9093 ;
  assign n9095 = ~n8913 & n9094 ;
  assign n9096 = n8913 & ~n9094 ;
  assign n9097 = ~n9095 & ~n9096 ;
  assign n9098 = ~n8912 & n9097 ;
  assign n9099 = n8912 & ~n9097 ;
  assign n9100 = ~n9098 & ~n9099 ;
  assign n9101 = ~n8646 & n9100 ;
  assign n9102 = n8646 & ~n9100 ;
  assign n9103 = ~n9101 & ~n9102 ;
  assign n9104 = x100 & n146 ;
  assign n9105 = x98 & n182 ;
  assign n9106 = x99 & n141 ;
  assign n9107 = ~n9105 & ~n9106 ;
  assign n9108 = ~n9104 & n9107 ;
  assign n9109 = ~n8656 & ~n8658 ;
  assign n9110 = ~x99 & ~x100 ;
  assign n9111 = x99 & x100 ;
  assign n9112 = ~n9110 & ~n9111 ;
  assign n9113 = ~n9109 & n9112 ;
  assign n9114 = n9109 & ~n9112 ;
  assign n9115 = ~n9113 & ~n9114 ;
  assign n9116 = n149 & n9115 ;
  assign n9117 = n9108 & ~n9116 ;
  assign n9118 = x2 & ~n9117 ;
  assign n9119 = x2 & ~n9118 ;
  assign n9120 = ~n9117 & ~n9118 ;
  assign n9121 = ~n9119 & ~n9120 ;
  assign n9122 = n9103 & ~n9121 ;
  assign n9123 = n9103 & ~n9122 ;
  assign n9124 = ~n9121 & ~n9122 ;
  assign n9125 = ~n9123 & ~n9124 ;
  assign n9126 = ~n8648 & ~n8666 ;
  assign n9127 = ~n8670 & ~n9126 ;
  assign n9128 = ~n9125 & ~n9127 ;
  assign n9129 = n9125 & n9127 ;
  assign n9130 = ~n9128 & ~n9129 ;
  assign n9355 = n9130 & x164 ;
  assign n9131 = ~x97 & n293 ;
  assign n9132 = ~x95 & n373 ;
  assign n9133 = ~x96 & n288 ;
  assign n9134 = ~n9132 & ~n9133 ;
  assign n9135 = ~n9131 & n9134 ;
  assign n9136 = n296 & n7949 ;
  assign n9137 = n9135 & ~n9136 ;
  assign n9138 = ~x5 & ~n9137 ;
  assign n9139 = ~x5 & ~n9138 ;
  assign n9140 = ~n9137 & ~n9138 ;
  assign n9141 = ~n9139 & ~n9140 ;
  assign n9142 = ~n8850 & ~n8856 ;
  assign n9143 = ~n8834 & ~n8836 ;
  assign n9144 = ~n8828 & ~n8830 ;
  assign n9145 = ~n8789 & ~n8795 ;
  assign n9146 = ~n8773 & ~n8775 ;
  assign n9147 = ~n8746 & ~n8750 ;
  assign n9148 = ~x64 & ~n8921 ;
  assign n9149 = ~n8714 & n9148 ;
  assign n9150 = n8714 & ~n9148 ;
  assign n9151 = ~n9149 & ~n9150 ;
  assign n9152 = ~x67 & n8006 ;
  assign n9153 = ~x65 & n8474 ;
  assign n9154 = ~x66 & n8001 ;
  assign n9155 = ~n9153 & ~n9154 ;
  assign n9156 = ~n9152 & n9155 ;
  assign n9157 = n266 & n8009 ;
  assign n9158 = n9156 & ~n9157 ;
  assign n9159 = ~x35 & ~n9158 ;
  assign n9160 = ~x35 & ~n9159 ;
  assign n9161 = ~n9158 & ~n9159 ;
  assign n9162 = ~n9160 & ~n9161 ;
  assign n9163 = ~n9151 & ~n9162 ;
  assign n9164 = n9151 & n9162 ;
  assign n9165 = ~n9163 & ~n9164 ;
  assign n9166 = ~x70 & n6725 ;
  assign n9167 = ~x68 & n7129 ;
  assign n9168 = ~x69 & n6720 ;
  assign n9169 = ~n9167 & ~n9168 ;
  assign n9170 = ~n9166 & n9169 ;
  assign n9171 = n529 & n6728 ;
  assign n9172 = n9170 & ~n9171 ;
  assign n9173 = ~x32 & ~n9172 ;
  assign n9174 = ~x32 & ~n9173 ;
  assign n9175 = ~n9172 & ~n9173 ;
  assign n9176 = ~n9174 & ~n9175 ;
  assign n9177 = n9165 & ~n9176 ;
  assign n9178 = n9165 & ~n9177 ;
  assign n9179 = ~n9176 & ~n9177 ;
  assign n9180 = ~n9178 & ~n9179 ;
  assign n9181 = ~n8732 & n9180 ;
  assign n9182 = n8732 & ~n9180 ;
  assign n9183 = ~n9181 & ~n9182 ;
  assign n9184 = ~x73 & n5560 ;
  assign n9185 = ~x71 & n5943 ;
  assign n9186 = ~x72 & n5555 ;
  assign n9187 = ~n9185 & ~n9186 ;
  assign n9188 = ~n9184 & n9187 ;
  assign n9189 = n903 & n5563 ;
  assign n9190 = n9188 & ~n9189 ;
  assign n9191 = ~x29 & ~n9190 ;
  assign n9192 = ~x29 & ~n9191 ;
  assign n9193 = ~n9190 & ~n9191 ;
  assign n9194 = ~n9192 & ~n9193 ;
  assign n9195 = ~n9183 & ~n9194 ;
  assign n9196 = n9183 & n9194 ;
  assign n9197 = ~n9195 & ~n9196 ;
  assign n9198 = n9147 & ~n9197 ;
  assign n9199 = ~n9147 & n9197 ;
  assign n9200 = ~n9198 & ~n9199 ;
  assign n9201 = ~x76 & n4531 ;
  assign n9202 = ~x74 & n4847 ;
  assign n9203 = ~x75 & n4526 ;
  assign n9204 = ~n9202 & ~n9203 ;
  assign n9205 = ~n9201 & n9204 ;
  assign n9206 = n1390 & n4534 ;
  assign n9207 = n9205 & ~n9206 ;
  assign n9208 = ~x26 & ~n9207 ;
  assign n9209 = ~x26 & ~n9208 ;
  assign n9210 = ~n9207 & ~n9208 ;
  assign n9211 = ~n9209 & ~n9210 ;
  assign n9212 = ~n9200 & n9211 ;
  assign n9213 = n9200 & ~n9211 ;
  assign n9214 = ~n9212 & ~n9213 ;
  assign n9215 = ~n8753 & ~n8757 ;
  assign n9216 = n9214 & ~n9215 ;
  assign n9217 = ~n9214 & n9215 ;
  assign n9218 = ~n9216 & ~n9217 ;
  assign n9219 = ~x79 & n3589 ;
  assign n9220 = ~x77 & n3878 ;
  assign n9221 = ~x78 & n3584 ;
  assign n9222 = ~n9220 & ~n9221 ;
  assign n9223 = ~n9219 & n9222 ;
  assign n9224 = n1921 & n3592 ;
  assign n9225 = n9223 & ~n9224 ;
  assign n9226 = ~x23 & ~n9225 ;
  assign n9227 = ~x23 & ~n9226 ;
  assign n9228 = ~n9225 & ~n9226 ;
  assign n9229 = ~n9227 & ~n9228 ;
  assign n9230 = n9218 & ~n9229 ;
  assign n9231 = n9218 & ~n9230 ;
  assign n9232 = ~n9229 & ~n9230 ;
  assign n9233 = ~n9231 & ~n9232 ;
  assign n9234 = ~n9146 & n9233 ;
  assign n9235 = n9146 & ~n9233 ;
  assign n9236 = ~n9234 & ~n9235 ;
  assign n9237 = ~x82 & n2751 ;
  assign n9238 = ~x80 & n3020 ;
  assign n9239 = ~x81 & n2746 ;
  assign n9240 = ~n9238 & ~n9239 ;
  assign n9241 = ~n9237 & n9240 ;
  assign n9242 = n2697 & n2754 ;
  assign n9243 = n9241 & ~n9242 ;
  assign n9244 = ~x20 & ~n9243 ;
  assign n9245 = ~x20 & ~n9244 ;
  assign n9246 = ~n9243 & ~n9244 ;
  assign n9247 = ~n9245 & ~n9246 ;
  assign n9248 = ~n9236 & ~n9247 ;
  assign n9249 = n9236 & n9247 ;
  assign n9250 = ~n9248 & ~n9249 ;
  assign n9251 = n9145 & ~n9250 ;
  assign n9252 = ~n9145 & n9250 ;
  assign n9253 = ~n9251 & ~n9252 ;
  assign n9254 = ~x85 & n2093 ;
  assign n9255 = ~x83 & n2275 ;
  assign n9256 = ~x84 & n2088 ;
  assign n9257 = ~n9255 & ~n9256 ;
  assign n9258 = ~n9254 & n9257 ;
  assign n9259 = n2096 & n3521 ;
  assign n9260 = n9258 & ~n9259 ;
  assign n9261 = ~x17 & ~n9260 ;
  assign n9262 = ~x17 & ~n9261 ;
  assign n9263 = ~n9260 & ~n9261 ;
  assign n9264 = ~n9262 & ~n9263 ;
  assign n9265 = n9253 & ~n9264 ;
  assign n9266 = n9253 & ~n9265 ;
  assign n9267 = ~n9264 & ~n9265 ;
  assign n9268 = ~n9266 & ~n9267 ;
  assign n9269 = ~n8813 & n9268 ;
  assign n9270 = n8813 & ~n9268 ;
  assign n9271 = ~n9269 & ~n9270 ;
  assign n9272 = ~x88 & n1434 ;
  assign n9273 = ~x86 & n1646 ;
  assign n9274 = ~x87 & n1429 ;
  assign n9275 = ~n9273 & ~n9274 ;
  assign n9276 = ~n9272 & n9275 ;
  assign n9277 = n1437 & n4457 ;
  assign n9278 = n9276 & ~n9277 ;
  assign n9279 = ~x14 & ~n9278 ;
  assign n9280 = ~x14 & ~n9279 ;
  assign n9281 = ~n9278 & ~n9279 ;
  assign n9282 = ~n9280 & ~n9281 ;
  assign n9283 = n9271 & n9282 ;
  assign n9284 = ~n9271 & ~n9282 ;
  assign n9285 = ~n9283 & ~n9284 ;
  assign n9286 = ~n9144 & n9285 ;
  assign n9287 = n9144 & ~n9285 ;
  assign n9288 = ~n9286 & ~n9287 ;
  assign n9289 = ~x91 & n945 ;
  assign n9290 = ~x89 & n1099 ;
  assign n9291 = ~x90 & n940 ;
  assign n9292 = ~n9290 & ~n9291 ;
  assign n9293 = ~n9289 & n9292 ;
  assign n9294 = n948 & n5507 ;
  assign n9295 = n9293 & ~n9294 ;
  assign n9296 = ~x11 & ~n9295 ;
  assign n9297 = ~x11 & ~n9296 ;
  assign n9298 = ~n9295 & ~n9296 ;
  assign n9299 = ~n9297 & ~n9298 ;
  assign n9300 = n9288 & ~n9299 ;
  assign n9301 = n9288 & ~n9300 ;
  assign n9302 = ~n9299 & ~n9300 ;
  assign n9303 = ~n9301 & ~n9302 ;
  assign n9304 = ~n9143 & n9303 ;
  assign n9305 = n9143 & ~n9303 ;
  assign n9306 = ~n9304 & ~n9305 ;
  assign n9307 = ~x94 & n574 ;
  assign n9308 = ~x92 & n673 ;
  assign n9309 = ~x93 & n569 ;
  assign n9310 = ~n9308 & ~n9309 ;
  assign n9311 = ~n9307 & n9310 ;
  assign n9312 = n577 & n6671 ;
  assign n9313 = n9311 & ~n9312 ;
  assign n9314 = ~x8 & ~n9313 ;
  assign n9315 = ~x8 & ~n9314 ;
  assign n9316 = ~n9313 & ~n9314 ;
  assign n9317 = ~n9315 & ~n9316 ;
  assign n9318 = n9306 & n9317 ;
  assign n9319 = ~n9306 & ~n9317 ;
  assign n9320 = ~n9318 & ~n9319 ;
  assign n9321 = ~n9142 & n9320 ;
  assign n9322 = n9142 & ~n9320 ;
  assign n9323 = ~n9321 & ~n9322 ;
  assign n9324 = ~n9141 & n9323 ;
  assign n9325 = n9141 & ~n9323 ;
  assign n9326 = ~n9324 & ~n9325 ;
  assign n9327 = ~n8874 & n9326 ;
  assign n9328 = n8874 & ~n9326 ;
  assign n9329 = ~n9327 & ~n9328 ;
  assign n9330 = ~x100 & n164 ;
  assign n9331 = ~x98 & n205 ;
  assign n9332 = ~x99 & n162 ;
  assign n9333 = ~n9331 & ~n9332 ;
  assign n9334 = ~n9330 & n9333 ;
  assign n9335 = ~n8655 & ~n8883 ;
  assign n9336 = n9112 & ~n9335 ;
  assign n9337 = ~n9112 & n9335 ;
  assign n9338 = ~n9336 & ~n9337 ;
  assign n9339 = n167 & n9338 ;
  assign n9340 = n9334 & ~n9339 ;
  assign n9341 = ~x2 & ~n9340 ;
  assign n9342 = ~x2 & ~n9341 ;
  assign n9343 = ~n9340 & ~n9341 ;
  assign n9344 = ~n9342 & ~n9343 ;
  assign n9345 = n9329 & ~n9344 ;
  assign n9346 = n9329 & ~n9345 ;
  assign n9347 = ~n9344 & ~n9345 ;
  assign n9348 = ~n9346 & ~n9347 ;
  assign n9349 = ~n8876 & ~n8891 ;
  assign n9350 = ~n8895 & ~n9349 ;
  assign n9351 = ~n9348 & ~n9350 ;
  assign n9352 = n9348 & n9350 ;
  assign n9353 = ~n9351 & ~n9352 ;
  assign n9356 = ~n9353 & ~x164 ;
  assign n9357 = ~n9355 & ~n9356 ;
  assign n9358 = ~n9122 & ~n9128 ;
  assign n9359 = ~n9093 & ~n9095 ;
  assign n9360 = x95 & n574 ;
  assign n9361 = x93 & n673 ;
  assign n9362 = x94 & n569 ;
  assign n9363 = ~n9361 & ~n9362 ;
  assign n9364 = ~n9360 & n9363 ;
  assign n9365 = n577 & n6894 ;
  assign n9366 = n9364 & ~n9365 ;
  assign n9367 = x8 & ~n9366 ;
  assign n9368 = x8 & ~n9367 ;
  assign n9369 = ~n9366 & ~n9367 ;
  assign n9370 = ~n9368 & ~n9369 ;
  assign n9371 = ~n8914 & ~n9077 ;
  assign n9372 = ~n9074 & ~n9371 ;
  assign n9373 = ~n9058 & ~n9060 ;
  assign n9374 = ~n8987 & ~n8990 ;
  assign n9375 = x77 & n4531 ;
  assign n9376 = x75 & n4847 ;
  assign n9377 = x76 & n4526 ;
  assign n9378 = ~n9376 & ~n9377 ;
  assign n9379 = ~n9375 & n9378 ;
  assign n9380 = n1502 & n4534 ;
  assign n9381 = n9379 & ~n9380 ;
  assign n9382 = x26 & ~n9381 ;
  assign n9383 = x26 & ~n9382 ;
  assign n9384 = ~n9381 & ~n9382 ;
  assign n9385 = ~n9383 & ~n9384 ;
  assign n9386 = ~n8969 & ~n8973 ;
  assign n9387 = x74 & n5560 ;
  assign n9388 = x72 & n5943 ;
  assign n9389 = x73 & n5555 ;
  assign n9390 = ~n9388 & ~n9389 ;
  assign n9391 = ~n9387 & n9390 ;
  assign n9392 = n994 & n5563 ;
  assign n9393 = n9391 & ~n9392 ;
  assign n9394 = x29 & ~n9393 ;
  assign n9395 = x29 & ~n9394 ;
  assign n9396 = ~n9393 & ~n9394 ;
  assign n9397 = ~n9395 & ~n9396 ;
  assign n9398 = ~n8504 & ~n8954 ;
  assign n9399 = ~n8951 & ~n9398 ;
  assign n9400 = x71 & n6725 ;
  assign n9401 = x69 & n7129 ;
  assign n9402 = x70 & n6720 ;
  assign n9403 = ~n9401 & ~n9402 ;
  assign n9404 = ~n9400 & n9403 ;
  assign n9405 = n558 & n6728 ;
  assign n9406 = n9404 & ~n9405 ;
  assign n9407 = x32 & ~n9406 ;
  assign n9408 = x32 & ~n9407 ;
  assign n9409 = ~n9406 & ~n9407 ;
  assign n9410 = ~n9408 & ~n9409 ;
  assign n9411 = n8486 & n8922 ;
  assign n9412 = ~n8937 & ~n9411 ;
  assign n9413 = x68 & n8006 ;
  assign n9414 = x66 & n8474 ;
  assign n9415 = x67 & n8001 ;
  assign n9416 = ~n9414 & ~n9415 ;
  assign n9417 = ~n9413 & n9416 ;
  assign n9418 = n317 & n8009 ;
  assign n9419 = n9417 & ~n9418 ;
  assign n9420 = x35 & ~n9419 ;
  assign n9421 = x35 & ~n9420 ;
  assign n9422 = ~n9419 & ~n9420 ;
  assign n9423 = ~n9421 & ~n9422 ;
  assign n9424 = x38 & ~n8922 ;
  assign n9425 = ~x36 & x37 ;
  assign n9426 = x36 & ~x37 ;
  assign n9427 = ~n9425 & ~n9426 ;
  assign n9428 = n8921 & ~n9427 ;
  assign n9429 = x64 & n9428 ;
  assign n9430 = ~x37 & x38 ;
  assign n9431 = x37 & ~x38 ;
  assign n9432 = ~n9430 & ~n9431 ;
  assign n9433 = ~n8921 & n9432 ;
  assign n9434 = x65 & n9433 ;
  assign n9435 = ~n9429 & ~n9434 ;
  assign n9436 = ~n8921 & ~n9432 ;
  assign n9437 = ~n152 & n9436 ;
  assign n9438 = n9435 & ~n9437 ;
  assign n9439 = x38 & ~n9438 ;
  assign n9440 = x38 & ~n9439 ;
  assign n9441 = ~n9438 & ~n9439 ;
  assign n9442 = ~n9440 & ~n9441 ;
  assign n9443 = n9424 & ~n9442 ;
  assign n9444 = ~n9424 & n9442 ;
  assign n9445 = ~n9443 & ~n9444 ;
  assign n9446 = n9423 & ~n9445 ;
  assign n9447 = ~n9423 & n9445 ;
  assign n9448 = ~n9446 & ~n9447 ;
  assign n9449 = ~n9412 & n9448 ;
  assign n9450 = n9412 & ~n9448 ;
  assign n9451 = ~n9449 & ~n9450 ;
  assign n9452 = n9410 & ~n9451 ;
  assign n9453 = ~n9410 & n9451 ;
  assign n9454 = ~n9452 & ~n9453 ;
  assign n9455 = ~n9399 & n9454 ;
  assign n9456 = n9399 & ~n9454 ;
  assign n9457 = ~n9455 & ~n9456 ;
  assign n9458 = n9397 & ~n9457 ;
  assign n9459 = ~n9397 & n9457 ;
  assign n9460 = ~n9458 & ~n9459 ;
  assign n9461 = ~n9386 & n9460 ;
  assign n9462 = n9386 & ~n9460 ;
  assign n9463 = ~n9461 & ~n9462 ;
  assign n9464 = n9385 & ~n9463 ;
  assign n9465 = ~n9385 & n9463 ;
  assign n9466 = ~n9464 & ~n9465 ;
  assign n9467 = ~n9374 & n9466 ;
  assign n9468 = n9374 & ~n9466 ;
  assign n9469 = ~n9467 & ~n9468 ;
  assign n9470 = x80 & n3589 ;
  assign n9471 = x78 & n3878 ;
  assign n9472 = x79 & n3584 ;
  assign n9473 = ~n9471 & ~n9472 ;
  assign n9474 = ~n9470 & n9473 ;
  assign n9475 = n2028 & n3592 ;
  assign n9476 = n9474 & ~n9475 ;
  assign n9477 = x23 & ~n9476 ;
  assign n9478 = x23 & ~n9477 ;
  assign n9479 = ~n9476 & ~n9477 ;
  assign n9480 = ~n9478 & ~n9479 ;
  assign n9481 = n9469 & ~n9480 ;
  assign n9482 = n9469 & ~n9481 ;
  assign n9483 = ~n9480 & ~n9481 ;
  assign n9484 = ~n9482 & ~n9483 ;
  assign n9485 = ~n8917 & ~n9007 ;
  assign n9486 = ~n9004 & ~n9485 ;
  assign n9487 = n9484 & n9486 ;
  assign n9488 = ~n9484 & ~n9486 ;
  assign n9489 = ~n9487 & ~n9488 ;
  assign n9490 = x83 & n2751 ;
  assign n9491 = x81 & n3020 ;
  assign n9492 = x82 & n2746 ;
  assign n9493 = ~n9491 & ~n9492 ;
  assign n9494 = ~n9490 & n9493 ;
  assign n9495 = n2754 & n2843 ;
  assign n9496 = n9494 & ~n9495 ;
  assign n9497 = x20 & ~n9496 ;
  assign n9498 = x20 & ~n9497 ;
  assign n9499 = ~n9496 & ~n9497 ;
  assign n9500 = ~n9498 & ~n9499 ;
  assign n9501 = n9489 & ~n9500 ;
  assign n9502 = n9489 & ~n9501 ;
  assign n9503 = ~n9500 & ~n9501 ;
  assign n9504 = ~n9502 & ~n9503 ;
  assign n9505 = ~n9022 & ~n9026 ;
  assign n9506 = n9504 & n9505 ;
  assign n9507 = ~n9504 & ~n9505 ;
  assign n9508 = ~n9506 & ~n9507 ;
  assign n9509 = x86 & n2093 ;
  assign n9510 = x84 & n2275 ;
  assign n9511 = x85 & n2088 ;
  assign n9512 = ~n9510 & ~n9511 ;
  assign n9513 = ~n9509 & n9512 ;
  assign n9514 = n2096 & n3686 ;
  assign n9515 = n9513 & ~n9514 ;
  assign n9516 = x17 & ~n9515 ;
  assign n9517 = x17 & ~n9516 ;
  assign n9518 = ~n9515 & ~n9516 ;
  assign n9519 = ~n9517 & ~n9518 ;
  assign n9520 = n9508 & ~n9519 ;
  assign n9521 = n9508 & ~n9520 ;
  assign n9522 = ~n9519 & ~n9520 ;
  assign n9523 = ~n9521 & ~n9522 ;
  assign n9524 = ~n8585 & ~n9042 ;
  assign n9525 = ~n9039 & ~n9524 ;
  assign n9526 = n9523 & n9525 ;
  assign n9527 = ~n9523 & ~n9525 ;
  assign n9528 = ~n9526 & ~n9527 ;
  assign n9529 = x89 & n1434 ;
  assign n9530 = x87 & n1646 ;
  assign n9531 = x88 & n1429 ;
  assign n9532 = ~n9530 & ~n9531 ;
  assign n9533 = ~n9529 & n9532 ;
  assign n9534 = n1437 & n4488 ;
  assign n9535 = n9533 & ~n9534 ;
  assign n9536 = x14 & ~n9535 ;
  assign n9537 = x14 & ~n9536 ;
  assign n9538 = ~n9535 & ~n9536 ;
  assign n9539 = ~n9537 & ~n9538 ;
  assign n9540 = n9528 & ~n9539 ;
  assign n9541 = ~n9528 & n9539 ;
  assign n9542 = ~n9373 & ~n9541 ;
  assign n9543 = ~n9540 & n9542 ;
  assign n9544 = ~n9373 & ~n9543 ;
  assign n9545 = ~n9540 & ~n9543 ;
  assign n9546 = ~n9541 & n9545 ;
  assign n9547 = ~n9544 & ~n9546 ;
  assign n9548 = x92 & n945 ;
  assign n9549 = x90 & n1099 ;
  assign n9550 = x91 & n940 ;
  assign n9551 = ~n9549 & ~n9550 ;
  assign n9552 = ~n9548 & n9551 ;
  assign n9553 = n948 & n5710 ;
  assign n9554 = n9552 & ~n9553 ;
  assign n9555 = x11 & ~n9554 ;
  assign n9556 = x11 & ~n9555 ;
  assign n9557 = ~n9554 & ~n9555 ;
  assign n9558 = ~n9556 & ~n9557 ;
  assign n9559 = n9547 & n9558 ;
  assign n9560 = ~n9547 & ~n9558 ;
  assign n9561 = ~n9559 & ~n9560 ;
  assign n9562 = ~n9372 & n9561 ;
  assign n9563 = n9372 & ~n9561 ;
  assign n9564 = ~n9562 & ~n9563 ;
  assign n9565 = n9370 & ~n9564 ;
  assign n9566 = ~n9370 & n9564 ;
  assign n9567 = ~n9565 & ~n9566 ;
  assign n9568 = ~n9359 & n9567 ;
  assign n9569 = n9359 & ~n9567 ;
  assign n9570 = ~n9568 & ~n9569 ;
  assign n9571 = x98 & n293 ;
  assign n9572 = x96 & n373 ;
  assign n9573 = x97 & n288 ;
  assign n9574 = ~n9572 & ~n9573 ;
  assign n9575 = ~n9571 & n9574 ;
  assign n9576 = n296 & n8196 ;
  assign n9577 = n9575 & ~n9576 ;
  assign n9578 = x5 & ~n9577 ;
  assign n9579 = x5 & ~n9578 ;
  assign n9580 = ~n9577 & ~n9578 ;
  assign n9581 = ~n9579 & ~n9580 ;
  assign n9582 = n9570 & ~n9581 ;
  assign n9583 = n9570 & ~n9582 ;
  assign n9584 = ~n9581 & ~n9582 ;
  assign n9585 = ~n9583 & ~n9584 ;
  assign n9586 = ~n9098 & ~n9101 ;
  assign n9587 = n9585 & n9586 ;
  assign n9588 = ~n9585 & ~n9586 ;
  assign n9589 = ~n9587 & ~n9588 ;
  assign n9590 = x101 & n146 ;
  assign n9591 = x99 & n182 ;
  assign n9592 = x100 & n141 ;
  assign n9593 = ~n9591 & ~n9592 ;
  assign n9594 = ~n9590 & n9593 ;
  assign n9595 = ~n9111 & ~n9113 ;
  assign n9596 = ~x100 & ~x101 ;
  assign n9597 = x100 & x101 ;
  assign n9598 = ~n9596 & ~n9597 ;
  assign n9599 = ~n9595 & n9598 ;
  assign n9600 = n9595 & ~n9598 ;
  assign n9601 = ~n9599 & ~n9600 ;
  assign n9602 = n149 & n9601 ;
  assign n9603 = n9594 & ~n9602 ;
  assign n9604 = x2 & ~n9603 ;
  assign n9605 = x2 & ~n9604 ;
  assign n9606 = ~n9603 & ~n9604 ;
  assign n9607 = ~n9605 & ~n9606 ;
  assign n9608 = ~n9589 & n9607 ;
  assign n9609 = n9589 & ~n9607 ;
  assign n9610 = ~n9608 & ~n9609 ;
  assign n9611 = ~n9358 & n9610 ;
  assign n9612 = n9358 & ~n9610 ;
  assign n9613 = ~n9611 & ~n9612 ;
  assign n9858 = n9613 & x165 ;
  assign n9614 = ~n9345 & ~n9351 ;
  assign n9615 = ~n9319 & ~n9321 ;
  assign n9616 = ~x95 & n574 ;
  assign n9617 = ~x93 & n673 ;
  assign n9618 = ~x94 & n569 ;
  assign n9619 = ~n9617 & ~n9618 ;
  assign n9620 = ~n9616 & n9619 ;
  assign n9621 = n577 & n7100 ;
  assign n9622 = n9620 & ~n9621 ;
  assign n9623 = ~x8 & ~n9622 ;
  assign n9624 = ~x8 & ~n9623 ;
  assign n9625 = ~n9622 & ~n9623 ;
  assign n9626 = ~n9624 & ~n9625 ;
  assign n9627 = ~n9143 & ~n9303 ;
  assign n9628 = ~n9300 & ~n9627 ;
  assign n9629 = ~n9284 & ~n9286 ;
  assign n9630 = ~n9213 & ~n9216 ;
  assign n9631 = ~x77 & n4531 ;
  assign n9632 = ~x75 & n4847 ;
  assign n9633 = ~x76 & n4526 ;
  assign n9634 = ~n9632 & ~n9633 ;
  assign n9635 = ~n9631 & n9634 ;
  assign n9636 = n1594 & n4534 ;
  assign n9637 = n9635 & ~n9636 ;
  assign n9638 = ~x26 & ~n9637 ;
  assign n9639 = ~x26 & ~n9638 ;
  assign n9640 = ~n9637 & ~n9638 ;
  assign n9641 = ~n9639 & ~n9640 ;
  assign n9642 = ~n9195 & ~n9199 ;
  assign n9643 = ~x74 & n5560 ;
  assign n9644 = ~x72 & n5943 ;
  assign n9645 = ~x73 & n5555 ;
  assign n9646 = ~n9644 & ~n9645 ;
  assign n9647 = ~n9643 & n9646 ;
  assign n9648 = n1066 & n5563 ;
  assign n9649 = n9647 & ~n9648 ;
  assign n9650 = ~x29 & ~n9649 ;
  assign n9651 = ~x29 & ~n9650 ;
  assign n9652 = ~n9649 & ~n9650 ;
  assign n9653 = ~n9651 & ~n9652 ;
  assign n9654 = ~n8732 & ~n9180 ;
  assign n9655 = ~n9177 & ~n9654 ;
  assign n9656 = ~x71 & n6725 ;
  assign n9657 = ~x69 & n7129 ;
  assign n9658 = ~x70 & n6720 ;
  assign n9659 = ~n9657 & ~n9658 ;
  assign n9660 = ~n9656 & n9659 ;
  assign n9661 = n622 & n6728 ;
  assign n9662 = n9660 & ~n9661 ;
  assign n9663 = ~x32 & ~n9662 ;
  assign n9664 = ~x32 & ~n9663 ;
  assign n9665 = ~n9662 & ~n9663 ;
  assign n9666 = ~n9664 & ~n9665 ;
  assign n9667 = n8714 & n9148 ;
  assign n9668 = ~n9163 & ~n9667 ;
  assign n9669 = ~x68 & n8006 ;
  assign n9670 = ~x66 & n8474 ;
  assign n9671 = ~x67 & n8001 ;
  assign n9672 = ~n9670 & ~n9671 ;
  assign n9673 = ~n9669 & n9672 ;
  assign n9674 = n352 & n8009 ;
  assign n9675 = n9673 & ~n9674 ;
  assign n9676 = ~x35 & ~n9675 ;
  assign n9677 = ~x35 & ~n9676 ;
  assign n9678 = ~n9675 & ~n9676 ;
  assign n9679 = ~n9677 & ~n9678 ;
  assign n9680 = ~x38 & ~n9148 ;
  assign n9681 = ~x64 & n9428 ;
  assign n9682 = ~x65 & n9433 ;
  assign n9683 = ~n9681 & ~n9682 ;
  assign n9684 = ~n9437 & n9683 ;
  assign n9685 = ~x38 & ~n9684 ;
  assign n9686 = ~x38 & ~n9685 ;
  assign n9687 = ~n9684 & ~n9685 ;
  assign n9688 = ~n9686 & ~n9687 ;
  assign n9689 = n9680 & ~n9688 ;
  assign n9690 = ~n9680 & n9688 ;
  assign n9691 = ~n9689 & ~n9690 ;
  assign n9692 = n9679 & ~n9691 ;
  assign n9693 = ~n9679 & n9691 ;
  assign n9694 = ~n9692 & ~n9693 ;
  assign n9695 = ~n9668 & n9694 ;
  assign n9696 = n9668 & ~n9694 ;
  assign n9697 = ~n9695 & ~n9696 ;
  assign n9698 = n9666 & ~n9697 ;
  assign n9699 = ~n9666 & n9697 ;
  assign n9700 = ~n9698 & ~n9699 ;
  assign n9701 = ~n9655 & n9700 ;
  assign n9702 = n9655 & ~n9700 ;
  assign n9703 = ~n9701 & ~n9702 ;
  assign n9704 = n9653 & ~n9703 ;
  assign n9705 = ~n9653 & n9703 ;
  assign n9706 = ~n9704 & ~n9705 ;
  assign n9707 = ~n9642 & n9706 ;
  assign n9708 = n9642 & ~n9706 ;
  assign n9709 = ~n9707 & ~n9708 ;
  assign n9710 = n9641 & ~n9709 ;
  assign n9711 = ~n9641 & n9709 ;
  assign n9712 = ~n9710 & ~n9711 ;
  assign n9713 = ~n9630 & n9712 ;
  assign n9714 = n9630 & ~n9712 ;
  assign n9715 = ~n9713 & ~n9714 ;
  assign n9716 = ~x80 & n3589 ;
  assign n9717 = ~x78 & n3878 ;
  assign n9718 = ~x79 & n3584 ;
  assign n9719 = ~n9717 & ~n9718 ;
  assign n9720 = ~n9716 & n9719 ;
  assign n9721 = n2145 & n3592 ;
  assign n9722 = n9720 & ~n9721 ;
  assign n9723 = ~x23 & ~n9722 ;
  assign n9724 = ~x23 & ~n9723 ;
  assign n9725 = ~n9722 & ~n9723 ;
  assign n9726 = ~n9724 & ~n9725 ;
  assign n9727 = n9715 & ~n9726 ;
  assign n9728 = n9715 & ~n9727 ;
  assign n9729 = ~n9726 & ~n9727 ;
  assign n9730 = ~n9728 & ~n9729 ;
  assign n9731 = ~n9146 & ~n9233 ;
  assign n9732 = ~n9230 & ~n9731 ;
  assign n9733 = n9730 & n9732 ;
  assign n9734 = ~n9730 & ~n9732 ;
  assign n9735 = ~n9733 & ~n9734 ;
  assign n9736 = ~x83 & n2751 ;
  assign n9737 = ~x81 & n3020 ;
  assign n9738 = ~x82 & n2746 ;
  assign n9739 = ~n9737 & ~n9738 ;
  assign n9740 = ~n9736 & n9739 ;
  assign n9741 = n2754 & n2972 ;
  assign n9742 = n9740 & ~n9741 ;
  assign n9743 = ~x20 & ~n9742 ;
  assign n9744 = ~x20 & ~n9743 ;
  assign n9745 = ~n9742 & ~n9743 ;
  assign n9746 = ~n9744 & ~n9745 ;
  assign n9747 = n9735 & ~n9746 ;
  assign n9748 = n9735 & ~n9747 ;
  assign n9749 = ~n9746 & ~n9747 ;
  assign n9750 = ~n9748 & ~n9749 ;
  assign n9751 = ~n9248 & ~n9252 ;
  assign n9752 = n9750 & n9751 ;
  assign n9753 = ~n9750 & ~n9751 ;
  assign n9754 = ~n9752 & ~n9753 ;
  assign n9755 = ~x86 & n2093 ;
  assign n9756 = ~x84 & n2275 ;
  assign n9757 = ~x85 & n2088 ;
  assign n9758 = ~n9756 & ~n9757 ;
  assign n9759 = ~n9755 & n9758 ;
  assign n9760 = n2096 & n3832 ;
  assign n9761 = n9759 & ~n9760 ;
  assign n9762 = ~x17 & ~n9761 ;
  assign n9763 = ~x17 & ~n9762 ;
  assign n9764 = ~n9761 & ~n9762 ;
  assign n9765 = ~n9763 & ~n9764 ;
  assign n9766 = n9754 & ~n9765 ;
  assign n9767 = n9754 & ~n9766 ;
  assign n9768 = ~n9765 & ~n9766 ;
  assign n9769 = ~n9767 & ~n9768 ;
  assign n9770 = ~n8813 & ~n9268 ;
  assign n9771 = ~n9265 & ~n9770 ;
  assign n9772 = n9769 & n9771 ;
  assign n9773 = ~n9769 & ~n9771 ;
  assign n9774 = ~n9772 & ~n9773 ;
  assign n9775 = ~x89 & n1434 ;
  assign n9776 = ~x87 & n1646 ;
  assign n9777 = ~x88 & n1429 ;
  assign n9778 = ~n9776 & ~n9777 ;
  assign n9779 = ~n9775 & n9778 ;
  assign n9780 = n1437 & n4664 ;
  assign n9781 = n9779 & ~n9780 ;
  assign n9782 = ~x14 & ~n9781 ;
  assign n9783 = ~x14 & ~n9782 ;
  assign n9784 = ~n9781 & ~n9782 ;
  assign n9785 = ~n9783 & ~n9784 ;
  assign n9786 = n9774 & ~n9785 ;
  assign n9787 = ~n9774 & n9785 ;
  assign n9788 = ~n9629 & ~n9787 ;
  assign n9789 = ~n9786 & n9788 ;
  assign n9790 = ~n9629 & ~n9789 ;
  assign n9791 = ~n9786 & ~n9789 ;
  assign n9792 = ~n9787 & n9791 ;
  assign n9793 = ~n9790 & ~n9792 ;
  assign n9794 = ~x92 & n945 ;
  assign n9795 = ~x90 & n1099 ;
  assign n9796 = ~x91 & n940 ;
  assign n9797 = ~n9795 & ~n9796 ;
  assign n9798 = ~n9794 & n9797 ;
  assign n9799 = n948 & n5896 ;
  assign n9800 = n9798 & ~n9799 ;
  assign n9801 = ~x11 & ~n9800 ;
  assign n9802 = ~x11 & ~n9801 ;
  assign n9803 = ~n9800 & ~n9801 ;
  assign n9804 = ~n9802 & ~n9803 ;
  assign n9805 = n9793 & n9804 ;
  assign n9806 = ~n9793 & ~n9804 ;
  assign n9807 = ~n9805 & ~n9806 ;
  assign n9808 = ~n9628 & n9807 ;
  assign n9809 = n9628 & ~n9807 ;
  assign n9810 = ~n9808 & ~n9809 ;
  assign n9811 = n9626 & ~n9810 ;
  assign n9812 = ~n9626 & n9810 ;
  assign n9813 = ~n9811 & ~n9812 ;
  assign n9814 = ~n9615 & n9813 ;
  assign n9815 = n9615 & ~n9813 ;
  assign n9816 = ~n9814 & ~n9815 ;
  assign n9817 = ~x98 & n293 ;
  assign n9818 = ~x96 & n373 ;
  assign n9819 = ~x97 & n288 ;
  assign n9820 = ~n9818 & ~n9819 ;
  assign n9821 = ~n9817 & n9820 ;
  assign n9822 = n296 & n8426 ;
  assign n9823 = n9821 & ~n9822 ;
  assign n9824 = ~x5 & ~n9823 ;
  assign n9825 = ~x5 & ~n9824 ;
  assign n9826 = ~n9823 & ~n9824 ;
  assign n9827 = ~n9825 & ~n9826 ;
  assign n9828 = n9816 & ~n9827 ;
  assign n9829 = n9816 & ~n9828 ;
  assign n9830 = ~n9827 & ~n9828 ;
  assign n9831 = ~n9829 & ~n9830 ;
  assign n9832 = ~n9324 & ~n9327 ;
  assign n9833 = n9831 & n9832 ;
  assign n9834 = ~n9831 & ~n9832 ;
  assign n9835 = ~n9833 & ~n9834 ;
  assign n9836 = ~x101 & n164 ;
  assign n9837 = ~x99 & n205 ;
  assign n9838 = ~x100 & n162 ;
  assign n9839 = ~n9837 & ~n9838 ;
  assign n9840 = ~n9836 & n9839 ;
  assign n9841 = ~n9110 & ~n9336 ;
  assign n9842 = n9598 & ~n9841 ;
  assign n9843 = ~n9598 & n9841 ;
  assign n9844 = ~n9842 & ~n9843 ;
  assign n9845 = n167 & n9844 ;
  assign n9846 = n9840 & ~n9845 ;
  assign n9847 = ~x2 & ~n9846 ;
  assign n9848 = ~x2 & ~n9847 ;
  assign n9849 = ~n9846 & ~n9847 ;
  assign n9850 = ~n9848 & ~n9849 ;
  assign n9851 = ~n9835 & n9850 ;
  assign n9852 = n9835 & ~n9850 ;
  assign n9853 = ~n9851 & ~n9852 ;
  assign n9854 = ~n9614 & n9853 ;
  assign n9855 = n9614 & ~n9853 ;
  assign n9856 = ~n9854 & ~n9855 ;
  assign n9859 = ~n9856 & ~x165 ;
  assign n9860 = ~n9858 & ~n9859 ;
  assign n9861 = ~n9582 & ~n9588 ;
  assign n9862 = x99 & n293 ;
  assign n9863 = x97 & n373 ;
  assign n9864 = x98 & n288 ;
  assign n9865 = ~n9863 & ~n9864 ;
  assign n9866 = ~n9862 & n9865 ;
  assign n9867 = n296 & n8660 ;
  assign n9868 = n9866 & ~n9867 ;
  assign n9869 = x5 & ~n9868 ;
  assign n9870 = x5 & ~n9869 ;
  assign n9871 = ~n9868 & ~n9869 ;
  assign n9872 = ~n9870 & ~n9871 ;
  assign n9873 = ~n9566 & ~n9568 ;
  assign n9874 = x96 & n574 ;
  assign n9875 = x94 & n673 ;
  assign n9876 = x95 & n569 ;
  assign n9877 = ~n9875 & ~n9876 ;
  assign n9878 = ~n9874 & n9877 ;
  assign n9879 = n577 & n7321 ;
  assign n9880 = n9878 & ~n9879 ;
  assign n9881 = x8 & ~n9880 ;
  assign n9882 = x8 & ~n9881 ;
  assign n9883 = ~n9880 & ~n9881 ;
  assign n9884 = ~n9882 & ~n9883 ;
  assign n9885 = ~n9560 & ~n9562 ;
  assign n9886 = x93 & n945 ;
  assign n9887 = x91 & n1099 ;
  assign n9888 = x92 & n940 ;
  assign n9889 = ~n9887 & ~n9888 ;
  assign n9890 = ~n9886 & n9889 ;
  assign n9891 = n948 & n6094 ;
  assign n9892 = n9890 & ~n9891 ;
  assign n9893 = x11 & ~n9892 ;
  assign n9894 = x11 & ~n9893 ;
  assign n9895 = ~n9892 & ~n9893 ;
  assign n9896 = ~n9894 & ~n9895 ;
  assign n9897 = ~n9520 & ~n9527 ;
  assign n9898 = ~n9465 & ~n9467 ;
  assign n9899 = ~n9459 & ~n9461 ;
  assign n9900 = x75 & n5560 ;
  assign n9901 = x73 & n5943 ;
  assign n9902 = x74 & n5555 ;
  assign n9903 = ~n9901 & ~n9902 ;
  assign n9904 = ~n9900 & n9903 ;
  assign n9905 = n1150 & n5563 ;
  assign n9906 = n9904 & ~n9905 ;
  assign n9907 = x29 & ~n9906 ;
  assign n9908 = x29 & ~n9907 ;
  assign n9909 = ~n9906 & ~n9907 ;
  assign n9910 = ~n9908 & ~n9909 ;
  assign n9911 = ~n9453 & ~n9455 ;
  assign n9912 = ~n9447 & ~n9449 ;
  assign n9913 = x66 & n9433 ;
  assign n9914 = n8921 & ~n9432 ;
  assign n9915 = n9427 & n9914 ;
  assign n9916 = x64 & n9915 ;
  assign n9917 = x65 & n9428 ;
  assign n9918 = ~n9916 & ~n9917 ;
  assign n9919 = ~n9913 & n9918 ;
  assign n9920 = n194 & n9436 ;
  assign n9921 = n9919 & ~n9920 ;
  assign n9922 = x38 & ~n9921 ;
  assign n9923 = x38 & ~n9922 ;
  assign n9924 = ~n9921 & ~n9922 ;
  assign n9925 = ~n9923 & ~n9924 ;
  assign n9926 = ~n9443 & n9925 ;
  assign n9927 = n9443 & ~n9925 ;
  assign n9928 = ~n9926 & ~n9927 ;
  assign n9929 = x69 & n8006 ;
  assign n9930 = x67 & n8474 ;
  assign n9931 = x68 & n8001 ;
  assign n9932 = ~n9930 & ~n9931 ;
  assign n9933 = ~n9929 & n9932 ;
  assign n9934 = n398 & n8009 ;
  assign n9935 = n9933 & ~n9934 ;
  assign n9936 = x35 & ~n9935 ;
  assign n9937 = x35 & ~n9936 ;
  assign n9938 = ~n9935 & ~n9936 ;
  assign n9939 = ~n9937 & ~n9938 ;
  assign n9940 = n9928 & ~n9939 ;
  assign n9941 = n9928 & ~n9940 ;
  assign n9942 = ~n9939 & ~n9940 ;
  assign n9943 = ~n9941 & ~n9942 ;
  assign n9944 = ~n9912 & n9943 ;
  assign n9945 = n9912 & ~n9943 ;
  assign n9946 = ~n9944 & ~n9945 ;
  assign n9947 = x72 & n6725 ;
  assign n9948 = x70 & n7129 ;
  assign n9949 = x71 & n6720 ;
  assign n9950 = ~n9948 & ~n9949 ;
  assign n9951 = ~n9947 & n9950 ;
  assign n9952 = n717 & n6728 ;
  assign n9953 = n9951 & ~n9952 ;
  assign n9954 = x32 & ~n9953 ;
  assign n9955 = x32 & ~n9954 ;
  assign n9956 = ~n9953 & ~n9954 ;
  assign n9957 = ~n9955 & ~n9956 ;
  assign n9958 = ~n9946 & ~n9957 ;
  assign n9959 = n9946 & n9957 ;
  assign n9960 = ~n9958 & ~n9959 ;
  assign n9961 = ~n9911 & n9960 ;
  assign n9962 = n9911 & ~n9960 ;
  assign n9963 = ~n9961 & ~n9962 ;
  assign n9964 = ~n9910 & n9963 ;
  assign n9965 = ~n9910 & ~n9964 ;
  assign n9966 = n9963 & ~n9964 ;
  assign n9967 = ~n9965 & ~n9966 ;
  assign n9968 = ~n9899 & ~n9967 ;
  assign n9969 = ~n9899 & ~n9968 ;
  assign n9970 = ~n9967 & ~n9968 ;
  assign n9971 = ~n9969 & ~n9970 ;
  assign n9972 = x78 & n4531 ;
  assign n9973 = x76 & n4847 ;
  assign n9974 = x77 & n4526 ;
  assign n9975 = ~n9973 & ~n9974 ;
  assign n9976 = ~n9972 & n9975 ;
  assign n9977 = n1624 & n4534 ;
  assign n9978 = n9976 & ~n9977 ;
  assign n9979 = x26 & ~n9978 ;
  assign n9980 = x26 & ~n9979 ;
  assign n9981 = ~n9978 & ~n9979 ;
  assign n9982 = ~n9980 & ~n9981 ;
  assign n9983 = n9971 & n9982 ;
  assign n9984 = ~n9971 & ~n9982 ;
  assign n9985 = ~n9983 & ~n9984 ;
  assign n9986 = ~n9898 & n9985 ;
  assign n9987 = n9898 & ~n9985 ;
  assign n9988 = ~n9986 & ~n9987 ;
  assign n9989 = x81 & n3589 ;
  assign n9990 = x79 & n3878 ;
  assign n9991 = x80 & n3584 ;
  assign n9992 = ~n9990 & ~n9991 ;
  assign n9993 = ~n9989 & n9992 ;
  assign n9994 = n2348 & n3592 ;
  assign n9995 = n9993 & ~n9994 ;
  assign n9996 = x23 & ~n9995 ;
  assign n9997 = x23 & ~n9996 ;
  assign n9998 = ~n9995 & ~n9996 ;
  assign n9999 = ~n9997 & ~n9998 ;
  assign n10000 = n9988 & ~n9999 ;
  assign n10001 = n9988 & ~n10000 ;
  assign n10002 = ~n9999 & ~n10000 ;
  assign n10003 = ~n10001 & ~n10002 ;
  assign n10004 = ~n9481 & ~n9488 ;
  assign n10005 = n10003 & n10004 ;
  assign n10006 = ~n10003 & ~n10004 ;
  assign n10007 = ~n10005 & ~n10006 ;
  assign n10008 = x84 & n2751 ;
  assign n10009 = x82 & n3020 ;
  assign n10010 = x83 & n2746 ;
  assign n10011 = ~n10009 & ~n10010 ;
  assign n10012 = ~n10008 & n10011 ;
  assign n10013 = n2754 & n3114 ;
  assign n10014 = n10012 & ~n10013 ;
  assign n10015 = x20 & ~n10014 ;
  assign n10016 = x20 & ~n10015 ;
  assign n10017 = ~n10014 & ~n10015 ;
  assign n10018 = ~n10016 & ~n10017 ;
  assign n10019 = n10007 & ~n10018 ;
  assign n10020 = n10007 & ~n10019 ;
  assign n10021 = ~n10018 & ~n10019 ;
  assign n10022 = ~n10020 & ~n10021 ;
  assign n10023 = ~n9501 & ~n9507 ;
  assign n10024 = n10022 & n10023 ;
  assign n10025 = ~n10022 & ~n10023 ;
  assign n10026 = ~n10024 & ~n10025 ;
  assign n10027 = x87 & n2093 ;
  assign n10028 = x85 & n2275 ;
  assign n10029 = x86 & n2088 ;
  assign n10030 = ~n10028 & ~n10029 ;
  assign n10031 = ~n10027 & n10030 ;
  assign n10032 = n2096 & n3991 ;
  assign n10033 = n10031 & ~n10032 ;
  assign n10034 = x17 & ~n10033 ;
  assign n10035 = x17 & ~n10034 ;
  assign n10036 = ~n10033 & ~n10034 ;
  assign n10037 = ~n10035 & ~n10036 ;
  assign n10038 = n10026 & ~n10037 ;
  assign n10039 = ~n10026 & n10037 ;
  assign n10040 = ~n9897 & ~n10039 ;
  assign n10041 = ~n10038 & n10040 ;
  assign n10042 = ~n9897 & ~n10041 ;
  assign n10043 = ~n10038 & ~n10041 ;
  assign n10044 = ~n10039 & n10043 ;
  assign n10045 = ~n10042 & ~n10044 ;
  assign n10046 = x90 & n1434 ;
  assign n10047 = x88 & n1646 ;
  assign n10048 = x89 & n1429 ;
  assign n10049 = ~n10047 & ~n10048 ;
  assign n10050 = ~n10046 & n10049 ;
  assign n10051 = n1437 & n4986 ;
  assign n10052 = n10050 & ~n10051 ;
  assign n10053 = x14 & ~n10052 ;
  assign n10054 = x14 & ~n10053 ;
  assign n10055 = ~n10052 & ~n10053 ;
  assign n10056 = ~n10054 & ~n10055 ;
  assign n10057 = n10045 & n10056 ;
  assign n10058 = ~n10045 & ~n10056 ;
  assign n10059 = ~n10057 & ~n10058 ;
  assign n10060 = ~n9545 & n10059 ;
  assign n10061 = n9545 & ~n10059 ;
  assign n10062 = ~n10060 & ~n10061 ;
  assign n10063 = n9896 & ~n10062 ;
  assign n10064 = ~n9896 & n10062 ;
  assign n10065 = ~n10063 & ~n10064 ;
  assign n10066 = ~n9885 & n10065 ;
  assign n10067 = n9885 & ~n10065 ;
  assign n10068 = ~n10066 & ~n10067 ;
  assign n10069 = n9884 & ~n10068 ;
  assign n10070 = ~n9884 & n10068 ;
  assign n10071 = ~n10069 & ~n10070 ;
  assign n10072 = ~n9873 & n10071 ;
  assign n10073 = n9873 & ~n10071 ;
  assign n10074 = ~n10072 & ~n10073 ;
  assign n10075 = n9872 & ~n10074 ;
  assign n10076 = ~n9872 & n10074 ;
  assign n10077 = ~n10075 & ~n10076 ;
  assign n10078 = ~n9861 & n10077 ;
  assign n10079 = n9861 & ~n10077 ;
  assign n10080 = ~n10078 & ~n10079 ;
  assign n10081 = x102 & n146 ;
  assign n10082 = x100 & n182 ;
  assign n10083 = x101 & n141 ;
  assign n10084 = ~n10082 & ~n10083 ;
  assign n10085 = ~n10081 & n10084 ;
  assign n10086 = ~n9597 & ~n9599 ;
  assign n10087 = ~x101 & ~x102 ;
  assign n10088 = x101 & x102 ;
  assign n10089 = ~n10087 & ~n10088 ;
  assign n10090 = ~n10086 & n10089 ;
  assign n10091 = n10086 & ~n10089 ;
  assign n10092 = ~n10090 & ~n10091 ;
  assign n10093 = n149 & n10092 ;
  assign n10094 = n10085 & ~n10093 ;
  assign n10095 = x2 & ~n10094 ;
  assign n10096 = x2 & ~n10095 ;
  assign n10097 = ~n10094 & ~n10095 ;
  assign n10098 = ~n10096 & ~n10097 ;
  assign n10099 = n10080 & ~n10098 ;
  assign n10100 = n10080 & ~n10099 ;
  assign n10101 = ~n10098 & ~n10099 ;
  assign n10102 = ~n10100 & ~n10101 ;
  assign n10103 = ~n9609 & ~n9611 ;
  assign n10104 = ~n10102 & ~n10103 ;
  assign n10105 = n10102 & n10103 ;
  assign n10106 = ~n10104 & ~n10105 ;
  assign n10349 = n10106 & x166 ;
  assign n10107 = ~n9828 & ~n9834 ;
  assign n10108 = ~x99 & n293 ;
  assign n10109 = ~x97 & n373 ;
  assign n10110 = ~x98 & n288 ;
  assign n10111 = ~n10109 & ~n10110 ;
  assign n10112 = ~n10108 & n10111 ;
  assign n10113 = n296 & n8885 ;
  assign n10114 = n10112 & ~n10113 ;
  assign n10115 = ~x5 & ~n10114 ;
  assign n10116 = ~x5 & ~n10115 ;
  assign n10117 = ~n10114 & ~n10115 ;
  assign n10118 = ~n10116 & ~n10117 ;
  assign n10119 = ~n9812 & ~n9814 ;
  assign n10120 = ~x96 & n574 ;
  assign n10121 = ~x94 & n673 ;
  assign n10122 = ~x95 & n569 ;
  assign n10123 = ~n10121 & ~n10122 ;
  assign n10124 = ~n10120 & n10123 ;
  assign n10125 = n577 & n7531 ;
  assign n10126 = n10124 & ~n10125 ;
  assign n10127 = ~x8 & ~n10126 ;
  assign n10128 = ~x8 & ~n10127 ;
  assign n10129 = ~n10126 & ~n10127 ;
  assign n10130 = ~n10128 & ~n10129 ;
  assign n10131 = ~n9806 & ~n9808 ;
  assign n10132 = ~x93 & n945 ;
  assign n10133 = ~x91 & n1099 ;
  assign n10134 = ~x92 & n940 ;
  assign n10135 = ~n10133 & ~n10134 ;
  assign n10136 = ~n10132 & n10135 ;
  assign n10137 = n948 & n6285 ;
  assign n10138 = n10136 & ~n10137 ;
  assign n10139 = ~x11 & ~n10138 ;
  assign n10140 = ~x11 & ~n10139 ;
  assign n10141 = ~n10138 & ~n10139 ;
  assign n10142 = ~n10140 & ~n10141 ;
  assign n10143 = ~n9766 & ~n9773 ;
  assign n10144 = ~n9711 & ~n9713 ;
  assign n10145 = ~n9705 & ~n9707 ;
  assign n10146 = ~x75 & n5560 ;
  assign n10147 = ~x73 & n5943 ;
  assign n10148 = ~x74 & n5555 ;
  assign n10149 = ~n10147 & ~n10148 ;
  assign n10150 = ~n10146 & n10149 ;
  assign n10151 = n1225 & n5563 ;
  assign n10152 = n10150 & ~n10151 ;
  assign n10153 = ~x29 & ~n10152 ;
  assign n10154 = ~x29 & ~n10153 ;
  assign n10155 = ~n10152 & ~n10153 ;
  assign n10156 = ~n10154 & ~n10155 ;
  assign n10157 = ~n9699 & ~n9701 ;
  assign n10158 = ~n9693 & ~n9695 ;
  assign n10159 = ~x66 & n9433 ;
  assign n10160 = ~x64 & n9915 ;
  assign n10161 = ~x65 & n9428 ;
  assign n10162 = ~n10160 & ~n10161 ;
  assign n10163 = ~n10159 & n10162 ;
  assign n10164 = n214 & n9436 ;
  assign n10165 = n10163 & ~n10164 ;
  assign n10166 = ~x38 & ~n10165 ;
  assign n10167 = ~x38 & ~n10166 ;
  assign n10168 = ~n10165 & ~n10166 ;
  assign n10169 = ~n10167 & ~n10168 ;
  assign n10170 = ~n9689 & n10169 ;
  assign n10171 = n9689 & ~n10169 ;
  assign n10172 = ~n10170 & ~n10171 ;
  assign n10173 = ~x69 & n8006 ;
  assign n10174 = ~x67 & n8474 ;
  assign n10175 = ~x68 & n8001 ;
  assign n10176 = ~n10174 & ~n10175 ;
  assign n10177 = ~n10173 & n10176 ;
  assign n10178 = n435 & n8009 ;
  assign n10179 = n10177 & ~n10178 ;
  assign n10180 = ~x35 & ~n10179 ;
  assign n10181 = ~x35 & ~n10180 ;
  assign n10182 = ~n10179 & ~n10180 ;
  assign n10183 = ~n10181 & ~n10182 ;
  assign n10184 = n10172 & ~n10183 ;
  assign n10185 = n10172 & ~n10184 ;
  assign n10186 = ~n10183 & ~n10184 ;
  assign n10187 = ~n10185 & ~n10186 ;
  assign n10188 = ~n10158 & n10187 ;
  assign n10189 = n10158 & ~n10187 ;
  assign n10190 = ~n10188 & ~n10189 ;
  assign n10191 = ~x72 & n6725 ;
  assign n10192 = ~x70 & n7129 ;
  assign n10193 = ~x71 & n6720 ;
  assign n10194 = ~n10192 & ~n10193 ;
  assign n10195 = ~n10191 & n10194 ;
  assign n10196 = n773 & n6728 ;
  assign n10197 = n10195 & ~n10196 ;
  assign n10198 = ~x32 & ~n10197 ;
  assign n10199 = ~x32 & ~n10198 ;
  assign n10200 = ~n10197 & ~n10198 ;
  assign n10201 = ~n10199 & ~n10200 ;
  assign n10202 = ~n10190 & ~n10201 ;
  assign n10203 = n10190 & n10201 ;
  assign n10204 = ~n10202 & ~n10203 ;
  assign n10205 = ~n10157 & n10204 ;
  assign n10206 = n10157 & ~n10204 ;
  assign n10207 = ~n10205 & ~n10206 ;
  assign n10208 = ~n10156 & n10207 ;
  assign n10209 = ~n10156 & ~n10208 ;
  assign n10210 = n10207 & ~n10208 ;
  assign n10211 = ~n10209 & ~n10210 ;
  assign n10212 = ~n10145 & ~n10211 ;
  assign n10213 = ~n10145 & ~n10212 ;
  assign n10214 = ~n10211 & ~n10212 ;
  assign n10215 = ~n10213 & ~n10214 ;
  assign n10216 = ~x78 & n4531 ;
  assign n10217 = ~x76 & n4847 ;
  assign n10218 = ~x77 & n4526 ;
  assign n10219 = ~n10217 & ~n10218 ;
  assign n10220 = ~n10216 & n10219 ;
  assign n10221 = n1718 & n4534 ;
  assign n10222 = n10220 & ~n10221 ;
  assign n10223 = ~x26 & ~n10222 ;
  assign n10224 = ~x26 & ~n10223 ;
  assign n10225 = ~n10222 & ~n10223 ;
  assign n10226 = ~n10224 & ~n10225 ;
  assign n10227 = n10215 & n10226 ;
  assign n10228 = ~n10215 & ~n10226 ;
  assign n10229 = ~n10227 & ~n10228 ;
  assign n10230 = ~n10144 & n10229 ;
  assign n10231 = n10144 & ~n10229 ;
  assign n10232 = ~n10230 & ~n10231 ;
  assign n10233 = ~x81 & n3589 ;
  assign n10234 = ~x79 & n3878 ;
  assign n10235 = ~x80 & n3584 ;
  assign n10236 = ~n10234 & ~n10235 ;
  assign n10237 = ~n10233 & n10236 ;
  assign n10238 = n2460 & n3592 ;
  assign n10239 = n10237 & ~n10238 ;
  assign n10240 = ~x23 & ~n10239 ;
  assign n10241 = ~x23 & ~n10240 ;
  assign n10242 = ~n10239 & ~n10240 ;
  assign n10243 = ~n10241 & ~n10242 ;
  assign n10244 = n10232 & ~n10243 ;
  assign n10245 = n10232 & ~n10244 ;
  assign n10246 = ~n10243 & ~n10244 ;
  assign n10247 = ~n10245 & ~n10246 ;
  assign n10248 = ~n9727 & ~n9734 ;
  assign n10249 = n10247 & n10248 ;
  assign n10250 = ~n10247 & ~n10248 ;
  assign n10251 = ~n10249 & ~n10250 ;
  assign n10252 = ~x84 & n2751 ;
  assign n10253 = ~x82 & n3020 ;
  assign n10254 = ~x83 & n2746 ;
  assign n10255 = ~n10253 & ~n10254 ;
  assign n10256 = ~n10252 & n10255 ;
  assign n10257 = n2754 & n3247 ;
  assign n10258 = n10256 & ~n10257 ;
  assign n10259 = ~x20 & ~n10258 ;
  assign n10260 = ~x20 & ~n10259 ;
  assign n10261 = ~n10258 & ~n10259 ;
  assign n10262 = ~n10260 & ~n10261 ;
  assign n10263 = n10251 & ~n10262 ;
  assign n10264 = n10251 & ~n10263 ;
  assign n10265 = ~n10262 & ~n10263 ;
  assign n10266 = ~n10264 & ~n10265 ;
  assign n10267 = ~n9747 & ~n9753 ;
  assign n10268 = n10266 & n10267 ;
  assign n10269 = ~n10266 & ~n10267 ;
  assign n10270 = ~n10268 & ~n10269 ;
  assign n10271 = ~x87 & n2093 ;
  assign n10272 = ~x85 & n2275 ;
  assign n10273 = ~x86 & n2088 ;
  assign n10274 = ~n10272 & ~n10273 ;
  assign n10275 = ~n10271 & n10274 ;
  assign n10276 = n2096 & n4143 ;
  assign n10277 = n10275 & ~n10276 ;
  assign n10278 = ~x17 & ~n10277 ;
  assign n10279 = ~x17 & ~n10278 ;
  assign n10280 = ~n10277 & ~n10278 ;
  assign n10281 = ~n10279 & ~n10280 ;
  assign n10282 = n10270 & ~n10281 ;
  assign n10283 = ~n10270 & n10281 ;
  assign n10284 = ~n10143 & ~n10283 ;
  assign n10285 = ~n10282 & n10284 ;
  assign n10286 = ~n10143 & ~n10285 ;
  assign n10287 = ~n10282 & ~n10285 ;
  assign n10288 = ~n10283 & n10287 ;
  assign n10289 = ~n10286 & ~n10288 ;
  assign n10290 = ~x90 & n1434 ;
  assign n10291 = ~x88 & n1646 ;
  assign n10292 = ~x89 & n1429 ;
  assign n10293 = ~n10291 & ~n10292 ;
  assign n10294 = ~n10290 & n10293 ;
  assign n10295 = n1437 & n5155 ;
  assign n10296 = n10294 & ~n10295 ;
  assign n10297 = ~x14 & ~n10296 ;
  assign n10298 = ~x14 & ~n10297 ;
  assign n10299 = ~n10296 & ~n10297 ;
  assign n10300 = ~n10298 & ~n10299 ;
  assign n10301 = n10289 & n10300 ;
  assign n10302 = ~n10289 & ~n10300 ;
  assign n10303 = ~n10301 & ~n10302 ;
  assign n10304 = ~n9791 & n10303 ;
  assign n10305 = n9791 & ~n10303 ;
  assign n10306 = ~n10304 & ~n10305 ;
  assign n10307 = n10142 & ~n10306 ;
  assign n10308 = ~n10142 & n10306 ;
  assign n10309 = ~n10307 & ~n10308 ;
  assign n10310 = ~n10131 & n10309 ;
  assign n10311 = n10131 & ~n10309 ;
  assign n10312 = ~n10310 & ~n10311 ;
  assign n10313 = n10130 & ~n10312 ;
  assign n10314 = ~n10130 & n10312 ;
  assign n10315 = ~n10313 & ~n10314 ;
  assign n10316 = ~n10119 & n10315 ;
  assign n10317 = n10119 & ~n10315 ;
  assign n10318 = ~n10316 & ~n10317 ;
  assign n10319 = n10118 & ~n10318 ;
  assign n10320 = ~n10118 & n10318 ;
  assign n10321 = ~n10319 & ~n10320 ;
  assign n10322 = ~n10107 & n10321 ;
  assign n10323 = n10107 & ~n10321 ;
  assign n10324 = ~n10322 & ~n10323 ;
  assign n10325 = ~x102 & n164 ;
  assign n10326 = ~x100 & n205 ;
  assign n10327 = ~x101 & n162 ;
  assign n10328 = ~n10326 & ~n10327 ;
  assign n10329 = ~n10325 & n10328 ;
  assign n10330 = ~n9596 & ~n9842 ;
  assign n10331 = n10089 & ~n10330 ;
  assign n10332 = ~n10089 & n10330 ;
  assign n10333 = ~n10331 & ~n10332 ;
  assign n10334 = n167 & n10333 ;
  assign n10335 = n10329 & ~n10334 ;
  assign n10336 = ~x2 & ~n10335 ;
  assign n10337 = ~x2 & ~n10336 ;
  assign n10338 = ~n10335 & ~n10336 ;
  assign n10339 = ~n10337 & ~n10338 ;
  assign n10340 = n10324 & ~n10339 ;
  assign n10341 = n10324 & ~n10340 ;
  assign n10342 = ~n10339 & ~n10340 ;
  assign n10343 = ~n10341 & ~n10342 ;
  assign n10344 = ~n9852 & ~n9854 ;
  assign n10345 = ~n10343 & ~n10344 ;
  assign n10346 = n10343 & n10344 ;
  assign n10347 = ~n10345 & ~n10346 ;
  assign n10350 = ~n10347 & ~x166 ;
  assign n10351 = ~n10349 & ~n10350 ;
  assign n10352 = ~n10076 & ~n10078 ;
  assign n10353 = ~n10070 & ~n10072 ;
  assign n10354 = ~n10064 & ~n10066 ;
  assign n10355 = ~n10058 & ~n10060 ;
  assign n10356 = ~n10000 & ~n10006 ;
  assign n10357 = ~n9984 & ~n9986 ;
  assign n10358 = x38 & ~x39 ;
  assign n10359 = ~x38 & x39 ;
  assign n10360 = ~n10358 & ~n10359 ;
  assign n10361 = x64 & ~n10360 ;
  assign n10362 = ~n9927 & n10361 ;
  assign n10363 = n9927 & ~n10361 ;
  assign n10364 = ~n10362 & ~n10363 ;
  assign n10365 = x67 & n9433 ;
  assign n10366 = x65 & n9915 ;
  assign n10367 = x66 & n9428 ;
  assign n10368 = ~n10366 & ~n10367 ;
  assign n10369 = ~n10365 & n10368 ;
  assign n10370 = n240 & n9436 ;
  assign n10371 = n10369 & ~n10370 ;
  assign n10372 = x38 & ~n10371 ;
  assign n10373 = x38 & ~n10372 ;
  assign n10374 = ~n10371 & ~n10372 ;
  assign n10375 = ~n10373 & ~n10374 ;
  assign n10376 = ~n10364 & ~n10375 ;
  assign n10377 = n10364 & n10375 ;
  assign n10378 = ~n10376 & ~n10377 ;
  assign n10379 = x70 & n8006 ;
  assign n10380 = x68 & n8474 ;
  assign n10381 = x69 & n8001 ;
  assign n10382 = ~n10380 & ~n10381 ;
  assign n10383 = ~n10379 & n10382 ;
  assign n10384 = n488 & n8009 ;
  assign n10385 = n10383 & ~n10384 ;
  assign n10386 = x35 & ~n10385 ;
  assign n10387 = x35 & ~n10386 ;
  assign n10388 = ~n10385 & ~n10386 ;
  assign n10389 = ~n10387 & ~n10388 ;
  assign n10390 = n10378 & ~n10389 ;
  assign n10391 = n10378 & ~n10390 ;
  assign n10392 = ~n10389 & ~n10390 ;
  assign n10393 = ~n10391 & ~n10392 ;
  assign n10394 = ~n9912 & ~n9943 ;
  assign n10395 = ~n9940 & ~n10394 ;
  assign n10396 = n10393 & n10395 ;
  assign n10397 = ~n10393 & ~n10395 ;
  assign n10398 = ~n10396 & ~n10397 ;
  assign n10399 = x73 & n6725 ;
  assign n10400 = x71 & n7129 ;
  assign n10401 = x72 & n6720 ;
  assign n10402 = ~n10400 & ~n10401 ;
  assign n10403 = ~n10399 & n10402 ;
  assign n10404 = n843 & n6728 ;
  assign n10405 = n10403 & ~n10404 ;
  assign n10406 = x32 & ~n10405 ;
  assign n10407 = x32 & ~n10406 ;
  assign n10408 = ~n10405 & ~n10406 ;
  assign n10409 = ~n10407 & ~n10408 ;
  assign n10410 = n10398 & ~n10409 ;
  assign n10411 = n10398 & ~n10410 ;
  assign n10412 = ~n10409 & ~n10410 ;
  assign n10413 = ~n10411 & ~n10412 ;
  assign n10414 = ~n9958 & ~n9961 ;
  assign n10415 = n10413 & n10414 ;
  assign n10416 = ~n10413 & ~n10414 ;
  assign n10417 = ~n10415 & ~n10416 ;
  assign n10418 = x76 & n5560 ;
  assign n10419 = x74 & n5943 ;
  assign n10420 = x75 & n5555 ;
  assign n10421 = ~n10419 & ~n10420 ;
  assign n10422 = ~n10418 & n10421 ;
  assign n10423 = n1311 & n5563 ;
  assign n10424 = n10422 & ~n10423 ;
  assign n10425 = x29 & ~n10424 ;
  assign n10426 = x29 & ~n10425 ;
  assign n10427 = ~n10424 & ~n10425 ;
  assign n10428 = ~n10426 & ~n10427 ;
  assign n10429 = ~n10417 & n10428 ;
  assign n10430 = n10417 & ~n10428 ;
  assign n10431 = ~n10429 & ~n10430 ;
  assign n10432 = ~n9964 & ~n9968 ;
  assign n10433 = n10431 & ~n10432 ;
  assign n10434 = ~n10431 & n10432 ;
  assign n10435 = ~n10433 & ~n10434 ;
  assign n10436 = x79 & n4531 ;
  assign n10437 = x77 & n4847 ;
  assign n10438 = x78 & n4526 ;
  assign n10439 = ~n10437 & ~n10438 ;
  assign n10440 = ~n10436 & n10439 ;
  assign n10441 = n1817 & n4534 ;
  assign n10442 = n10440 & ~n10441 ;
  assign n10443 = x26 & ~n10442 ;
  assign n10444 = x26 & ~n10443 ;
  assign n10445 = ~n10442 & ~n10443 ;
  assign n10446 = ~n10444 & ~n10445 ;
  assign n10447 = n10435 & ~n10446 ;
  assign n10448 = n10435 & ~n10447 ;
  assign n10449 = ~n10446 & ~n10447 ;
  assign n10450 = ~n10448 & ~n10449 ;
  assign n10451 = ~n10357 & n10450 ;
  assign n10452 = n10357 & ~n10450 ;
  assign n10453 = ~n10451 & ~n10452 ;
  assign n10454 = x82 & n3589 ;
  assign n10455 = x80 & n3878 ;
  assign n10456 = x81 & n3584 ;
  assign n10457 = ~n10455 & ~n10456 ;
  assign n10458 = ~n10454 & n10457 ;
  assign n10459 = n2584 & n3592 ;
  assign n10460 = n10458 & ~n10459 ;
  assign n10461 = x23 & ~n10460 ;
  assign n10462 = x23 & ~n10461 ;
  assign n10463 = ~n10460 & ~n10461 ;
  assign n10464 = ~n10462 & ~n10463 ;
  assign n10465 = ~n10453 & ~n10464 ;
  assign n10466 = n10453 & n10464 ;
  assign n10467 = ~n10465 & ~n10466 ;
  assign n10468 = n10356 & ~n10467 ;
  assign n10469 = ~n10356 & n10467 ;
  assign n10470 = ~n10468 & ~n10469 ;
  assign n10471 = x85 & n2751 ;
  assign n10472 = x83 & n3020 ;
  assign n10473 = x84 & n2746 ;
  assign n10474 = ~n10472 & ~n10473 ;
  assign n10475 = ~n10471 & n10474 ;
  assign n10476 = n2754 & n3389 ;
  assign n10477 = n10475 & ~n10476 ;
  assign n10478 = x20 & ~n10477 ;
  assign n10479 = x20 & ~n10478 ;
  assign n10480 = ~n10477 & ~n10478 ;
  assign n10481 = ~n10479 & ~n10480 ;
  assign n10482 = n10470 & ~n10481 ;
  assign n10483 = n10470 & ~n10482 ;
  assign n10484 = ~n10481 & ~n10482 ;
  assign n10485 = ~n10483 & ~n10484 ;
  assign n10486 = ~n10019 & ~n10025 ;
  assign n10487 = n10485 & n10486 ;
  assign n10488 = ~n10485 & ~n10486 ;
  assign n10489 = ~n10487 & ~n10488 ;
  assign n10490 = x88 & n2093 ;
  assign n10491 = x86 & n2275 ;
  assign n10492 = x87 & n2088 ;
  assign n10493 = ~n10491 & ~n10492 ;
  assign n10494 = ~n10490 & n10493 ;
  assign n10495 = n2096 & n4305 ;
  assign n10496 = n10494 & ~n10495 ;
  assign n10497 = x17 & ~n10496 ;
  assign n10498 = x17 & ~n10497 ;
  assign n10499 = ~n10496 & ~n10497 ;
  assign n10500 = ~n10498 & ~n10499 ;
  assign n10501 = ~n10489 & n10500 ;
  assign n10502 = n10489 & ~n10500 ;
  assign n10503 = ~n10501 & ~n10502 ;
  assign n10504 = ~n10043 & n10503 ;
  assign n10505 = n10043 & ~n10503 ;
  assign n10506 = ~n10504 & ~n10505 ;
  assign n10507 = x91 & n1434 ;
  assign n10508 = x89 & n1646 ;
  assign n10509 = x90 & n1429 ;
  assign n10510 = ~n10508 & ~n10509 ;
  assign n10511 = ~n10507 & n10510 ;
  assign n10512 = n1437 & n5336 ;
  assign n10513 = n10511 & ~n10512 ;
  assign n10514 = x14 & ~n10513 ;
  assign n10515 = x14 & ~n10514 ;
  assign n10516 = ~n10513 & ~n10514 ;
  assign n10517 = ~n10515 & ~n10516 ;
  assign n10518 = n10506 & ~n10517 ;
  assign n10519 = n10506 & ~n10518 ;
  assign n10520 = ~n10517 & ~n10518 ;
  assign n10521 = ~n10519 & ~n10520 ;
  assign n10522 = ~n10355 & n10521 ;
  assign n10523 = n10355 & ~n10521 ;
  assign n10524 = ~n10522 & ~n10523 ;
  assign n10525 = x94 & n945 ;
  assign n10526 = x92 & n1099 ;
  assign n10527 = x93 & n940 ;
  assign n10528 = ~n10526 & ~n10527 ;
  assign n10529 = ~n10525 & n10528 ;
  assign n10530 = n948 & n6483 ;
  assign n10531 = n10529 & ~n10530 ;
  assign n10532 = x11 & ~n10531 ;
  assign n10533 = x11 & ~n10532 ;
  assign n10534 = ~n10531 & ~n10532 ;
  assign n10535 = ~n10533 & ~n10534 ;
  assign n10536 = ~n10524 & ~n10535 ;
  assign n10537 = n10524 & n10535 ;
  assign n10538 = ~n10536 & ~n10537 ;
  assign n10539 = ~n10354 & n10538 ;
  assign n10540 = n10354 & ~n10538 ;
  assign n10541 = ~n10539 & ~n10540 ;
  assign n10542 = x97 & n574 ;
  assign n10543 = x95 & n673 ;
  assign n10544 = x96 & n569 ;
  assign n10545 = ~n10543 & ~n10544 ;
  assign n10546 = ~n10542 & n10545 ;
  assign n10547 = n577 & n7745 ;
  assign n10548 = n10546 & ~n10547 ;
  assign n10549 = x8 & ~n10548 ;
  assign n10550 = x8 & ~n10549 ;
  assign n10551 = ~n10548 & ~n10549 ;
  assign n10552 = ~n10550 & ~n10551 ;
  assign n10553 = n10541 & ~n10552 ;
  assign n10554 = n10541 & ~n10553 ;
  assign n10555 = ~n10552 & ~n10553 ;
  assign n10556 = ~n10554 & ~n10555 ;
  assign n10557 = ~n10353 & n10556 ;
  assign n10558 = n10353 & ~n10556 ;
  assign n10559 = ~n10557 & ~n10558 ;
  assign n10560 = x100 & n293 ;
  assign n10561 = x98 & n373 ;
  assign n10562 = x99 & n288 ;
  assign n10563 = ~n10561 & ~n10562 ;
  assign n10564 = ~n10560 & n10563 ;
  assign n10565 = n296 & n9115 ;
  assign n10566 = n10564 & ~n10565 ;
  assign n10567 = x5 & ~n10566 ;
  assign n10568 = x5 & ~n10567 ;
  assign n10569 = ~n10566 & ~n10567 ;
  assign n10570 = ~n10568 & ~n10569 ;
  assign n10571 = n10559 & n10570 ;
  assign n10572 = ~n10559 & ~n10570 ;
  assign n10573 = ~n10571 & ~n10572 ;
  assign n10574 = ~n10352 & n10573 ;
  assign n10575 = n10352 & ~n10573 ;
  assign n10576 = ~n10574 & ~n10575 ;
  assign n10577 = x103 & n146 ;
  assign n10578 = x101 & n182 ;
  assign n10579 = x102 & n141 ;
  assign n10580 = ~n10578 & ~n10579 ;
  assign n10581 = ~n10577 & n10580 ;
  assign n10582 = ~n10088 & ~n10090 ;
  assign n10583 = ~x102 & ~x103 ;
  assign n10584 = x102 & x103 ;
  assign n10585 = ~n10583 & ~n10584 ;
  assign n10586 = ~n10582 & n10585 ;
  assign n10587 = n10582 & ~n10585 ;
  assign n10588 = ~n10586 & ~n10587 ;
  assign n10589 = n149 & n10588 ;
  assign n10590 = n10581 & ~n10589 ;
  assign n10591 = x2 & ~n10590 ;
  assign n10592 = x2 & ~n10591 ;
  assign n10593 = ~n10590 & ~n10591 ;
  assign n10594 = ~n10592 & ~n10593 ;
  assign n10595 = n10576 & ~n10594 ;
  assign n10596 = n10576 & ~n10595 ;
  assign n10597 = ~n10594 & ~n10595 ;
  assign n10598 = ~n10596 & ~n10597 ;
  assign n10599 = ~n10099 & ~n10104 ;
  assign n10600 = ~n10598 & ~n10599 ;
  assign n10601 = n10598 & n10599 ;
  assign n10602 = ~n10600 & ~n10601 ;
  assign n10849 = n10602 & x167 ;
  assign n10603 = ~n10320 & ~n10322 ;
  assign n10604 = ~n10314 & ~n10316 ;
  assign n10605 = ~n10308 & ~n10310 ;
  assign n10606 = ~n10302 & ~n10304 ;
  assign n10607 = ~n10244 & ~n10250 ;
  assign n10608 = ~n10228 & ~n10230 ;
  assign n10609 = ~x64 & ~n10360 ;
  assign n10610 = ~n10171 & n10609 ;
  assign n10611 = n10171 & ~n10609 ;
  assign n10612 = ~n10610 & ~n10611 ;
  assign n10613 = ~x67 & n9433 ;
  assign n10614 = ~x65 & n9915 ;
  assign n10615 = ~x66 & n9428 ;
  assign n10616 = ~n10614 & ~n10615 ;
  assign n10617 = ~n10613 & n10616 ;
  assign n10618 = n266 & n9436 ;
  assign n10619 = n10617 & ~n10618 ;
  assign n10620 = ~x38 & ~n10619 ;
  assign n10621 = ~x38 & ~n10620 ;
  assign n10622 = ~n10619 & ~n10620 ;
  assign n10623 = ~n10621 & ~n10622 ;
  assign n10624 = ~n10612 & ~n10623 ;
  assign n10625 = n10612 & n10623 ;
  assign n10626 = ~n10624 & ~n10625 ;
  assign n10627 = ~x70 & n8006 ;
  assign n10628 = ~x68 & n8474 ;
  assign n10629 = ~x69 & n8001 ;
  assign n10630 = ~n10628 & ~n10629 ;
  assign n10631 = ~n10627 & n10630 ;
  assign n10632 = n529 & n8009 ;
  assign n10633 = n10631 & ~n10632 ;
  assign n10634 = ~x35 & ~n10633 ;
  assign n10635 = ~x35 & ~n10634 ;
  assign n10636 = ~n10633 & ~n10634 ;
  assign n10637 = ~n10635 & ~n10636 ;
  assign n10638 = n10626 & ~n10637 ;
  assign n10639 = n10626 & ~n10638 ;
  assign n10640 = ~n10637 & ~n10638 ;
  assign n10641 = ~n10639 & ~n10640 ;
  assign n10642 = ~n10158 & ~n10187 ;
  assign n10643 = ~n10184 & ~n10642 ;
  assign n10644 = n10641 & n10643 ;
  assign n10645 = ~n10641 & ~n10643 ;
  assign n10646 = ~n10644 & ~n10645 ;
  assign n10647 = ~x73 & n6725 ;
  assign n10648 = ~x71 & n7129 ;
  assign n10649 = ~x72 & n6720 ;
  assign n10650 = ~n10648 & ~n10649 ;
  assign n10651 = ~n10647 & n10650 ;
  assign n10652 = n903 & n6728 ;
  assign n10653 = n10651 & ~n10652 ;
  assign n10654 = ~x32 & ~n10653 ;
  assign n10655 = ~x32 & ~n10654 ;
  assign n10656 = ~n10653 & ~n10654 ;
  assign n10657 = ~n10655 & ~n10656 ;
  assign n10658 = n10646 & ~n10657 ;
  assign n10659 = n10646 & ~n10658 ;
  assign n10660 = ~n10657 & ~n10658 ;
  assign n10661 = ~n10659 & ~n10660 ;
  assign n10662 = ~n10202 & ~n10205 ;
  assign n10663 = n10661 & n10662 ;
  assign n10664 = ~n10661 & ~n10662 ;
  assign n10665 = ~n10663 & ~n10664 ;
  assign n10666 = ~x76 & n5560 ;
  assign n10667 = ~x74 & n5943 ;
  assign n10668 = ~x75 & n5555 ;
  assign n10669 = ~n10667 & ~n10668 ;
  assign n10670 = ~n10666 & n10669 ;
  assign n10671 = n1390 & n5563 ;
  assign n10672 = n10670 & ~n10671 ;
  assign n10673 = ~x29 & ~n10672 ;
  assign n10674 = ~x29 & ~n10673 ;
  assign n10675 = ~n10672 & ~n10673 ;
  assign n10676 = ~n10674 & ~n10675 ;
  assign n10677 = ~n10665 & n10676 ;
  assign n10678 = n10665 & ~n10676 ;
  assign n10679 = ~n10677 & ~n10678 ;
  assign n10680 = ~n10208 & ~n10212 ;
  assign n10681 = n10679 & ~n10680 ;
  assign n10682 = ~n10679 & n10680 ;
  assign n10683 = ~n10681 & ~n10682 ;
  assign n10684 = ~x79 & n4531 ;
  assign n10685 = ~x77 & n4847 ;
  assign n10686 = ~x78 & n4526 ;
  assign n10687 = ~n10685 & ~n10686 ;
  assign n10688 = ~n10684 & n10687 ;
  assign n10689 = n1921 & n4534 ;
  assign n10690 = n10688 & ~n10689 ;
  assign n10691 = ~x26 & ~n10690 ;
  assign n10692 = ~x26 & ~n10691 ;
  assign n10693 = ~n10690 & ~n10691 ;
  assign n10694 = ~n10692 & ~n10693 ;
  assign n10695 = n10683 & ~n10694 ;
  assign n10696 = n10683 & ~n10695 ;
  assign n10697 = ~n10694 & ~n10695 ;
  assign n10698 = ~n10696 & ~n10697 ;
  assign n10699 = ~n10608 & n10698 ;
  assign n10700 = n10608 & ~n10698 ;
  assign n10701 = ~n10699 & ~n10700 ;
  assign n10702 = ~x82 & n3589 ;
  assign n10703 = ~x80 & n3878 ;
  assign n10704 = ~x81 & n3584 ;
  assign n10705 = ~n10703 & ~n10704 ;
  assign n10706 = ~n10702 & n10705 ;
  assign n10707 = n2697 & n3592 ;
  assign n10708 = n10706 & ~n10707 ;
  assign n10709 = ~x23 & ~n10708 ;
  assign n10710 = ~x23 & ~n10709 ;
  assign n10711 = ~n10708 & ~n10709 ;
  assign n10712 = ~n10710 & ~n10711 ;
  assign n10713 = ~n10701 & ~n10712 ;
  assign n10714 = n10701 & n10712 ;
  assign n10715 = ~n10713 & ~n10714 ;
  assign n10716 = n10607 & ~n10715 ;
  assign n10717 = ~n10607 & n10715 ;
  assign n10718 = ~n10716 & ~n10717 ;
  assign n10719 = ~x85 & n2751 ;
  assign n10720 = ~x83 & n3020 ;
  assign n10721 = ~x84 & n2746 ;
  assign n10722 = ~n10720 & ~n10721 ;
  assign n10723 = ~n10719 & n10722 ;
  assign n10724 = n2754 & n3521 ;
  assign n10725 = n10723 & ~n10724 ;
  assign n10726 = ~x20 & ~n10725 ;
  assign n10727 = ~x20 & ~n10726 ;
  assign n10728 = ~n10725 & ~n10726 ;
  assign n10729 = ~n10727 & ~n10728 ;
  assign n10730 = n10718 & ~n10729 ;
  assign n10731 = n10718 & ~n10730 ;
  assign n10732 = ~n10729 & ~n10730 ;
  assign n10733 = ~n10731 & ~n10732 ;
  assign n10734 = ~n10263 & ~n10269 ;
  assign n10735 = n10733 & n10734 ;
  assign n10736 = ~n10733 & ~n10734 ;
  assign n10737 = ~n10735 & ~n10736 ;
  assign n10738 = ~x88 & n2093 ;
  assign n10739 = ~x86 & n2275 ;
  assign n10740 = ~x87 & n2088 ;
  assign n10741 = ~n10739 & ~n10740 ;
  assign n10742 = ~n10738 & n10741 ;
  assign n10743 = n2096 & n4457 ;
  assign n10744 = n10742 & ~n10743 ;
  assign n10745 = ~x17 & ~n10744 ;
  assign n10746 = ~x17 & ~n10745 ;
  assign n10747 = ~n10744 & ~n10745 ;
  assign n10748 = ~n10746 & ~n10747 ;
  assign n10749 = ~n10737 & n10748 ;
  assign n10750 = n10737 & ~n10748 ;
  assign n10751 = ~n10749 & ~n10750 ;
  assign n10752 = ~n10287 & n10751 ;
  assign n10753 = n10287 & ~n10751 ;
  assign n10754 = ~n10752 & ~n10753 ;
  assign n10755 = ~x91 & n1434 ;
  assign n10756 = ~x89 & n1646 ;
  assign n10757 = ~x90 & n1429 ;
  assign n10758 = ~n10756 & ~n10757 ;
  assign n10759 = ~n10755 & n10758 ;
  assign n10760 = n1437 & n5507 ;
  assign n10761 = n10759 & ~n10760 ;
  assign n10762 = ~x14 & ~n10761 ;
  assign n10763 = ~x14 & ~n10762 ;
  assign n10764 = ~n10761 & ~n10762 ;
  assign n10765 = ~n10763 & ~n10764 ;
  assign n10766 = n10754 & ~n10765 ;
  assign n10767 = n10754 & ~n10766 ;
  assign n10768 = ~n10765 & ~n10766 ;
  assign n10769 = ~n10767 & ~n10768 ;
  assign n10770 = ~n10606 & n10769 ;
  assign n10771 = n10606 & ~n10769 ;
  assign n10772 = ~n10770 & ~n10771 ;
  assign n10773 = ~x94 & n945 ;
  assign n10774 = ~x92 & n1099 ;
  assign n10775 = ~x93 & n940 ;
  assign n10776 = ~n10774 & ~n10775 ;
  assign n10777 = ~n10773 & n10776 ;
  assign n10778 = n948 & n6671 ;
  assign n10779 = n10777 & ~n10778 ;
  assign n10780 = ~x11 & ~n10779 ;
  assign n10781 = ~x11 & ~n10780 ;
  assign n10782 = ~n10779 & ~n10780 ;
  assign n10783 = ~n10781 & ~n10782 ;
  assign n10784 = ~n10772 & ~n10783 ;
  assign n10785 = n10772 & n10783 ;
  assign n10786 = ~n10784 & ~n10785 ;
  assign n10787 = ~n10605 & n10786 ;
  assign n10788 = n10605 & ~n10786 ;
  assign n10789 = ~n10787 & ~n10788 ;
  assign n10790 = ~x97 & n574 ;
  assign n10791 = ~x95 & n673 ;
  assign n10792 = ~x96 & n569 ;
  assign n10793 = ~n10791 & ~n10792 ;
  assign n10794 = ~n10790 & n10793 ;
  assign n10795 = n577 & n7949 ;
  assign n10796 = n10794 & ~n10795 ;
  assign n10797 = ~x8 & ~n10796 ;
  assign n10798 = ~x8 & ~n10797 ;
  assign n10799 = ~n10796 & ~n10797 ;
  assign n10800 = ~n10798 & ~n10799 ;
  assign n10801 = n10789 & ~n10800 ;
  assign n10802 = n10789 & ~n10801 ;
  assign n10803 = ~n10800 & ~n10801 ;
  assign n10804 = ~n10802 & ~n10803 ;
  assign n10805 = ~n10604 & n10804 ;
  assign n10806 = n10604 & ~n10804 ;
  assign n10807 = ~n10805 & ~n10806 ;
  assign n10808 = ~x100 & n293 ;
  assign n10809 = ~x98 & n373 ;
  assign n10810 = ~x99 & n288 ;
  assign n10811 = ~n10809 & ~n10810 ;
  assign n10812 = ~n10808 & n10811 ;
  assign n10813 = n296 & n9338 ;
  assign n10814 = n10812 & ~n10813 ;
  assign n10815 = ~x5 & ~n10814 ;
  assign n10816 = ~x5 & ~n10815 ;
  assign n10817 = ~n10814 & ~n10815 ;
  assign n10818 = ~n10816 & ~n10817 ;
  assign n10819 = n10807 & n10818 ;
  assign n10820 = ~n10807 & ~n10818 ;
  assign n10821 = ~n10819 & ~n10820 ;
  assign n10822 = ~n10603 & n10821 ;
  assign n10823 = n10603 & ~n10821 ;
  assign n10824 = ~n10822 & ~n10823 ;
  assign n10825 = ~x103 & n164 ;
  assign n10826 = ~x101 & n205 ;
  assign n10827 = ~x102 & n162 ;
  assign n10828 = ~n10826 & ~n10827 ;
  assign n10829 = ~n10825 & n10828 ;
  assign n10830 = ~n10087 & ~n10331 ;
  assign n10831 = n10585 & ~n10830 ;
  assign n10832 = ~n10585 & n10830 ;
  assign n10833 = ~n10831 & ~n10832 ;
  assign n10834 = n167 & n10833 ;
  assign n10835 = n10829 & ~n10834 ;
  assign n10836 = ~x2 & ~n10835 ;
  assign n10837 = ~x2 & ~n10836 ;
  assign n10838 = ~n10835 & ~n10836 ;
  assign n10839 = ~n10837 & ~n10838 ;
  assign n10840 = n10824 & ~n10839 ;
  assign n10841 = n10824 & ~n10840 ;
  assign n10842 = ~n10839 & ~n10840 ;
  assign n10843 = ~n10841 & ~n10842 ;
  assign n10844 = ~n10340 & ~n10345 ;
  assign n10845 = ~n10843 & ~n10844 ;
  assign n10846 = n10843 & n10844 ;
  assign n10847 = ~n10845 & ~n10846 ;
  assign n10850 = ~n10847 & ~x167 ;
  assign n10851 = ~n10849 & ~n10850 ;
  assign n10852 = ~n10595 & ~n10600 ;
  assign n10853 = ~n10572 & ~n10574 ;
  assign n10854 = ~n10353 & ~n10556 ;
  assign n10855 = ~n10553 & ~n10854 ;
  assign n10856 = x98 & n574 ;
  assign n10857 = x96 & n673 ;
  assign n10858 = x97 & n569 ;
  assign n10859 = ~n10857 & ~n10858 ;
  assign n10860 = ~n10856 & n10859 ;
  assign n10861 = n577 & n8196 ;
  assign n10862 = n10860 & ~n10861 ;
  assign n10863 = x8 & ~n10862 ;
  assign n10864 = x8 & ~n10863 ;
  assign n10865 = ~n10862 & ~n10863 ;
  assign n10866 = ~n10864 & ~n10865 ;
  assign n10867 = ~n10536 & ~n10539 ;
  assign n10868 = ~n10355 & ~n10521 ;
  assign n10869 = ~n10518 & ~n10868 ;
  assign n10870 = x92 & n1434 ;
  assign n10871 = x90 & n1646 ;
  assign n10872 = x91 & n1429 ;
  assign n10873 = ~n10871 & ~n10872 ;
  assign n10874 = ~n10870 & n10873 ;
  assign n10875 = n1437 & n5710 ;
  assign n10876 = n10874 & ~n10875 ;
  assign n10877 = x14 & ~n10876 ;
  assign n10878 = x14 & ~n10877 ;
  assign n10879 = ~n10876 & ~n10877 ;
  assign n10880 = ~n10878 & ~n10879 ;
  assign n10881 = ~n10430 & ~n10433 ;
  assign n10882 = ~n10410 & ~n10416 ;
  assign n10883 = n9927 & n10361 ;
  assign n10884 = ~n10376 & ~n10883 ;
  assign n10885 = x68 & n9433 ;
  assign n10886 = x66 & n9915 ;
  assign n10887 = x67 & n9428 ;
  assign n10888 = ~n10886 & ~n10887 ;
  assign n10889 = ~n10885 & n10888 ;
  assign n10890 = n317 & n9436 ;
  assign n10891 = n10889 & ~n10890 ;
  assign n10892 = x38 & ~n10891 ;
  assign n10893 = x38 & ~n10892 ;
  assign n10894 = ~n10891 & ~n10892 ;
  assign n10895 = ~n10893 & ~n10894 ;
  assign n10896 = x41 & ~n10361 ;
  assign n10897 = ~x39 & x40 ;
  assign n10898 = x39 & ~x40 ;
  assign n10899 = ~n10897 & ~n10898 ;
  assign n10900 = n10360 & ~n10899 ;
  assign n10901 = x64 & n10900 ;
  assign n10902 = ~x40 & x41 ;
  assign n10903 = x40 & ~x41 ;
  assign n10904 = ~n10902 & ~n10903 ;
  assign n10905 = ~n10360 & n10904 ;
  assign n10906 = x65 & n10905 ;
  assign n10907 = ~n10901 & ~n10906 ;
  assign n10908 = ~n10360 & ~n10904 ;
  assign n10909 = ~n152 & n10908 ;
  assign n10910 = n10907 & ~n10909 ;
  assign n10911 = x41 & ~n10910 ;
  assign n10912 = x41 & ~n10911 ;
  assign n10913 = ~n10910 & ~n10911 ;
  assign n10914 = ~n10912 & ~n10913 ;
  assign n10915 = n10896 & ~n10914 ;
  assign n10916 = ~n10896 & n10914 ;
  assign n10917 = ~n10915 & ~n10916 ;
  assign n10918 = n10895 & ~n10917 ;
  assign n10919 = ~n10895 & n10917 ;
  assign n10920 = ~n10918 & ~n10919 ;
  assign n10921 = ~n10884 & n10920 ;
  assign n10922 = n10884 & ~n10920 ;
  assign n10923 = ~n10921 & ~n10922 ;
  assign n10924 = x71 & n8006 ;
  assign n10925 = x69 & n8474 ;
  assign n10926 = x70 & n8001 ;
  assign n10927 = ~n10925 & ~n10926 ;
  assign n10928 = ~n10924 & n10927 ;
  assign n10929 = n558 & n8009 ;
  assign n10930 = n10928 & ~n10929 ;
  assign n10931 = x35 & ~n10930 ;
  assign n10932 = x35 & ~n10931 ;
  assign n10933 = ~n10930 & ~n10931 ;
  assign n10934 = ~n10932 & ~n10933 ;
  assign n10935 = n10923 & ~n10934 ;
  assign n10936 = n10923 & ~n10935 ;
  assign n10937 = ~n10934 & ~n10935 ;
  assign n10938 = ~n10936 & ~n10937 ;
  assign n10939 = ~n10390 & ~n10397 ;
  assign n10940 = n10938 & n10939 ;
  assign n10941 = ~n10938 & ~n10939 ;
  assign n10942 = ~n10940 & ~n10941 ;
  assign n10943 = x74 & n6725 ;
  assign n10944 = x72 & n7129 ;
  assign n10945 = x73 & n6720 ;
  assign n10946 = ~n10944 & ~n10945 ;
  assign n10947 = ~n10943 & n10946 ;
  assign n10948 = n994 & n6728 ;
  assign n10949 = n10947 & ~n10948 ;
  assign n10950 = x32 & ~n10949 ;
  assign n10951 = x32 & ~n10950 ;
  assign n10952 = ~n10949 & ~n10950 ;
  assign n10953 = ~n10951 & ~n10952 ;
  assign n10954 = n10942 & ~n10953 ;
  assign n10955 = ~n10942 & n10953 ;
  assign n10956 = ~n10882 & ~n10955 ;
  assign n10957 = ~n10954 & n10956 ;
  assign n10958 = ~n10882 & ~n10957 ;
  assign n10959 = ~n10954 & ~n10957 ;
  assign n10960 = ~n10955 & n10959 ;
  assign n10961 = ~n10958 & ~n10960 ;
  assign n10962 = x77 & n5560 ;
  assign n10963 = x75 & n5943 ;
  assign n10964 = x76 & n5555 ;
  assign n10965 = ~n10963 & ~n10964 ;
  assign n10966 = ~n10962 & n10965 ;
  assign n10967 = n1502 & n5563 ;
  assign n10968 = n10966 & ~n10967 ;
  assign n10969 = x29 & ~n10968 ;
  assign n10970 = x29 & ~n10969 ;
  assign n10971 = ~n10968 & ~n10969 ;
  assign n10972 = ~n10970 & ~n10971 ;
  assign n10973 = n10961 & n10972 ;
  assign n10974 = ~n10961 & ~n10972 ;
  assign n10975 = ~n10973 & ~n10974 ;
  assign n10976 = ~n10881 & n10975 ;
  assign n10977 = n10881 & ~n10975 ;
  assign n10978 = ~n10976 & ~n10977 ;
  assign n10979 = x80 & n4531 ;
  assign n10980 = x78 & n4847 ;
  assign n10981 = x79 & n4526 ;
  assign n10982 = ~n10980 & ~n10981 ;
  assign n10983 = ~n10979 & n10982 ;
  assign n10984 = n2028 & n4534 ;
  assign n10985 = n10983 & ~n10984 ;
  assign n10986 = x26 & ~n10985 ;
  assign n10987 = x26 & ~n10986 ;
  assign n10988 = ~n10985 & ~n10986 ;
  assign n10989 = ~n10987 & ~n10988 ;
  assign n10990 = n10978 & ~n10989 ;
  assign n10991 = n10978 & ~n10990 ;
  assign n10992 = ~n10989 & ~n10990 ;
  assign n10993 = ~n10991 & ~n10992 ;
  assign n10994 = ~n10357 & ~n10450 ;
  assign n10995 = ~n10447 & ~n10994 ;
  assign n10996 = n10993 & n10995 ;
  assign n10997 = ~n10993 & ~n10995 ;
  assign n10998 = ~n10996 & ~n10997 ;
  assign n10999 = x83 & n3589 ;
  assign n11000 = x81 & n3878 ;
  assign n11001 = x82 & n3584 ;
  assign n11002 = ~n11000 & ~n11001 ;
  assign n11003 = ~n10999 & n11002 ;
  assign n11004 = n2843 & n3592 ;
  assign n11005 = n11003 & ~n11004 ;
  assign n11006 = x23 & ~n11005 ;
  assign n11007 = x23 & ~n11006 ;
  assign n11008 = ~n11005 & ~n11006 ;
  assign n11009 = ~n11007 & ~n11008 ;
  assign n11010 = n10998 & ~n11009 ;
  assign n11011 = n10998 & ~n11010 ;
  assign n11012 = ~n11009 & ~n11010 ;
  assign n11013 = ~n11011 & ~n11012 ;
  assign n11014 = ~n10465 & ~n10469 ;
  assign n11015 = n11013 & n11014 ;
  assign n11016 = ~n11013 & ~n11014 ;
  assign n11017 = ~n11015 & ~n11016 ;
  assign n11018 = x86 & n2751 ;
  assign n11019 = x84 & n3020 ;
  assign n11020 = x85 & n2746 ;
  assign n11021 = ~n11019 & ~n11020 ;
  assign n11022 = ~n11018 & n11021 ;
  assign n11023 = n2754 & n3686 ;
  assign n11024 = n11022 & ~n11023 ;
  assign n11025 = x20 & ~n11024 ;
  assign n11026 = x20 & ~n11025 ;
  assign n11027 = ~n11024 & ~n11025 ;
  assign n11028 = ~n11026 & ~n11027 ;
  assign n11029 = n11017 & ~n11028 ;
  assign n11030 = n11017 & ~n11029 ;
  assign n11031 = ~n11028 & ~n11029 ;
  assign n11032 = ~n11030 & ~n11031 ;
  assign n11033 = ~n10482 & ~n10488 ;
  assign n11034 = n11032 & n11033 ;
  assign n11035 = ~n11032 & ~n11033 ;
  assign n11036 = ~n11034 & ~n11035 ;
  assign n11037 = x89 & n2093 ;
  assign n11038 = x87 & n2275 ;
  assign n11039 = x88 & n2088 ;
  assign n11040 = ~n11038 & ~n11039 ;
  assign n11041 = ~n11037 & n11040 ;
  assign n11042 = n2096 & n4488 ;
  assign n11043 = n11041 & ~n11042 ;
  assign n11044 = x17 & ~n11043 ;
  assign n11045 = x17 & ~n11044 ;
  assign n11046 = ~n11043 & ~n11044 ;
  assign n11047 = ~n11045 & ~n11046 ;
  assign n11048 = n11036 & ~n11047 ;
  assign n11049 = n11036 & ~n11048 ;
  assign n11050 = ~n11047 & ~n11048 ;
  assign n11051 = ~n11049 & ~n11050 ;
  assign n11052 = ~n10502 & ~n10504 ;
  assign n11053 = ~n11051 & ~n11052 ;
  assign n11054 = n11051 & n11052 ;
  assign n11055 = ~n11053 & ~n11054 ;
  assign n11056 = ~n10880 & n11055 ;
  assign n11057 = ~n10880 & ~n11056 ;
  assign n11058 = n11055 & ~n11056 ;
  assign n11059 = ~n11057 & ~n11058 ;
  assign n11060 = ~n10869 & ~n11059 ;
  assign n11061 = ~n10869 & ~n11060 ;
  assign n11062 = ~n11059 & ~n11060 ;
  assign n11063 = ~n11061 & ~n11062 ;
  assign n11064 = x95 & n945 ;
  assign n11065 = x93 & n1099 ;
  assign n11066 = x94 & n940 ;
  assign n11067 = ~n11065 & ~n11066 ;
  assign n11068 = ~n11064 & n11067 ;
  assign n11069 = n948 & n6894 ;
  assign n11070 = n11068 & ~n11069 ;
  assign n11071 = x11 & ~n11070 ;
  assign n11072 = x11 & ~n11071 ;
  assign n11073 = ~n11070 & ~n11071 ;
  assign n11074 = ~n11072 & ~n11073 ;
  assign n11075 = n11063 & n11074 ;
  assign n11076 = ~n11063 & ~n11074 ;
  assign n11077 = ~n11075 & ~n11076 ;
  assign n11078 = ~n10867 & n11077 ;
  assign n11079 = n10867 & ~n11077 ;
  assign n11080 = ~n11078 & ~n11079 ;
  assign n11081 = n10866 & ~n11080 ;
  assign n11082 = ~n10866 & n11080 ;
  assign n11083 = ~n11081 & ~n11082 ;
  assign n11084 = ~n10855 & n11083 ;
  assign n11085 = n10855 & ~n11083 ;
  assign n11086 = ~n11084 & ~n11085 ;
  assign n11087 = x101 & n293 ;
  assign n11088 = x99 & n373 ;
  assign n11089 = x100 & n288 ;
  assign n11090 = ~n11088 & ~n11089 ;
  assign n11091 = ~n11087 & n11090 ;
  assign n11092 = n296 & n9601 ;
  assign n11093 = n11091 & ~n11092 ;
  assign n11094 = x5 & ~n11093 ;
  assign n11095 = x5 & ~n11094 ;
  assign n11096 = ~n11093 & ~n11094 ;
  assign n11097 = ~n11095 & ~n11096 ;
  assign n11098 = n11086 & ~n11097 ;
  assign n11099 = n11086 & ~n11098 ;
  assign n11100 = ~n11097 & ~n11098 ;
  assign n11101 = ~n11099 & ~n11100 ;
  assign n11102 = ~n10853 & n11101 ;
  assign n11103 = n10853 & ~n11101 ;
  assign n11104 = ~n11102 & ~n11103 ;
  assign n11105 = x104 & n146 ;
  assign n11106 = x102 & n182 ;
  assign n11107 = x103 & n141 ;
  assign n11108 = ~n11106 & ~n11107 ;
  assign n11109 = ~n11105 & n11108 ;
  assign n11110 = ~n10584 & ~n10586 ;
  assign n11111 = ~x103 & ~x104 ;
  assign n11112 = x103 & x104 ;
  assign n11113 = ~n11111 & ~n11112 ;
  assign n11114 = ~n11110 & n11113 ;
  assign n11115 = n11110 & ~n11113 ;
  assign n11116 = ~n11114 & ~n11115 ;
  assign n11117 = n149 & n11116 ;
  assign n11118 = n11109 & ~n11117 ;
  assign n11119 = x2 & ~n11118 ;
  assign n11120 = x2 & ~n11119 ;
  assign n11121 = ~n11118 & ~n11119 ;
  assign n11122 = ~n11120 & ~n11121 ;
  assign n11123 = ~n11104 & ~n11122 ;
  assign n11124 = n11104 & n11122 ;
  assign n11125 = ~n11123 & ~n11124 ;
  assign n11126 = ~n10852 & n11125 ;
  assign n11127 = n10852 & ~n11125 ;
  assign n11128 = ~n11126 & ~n11127 ;
  assign n11394 = n11128 & x168 ;
  assign n11129 = ~n10840 & ~n10845 ;
  assign n11130 = ~n10820 & ~n10822 ;
  assign n11131 = ~n10604 & ~n10804 ;
  assign n11132 = ~n10801 & ~n11131 ;
  assign n11133 = ~x98 & n574 ;
  assign n11134 = ~x96 & n673 ;
  assign n11135 = ~x97 & n569 ;
  assign n11136 = ~n11134 & ~n11135 ;
  assign n11137 = ~n11133 & n11136 ;
  assign n11138 = n577 & n8426 ;
  assign n11139 = n11137 & ~n11138 ;
  assign n11140 = ~x8 & ~n11139 ;
  assign n11141 = ~x8 & ~n11140 ;
  assign n11142 = ~n11139 & ~n11140 ;
  assign n11143 = ~n11141 & ~n11142 ;
  assign n11144 = ~n10784 & ~n10787 ;
  assign n11145 = ~n10606 & ~n10769 ;
  assign n11146 = ~n10766 & ~n11145 ;
  assign n11147 = ~x92 & n1434 ;
  assign n11148 = ~x90 & n1646 ;
  assign n11149 = ~x91 & n1429 ;
  assign n11150 = ~n11148 & ~n11149 ;
  assign n11151 = ~n11147 & n11150 ;
  assign n11152 = n1437 & n5896 ;
  assign n11153 = n11151 & ~n11152 ;
  assign n11154 = ~x14 & ~n11153 ;
  assign n11155 = ~x14 & ~n11154 ;
  assign n11156 = ~n11153 & ~n11154 ;
  assign n11157 = ~n11155 & ~n11156 ;
  assign n11158 = ~n10678 & ~n10681 ;
  assign n11159 = ~n10658 & ~n10664 ;
  assign n11160 = n10171 & n10609 ;
  assign n11161 = ~n10624 & ~n11160 ;
  assign n11162 = ~x68 & n9433 ;
  assign n11163 = ~x66 & n9915 ;
  assign n11164 = ~x67 & n9428 ;
  assign n11165 = ~n11163 & ~n11164 ;
  assign n11166 = ~n11162 & n11165 ;
  assign n11167 = n352 & n9436 ;
  assign n11168 = n11166 & ~n11167 ;
  assign n11169 = ~x38 & ~n11168 ;
  assign n11170 = ~x38 & ~n11169 ;
  assign n11171 = ~n11168 & ~n11169 ;
  assign n11172 = ~n11170 & ~n11171 ;
  assign n11173 = ~x41 & ~n10609 ;
  assign n11174 = ~x64 & n10900 ;
  assign n11175 = ~x65 & n10905 ;
  assign n11176 = ~n11174 & ~n11175 ;
  assign n11177 = ~n10909 & n11176 ;
  assign n11178 = ~x41 & ~n11177 ;
  assign n11179 = ~x41 & ~n11178 ;
  assign n11180 = ~n11177 & ~n11178 ;
  assign n11181 = ~n11179 & ~n11180 ;
  assign n11182 = n11173 & ~n11181 ;
  assign n11183 = ~n11173 & n11181 ;
  assign n11184 = ~n11182 & ~n11183 ;
  assign n11185 = n11172 & ~n11184 ;
  assign n11186 = ~n11172 & n11184 ;
  assign n11187 = ~n11185 & ~n11186 ;
  assign n11188 = ~n11161 & n11187 ;
  assign n11189 = n11161 & ~n11187 ;
  assign n11190 = ~n11188 & ~n11189 ;
  assign n11191 = ~x71 & n8006 ;
  assign n11192 = ~x69 & n8474 ;
  assign n11193 = ~x70 & n8001 ;
  assign n11194 = ~n11192 & ~n11193 ;
  assign n11195 = ~n11191 & n11194 ;
  assign n11196 = n622 & n8009 ;
  assign n11197 = n11195 & ~n11196 ;
  assign n11198 = ~x35 & ~n11197 ;
  assign n11199 = ~x35 & ~n11198 ;
  assign n11200 = ~n11197 & ~n11198 ;
  assign n11201 = ~n11199 & ~n11200 ;
  assign n11202 = n11190 & ~n11201 ;
  assign n11203 = n11190 & ~n11202 ;
  assign n11204 = ~n11201 & ~n11202 ;
  assign n11205 = ~n11203 & ~n11204 ;
  assign n11206 = ~n10638 & ~n10645 ;
  assign n11207 = n11205 & n11206 ;
  assign n11208 = ~n11205 & ~n11206 ;
  assign n11209 = ~n11207 & ~n11208 ;
  assign n11210 = ~x74 & n6725 ;
  assign n11211 = ~x72 & n7129 ;
  assign n11212 = ~x73 & n6720 ;
  assign n11213 = ~n11211 & ~n11212 ;
  assign n11214 = ~n11210 & n11213 ;
  assign n11215 = n1066 & n6728 ;
  assign n11216 = n11214 & ~n11215 ;
  assign n11217 = ~x32 & ~n11216 ;
  assign n11218 = ~x32 & ~n11217 ;
  assign n11219 = ~n11216 & ~n11217 ;
  assign n11220 = ~n11218 & ~n11219 ;
  assign n11221 = n11209 & ~n11220 ;
  assign n11222 = ~n11209 & n11220 ;
  assign n11223 = ~n11159 & ~n11222 ;
  assign n11224 = ~n11221 & n11223 ;
  assign n11225 = ~n11159 & ~n11224 ;
  assign n11226 = ~n11221 & ~n11224 ;
  assign n11227 = ~n11222 & n11226 ;
  assign n11228 = ~n11225 & ~n11227 ;
  assign n11229 = ~x77 & n5560 ;
  assign n11230 = ~x75 & n5943 ;
  assign n11231 = ~x76 & n5555 ;
  assign n11232 = ~n11230 & ~n11231 ;
  assign n11233 = ~n11229 & n11232 ;
  assign n11234 = n1594 & n5563 ;
  assign n11235 = n11233 & ~n11234 ;
  assign n11236 = ~x29 & ~n11235 ;
  assign n11237 = ~x29 & ~n11236 ;
  assign n11238 = ~n11235 & ~n11236 ;
  assign n11239 = ~n11237 & ~n11238 ;
  assign n11240 = n11228 & n11239 ;
  assign n11241 = ~n11228 & ~n11239 ;
  assign n11242 = ~n11240 & ~n11241 ;
  assign n11243 = ~n11158 & n11242 ;
  assign n11244 = n11158 & ~n11242 ;
  assign n11245 = ~n11243 & ~n11244 ;
  assign n11246 = ~x80 & n4531 ;
  assign n11247 = ~x78 & n4847 ;
  assign n11248 = ~x79 & n4526 ;
  assign n11249 = ~n11247 & ~n11248 ;
  assign n11250 = ~n11246 & n11249 ;
  assign n11251 = n2145 & n4534 ;
  assign n11252 = n11250 & ~n11251 ;
  assign n11253 = ~x26 & ~n11252 ;
  assign n11254 = ~x26 & ~n11253 ;
  assign n11255 = ~n11252 & ~n11253 ;
  assign n11256 = ~n11254 & ~n11255 ;
  assign n11257 = n11245 & ~n11256 ;
  assign n11258 = n11245 & ~n11257 ;
  assign n11259 = ~n11256 & ~n11257 ;
  assign n11260 = ~n11258 & ~n11259 ;
  assign n11261 = ~n10608 & ~n10698 ;
  assign n11262 = ~n10695 & ~n11261 ;
  assign n11263 = n11260 & n11262 ;
  assign n11264 = ~n11260 & ~n11262 ;
  assign n11265 = ~n11263 & ~n11264 ;
  assign n11266 = ~x83 & n3589 ;
  assign n11267 = ~x81 & n3878 ;
  assign n11268 = ~x82 & n3584 ;
  assign n11269 = ~n11267 & ~n11268 ;
  assign n11270 = ~n11266 & n11269 ;
  assign n11271 = n2972 & n3592 ;
  assign n11272 = n11270 & ~n11271 ;
  assign n11273 = ~x23 & ~n11272 ;
  assign n11274 = ~x23 & ~n11273 ;
  assign n11275 = ~n11272 & ~n11273 ;
  assign n11276 = ~n11274 & ~n11275 ;
  assign n11277 = n11265 & ~n11276 ;
  assign n11278 = n11265 & ~n11277 ;
  assign n11279 = ~n11276 & ~n11277 ;
  assign n11280 = ~n11278 & ~n11279 ;
  assign n11281 = ~n10713 & ~n10717 ;
  assign n11282 = n11280 & n11281 ;
  assign n11283 = ~n11280 & ~n11281 ;
  assign n11284 = ~n11282 & ~n11283 ;
  assign n11285 = ~x86 & n2751 ;
  assign n11286 = ~x84 & n3020 ;
  assign n11287 = ~x85 & n2746 ;
  assign n11288 = ~n11286 & ~n11287 ;
  assign n11289 = ~n11285 & n11288 ;
  assign n11290 = n2754 & n3832 ;
  assign n11291 = n11289 & ~n11290 ;
  assign n11292 = ~x20 & ~n11291 ;
  assign n11293 = ~x20 & ~n11292 ;
  assign n11294 = ~n11291 & ~n11292 ;
  assign n11295 = ~n11293 & ~n11294 ;
  assign n11296 = n11284 & ~n11295 ;
  assign n11297 = n11284 & ~n11296 ;
  assign n11298 = ~n11295 & ~n11296 ;
  assign n11299 = ~n11297 & ~n11298 ;
  assign n11300 = ~n10730 & ~n10736 ;
  assign n11301 = n11299 & n11300 ;
  assign n11302 = ~n11299 & ~n11300 ;
  assign n11303 = ~n11301 & ~n11302 ;
  assign n11304 = ~x89 & n2093 ;
  assign n11305 = ~x87 & n2275 ;
  assign n11306 = ~x88 & n2088 ;
  assign n11307 = ~n11305 & ~n11306 ;
  assign n11308 = ~n11304 & n11307 ;
  assign n11309 = n2096 & n4664 ;
  assign n11310 = n11308 & ~n11309 ;
  assign n11311 = ~x17 & ~n11310 ;
  assign n11312 = ~x17 & ~n11311 ;
  assign n11313 = ~n11310 & ~n11311 ;
  assign n11314 = ~n11312 & ~n11313 ;
  assign n11315 = n11303 & ~n11314 ;
  assign n11316 = n11303 & ~n11315 ;
  assign n11317 = ~n11314 & ~n11315 ;
  assign n11318 = ~n11316 & ~n11317 ;
  assign n11319 = ~n10750 & ~n10752 ;
  assign n11320 = ~n11318 & ~n11319 ;
  assign n11321 = n11318 & n11319 ;
  assign n11322 = ~n11320 & ~n11321 ;
  assign n11323 = ~n11157 & n11322 ;
  assign n11324 = ~n11157 & ~n11323 ;
  assign n11325 = n11322 & ~n11323 ;
  assign n11326 = ~n11324 & ~n11325 ;
  assign n11327 = ~n11146 & ~n11326 ;
  assign n11328 = ~n11146 & ~n11327 ;
  assign n11329 = ~n11326 & ~n11327 ;
  assign n11330 = ~n11328 & ~n11329 ;
  assign n11331 = ~x95 & n945 ;
  assign n11332 = ~x93 & n1099 ;
  assign n11333 = ~x94 & n940 ;
  assign n11334 = ~n11332 & ~n11333 ;
  assign n11335 = ~n11331 & n11334 ;
  assign n11336 = n948 & n7100 ;
  assign n11337 = n11335 & ~n11336 ;
  assign n11338 = ~x11 & ~n11337 ;
  assign n11339 = ~x11 & ~n11338 ;
  assign n11340 = ~n11337 & ~n11338 ;
  assign n11341 = ~n11339 & ~n11340 ;
  assign n11342 = n11330 & n11341 ;
  assign n11343 = ~n11330 & ~n11341 ;
  assign n11344 = ~n11342 & ~n11343 ;
  assign n11345 = ~n11144 & n11344 ;
  assign n11346 = n11144 & ~n11344 ;
  assign n11347 = ~n11345 & ~n11346 ;
  assign n11348 = n11143 & ~n11347 ;
  assign n11349 = ~n11143 & n11347 ;
  assign n11350 = ~n11348 & ~n11349 ;
  assign n11351 = ~n11132 & n11350 ;
  assign n11352 = n11132 & ~n11350 ;
  assign n11353 = ~n11351 & ~n11352 ;
  assign n11354 = ~x101 & n293 ;
  assign n11355 = ~x99 & n373 ;
  assign n11356 = ~x100 & n288 ;
  assign n11357 = ~n11355 & ~n11356 ;
  assign n11358 = ~n11354 & n11357 ;
  assign n11359 = n296 & n9844 ;
  assign n11360 = n11358 & ~n11359 ;
  assign n11361 = ~x5 & ~n11360 ;
  assign n11362 = ~x5 & ~n11361 ;
  assign n11363 = ~n11360 & ~n11361 ;
  assign n11364 = ~n11362 & ~n11363 ;
  assign n11365 = n11353 & ~n11364 ;
  assign n11366 = n11353 & ~n11365 ;
  assign n11367 = ~n11364 & ~n11365 ;
  assign n11368 = ~n11366 & ~n11367 ;
  assign n11369 = ~n11130 & n11368 ;
  assign n11370 = n11130 & ~n11368 ;
  assign n11371 = ~n11369 & ~n11370 ;
  assign n11372 = ~x104 & n164 ;
  assign n11373 = ~x102 & n205 ;
  assign n11374 = ~x103 & n162 ;
  assign n11375 = ~n11373 & ~n11374 ;
  assign n11376 = ~n11372 & n11375 ;
  assign n11377 = ~n10583 & ~n10831 ;
  assign n11378 = n11113 & ~n11377 ;
  assign n11379 = ~n11113 & n11377 ;
  assign n11380 = ~n11378 & ~n11379 ;
  assign n11381 = n167 & n11380 ;
  assign n11382 = n11376 & ~n11381 ;
  assign n11383 = ~x2 & ~n11382 ;
  assign n11384 = ~x2 & ~n11383 ;
  assign n11385 = ~n11382 & ~n11383 ;
  assign n11386 = ~n11384 & ~n11385 ;
  assign n11387 = ~n11371 & ~n11386 ;
  assign n11388 = n11371 & n11386 ;
  assign n11389 = ~n11387 & ~n11388 ;
  assign n11390 = ~n11129 & n11389 ;
  assign n11391 = n11129 & ~n11389 ;
  assign n11392 = ~n11390 & ~n11391 ;
  assign n11395 = ~n11392 & ~x168 ;
  assign n11396 = ~n11394 & ~n11395 ;
  assign n11397 = ~n11123 & ~n11126 ;
  assign n11398 = ~n10853 & ~n11101 ;
  assign n11399 = ~n11098 & ~n11398 ;
  assign n11400 = ~n11082 & ~n11084 ;
  assign n11401 = ~n11076 & ~n11078 ;
  assign n11402 = x96 & n945 ;
  assign n11403 = x94 & n1099 ;
  assign n11404 = x95 & n940 ;
  assign n11405 = ~n11403 & ~n11404 ;
  assign n11406 = ~n11402 & n11405 ;
  assign n11407 = n948 & n7321 ;
  assign n11408 = n11406 & ~n11407 ;
  assign n11409 = x11 & ~n11408 ;
  assign n11410 = x11 & ~n11409 ;
  assign n11411 = ~n11408 & ~n11409 ;
  assign n11412 = ~n11410 & ~n11411 ;
  assign n11413 = ~n11056 & ~n11060 ;
  assign n11414 = x93 & n1434 ;
  assign n11415 = x91 & n1646 ;
  assign n11416 = x92 & n1429 ;
  assign n11417 = ~n11415 & ~n11416 ;
  assign n11418 = ~n11414 & n11417 ;
  assign n11419 = n1437 & n6094 ;
  assign n11420 = n11418 & ~n11419 ;
  assign n11421 = x14 & ~n11420 ;
  assign n11422 = x14 & ~n11421 ;
  assign n11423 = ~n11420 & ~n11421 ;
  assign n11424 = ~n11422 & ~n11423 ;
  assign n11425 = ~n11048 & ~n11053 ;
  assign n11426 = ~n11029 & ~n11035 ;
  assign n11427 = ~n10990 & ~n10997 ;
  assign n11428 = x81 & n4531 ;
  assign n11429 = x79 & n4847 ;
  assign n11430 = x80 & n4526 ;
  assign n11431 = ~n11429 & ~n11430 ;
  assign n11432 = ~n11428 & n11431 ;
  assign n11433 = n2348 & n4534 ;
  assign n11434 = n11432 & ~n11433 ;
  assign n11435 = x26 & ~n11434 ;
  assign n11436 = x26 & ~n11435 ;
  assign n11437 = ~n11434 & ~n11435 ;
  assign n11438 = ~n11436 & ~n11437 ;
  assign n11439 = ~n10974 & ~n10976 ;
  assign n11440 = x78 & n5560 ;
  assign n11441 = x76 & n5943 ;
  assign n11442 = x77 & n5555 ;
  assign n11443 = ~n11441 & ~n11442 ;
  assign n11444 = ~n11440 & n11443 ;
  assign n11445 = n1624 & n5563 ;
  assign n11446 = n11444 & ~n11445 ;
  assign n11447 = x29 & ~n11446 ;
  assign n11448 = x29 & ~n11447 ;
  assign n11449 = ~n11446 & ~n11447 ;
  assign n11450 = ~n11448 & ~n11449 ;
  assign n11451 = ~n10935 & ~n10941 ;
  assign n11452 = x72 & n8006 ;
  assign n11453 = x70 & n8474 ;
  assign n11454 = x71 & n8001 ;
  assign n11455 = ~n11453 & ~n11454 ;
  assign n11456 = ~n11452 & n11455 ;
  assign n11457 = n717 & n8009 ;
  assign n11458 = n11456 & ~n11457 ;
  assign n11459 = x35 & ~n11458 ;
  assign n11460 = x35 & ~n11459 ;
  assign n11461 = ~n11458 & ~n11459 ;
  assign n11462 = ~n11460 & ~n11461 ;
  assign n11463 = ~n10919 & ~n10921 ;
  assign n11464 = x66 & n10905 ;
  assign n11465 = n10360 & ~n10904 ;
  assign n11466 = n10899 & n11465 ;
  assign n11467 = x64 & n11466 ;
  assign n11468 = x65 & n10900 ;
  assign n11469 = ~n11467 & ~n11468 ;
  assign n11470 = ~n11464 & n11469 ;
  assign n11471 = n194 & n10908 ;
  assign n11472 = n11470 & ~n11471 ;
  assign n11473 = x41 & ~n11472 ;
  assign n11474 = x41 & ~n11473 ;
  assign n11475 = ~n11472 & ~n11473 ;
  assign n11476 = ~n11474 & ~n11475 ;
  assign n11477 = ~n10915 & n11476 ;
  assign n11478 = n10915 & ~n11476 ;
  assign n11479 = ~n11477 & ~n11478 ;
  assign n11480 = x69 & n9433 ;
  assign n11481 = x67 & n9915 ;
  assign n11482 = x68 & n9428 ;
  assign n11483 = ~n11481 & ~n11482 ;
  assign n11484 = ~n11480 & n11483 ;
  assign n11485 = n398 & n9436 ;
  assign n11486 = n11484 & ~n11485 ;
  assign n11487 = x38 & ~n11486 ;
  assign n11488 = x38 & ~n11487 ;
  assign n11489 = ~n11486 & ~n11487 ;
  assign n11490 = ~n11488 & ~n11489 ;
  assign n11491 = n11479 & ~n11490 ;
  assign n11492 = n11479 & ~n11491 ;
  assign n11493 = ~n11490 & ~n11491 ;
  assign n11494 = ~n11492 & ~n11493 ;
  assign n11495 = ~n11463 & ~n11494 ;
  assign n11496 = n11463 & n11494 ;
  assign n11497 = ~n11495 & ~n11496 ;
  assign n11498 = ~n11462 & n11497 ;
  assign n11499 = ~n11462 & ~n11498 ;
  assign n11500 = n11497 & ~n11498 ;
  assign n11501 = ~n11499 & ~n11500 ;
  assign n11502 = ~n11451 & ~n11501 ;
  assign n11503 = ~n11451 & ~n11502 ;
  assign n11504 = ~n11501 & ~n11502 ;
  assign n11505 = ~n11503 & ~n11504 ;
  assign n11506 = x75 & n6725 ;
  assign n11507 = x73 & n7129 ;
  assign n11508 = x74 & n6720 ;
  assign n11509 = ~n11507 & ~n11508 ;
  assign n11510 = ~n11506 & n11509 ;
  assign n11511 = n1150 & n6728 ;
  assign n11512 = n11510 & ~n11511 ;
  assign n11513 = x32 & ~n11512 ;
  assign n11514 = x32 & ~n11513 ;
  assign n11515 = ~n11512 & ~n11513 ;
  assign n11516 = ~n11514 & ~n11515 ;
  assign n11517 = n11505 & n11516 ;
  assign n11518 = ~n11505 & ~n11516 ;
  assign n11519 = ~n11517 & ~n11518 ;
  assign n11520 = ~n10959 & n11519 ;
  assign n11521 = n10959 & ~n11519 ;
  assign n11522 = ~n11520 & ~n11521 ;
  assign n11523 = n11450 & ~n11522 ;
  assign n11524 = ~n11450 & n11522 ;
  assign n11525 = ~n11523 & ~n11524 ;
  assign n11526 = ~n11439 & n11525 ;
  assign n11527 = n11439 & ~n11525 ;
  assign n11528 = ~n11526 & ~n11527 ;
  assign n11529 = n11438 & ~n11528 ;
  assign n11530 = ~n11438 & n11528 ;
  assign n11531 = ~n11529 & ~n11530 ;
  assign n11532 = ~n11427 & n11531 ;
  assign n11533 = n11427 & ~n11531 ;
  assign n11534 = ~n11532 & ~n11533 ;
  assign n11535 = x84 & n3589 ;
  assign n11536 = x82 & n3878 ;
  assign n11537 = x83 & n3584 ;
  assign n11538 = ~n11536 & ~n11537 ;
  assign n11539 = ~n11535 & n11538 ;
  assign n11540 = n3114 & n3592 ;
  assign n11541 = n11539 & ~n11540 ;
  assign n11542 = x23 & ~n11541 ;
  assign n11543 = x23 & ~n11542 ;
  assign n11544 = ~n11541 & ~n11542 ;
  assign n11545 = ~n11543 & ~n11544 ;
  assign n11546 = n11534 & ~n11545 ;
  assign n11547 = n11534 & ~n11546 ;
  assign n11548 = ~n11545 & ~n11546 ;
  assign n11549 = ~n11547 & ~n11548 ;
  assign n11550 = ~n11010 & ~n11016 ;
  assign n11551 = n11549 & n11550 ;
  assign n11552 = ~n11549 & ~n11550 ;
  assign n11553 = ~n11551 & ~n11552 ;
  assign n11554 = x87 & n2751 ;
  assign n11555 = x85 & n3020 ;
  assign n11556 = x86 & n2746 ;
  assign n11557 = ~n11555 & ~n11556 ;
  assign n11558 = ~n11554 & n11557 ;
  assign n11559 = n2754 & n3991 ;
  assign n11560 = n11558 & ~n11559 ;
  assign n11561 = x20 & ~n11560 ;
  assign n11562 = x20 & ~n11561 ;
  assign n11563 = ~n11560 & ~n11561 ;
  assign n11564 = ~n11562 & ~n11563 ;
  assign n11565 = n11553 & ~n11564 ;
  assign n11566 = ~n11553 & n11564 ;
  assign n11567 = ~n11426 & ~n11566 ;
  assign n11568 = ~n11565 & n11567 ;
  assign n11569 = ~n11426 & ~n11568 ;
  assign n11570 = ~n11565 & ~n11568 ;
  assign n11571 = ~n11566 & n11570 ;
  assign n11572 = ~n11569 & ~n11571 ;
  assign n11573 = x90 & n2093 ;
  assign n11574 = x88 & n2275 ;
  assign n11575 = x89 & n2088 ;
  assign n11576 = ~n11574 & ~n11575 ;
  assign n11577 = ~n11573 & n11576 ;
  assign n11578 = n2096 & n4986 ;
  assign n11579 = n11577 & ~n11578 ;
  assign n11580 = x17 & ~n11579 ;
  assign n11581 = x17 & ~n11580 ;
  assign n11582 = ~n11579 & ~n11580 ;
  assign n11583 = ~n11581 & ~n11582 ;
  assign n11584 = n11572 & n11583 ;
  assign n11585 = ~n11572 & ~n11583 ;
  assign n11586 = ~n11584 & ~n11585 ;
  assign n11587 = ~n11425 & n11586 ;
  assign n11588 = n11425 & ~n11586 ;
  assign n11589 = ~n11587 & ~n11588 ;
  assign n11590 = n11424 & ~n11589 ;
  assign n11591 = ~n11424 & n11589 ;
  assign n11592 = ~n11590 & ~n11591 ;
  assign n11593 = ~n11413 & n11592 ;
  assign n11594 = n11413 & ~n11592 ;
  assign n11595 = ~n11593 & ~n11594 ;
  assign n11596 = n11412 & ~n11595 ;
  assign n11597 = ~n11412 & n11595 ;
  assign n11598 = ~n11596 & ~n11597 ;
  assign n11599 = ~n11401 & n11598 ;
  assign n11600 = n11401 & ~n11598 ;
  assign n11601 = ~n11599 & ~n11600 ;
  assign n11602 = x99 & n574 ;
  assign n11603 = x97 & n673 ;
  assign n11604 = x98 & n569 ;
  assign n11605 = ~n11603 & ~n11604 ;
  assign n11606 = ~n11602 & n11605 ;
  assign n11607 = n577 & n8660 ;
  assign n11608 = n11606 & ~n11607 ;
  assign n11609 = x8 & ~n11608 ;
  assign n11610 = x8 & ~n11609 ;
  assign n11611 = ~n11608 & ~n11609 ;
  assign n11612 = ~n11610 & ~n11611 ;
  assign n11613 = n11601 & ~n11612 ;
  assign n11614 = n11601 & ~n11613 ;
  assign n11615 = ~n11612 & ~n11613 ;
  assign n11616 = ~n11614 & ~n11615 ;
  assign n11617 = ~n11400 & n11616 ;
  assign n11618 = n11400 & ~n11616 ;
  assign n11619 = ~n11617 & ~n11618 ;
  assign n11620 = x102 & n293 ;
  assign n11621 = x100 & n373 ;
  assign n11622 = x101 & n288 ;
  assign n11623 = ~n11621 & ~n11622 ;
  assign n11624 = ~n11620 & n11623 ;
  assign n11625 = n296 & n10092 ;
  assign n11626 = n11624 & ~n11625 ;
  assign n11627 = x5 & ~n11626 ;
  assign n11628 = x5 & ~n11627 ;
  assign n11629 = ~n11626 & ~n11627 ;
  assign n11630 = ~n11628 & ~n11629 ;
  assign n11631 = ~n11619 & ~n11630 ;
  assign n11632 = n11619 & n11630 ;
  assign n11633 = ~n11631 & ~n11632 ;
  assign n11634 = n11399 & ~n11633 ;
  assign n11635 = ~n11399 & n11633 ;
  assign n11636 = ~n11634 & ~n11635 ;
  assign n11637 = x105 & n146 ;
  assign n11638 = x103 & n182 ;
  assign n11639 = x104 & n141 ;
  assign n11640 = ~n11638 & ~n11639 ;
  assign n11641 = ~n11637 & n11640 ;
  assign n11642 = ~n11112 & ~n11114 ;
  assign n11643 = ~x104 & ~x105 ;
  assign n11644 = x104 & x105 ;
  assign n11645 = ~n11643 & ~n11644 ;
  assign n11646 = ~n11642 & n11645 ;
  assign n11647 = n11642 & ~n11645 ;
  assign n11648 = ~n11646 & ~n11647 ;
  assign n11649 = n149 & n11648 ;
  assign n11650 = n11641 & ~n11649 ;
  assign n11651 = x2 & ~n11650 ;
  assign n11652 = x2 & ~n11651 ;
  assign n11653 = ~n11650 & ~n11651 ;
  assign n11654 = ~n11652 & ~n11653 ;
  assign n11655 = ~n11636 & n11654 ;
  assign n11656 = n11636 & ~n11654 ;
  assign n11657 = ~n11655 & ~n11656 ;
  assign n11658 = ~n11397 & n11657 ;
  assign n11659 = n11397 & ~n11657 ;
  assign n11660 = ~n11658 & ~n11659 ;
  assign n11921 = n11660 & x169 ;
  assign n11661 = ~n11387 & ~n11390 ;
  assign n11662 = ~n11130 & ~n11368 ;
  assign n11663 = ~n11365 & ~n11662 ;
  assign n11664 = ~n11349 & ~n11351 ;
  assign n11665 = ~n11343 & ~n11345 ;
  assign n11666 = ~x96 & n945 ;
  assign n11667 = ~x94 & n1099 ;
  assign n11668 = ~x95 & n940 ;
  assign n11669 = ~n11667 & ~n11668 ;
  assign n11670 = ~n11666 & n11669 ;
  assign n11671 = n948 & n7531 ;
  assign n11672 = n11670 & ~n11671 ;
  assign n11673 = ~x11 & ~n11672 ;
  assign n11674 = ~x11 & ~n11673 ;
  assign n11675 = ~n11672 & ~n11673 ;
  assign n11676 = ~n11674 & ~n11675 ;
  assign n11677 = ~n11323 & ~n11327 ;
  assign n11678 = ~x93 & n1434 ;
  assign n11679 = ~x91 & n1646 ;
  assign n11680 = ~x92 & n1429 ;
  assign n11681 = ~n11679 & ~n11680 ;
  assign n11682 = ~n11678 & n11681 ;
  assign n11683 = n1437 & n6285 ;
  assign n11684 = n11682 & ~n11683 ;
  assign n11685 = ~x14 & ~n11684 ;
  assign n11686 = ~x14 & ~n11685 ;
  assign n11687 = ~n11684 & ~n11685 ;
  assign n11688 = ~n11686 & ~n11687 ;
  assign n11689 = ~n11315 & ~n11320 ;
  assign n11690 = ~n11296 & ~n11302 ;
  assign n11691 = ~n11257 & ~n11264 ;
  assign n11692 = ~x81 & n4531 ;
  assign n11693 = ~x79 & n4847 ;
  assign n11694 = ~x80 & n4526 ;
  assign n11695 = ~n11693 & ~n11694 ;
  assign n11696 = ~n11692 & n11695 ;
  assign n11697 = n2460 & n4534 ;
  assign n11698 = n11696 & ~n11697 ;
  assign n11699 = ~x26 & ~n11698 ;
  assign n11700 = ~x26 & ~n11699 ;
  assign n11701 = ~n11698 & ~n11699 ;
  assign n11702 = ~n11700 & ~n11701 ;
  assign n11703 = ~n11241 & ~n11243 ;
  assign n11704 = ~x78 & n5560 ;
  assign n11705 = ~x76 & n5943 ;
  assign n11706 = ~x77 & n5555 ;
  assign n11707 = ~n11705 & ~n11706 ;
  assign n11708 = ~n11704 & n11707 ;
  assign n11709 = n1718 & n5563 ;
  assign n11710 = n11708 & ~n11709 ;
  assign n11711 = ~x29 & ~n11710 ;
  assign n11712 = ~x29 & ~n11711 ;
  assign n11713 = ~n11710 & ~n11711 ;
  assign n11714 = ~n11712 & ~n11713 ;
  assign n11715 = ~n11202 & ~n11208 ;
  assign n11716 = ~x72 & n8006 ;
  assign n11717 = ~x70 & n8474 ;
  assign n11718 = ~x71 & n8001 ;
  assign n11719 = ~n11717 & ~n11718 ;
  assign n11720 = ~n11716 & n11719 ;
  assign n11721 = n773 & n8009 ;
  assign n11722 = n11720 & ~n11721 ;
  assign n11723 = ~x35 & ~n11722 ;
  assign n11724 = ~x35 & ~n11723 ;
  assign n11725 = ~n11722 & ~n11723 ;
  assign n11726 = ~n11724 & ~n11725 ;
  assign n11727 = ~n11186 & ~n11188 ;
  assign n11728 = ~x66 & n10905 ;
  assign n11729 = ~x64 & n11466 ;
  assign n11730 = ~x65 & n10900 ;
  assign n11731 = ~n11729 & ~n11730 ;
  assign n11732 = ~n11728 & n11731 ;
  assign n11733 = n214 & n10908 ;
  assign n11734 = n11732 & ~n11733 ;
  assign n11735 = ~x41 & ~n11734 ;
  assign n11736 = ~x41 & ~n11735 ;
  assign n11737 = ~n11734 & ~n11735 ;
  assign n11738 = ~n11736 & ~n11737 ;
  assign n11739 = ~n11182 & n11738 ;
  assign n11740 = n11182 & ~n11738 ;
  assign n11741 = ~n11739 & ~n11740 ;
  assign n11742 = ~x69 & n9433 ;
  assign n11743 = ~x67 & n9915 ;
  assign n11744 = ~x68 & n9428 ;
  assign n11745 = ~n11743 & ~n11744 ;
  assign n11746 = ~n11742 & n11745 ;
  assign n11747 = n435 & n9436 ;
  assign n11748 = n11746 & ~n11747 ;
  assign n11749 = ~x38 & ~n11748 ;
  assign n11750 = ~x38 & ~n11749 ;
  assign n11751 = ~n11748 & ~n11749 ;
  assign n11752 = ~n11750 & ~n11751 ;
  assign n11753 = n11741 & ~n11752 ;
  assign n11754 = n11741 & ~n11753 ;
  assign n11755 = ~n11752 & ~n11753 ;
  assign n11756 = ~n11754 & ~n11755 ;
  assign n11757 = ~n11727 & ~n11756 ;
  assign n11758 = n11727 & n11756 ;
  assign n11759 = ~n11757 & ~n11758 ;
  assign n11760 = ~n11726 & n11759 ;
  assign n11761 = ~n11726 & ~n11760 ;
  assign n11762 = n11759 & ~n11760 ;
  assign n11763 = ~n11761 & ~n11762 ;
  assign n11764 = ~n11715 & ~n11763 ;
  assign n11765 = ~n11715 & ~n11764 ;
  assign n11766 = ~n11763 & ~n11764 ;
  assign n11767 = ~n11765 & ~n11766 ;
  assign n11768 = ~x75 & n6725 ;
  assign n11769 = ~x73 & n7129 ;
  assign n11770 = ~x74 & n6720 ;
  assign n11771 = ~n11769 & ~n11770 ;
  assign n11772 = ~n11768 & n11771 ;
  assign n11773 = n1225 & n6728 ;
  assign n11774 = n11772 & ~n11773 ;
  assign n11775 = ~x32 & ~n11774 ;
  assign n11776 = ~x32 & ~n11775 ;
  assign n11777 = ~n11774 & ~n11775 ;
  assign n11778 = ~n11776 & ~n11777 ;
  assign n11779 = n11767 & n11778 ;
  assign n11780 = ~n11767 & ~n11778 ;
  assign n11781 = ~n11779 & ~n11780 ;
  assign n11782 = ~n11226 & n11781 ;
  assign n11783 = n11226 & ~n11781 ;
  assign n11784 = ~n11782 & ~n11783 ;
  assign n11785 = n11714 & ~n11784 ;
  assign n11786 = ~n11714 & n11784 ;
  assign n11787 = ~n11785 & ~n11786 ;
  assign n11788 = ~n11703 & n11787 ;
  assign n11789 = n11703 & ~n11787 ;
  assign n11790 = ~n11788 & ~n11789 ;
  assign n11791 = n11702 & ~n11790 ;
  assign n11792 = ~n11702 & n11790 ;
  assign n11793 = ~n11791 & ~n11792 ;
  assign n11794 = ~n11691 & n11793 ;
  assign n11795 = n11691 & ~n11793 ;
  assign n11796 = ~n11794 & ~n11795 ;
  assign n11797 = ~x84 & n3589 ;
  assign n11798 = ~x82 & n3878 ;
  assign n11799 = ~x83 & n3584 ;
  assign n11800 = ~n11798 & ~n11799 ;
  assign n11801 = ~n11797 & n11800 ;
  assign n11802 = n3247 & n3592 ;
  assign n11803 = n11801 & ~n11802 ;
  assign n11804 = ~x23 & ~n11803 ;
  assign n11805 = ~x23 & ~n11804 ;
  assign n11806 = ~n11803 & ~n11804 ;
  assign n11807 = ~n11805 & ~n11806 ;
  assign n11808 = n11796 & ~n11807 ;
  assign n11809 = n11796 & ~n11808 ;
  assign n11810 = ~n11807 & ~n11808 ;
  assign n11811 = ~n11809 & ~n11810 ;
  assign n11812 = ~n11277 & ~n11283 ;
  assign n11813 = n11811 & n11812 ;
  assign n11814 = ~n11811 & ~n11812 ;
  assign n11815 = ~n11813 & ~n11814 ;
  assign n11816 = ~x87 & n2751 ;
  assign n11817 = ~x85 & n3020 ;
  assign n11818 = ~x86 & n2746 ;
  assign n11819 = ~n11817 & ~n11818 ;
  assign n11820 = ~n11816 & n11819 ;
  assign n11821 = n2754 & n4143 ;
  assign n11822 = n11820 & ~n11821 ;
  assign n11823 = ~x20 & ~n11822 ;
  assign n11824 = ~x20 & ~n11823 ;
  assign n11825 = ~n11822 & ~n11823 ;
  assign n11826 = ~n11824 & ~n11825 ;
  assign n11827 = n11815 & ~n11826 ;
  assign n11828 = ~n11815 & n11826 ;
  assign n11829 = ~n11690 & ~n11828 ;
  assign n11830 = ~n11827 & n11829 ;
  assign n11831 = ~n11690 & ~n11830 ;
  assign n11832 = ~n11827 & ~n11830 ;
  assign n11833 = ~n11828 & n11832 ;
  assign n11834 = ~n11831 & ~n11833 ;
  assign n11835 = ~x90 & n2093 ;
  assign n11836 = ~x88 & n2275 ;
  assign n11837 = ~x89 & n2088 ;
  assign n11838 = ~n11836 & ~n11837 ;
  assign n11839 = ~n11835 & n11838 ;
  assign n11840 = n2096 & n5155 ;
  assign n11841 = n11839 & ~n11840 ;
  assign n11842 = ~x17 & ~n11841 ;
  assign n11843 = ~x17 & ~n11842 ;
  assign n11844 = ~n11841 & ~n11842 ;
  assign n11845 = ~n11843 & ~n11844 ;
  assign n11846 = n11834 & n11845 ;
  assign n11847 = ~n11834 & ~n11845 ;
  assign n11848 = ~n11846 & ~n11847 ;
  assign n11849 = ~n11689 & n11848 ;
  assign n11850 = n11689 & ~n11848 ;
  assign n11851 = ~n11849 & ~n11850 ;
  assign n11852 = n11688 & ~n11851 ;
  assign n11853 = ~n11688 & n11851 ;
  assign n11854 = ~n11852 & ~n11853 ;
  assign n11855 = ~n11677 & n11854 ;
  assign n11856 = n11677 & ~n11854 ;
  assign n11857 = ~n11855 & ~n11856 ;
  assign n11858 = n11676 & ~n11857 ;
  assign n11859 = ~n11676 & n11857 ;
  assign n11860 = ~n11858 & ~n11859 ;
  assign n11861 = ~n11665 & n11860 ;
  assign n11862 = n11665 & ~n11860 ;
  assign n11863 = ~n11861 & ~n11862 ;
  assign n11864 = ~x99 & n574 ;
  assign n11865 = ~x97 & n673 ;
  assign n11866 = ~x98 & n569 ;
  assign n11867 = ~n11865 & ~n11866 ;
  assign n11868 = ~n11864 & n11867 ;
  assign n11869 = n577 & n8885 ;
  assign n11870 = n11868 & ~n11869 ;
  assign n11871 = ~x8 & ~n11870 ;
  assign n11872 = ~x8 & ~n11871 ;
  assign n11873 = ~n11870 & ~n11871 ;
  assign n11874 = ~n11872 & ~n11873 ;
  assign n11875 = n11863 & ~n11874 ;
  assign n11876 = n11863 & ~n11875 ;
  assign n11877 = ~n11874 & ~n11875 ;
  assign n11878 = ~n11876 & ~n11877 ;
  assign n11879 = ~n11664 & n11878 ;
  assign n11880 = n11664 & ~n11878 ;
  assign n11881 = ~n11879 & ~n11880 ;
  assign n11882 = ~x102 & n293 ;
  assign n11883 = ~x100 & n373 ;
  assign n11884 = ~x101 & n288 ;
  assign n11885 = ~n11883 & ~n11884 ;
  assign n11886 = ~n11882 & n11885 ;
  assign n11887 = n296 & n10333 ;
  assign n11888 = n11886 & ~n11887 ;
  assign n11889 = ~x5 & ~n11888 ;
  assign n11890 = ~x5 & ~n11889 ;
  assign n11891 = ~n11888 & ~n11889 ;
  assign n11892 = ~n11890 & ~n11891 ;
  assign n11893 = ~n11881 & ~n11892 ;
  assign n11894 = n11881 & n11892 ;
  assign n11895 = ~n11893 & ~n11894 ;
  assign n11896 = n11663 & ~n11895 ;
  assign n11897 = ~n11663 & n11895 ;
  assign n11898 = ~n11896 & ~n11897 ;
  assign n11899 = ~x105 & n164 ;
  assign n11900 = ~x103 & n205 ;
  assign n11901 = ~x104 & n162 ;
  assign n11902 = ~n11900 & ~n11901 ;
  assign n11903 = ~n11899 & n11902 ;
  assign n11904 = ~n11111 & ~n11378 ;
  assign n11905 = n11645 & ~n11904 ;
  assign n11906 = ~n11645 & n11904 ;
  assign n11907 = ~n11905 & ~n11906 ;
  assign n11908 = n167 & n11907 ;
  assign n11909 = n11903 & ~n11908 ;
  assign n11910 = ~x2 & ~n11909 ;
  assign n11911 = ~x2 & ~n11910 ;
  assign n11912 = ~n11909 & ~n11910 ;
  assign n11913 = ~n11911 & ~n11912 ;
  assign n11914 = ~n11898 & n11913 ;
  assign n11915 = n11898 & ~n11913 ;
  assign n11916 = ~n11914 & ~n11915 ;
  assign n11917 = ~n11661 & n11916 ;
  assign n11918 = n11661 & ~n11916 ;
  assign n11919 = ~n11917 & ~n11918 ;
  assign n11922 = ~n11919 & ~x169 ;
  assign n11923 = ~n11921 & ~n11922 ;
  assign n11924 = ~n11631 & ~n11635 ;
  assign n11925 = x103 & n293 ;
  assign n11926 = x101 & n373 ;
  assign n11927 = x102 & n288 ;
  assign n11928 = ~n11926 & ~n11927 ;
  assign n11929 = ~n11925 & n11928 ;
  assign n11930 = n296 & n10588 ;
  assign n11931 = n11929 & ~n11930 ;
  assign n11932 = x5 & ~n11931 ;
  assign n11933 = x5 & ~n11932 ;
  assign n11934 = ~n11931 & ~n11932 ;
  assign n11935 = ~n11933 & ~n11934 ;
  assign n11936 = ~n11400 & ~n11616 ;
  assign n11937 = ~n11613 & ~n11936 ;
  assign n11938 = ~n11597 & ~n11599 ;
  assign n11939 = ~n11591 & ~n11593 ;
  assign n11940 = ~n11585 & ~n11587 ;
  assign n11941 = ~n11530 & ~n11532 ;
  assign n11942 = ~n11524 & ~n11526 ;
  assign n11943 = ~n11518 & ~n11520 ;
  assign n11944 = x76 & n6725 ;
  assign n11945 = x74 & n7129 ;
  assign n11946 = x75 & n6720 ;
  assign n11947 = ~n11945 & ~n11946 ;
  assign n11948 = ~n11944 & n11947 ;
  assign n11949 = n1311 & n6728 ;
  assign n11950 = n11948 & ~n11949 ;
  assign n11951 = x32 & ~n11950 ;
  assign n11952 = x32 & ~n11951 ;
  assign n11953 = ~n11950 & ~n11951 ;
  assign n11954 = ~n11952 & ~n11953 ;
  assign n11955 = ~n11498 & ~n11502 ;
  assign n11956 = x41 & ~x42 ;
  assign n11957 = ~x41 & x42 ;
  assign n11958 = ~n11956 & ~n11957 ;
  assign n11959 = x64 & ~n11958 ;
  assign n11960 = ~n11478 & n11959 ;
  assign n11961 = n11478 & ~n11959 ;
  assign n11962 = ~n11960 & ~n11961 ;
  assign n11963 = x67 & n10905 ;
  assign n11964 = x65 & n11466 ;
  assign n11965 = x66 & n10900 ;
  assign n11966 = ~n11964 & ~n11965 ;
  assign n11967 = ~n11963 & n11966 ;
  assign n11968 = n240 & n10908 ;
  assign n11969 = n11967 & ~n11968 ;
  assign n11970 = x41 & ~n11969 ;
  assign n11971 = x41 & ~n11970 ;
  assign n11972 = ~n11969 & ~n11970 ;
  assign n11973 = ~n11971 & ~n11972 ;
  assign n11974 = ~n11962 & ~n11973 ;
  assign n11975 = n11962 & n11973 ;
  assign n11976 = ~n11974 & ~n11975 ;
  assign n11977 = x70 & n9433 ;
  assign n11978 = x68 & n9915 ;
  assign n11979 = x69 & n9428 ;
  assign n11980 = ~n11978 & ~n11979 ;
  assign n11981 = ~n11977 & n11980 ;
  assign n11982 = n488 & n9436 ;
  assign n11983 = n11981 & ~n11982 ;
  assign n11984 = x38 & ~n11983 ;
  assign n11985 = x38 & ~n11984 ;
  assign n11986 = ~n11983 & ~n11984 ;
  assign n11987 = ~n11985 & ~n11986 ;
  assign n11988 = n11976 & ~n11987 ;
  assign n11989 = n11976 & ~n11988 ;
  assign n11990 = ~n11987 & ~n11988 ;
  assign n11991 = ~n11989 & ~n11990 ;
  assign n11992 = ~n11491 & ~n11495 ;
  assign n11993 = n11991 & n11992 ;
  assign n11994 = ~n11991 & ~n11992 ;
  assign n11995 = ~n11993 & ~n11994 ;
  assign n11996 = x73 & n8006 ;
  assign n11997 = x71 & n8474 ;
  assign n11998 = x72 & n8001 ;
  assign n11999 = ~n11997 & ~n11998 ;
  assign n12000 = ~n11996 & n11999 ;
  assign n12001 = n843 & n8009 ;
  assign n12002 = n12000 & ~n12001 ;
  assign n12003 = x35 & ~n12002 ;
  assign n12004 = x35 & ~n12003 ;
  assign n12005 = ~n12002 & ~n12003 ;
  assign n12006 = ~n12004 & ~n12005 ;
  assign n12007 = ~n11995 & n12006 ;
  assign n12008 = n11995 & ~n12006 ;
  assign n12009 = ~n12007 & ~n12008 ;
  assign n12010 = ~n11955 & n12009 ;
  assign n12011 = n11955 & ~n12009 ;
  assign n12012 = ~n12010 & ~n12011 ;
  assign n12013 = ~n11954 & n12012 ;
  assign n12014 = ~n11954 & ~n12013 ;
  assign n12015 = n12012 & ~n12013 ;
  assign n12016 = ~n12014 & ~n12015 ;
  assign n12017 = ~n11943 & ~n12016 ;
  assign n12018 = ~n11943 & ~n12017 ;
  assign n12019 = ~n12016 & ~n12017 ;
  assign n12020 = ~n12018 & ~n12019 ;
  assign n12021 = x79 & n5560 ;
  assign n12022 = x77 & n5943 ;
  assign n12023 = x78 & n5555 ;
  assign n12024 = ~n12022 & ~n12023 ;
  assign n12025 = ~n12021 & n12024 ;
  assign n12026 = n1817 & n5563 ;
  assign n12027 = n12025 & ~n12026 ;
  assign n12028 = x29 & ~n12027 ;
  assign n12029 = x29 & ~n12028 ;
  assign n12030 = ~n12027 & ~n12028 ;
  assign n12031 = ~n12029 & ~n12030 ;
  assign n12032 = ~n12020 & ~n12031 ;
  assign n12033 = ~n12020 & ~n12032 ;
  assign n12034 = ~n12031 & ~n12032 ;
  assign n12035 = ~n12033 & ~n12034 ;
  assign n12036 = ~n11942 & n12035 ;
  assign n12037 = n11942 & ~n12035 ;
  assign n12038 = ~n12036 & ~n12037 ;
  assign n12039 = x82 & n4531 ;
  assign n12040 = x80 & n4847 ;
  assign n12041 = x81 & n4526 ;
  assign n12042 = ~n12040 & ~n12041 ;
  assign n12043 = ~n12039 & n12042 ;
  assign n12044 = n2584 & n4534 ;
  assign n12045 = n12043 & ~n12044 ;
  assign n12046 = x26 & ~n12045 ;
  assign n12047 = x26 & ~n12046 ;
  assign n12048 = ~n12045 & ~n12046 ;
  assign n12049 = ~n12047 & ~n12048 ;
  assign n12050 = ~n12038 & ~n12049 ;
  assign n12051 = n12038 & n12049 ;
  assign n12052 = ~n12050 & ~n12051 ;
  assign n12053 = ~n11941 & n12052 ;
  assign n12054 = n11941 & ~n12052 ;
  assign n12055 = ~n12053 & ~n12054 ;
  assign n12056 = x85 & n3589 ;
  assign n12057 = x83 & n3878 ;
  assign n12058 = x84 & n3584 ;
  assign n12059 = ~n12057 & ~n12058 ;
  assign n12060 = ~n12056 & n12059 ;
  assign n12061 = n3389 & n3592 ;
  assign n12062 = n12060 & ~n12061 ;
  assign n12063 = x23 & ~n12062 ;
  assign n12064 = x23 & ~n12063 ;
  assign n12065 = ~n12062 & ~n12063 ;
  assign n12066 = ~n12064 & ~n12065 ;
  assign n12067 = n12055 & ~n12066 ;
  assign n12068 = n12055 & ~n12067 ;
  assign n12069 = ~n12066 & ~n12067 ;
  assign n12070 = ~n12068 & ~n12069 ;
  assign n12071 = ~n11546 & ~n11552 ;
  assign n12072 = n12070 & n12071 ;
  assign n12073 = ~n12070 & ~n12071 ;
  assign n12074 = ~n12072 & ~n12073 ;
  assign n12075 = x88 & n2751 ;
  assign n12076 = x86 & n3020 ;
  assign n12077 = x87 & n2746 ;
  assign n12078 = ~n12076 & ~n12077 ;
  assign n12079 = ~n12075 & n12078 ;
  assign n12080 = n2754 & n4305 ;
  assign n12081 = n12079 & ~n12080 ;
  assign n12082 = x20 & ~n12081 ;
  assign n12083 = x20 & ~n12082 ;
  assign n12084 = ~n12081 & ~n12082 ;
  assign n12085 = ~n12083 & ~n12084 ;
  assign n12086 = ~n12074 & n12085 ;
  assign n12087 = n12074 & ~n12085 ;
  assign n12088 = ~n12086 & ~n12087 ;
  assign n12089 = ~n11570 & n12088 ;
  assign n12090 = n11570 & ~n12088 ;
  assign n12091 = ~n12089 & ~n12090 ;
  assign n12092 = x91 & n2093 ;
  assign n12093 = x89 & n2275 ;
  assign n12094 = x90 & n2088 ;
  assign n12095 = ~n12093 & ~n12094 ;
  assign n12096 = ~n12092 & n12095 ;
  assign n12097 = n2096 & n5336 ;
  assign n12098 = n12096 & ~n12097 ;
  assign n12099 = x17 & ~n12098 ;
  assign n12100 = x17 & ~n12099 ;
  assign n12101 = ~n12098 & ~n12099 ;
  assign n12102 = ~n12100 & ~n12101 ;
  assign n12103 = n12091 & ~n12102 ;
  assign n12104 = n12091 & ~n12103 ;
  assign n12105 = ~n12102 & ~n12103 ;
  assign n12106 = ~n12104 & ~n12105 ;
  assign n12107 = ~n11940 & n12106 ;
  assign n12108 = n11940 & ~n12106 ;
  assign n12109 = ~n12107 & ~n12108 ;
  assign n12110 = x94 & n1434 ;
  assign n12111 = x92 & n1646 ;
  assign n12112 = x93 & n1429 ;
  assign n12113 = ~n12111 & ~n12112 ;
  assign n12114 = ~n12110 & n12113 ;
  assign n12115 = n1437 & n6483 ;
  assign n12116 = n12114 & ~n12115 ;
  assign n12117 = x14 & ~n12116 ;
  assign n12118 = x14 & ~n12117 ;
  assign n12119 = ~n12116 & ~n12117 ;
  assign n12120 = ~n12118 & ~n12119 ;
  assign n12121 = ~n12109 & ~n12120 ;
  assign n12122 = n12109 & n12120 ;
  assign n12123 = ~n12121 & ~n12122 ;
  assign n12124 = ~n11939 & n12123 ;
  assign n12125 = n11939 & ~n12123 ;
  assign n12126 = ~n12124 & ~n12125 ;
  assign n12127 = x97 & n945 ;
  assign n12128 = x95 & n1099 ;
  assign n12129 = x96 & n940 ;
  assign n12130 = ~n12128 & ~n12129 ;
  assign n12131 = ~n12127 & n12130 ;
  assign n12132 = n948 & n7745 ;
  assign n12133 = n12131 & ~n12132 ;
  assign n12134 = x11 & ~n12133 ;
  assign n12135 = x11 & ~n12134 ;
  assign n12136 = ~n12133 & ~n12134 ;
  assign n12137 = ~n12135 & ~n12136 ;
  assign n12138 = n12126 & ~n12137 ;
  assign n12139 = n12126 & ~n12138 ;
  assign n12140 = ~n12137 & ~n12138 ;
  assign n12141 = ~n12139 & ~n12140 ;
  assign n12142 = ~n11938 & n12141 ;
  assign n12143 = n11938 & ~n12141 ;
  assign n12144 = ~n12142 & ~n12143 ;
  assign n12145 = x100 & n574 ;
  assign n12146 = x98 & n673 ;
  assign n12147 = x99 & n569 ;
  assign n12148 = ~n12146 & ~n12147 ;
  assign n12149 = ~n12145 & n12148 ;
  assign n12150 = n577 & n9115 ;
  assign n12151 = n12149 & ~n12150 ;
  assign n12152 = x8 & ~n12151 ;
  assign n12153 = x8 & ~n12152 ;
  assign n12154 = ~n12151 & ~n12152 ;
  assign n12155 = ~n12153 & ~n12154 ;
  assign n12156 = n12144 & n12155 ;
  assign n12157 = ~n12144 & ~n12155 ;
  assign n12158 = ~n12156 & ~n12157 ;
  assign n12159 = ~n11937 & n12158 ;
  assign n12160 = n11937 & ~n12158 ;
  assign n12161 = ~n12159 & ~n12160 ;
  assign n12162 = ~n11935 & n12161 ;
  assign n12163 = ~n11935 & ~n12162 ;
  assign n12164 = n12161 & ~n12162 ;
  assign n12165 = ~n12163 & ~n12164 ;
  assign n12166 = ~n11924 & ~n12165 ;
  assign n12167 = ~n11924 & ~n12166 ;
  assign n12168 = ~n12165 & ~n12166 ;
  assign n12169 = ~n12167 & ~n12168 ;
  assign n12170 = x106 & n146 ;
  assign n12171 = x104 & n182 ;
  assign n12172 = x105 & n141 ;
  assign n12173 = ~n12171 & ~n12172 ;
  assign n12174 = ~n12170 & n12173 ;
  assign n12175 = ~n11644 & ~n11646 ;
  assign n12176 = ~x105 & ~x106 ;
  assign n12177 = x105 & x106 ;
  assign n12178 = ~n12176 & ~n12177 ;
  assign n12179 = ~n12175 & n12178 ;
  assign n12180 = n12175 & ~n12178 ;
  assign n12181 = ~n12179 & ~n12180 ;
  assign n12182 = n149 & n12181 ;
  assign n12183 = n12174 & ~n12182 ;
  assign n12184 = x2 & ~n12183 ;
  assign n12185 = x2 & ~n12184 ;
  assign n12186 = ~n12183 & ~n12184 ;
  assign n12187 = ~n12185 & ~n12186 ;
  assign n12188 = ~n12169 & ~n12187 ;
  assign n12189 = ~n12169 & ~n12188 ;
  assign n12190 = ~n12187 & ~n12188 ;
  assign n12191 = ~n12189 & ~n12190 ;
  assign n12192 = ~n11656 & ~n11658 ;
  assign n12193 = ~n12191 & ~n12192 ;
  assign n12194 = n12191 & n12192 ;
  assign n12195 = ~n12193 & ~n12194 ;
  assign n12463 = n12195 & x170 ;
  assign n12196 = ~n11893 & ~n11897 ;
  assign n12197 = ~x103 & n293 ;
  assign n12198 = ~x101 & n373 ;
  assign n12199 = ~x102 & n288 ;
  assign n12200 = ~n12198 & ~n12199 ;
  assign n12201 = ~n12197 & n12200 ;
  assign n12202 = n296 & n10833 ;
  assign n12203 = n12201 & ~n12202 ;
  assign n12204 = ~x5 & ~n12203 ;
  assign n12205 = ~x5 & ~n12204 ;
  assign n12206 = ~n12203 & ~n12204 ;
  assign n12207 = ~n12205 & ~n12206 ;
  assign n12208 = ~n11664 & ~n11878 ;
  assign n12209 = ~n11875 & ~n12208 ;
  assign n12210 = ~n11859 & ~n11861 ;
  assign n12211 = ~n11853 & ~n11855 ;
  assign n12212 = ~n11847 & ~n11849 ;
  assign n12213 = ~n11792 & ~n11794 ;
  assign n12214 = ~n11786 & ~n11788 ;
  assign n12215 = ~n11780 & ~n11782 ;
  assign n12216 = ~x76 & n6725 ;
  assign n12217 = ~x74 & n7129 ;
  assign n12218 = ~x75 & n6720 ;
  assign n12219 = ~n12217 & ~n12218 ;
  assign n12220 = ~n12216 & n12219 ;
  assign n12221 = n1390 & n6728 ;
  assign n12222 = n12220 & ~n12221 ;
  assign n12223 = ~x32 & ~n12222 ;
  assign n12224 = ~x32 & ~n12223 ;
  assign n12225 = ~n12222 & ~n12223 ;
  assign n12226 = ~n12224 & ~n12225 ;
  assign n12227 = ~n11760 & ~n11764 ;
  assign n12228 = ~x64 & ~n11958 ;
  assign n12229 = ~n11740 & n12228 ;
  assign n12230 = n11740 & ~n12228 ;
  assign n12231 = ~n12229 & ~n12230 ;
  assign n12232 = ~x67 & n10905 ;
  assign n12233 = ~x65 & n11466 ;
  assign n12234 = ~x66 & n10900 ;
  assign n12235 = ~n12233 & ~n12234 ;
  assign n12236 = ~n12232 & n12235 ;
  assign n12237 = n266 & n10908 ;
  assign n12238 = n12236 & ~n12237 ;
  assign n12239 = ~x41 & ~n12238 ;
  assign n12240 = ~x41 & ~n12239 ;
  assign n12241 = ~n12238 & ~n12239 ;
  assign n12242 = ~n12240 & ~n12241 ;
  assign n12243 = ~n12231 & ~n12242 ;
  assign n12244 = n12231 & n12242 ;
  assign n12245 = ~n12243 & ~n12244 ;
  assign n12246 = ~x70 & n9433 ;
  assign n12247 = ~x68 & n9915 ;
  assign n12248 = ~x69 & n9428 ;
  assign n12249 = ~n12247 & ~n12248 ;
  assign n12250 = ~n12246 & n12249 ;
  assign n12251 = n529 & n9436 ;
  assign n12252 = n12250 & ~n12251 ;
  assign n12253 = ~x38 & ~n12252 ;
  assign n12254 = ~x38 & ~n12253 ;
  assign n12255 = ~n12252 & ~n12253 ;
  assign n12256 = ~n12254 & ~n12255 ;
  assign n12257 = n12245 & ~n12256 ;
  assign n12258 = n12245 & ~n12257 ;
  assign n12259 = ~n12256 & ~n12257 ;
  assign n12260 = ~n12258 & ~n12259 ;
  assign n12261 = ~n11753 & ~n11757 ;
  assign n12262 = n12260 & n12261 ;
  assign n12263 = ~n12260 & ~n12261 ;
  assign n12264 = ~n12262 & ~n12263 ;
  assign n12265 = ~x73 & n8006 ;
  assign n12266 = ~x71 & n8474 ;
  assign n12267 = ~x72 & n8001 ;
  assign n12268 = ~n12266 & ~n12267 ;
  assign n12269 = ~n12265 & n12268 ;
  assign n12270 = n903 & n8009 ;
  assign n12271 = n12269 & ~n12270 ;
  assign n12272 = ~x35 & ~n12271 ;
  assign n12273 = ~x35 & ~n12272 ;
  assign n12274 = ~n12271 & ~n12272 ;
  assign n12275 = ~n12273 & ~n12274 ;
  assign n12276 = ~n12264 & n12275 ;
  assign n12277 = n12264 & ~n12275 ;
  assign n12278 = ~n12276 & ~n12277 ;
  assign n12279 = ~n12227 & n12278 ;
  assign n12280 = n12227 & ~n12278 ;
  assign n12281 = ~n12279 & ~n12280 ;
  assign n12282 = ~n12226 & n12281 ;
  assign n12283 = ~n12226 & ~n12282 ;
  assign n12284 = n12281 & ~n12282 ;
  assign n12285 = ~n12283 & ~n12284 ;
  assign n12286 = ~n12215 & ~n12285 ;
  assign n12287 = ~n12215 & ~n12286 ;
  assign n12288 = ~n12285 & ~n12286 ;
  assign n12289 = ~n12287 & ~n12288 ;
  assign n12290 = ~x79 & n5560 ;
  assign n12291 = ~x77 & n5943 ;
  assign n12292 = ~x78 & n5555 ;
  assign n12293 = ~n12291 & ~n12292 ;
  assign n12294 = ~n12290 & n12293 ;
  assign n12295 = n1921 & n5563 ;
  assign n12296 = n12294 & ~n12295 ;
  assign n12297 = ~x29 & ~n12296 ;
  assign n12298 = ~x29 & ~n12297 ;
  assign n12299 = ~n12296 & ~n12297 ;
  assign n12300 = ~n12298 & ~n12299 ;
  assign n12301 = ~n12289 & ~n12300 ;
  assign n12302 = ~n12289 & ~n12301 ;
  assign n12303 = ~n12300 & ~n12301 ;
  assign n12304 = ~n12302 & ~n12303 ;
  assign n12305 = ~n12214 & n12304 ;
  assign n12306 = n12214 & ~n12304 ;
  assign n12307 = ~n12305 & ~n12306 ;
  assign n12308 = ~x82 & n4531 ;
  assign n12309 = ~x80 & n4847 ;
  assign n12310 = ~x81 & n4526 ;
  assign n12311 = ~n12309 & ~n12310 ;
  assign n12312 = ~n12308 & n12311 ;
  assign n12313 = n2697 & n4534 ;
  assign n12314 = n12312 & ~n12313 ;
  assign n12315 = ~x26 & ~n12314 ;
  assign n12316 = ~x26 & ~n12315 ;
  assign n12317 = ~n12314 & ~n12315 ;
  assign n12318 = ~n12316 & ~n12317 ;
  assign n12319 = ~n12307 & ~n12318 ;
  assign n12320 = n12307 & n12318 ;
  assign n12321 = ~n12319 & ~n12320 ;
  assign n12322 = ~n12213 & n12321 ;
  assign n12323 = n12213 & ~n12321 ;
  assign n12324 = ~n12322 & ~n12323 ;
  assign n12325 = ~x85 & n3589 ;
  assign n12326 = ~x83 & n3878 ;
  assign n12327 = ~x84 & n3584 ;
  assign n12328 = ~n12326 & ~n12327 ;
  assign n12329 = ~n12325 & n12328 ;
  assign n12330 = n3521 & n3592 ;
  assign n12331 = n12329 & ~n12330 ;
  assign n12332 = ~x23 & ~n12331 ;
  assign n12333 = ~x23 & ~n12332 ;
  assign n12334 = ~n12331 & ~n12332 ;
  assign n12335 = ~n12333 & ~n12334 ;
  assign n12336 = n12324 & ~n12335 ;
  assign n12337 = n12324 & ~n12336 ;
  assign n12338 = ~n12335 & ~n12336 ;
  assign n12339 = ~n12337 & ~n12338 ;
  assign n12340 = ~n11808 & ~n11814 ;
  assign n12341 = n12339 & n12340 ;
  assign n12342 = ~n12339 & ~n12340 ;
  assign n12343 = ~n12341 & ~n12342 ;
  assign n12344 = ~x88 & n2751 ;
  assign n12345 = ~x86 & n3020 ;
  assign n12346 = ~x87 & n2746 ;
  assign n12347 = ~n12345 & ~n12346 ;
  assign n12348 = ~n12344 & n12347 ;
  assign n12349 = n2754 & n4457 ;
  assign n12350 = n12348 & ~n12349 ;
  assign n12351 = ~x20 & ~n12350 ;
  assign n12352 = ~x20 & ~n12351 ;
  assign n12353 = ~n12350 & ~n12351 ;
  assign n12354 = ~n12352 & ~n12353 ;
  assign n12355 = ~n12343 & n12354 ;
  assign n12356 = n12343 & ~n12354 ;
  assign n12357 = ~n12355 & ~n12356 ;
  assign n12358 = ~n11832 & n12357 ;
  assign n12359 = n11832 & ~n12357 ;
  assign n12360 = ~n12358 & ~n12359 ;
  assign n12361 = ~x91 & n2093 ;
  assign n12362 = ~x89 & n2275 ;
  assign n12363 = ~x90 & n2088 ;
  assign n12364 = ~n12362 & ~n12363 ;
  assign n12365 = ~n12361 & n12364 ;
  assign n12366 = n2096 & n5507 ;
  assign n12367 = n12365 & ~n12366 ;
  assign n12368 = ~x17 & ~n12367 ;
  assign n12369 = ~x17 & ~n12368 ;
  assign n12370 = ~n12367 & ~n12368 ;
  assign n12371 = ~n12369 & ~n12370 ;
  assign n12372 = n12360 & ~n12371 ;
  assign n12373 = n12360 & ~n12372 ;
  assign n12374 = ~n12371 & ~n12372 ;
  assign n12375 = ~n12373 & ~n12374 ;
  assign n12376 = ~n12212 & n12375 ;
  assign n12377 = n12212 & ~n12375 ;
  assign n12378 = ~n12376 & ~n12377 ;
  assign n12379 = ~x94 & n1434 ;
  assign n12380 = ~x92 & n1646 ;
  assign n12381 = ~x93 & n1429 ;
  assign n12382 = ~n12380 & ~n12381 ;
  assign n12383 = ~n12379 & n12382 ;
  assign n12384 = n1437 & n6671 ;
  assign n12385 = n12383 & ~n12384 ;
  assign n12386 = ~x14 & ~n12385 ;
  assign n12387 = ~x14 & ~n12386 ;
  assign n12388 = ~n12385 & ~n12386 ;
  assign n12389 = ~n12387 & ~n12388 ;
  assign n12390 = ~n12378 & ~n12389 ;
  assign n12391 = n12378 & n12389 ;
  assign n12392 = ~n12390 & ~n12391 ;
  assign n12393 = ~n12211 & n12392 ;
  assign n12394 = n12211 & ~n12392 ;
  assign n12395 = ~n12393 & ~n12394 ;
  assign n12396 = ~x97 & n945 ;
  assign n12397 = ~x95 & n1099 ;
  assign n12398 = ~x96 & n940 ;
  assign n12399 = ~n12397 & ~n12398 ;
  assign n12400 = ~n12396 & n12399 ;
  assign n12401 = n948 & n7949 ;
  assign n12402 = n12400 & ~n12401 ;
  assign n12403 = ~x11 & ~n12402 ;
  assign n12404 = ~x11 & ~n12403 ;
  assign n12405 = ~n12402 & ~n12403 ;
  assign n12406 = ~n12404 & ~n12405 ;
  assign n12407 = n12395 & ~n12406 ;
  assign n12408 = n12395 & ~n12407 ;
  assign n12409 = ~n12406 & ~n12407 ;
  assign n12410 = ~n12408 & ~n12409 ;
  assign n12411 = ~n12210 & n12410 ;
  assign n12412 = n12210 & ~n12410 ;
  assign n12413 = ~n12411 & ~n12412 ;
  assign n12414 = ~x100 & n574 ;
  assign n12415 = ~x98 & n673 ;
  assign n12416 = ~x99 & n569 ;
  assign n12417 = ~n12415 & ~n12416 ;
  assign n12418 = ~n12414 & n12417 ;
  assign n12419 = n577 & n9338 ;
  assign n12420 = n12418 & ~n12419 ;
  assign n12421 = ~x8 & ~n12420 ;
  assign n12422 = ~x8 & ~n12421 ;
  assign n12423 = ~n12420 & ~n12421 ;
  assign n12424 = ~n12422 & ~n12423 ;
  assign n12425 = n12413 & n12424 ;
  assign n12426 = ~n12413 & ~n12424 ;
  assign n12427 = ~n12425 & ~n12426 ;
  assign n12428 = ~n12209 & n12427 ;
  assign n12429 = n12209 & ~n12427 ;
  assign n12430 = ~n12428 & ~n12429 ;
  assign n12431 = ~n12207 & n12430 ;
  assign n12432 = ~n12207 & ~n12431 ;
  assign n12433 = n12430 & ~n12431 ;
  assign n12434 = ~n12432 & ~n12433 ;
  assign n12435 = ~n12196 & ~n12434 ;
  assign n12436 = ~n12196 & ~n12435 ;
  assign n12437 = ~n12434 & ~n12435 ;
  assign n12438 = ~n12436 & ~n12437 ;
  assign n12439 = ~x106 & n164 ;
  assign n12440 = ~x104 & n205 ;
  assign n12441 = ~x105 & n162 ;
  assign n12442 = ~n12440 & ~n12441 ;
  assign n12443 = ~n12439 & n12442 ;
  assign n12444 = ~n11643 & ~n11905 ;
  assign n12445 = n12178 & ~n12444 ;
  assign n12446 = ~n12178 & n12444 ;
  assign n12447 = ~n12445 & ~n12446 ;
  assign n12448 = n167 & n12447 ;
  assign n12449 = n12443 & ~n12448 ;
  assign n12450 = ~x2 & ~n12449 ;
  assign n12451 = ~x2 & ~n12450 ;
  assign n12452 = ~n12449 & ~n12450 ;
  assign n12453 = ~n12451 & ~n12452 ;
  assign n12454 = ~n12438 & ~n12453 ;
  assign n12455 = ~n12438 & ~n12454 ;
  assign n12456 = ~n12453 & ~n12454 ;
  assign n12457 = ~n12455 & ~n12456 ;
  assign n12458 = ~n11915 & ~n11917 ;
  assign n12459 = ~n12457 & ~n12458 ;
  assign n12460 = n12457 & n12458 ;
  assign n12461 = ~n12459 & ~n12460 ;
  assign n12464 = ~n12461 & ~x170 ;
  assign n12465 = ~n12463 & ~n12464 ;
  assign n12466 = ~n12162 & ~n12166 ;
  assign n12467 = ~n12157 & ~n12159 ;
  assign n12468 = ~n12121 & ~n12124 ;
  assign n12469 = ~n11940 & ~n12106 ;
  assign n12470 = ~n12103 & ~n12469 ;
  assign n12471 = x92 & n2093 ;
  assign n12472 = x90 & n2275 ;
  assign n12473 = x91 & n2088 ;
  assign n12474 = ~n12472 & ~n12473 ;
  assign n12475 = ~n12471 & n12474 ;
  assign n12476 = n2096 & n5710 ;
  assign n12477 = n12475 & ~n12476 ;
  assign n12478 = x17 & ~n12477 ;
  assign n12479 = x17 & ~n12478 ;
  assign n12480 = ~n12477 & ~n12478 ;
  assign n12481 = ~n12479 & ~n12480 ;
  assign n12482 = ~n12013 & ~n12017 ;
  assign n12483 = ~n12008 & ~n12010 ;
  assign n12484 = n11478 & n11959 ;
  assign n12485 = ~n11974 & ~n12484 ;
  assign n12486 = x68 & n10905 ;
  assign n12487 = x66 & n11466 ;
  assign n12488 = x67 & n10900 ;
  assign n12489 = ~n12487 & ~n12488 ;
  assign n12490 = ~n12486 & n12489 ;
  assign n12491 = n317 & n10908 ;
  assign n12492 = n12490 & ~n12491 ;
  assign n12493 = x41 & ~n12492 ;
  assign n12494 = x41 & ~n12493 ;
  assign n12495 = ~n12492 & ~n12493 ;
  assign n12496 = ~n12494 & ~n12495 ;
  assign n12497 = x44 & ~n11959 ;
  assign n12498 = ~x42 & x43 ;
  assign n12499 = x42 & ~x43 ;
  assign n12500 = ~n12498 & ~n12499 ;
  assign n12501 = n11958 & ~n12500 ;
  assign n12502 = x64 & n12501 ;
  assign n12503 = ~x43 & x44 ;
  assign n12504 = x43 & ~x44 ;
  assign n12505 = ~n12503 & ~n12504 ;
  assign n12506 = ~n11958 & n12505 ;
  assign n12507 = x65 & n12506 ;
  assign n12508 = ~n12502 & ~n12507 ;
  assign n12509 = ~n11958 & ~n12505 ;
  assign n12510 = ~n152 & n12509 ;
  assign n12511 = n12508 & ~n12510 ;
  assign n12512 = x44 & ~n12511 ;
  assign n12513 = x44 & ~n12512 ;
  assign n12514 = ~n12511 & ~n12512 ;
  assign n12515 = ~n12513 & ~n12514 ;
  assign n12516 = n12497 & ~n12515 ;
  assign n12517 = ~n12497 & n12515 ;
  assign n12518 = ~n12516 & ~n12517 ;
  assign n12519 = n12496 & ~n12518 ;
  assign n12520 = ~n12496 & n12518 ;
  assign n12521 = ~n12519 & ~n12520 ;
  assign n12522 = ~n12485 & n12521 ;
  assign n12523 = n12485 & ~n12521 ;
  assign n12524 = ~n12522 & ~n12523 ;
  assign n12525 = x71 & n9433 ;
  assign n12526 = x69 & n9915 ;
  assign n12527 = x70 & n9428 ;
  assign n12528 = ~n12526 & ~n12527 ;
  assign n12529 = ~n12525 & n12528 ;
  assign n12530 = n558 & n9436 ;
  assign n12531 = n12529 & ~n12530 ;
  assign n12532 = x38 & ~n12531 ;
  assign n12533 = x38 & ~n12532 ;
  assign n12534 = ~n12531 & ~n12532 ;
  assign n12535 = ~n12533 & ~n12534 ;
  assign n12536 = n12524 & ~n12535 ;
  assign n12537 = n12524 & ~n12536 ;
  assign n12538 = ~n12535 & ~n12536 ;
  assign n12539 = ~n12537 & ~n12538 ;
  assign n12540 = ~n11988 & ~n11994 ;
  assign n12541 = n12539 & n12540 ;
  assign n12542 = ~n12539 & ~n12540 ;
  assign n12543 = ~n12541 & ~n12542 ;
  assign n12544 = x74 & n8006 ;
  assign n12545 = x72 & n8474 ;
  assign n12546 = x73 & n8001 ;
  assign n12547 = ~n12545 & ~n12546 ;
  assign n12548 = ~n12544 & n12547 ;
  assign n12549 = n994 & n8009 ;
  assign n12550 = n12548 & ~n12549 ;
  assign n12551 = x35 & ~n12550 ;
  assign n12552 = x35 & ~n12551 ;
  assign n12553 = ~n12550 & ~n12551 ;
  assign n12554 = ~n12552 & ~n12553 ;
  assign n12555 = n12543 & ~n12554 ;
  assign n12556 = ~n12543 & n12554 ;
  assign n12557 = ~n12483 & ~n12556 ;
  assign n12558 = ~n12555 & n12557 ;
  assign n12559 = ~n12483 & ~n12558 ;
  assign n12560 = ~n12555 & ~n12558 ;
  assign n12561 = ~n12556 & n12560 ;
  assign n12562 = ~n12559 & ~n12561 ;
  assign n12563 = x77 & n6725 ;
  assign n12564 = x75 & n7129 ;
  assign n12565 = x76 & n6720 ;
  assign n12566 = ~n12564 & ~n12565 ;
  assign n12567 = ~n12563 & n12566 ;
  assign n12568 = n1502 & n6728 ;
  assign n12569 = n12567 & ~n12568 ;
  assign n12570 = x32 & ~n12569 ;
  assign n12571 = x32 & ~n12570 ;
  assign n12572 = ~n12569 & ~n12570 ;
  assign n12573 = ~n12571 & ~n12572 ;
  assign n12574 = n12562 & n12573 ;
  assign n12575 = ~n12562 & ~n12573 ;
  assign n12576 = ~n12574 & ~n12575 ;
  assign n12577 = ~n12482 & n12576 ;
  assign n12578 = n12482 & ~n12576 ;
  assign n12579 = ~n12577 & ~n12578 ;
  assign n12580 = x80 & n5560 ;
  assign n12581 = x78 & n5943 ;
  assign n12582 = x79 & n5555 ;
  assign n12583 = ~n12581 & ~n12582 ;
  assign n12584 = ~n12580 & n12583 ;
  assign n12585 = n2028 & n5563 ;
  assign n12586 = n12584 & ~n12585 ;
  assign n12587 = x29 & ~n12586 ;
  assign n12588 = x29 & ~n12587 ;
  assign n12589 = ~n12586 & ~n12587 ;
  assign n12590 = ~n12588 & ~n12589 ;
  assign n12591 = n12579 & ~n12590 ;
  assign n12592 = n12579 & ~n12591 ;
  assign n12593 = ~n12590 & ~n12591 ;
  assign n12594 = ~n12592 & ~n12593 ;
  assign n12595 = ~n11942 & ~n12035 ;
  assign n12596 = ~n12032 & ~n12595 ;
  assign n12597 = n12594 & n12596 ;
  assign n12598 = ~n12594 & ~n12596 ;
  assign n12599 = ~n12597 & ~n12598 ;
  assign n12600 = x83 & n4531 ;
  assign n12601 = x81 & n4847 ;
  assign n12602 = x82 & n4526 ;
  assign n12603 = ~n12601 & ~n12602 ;
  assign n12604 = ~n12600 & n12603 ;
  assign n12605 = n2843 & n4534 ;
  assign n12606 = n12604 & ~n12605 ;
  assign n12607 = x26 & ~n12606 ;
  assign n12608 = x26 & ~n12607 ;
  assign n12609 = ~n12606 & ~n12607 ;
  assign n12610 = ~n12608 & ~n12609 ;
  assign n12611 = n12599 & ~n12610 ;
  assign n12612 = n12599 & ~n12611 ;
  assign n12613 = ~n12610 & ~n12611 ;
  assign n12614 = ~n12612 & ~n12613 ;
  assign n12615 = ~n12050 & ~n12053 ;
  assign n12616 = n12614 & n12615 ;
  assign n12617 = ~n12614 & ~n12615 ;
  assign n12618 = ~n12616 & ~n12617 ;
  assign n12619 = x86 & n3589 ;
  assign n12620 = x84 & n3878 ;
  assign n12621 = x85 & n3584 ;
  assign n12622 = ~n12620 & ~n12621 ;
  assign n12623 = ~n12619 & n12622 ;
  assign n12624 = n3592 & n3686 ;
  assign n12625 = n12623 & ~n12624 ;
  assign n12626 = x23 & ~n12625 ;
  assign n12627 = x23 & ~n12626 ;
  assign n12628 = ~n12625 & ~n12626 ;
  assign n12629 = ~n12627 & ~n12628 ;
  assign n12630 = n12618 & ~n12629 ;
  assign n12631 = n12618 & ~n12630 ;
  assign n12632 = ~n12629 & ~n12630 ;
  assign n12633 = ~n12631 & ~n12632 ;
  assign n12634 = ~n12067 & ~n12073 ;
  assign n12635 = n12633 & n12634 ;
  assign n12636 = ~n12633 & ~n12634 ;
  assign n12637 = ~n12635 & ~n12636 ;
  assign n12638 = x89 & n2751 ;
  assign n12639 = x87 & n3020 ;
  assign n12640 = x88 & n2746 ;
  assign n12641 = ~n12639 & ~n12640 ;
  assign n12642 = ~n12638 & n12641 ;
  assign n12643 = n2754 & n4488 ;
  assign n12644 = n12642 & ~n12643 ;
  assign n12645 = x20 & ~n12644 ;
  assign n12646 = x20 & ~n12645 ;
  assign n12647 = ~n12644 & ~n12645 ;
  assign n12648 = ~n12646 & ~n12647 ;
  assign n12649 = n12637 & ~n12648 ;
  assign n12650 = n12637 & ~n12649 ;
  assign n12651 = ~n12648 & ~n12649 ;
  assign n12652 = ~n12650 & ~n12651 ;
  assign n12653 = ~n12087 & ~n12089 ;
  assign n12654 = ~n12652 & ~n12653 ;
  assign n12655 = n12652 & n12653 ;
  assign n12656 = ~n12654 & ~n12655 ;
  assign n12657 = ~n12481 & n12656 ;
  assign n12658 = ~n12481 & ~n12657 ;
  assign n12659 = n12656 & ~n12657 ;
  assign n12660 = ~n12658 & ~n12659 ;
  assign n12661 = ~n12470 & ~n12660 ;
  assign n12662 = ~n12470 & ~n12661 ;
  assign n12663 = ~n12660 & ~n12661 ;
  assign n12664 = ~n12662 & ~n12663 ;
  assign n12665 = x95 & n1434 ;
  assign n12666 = x93 & n1646 ;
  assign n12667 = x94 & n1429 ;
  assign n12668 = ~n12666 & ~n12667 ;
  assign n12669 = ~n12665 & n12668 ;
  assign n12670 = n1437 & n6894 ;
  assign n12671 = n12669 & ~n12670 ;
  assign n12672 = x14 & ~n12671 ;
  assign n12673 = x14 & ~n12672 ;
  assign n12674 = ~n12671 & ~n12672 ;
  assign n12675 = ~n12673 & ~n12674 ;
  assign n12676 = n12664 & n12675 ;
  assign n12677 = ~n12664 & ~n12675 ;
  assign n12678 = ~n12676 & ~n12677 ;
  assign n12679 = ~n12468 & n12678 ;
  assign n12680 = n12468 & ~n12678 ;
  assign n12681 = ~n12679 & ~n12680 ;
  assign n12682 = x98 & n945 ;
  assign n12683 = x96 & n1099 ;
  assign n12684 = x97 & n940 ;
  assign n12685 = ~n12683 & ~n12684 ;
  assign n12686 = ~n12682 & n12685 ;
  assign n12687 = n948 & n8196 ;
  assign n12688 = n12686 & ~n12687 ;
  assign n12689 = x11 & ~n12688 ;
  assign n12690 = x11 & ~n12689 ;
  assign n12691 = ~n12688 & ~n12689 ;
  assign n12692 = ~n12690 & ~n12691 ;
  assign n12693 = n12681 & ~n12692 ;
  assign n12694 = n12681 & ~n12693 ;
  assign n12695 = ~n12692 & ~n12693 ;
  assign n12696 = ~n12694 & ~n12695 ;
  assign n12697 = ~n11938 & ~n12141 ;
  assign n12698 = ~n12138 & ~n12697 ;
  assign n12699 = n12696 & n12698 ;
  assign n12700 = ~n12696 & ~n12698 ;
  assign n12701 = ~n12699 & ~n12700 ;
  assign n12702 = x101 & n574 ;
  assign n12703 = x99 & n673 ;
  assign n12704 = x100 & n569 ;
  assign n12705 = ~n12703 & ~n12704 ;
  assign n12706 = ~n12702 & n12705 ;
  assign n12707 = n577 & n9601 ;
  assign n12708 = n12706 & ~n12707 ;
  assign n12709 = x8 & ~n12708 ;
  assign n12710 = x8 & ~n12709 ;
  assign n12711 = ~n12708 & ~n12709 ;
  assign n12712 = ~n12710 & ~n12711 ;
  assign n12713 = n12701 & ~n12712 ;
  assign n12714 = ~n12701 & n12712 ;
  assign n12715 = ~n12467 & ~n12714 ;
  assign n12716 = ~n12713 & n12715 ;
  assign n12717 = ~n12467 & ~n12716 ;
  assign n12718 = ~n12713 & ~n12716 ;
  assign n12719 = ~n12714 & n12718 ;
  assign n12720 = ~n12717 & ~n12719 ;
  assign n12721 = x104 & n293 ;
  assign n12722 = x102 & n373 ;
  assign n12723 = x103 & n288 ;
  assign n12724 = ~n12722 & ~n12723 ;
  assign n12725 = ~n12721 & n12724 ;
  assign n12726 = n296 & n11116 ;
  assign n12727 = n12725 & ~n12726 ;
  assign n12728 = x5 & ~n12727 ;
  assign n12729 = x5 & ~n12728 ;
  assign n12730 = ~n12727 & ~n12728 ;
  assign n12731 = ~n12729 & ~n12730 ;
  assign n12732 = n12720 & n12731 ;
  assign n12733 = ~n12720 & ~n12731 ;
  assign n12734 = ~n12732 & ~n12733 ;
  assign n12735 = ~n12466 & n12734 ;
  assign n12736 = n12466 & ~n12734 ;
  assign n12737 = ~n12735 & ~n12736 ;
  assign n12738 = x107 & n146 ;
  assign n12739 = x105 & n182 ;
  assign n12740 = x106 & n141 ;
  assign n12741 = ~n12739 & ~n12740 ;
  assign n12742 = ~n12738 & n12741 ;
  assign n12743 = ~n12177 & ~n12179 ;
  assign n12744 = ~x106 & ~x107 ;
  assign n12745 = x106 & x107 ;
  assign n12746 = ~n12744 & ~n12745 ;
  assign n12747 = ~n12743 & n12746 ;
  assign n12748 = n12743 & ~n12746 ;
  assign n12749 = ~n12747 & ~n12748 ;
  assign n12750 = n149 & n12749 ;
  assign n12751 = n12742 & ~n12750 ;
  assign n12752 = x2 & ~n12751 ;
  assign n12753 = x2 & ~n12752 ;
  assign n12754 = ~n12751 & ~n12752 ;
  assign n12755 = ~n12753 & ~n12754 ;
  assign n12756 = n12737 & ~n12755 ;
  assign n12757 = n12737 & ~n12756 ;
  assign n12758 = ~n12755 & ~n12756 ;
  assign n12759 = ~n12757 & ~n12758 ;
  assign n12760 = ~n12188 & ~n12193 ;
  assign n12761 = ~n12759 & ~n12760 ;
  assign n12762 = n12759 & n12760 ;
  assign n12763 = ~n12761 & ~n12762 ;
  assign n13050 = n12763 & x171 ;
  assign n12764 = ~n12431 & ~n12435 ;
  assign n12765 = ~n12426 & ~n12428 ;
  assign n12766 = ~n12390 & ~n12393 ;
  assign n12767 = ~n12212 & ~n12375 ;
  assign n12768 = ~n12372 & ~n12767 ;
  assign n12769 = ~x92 & n2093 ;
  assign n12770 = ~x90 & n2275 ;
  assign n12771 = ~x91 & n2088 ;
  assign n12772 = ~n12770 & ~n12771 ;
  assign n12773 = ~n12769 & n12772 ;
  assign n12774 = n2096 & n5896 ;
  assign n12775 = n12773 & ~n12774 ;
  assign n12776 = ~x17 & ~n12775 ;
  assign n12777 = ~x17 & ~n12776 ;
  assign n12778 = ~n12775 & ~n12776 ;
  assign n12779 = ~n12777 & ~n12778 ;
  assign n12780 = ~n12282 & ~n12286 ;
  assign n12781 = ~n12277 & ~n12279 ;
  assign n12782 = n11740 & n12228 ;
  assign n12783 = ~n12243 & ~n12782 ;
  assign n12784 = ~x68 & n10905 ;
  assign n12785 = ~x66 & n11466 ;
  assign n12786 = ~x67 & n10900 ;
  assign n12787 = ~n12785 & ~n12786 ;
  assign n12788 = ~n12784 & n12787 ;
  assign n12789 = n352 & n10908 ;
  assign n12790 = n12788 & ~n12789 ;
  assign n12791 = ~x41 & ~n12790 ;
  assign n12792 = ~x41 & ~n12791 ;
  assign n12793 = ~n12790 & ~n12791 ;
  assign n12794 = ~n12792 & ~n12793 ;
  assign n12795 = ~x44 & ~n12228 ;
  assign n12796 = ~x64 & n12501 ;
  assign n12797 = ~x65 & n12506 ;
  assign n12798 = ~n12796 & ~n12797 ;
  assign n12799 = ~n12510 & n12798 ;
  assign n12800 = ~x44 & ~n12799 ;
  assign n12801 = ~x44 & ~n12800 ;
  assign n12802 = ~n12799 & ~n12800 ;
  assign n12803 = ~n12801 & ~n12802 ;
  assign n12804 = n12795 & ~n12803 ;
  assign n12805 = ~n12795 & n12803 ;
  assign n12806 = ~n12804 & ~n12805 ;
  assign n12807 = n12794 & ~n12806 ;
  assign n12808 = ~n12794 & n12806 ;
  assign n12809 = ~n12807 & ~n12808 ;
  assign n12810 = ~n12783 & n12809 ;
  assign n12811 = n12783 & ~n12809 ;
  assign n12812 = ~n12810 & ~n12811 ;
  assign n12813 = ~x71 & n9433 ;
  assign n12814 = ~x69 & n9915 ;
  assign n12815 = ~x70 & n9428 ;
  assign n12816 = ~n12814 & ~n12815 ;
  assign n12817 = ~n12813 & n12816 ;
  assign n12818 = n622 & n9436 ;
  assign n12819 = n12817 & ~n12818 ;
  assign n12820 = ~x38 & ~n12819 ;
  assign n12821 = ~x38 & ~n12820 ;
  assign n12822 = ~n12819 & ~n12820 ;
  assign n12823 = ~n12821 & ~n12822 ;
  assign n12824 = n12812 & ~n12823 ;
  assign n12825 = n12812 & ~n12824 ;
  assign n12826 = ~n12823 & ~n12824 ;
  assign n12827 = ~n12825 & ~n12826 ;
  assign n12828 = ~n12257 & ~n12263 ;
  assign n12829 = n12827 & n12828 ;
  assign n12830 = ~n12827 & ~n12828 ;
  assign n12831 = ~n12829 & ~n12830 ;
  assign n12832 = ~x74 & n8006 ;
  assign n12833 = ~x72 & n8474 ;
  assign n12834 = ~x73 & n8001 ;
  assign n12835 = ~n12833 & ~n12834 ;
  assign n12836 = ~n12832 & n12835 ;
  assign n12837 = n1066 & n8009 ;
  assign n12838 = n12836 & ~n12837 ;
  assign n12839 = ~x35 & ~n12838 ;
  assign n12840 = ~x35 & ~n12839 ;
  assign n12841 = ~n12838 & ~n12839 ;
  assign n12842 = ~n12840 & ~n12841 ;
  assign n12843 = n12831 & ~n12842 ;
  assign n12844 = ~n12831 & n12842 ;
  assign n12845 = ~n12781 & ~n12844 ;
  assign n12846 = ~n12843 & n12845 ;
  assign n12847 = ~n12781 & ~n12846 ;
  assign n12848 = ~n12843 & ~n12846 ;
  assign n12849 = ~n12844 & n12848 ;
  assign n12850 = ~n12847 & ~n12849 ;
  assign n12851 = ~x77 & n6725 ;
  assign n12852 = ~x75 & n7129 ;
  assign n12853 = ~x76 & n6720 ;
  assign n12854 = ~n12852 & ~n12853 ;
  assign n12855 = ~n12851 & n12854 ;
  assign n12856 = n1594 & n6728 ;
  assign n12857 = n12855 & ~n12856 ;
  assign n12858 = ~x32 & ~n12857 ;
  assign n12859 = ~x32 & ~n12858 ;
  assign n12860 = ~n12857 & ~n12858 ;
  assign n12861 = ~n12859 & ~n12860 ;
  assign n12862 = n12850 & n12861 ;
  assign n12863 = ~n12850 & ~n12861 ;
  assign n12864 = ~n12862 & ~n12863 ;
  assign n12865 = ~n12780 & n12864 ;
  assign n12866 = n12780 & ~n12864 ;
  assign n12867 = ~n12865 & ~n12866 ;
  assign n12868 = ~x80 & n5560 ;
  assign n12869 = ~x78 & n5943 ;
  assign n12870 = ~x79 & n5555 ;
  assign n12871 = ~n12869 & ~n12870 ;
  assign n12872 = ~n12868 & n12871 ;
  assign n12873 = n2145 & n5563 ;
  assign n12874 = n12872 & ~n12873 ;
  assign n12875 = ~x29 & ~n12874 ;
  assign n12876 = ~x29 & ~n12875 ;
  assign n12877 = ~n12874 & ~n12875 ;
  assign n12878 = ~n12876 & ~n12877 ;
  assign n12879 = n12867 & ~n12878 ;
  assign n12880 = n12867 & ~n12879 ;
  assign n12881 = ~n12878 & ~n12879 ;
  assign n12882 = ~n12880 & ~n12881 ;
  assign n12883 = ~n12214 & ~n12304 ;
  assign n12884 = ~n12301 & ~n12883 ;
  assign n12885 = n12882 & n12884 ;
  assign n12886 = ~n12882 & ~n12884 ;
  assign n12887 = ~n12885 & ~n12886 ;
  assign n12888 = ~x83 & n4531 ;
  assign n12889 = ~x81 & n4847 ;
  assign n12890 = ~x82 & n4526 ;
  assign n12891 = ~n12889 & ~n12890 ;
  assign n12892 = ~n12888 & n12891 ;
  assign n12893 = n2972 & n4534 ;
  assign n12894 = n12892 & ~n12893 ;
  assign n12895 = ~x26 & ~n12894 ;
  assign n12896 = ~x26 & ~n12895 ;
  assign n12897 = ~n12894 & ~n12895 ;
  assign n12898 = ~n12896 & ~n12897 ;
  assign n12899 = n12887 & ~n12898 ;
  assign n12900 = n12887 & ~n12899 ;
  assign n12901 = ~n12898 & ~n12899 ;
  assign n12902 = ~n12900 & ~n12901 ;
  assign n12903 = ~n12319 & ~n12322 ;
  assign n12904 = n12902 & n12903 ;
  assign n12905 = ~n12902 & ~n12903 ;
  assign n12906 = ~n12904 & ~n12905 ;
  assign n12907 = ~x86 & n3589 ;
  assign n12908 = ~x84 & n3878 ;
  assign n12909 = ~x85 & n3584 ;
  assign n12910 = ~n12908 & ~n12909 ;
  assign n12911 = ~n12907 & n12910 ;
  assign n12912 = n3592 & n3832 ;
  assign n12913 = n12911 & ~n12912 ;
  assign n12914 = ~x23 & ~n12913 ;
  assign n12915 = ~x23 & ~n12914 ;
  assign n12916 = ~n12913 & ~n12914 ;
  assign n12917 = ~n12915 & ~n12916 ;
  assign n12918 = n12906 & ~n12917 ;
  assign n12919 = n12906 & ~n12918 ;
  assign n12920 = ~n12917 & ~n12918 ;
  assign n12921 = ~n12919 & ~n12920 ;
  assign n12922 = ~n12336 & ~n12342 ;
  assign n12923 = n12921 & n12922 ;
  assign n12924 = ~n12921 & ~n12922 ;
  assign n12925 = ~n12923 & ~n12924 ;
  assign n12926 = ~x89 & n2751 ;
  assign n12927 = ~x87 & n3020 ;
  assign n12928 = ~x88 & n2746 ;
  assign n12929 = ~n12927 & ~n12928 ;
  assign n12930 = ~n12926 & n12929 ;
  assign n12931 = n2754 & n4664 ;
  assign n12932 = n12930 & ~n12931 ;
  assign n12933 = ~x20 & ~n12932 ;
  assign n12934 = ~x20 & ~n12933 ;
  assign n12935 = ~n12932 & ~n12933 ;
  assign n12936 = ~n12934 & ~n12935 ;
  assign n12937 = n12925 & ~n12936 ;
  assign n12938 = n12925 & ~n12937 ;
  assign n12939 = ~n12936 & ~n12937 ;
  assign n12940 = ~n12938 & ~n12939 ;
  assign n12941 = ~n12356 & ~n12358 ;
  assign n12942 = ~n12940 & ~n12941 ;
  assign n12943 = n12940 & n12941 ;
  assign n12944 = ~n12942 & ~n12943 ;
  assign n12945 = ~n12779 & n12944 ;
  assign n12946 = ~n12779 & ~n12945 ;
  assign n12947 = n12944 & ~n12945 ;
  assign n12948 = ~n12946 & ~n12947 ;
  assign n12949 = ~n12768 & ~n12948 ;
  assign n12950 = ~n12768 & ~n12949 ;
  assign n12951 = ~n12948 & ~n12949 ;
  assign n12952 = ~n12950 & ~n12951 ;
  assign n12953 = ~x95 & n1434 ;
  assign n12954 = ~x93 & n1646 ;
  assign n12955 = ~x94 & n1429 ;
  assign n12956 = ~n12954 & ~n12955 ;
  assign n12957 = ~n12953 & n12956 ;
  assign n12958 = n1437 & n7100 ;
  assign n12959 = n12957 & ~n12958 ;
  assign n12960 = ~x14 & ~n12959 ;
  assign n12961 = ~x14 & ~n12960 ;
  assign n12962 = ~n12959 & ~n12960 ;
  assign n12963 = ~n12961 & ~n12962 ;
  assign n12964 = n12952 & n12963 ;
  assign n12965 = ~n12952 & ~n12963 ;
  assign n12966 = ~n12964 & ~n12965 ;
  assign n12967 = ~n12766 & n12966 ;
  assign n12968 = n12766 & ~n12966 ;
  assign n12969 = ~n12967 & ~n12968 ;
  assign n12970 = ~x98 & n945 ;
  assign n12971 = ~x96 & n1099 ;
  assign n12972 = ~x97 & n940 ;
  assign n12973 = ~n12971 & ~n12972 ;
  assign n12974 = ~n12970 & n12973 ;
  assign n12975 = n948 & n8426 ;
  assign n12976 = n12974 & ~n12975 ;
  assign n12977 = ~x11 & ~n12976 ;
  assign n12978 = ~x11 & ~n12977 ;
  assign n12979 = ~n12976 & ~n12977 ;
  assign n12980 = ~n12978 & ~n12979 ;
  assign n12981 = n12969 & ~n12980 ;
  assign n12982 = n12969 & ~n12981 ;
  assign n12983 = ~n12980 & ~n12981 ;
  assign n12984 = ~n12982 & ~n12983 ;
  assign n12985 = ~n12210 & ~n12410 ;
  assign n12986 = ~n12407 & ~n12985 ;
  assign n12987 = n12984 & n12986 ;
  assign n12988 = ~n12984 & ~n12986 ;
  assign n12989 = ~n12987 & ~n12988 ;
  assign n12990 = ~x101 & n574 ;
  assign n12991 = ~x99 & n673 ;
  assign n12992 = ~x100 & n569 ;
  assign n12993 = ~n12991 & ~n12992 ;
  assign n12994 = ~n12990 & n12993 ;
  assign n12995 = n577 & n9844 ;
  assign n12996 = n12994 & ~n12995 ;
  assign n12997 = ~x8 & ~n12996 ;
  assign n12998 = ~x8 & ~n12997 ;
  assign n12999 = ~n12996 & ~n12997 ;
  assign n13000 = ~n12998 & ~n12999 ;
  assign n13001 = n12989 & ~n13000 ;
  assign n13002 = ~n12989 & n13000 ;
  assign n13003 = ~n12765 & ~n13002 ;
  assign n13004 = ~n13001 & n13003 ;
  assign n13005 = ~n12765 & ~n13004 ;
  assign n13006 = ~n13001 & ~n13004 ;
  assign n13007 = ~n13002 & n13006 ;
  assign n13008 = ~n13005 & ~n13007 ;
  assign n13009 = ~x104 & n293 ;
  assign n13010 = ~x102 & n373 ;
  assign n13011 = ~x103 & n288 ;
  assign n13012 = ~n13010 & ~n13011 ;
  assign n13013 = ~n13009 & n13012 ;
  assign n13014 = n296 & n11380 ;
  assign n13015 = n13013 & ~n13014 ;
  assign n13016 = ~x5 & ~n13015 ;
  assign n13017 = ~x5 & ~n13016 ;
  assign n13018 = ~n13015 & ~n13016 ;
  assign n13019 = ~n13017 & ~n13018 ;
  assign n13020 = n13008 & n13019 ;
  assign n13021 = ~n13008 & ~n13019 ;
  assign n13022 = ~n13020 & ~n13021 ;
  assign n13023 = ~n12764 & n13022 ;
  assign n13024 = n12764 & ~n13022 ;
  assign n13025 = ~n13023 & ~n13024 ;
  assign n13026 = ~x107 & n164 ;
  assign n13027 = ~x105 & n205 ;
  assign n13028 = ~x106 & n162 ;
  assign n13029 = ~n13027 & ~n13028 ;
  assign n13030 = ~n13026 & n13029 ;
  assign n13031 = ~n12176 & ~n12445 ;
  assign n13032 = n12746 & ~n13031 ;
  assign n13033 = ~n12746 & n13031 ;
  assign n13034 = ~n13032 & ~n13033 ;
  assign n13035 = n167 & n13034 ;
  assign n13036 = n13030 & ~n13035 ;
  assign n13037 = ~x2 & ~n13036 ;
  assign n13038 = ~x2 & ~n13037 ;
  assign n13039 = ~n13036 & ~n13037 ;
  assign n13040 = ~n13038 & ~n13039 ;
  assign n13041 = n13025 & ~n13040 ;
  assign n13042 = n13025 & ~n13041 ;
  assign n13043 = ~n13040 & ~n13041 ;
  assign n13044 = ~n13042 & ~n13043 ;
  assign n13045 = ~n12454 & ~n12459 ;
  assign n13046 = ~n13044 & ~n13045 ;
  assign n13047 = n13044 & n13045 ;
  assign n13048 = ~n13046 & ~n13047 ;
  assign n13051 = ~n13048 & ~x171 ;
  assign n13052 = ~n13050 & ~n13051 ;
  assign n13053 = ~n12756 & ~n12761 ;
  assign n13054 = ~n12733 & ~n12735 ;
  assign n13055 = x105 & n293 ;
  assign n13056 = x103 & n373 ;
  assign n13057 = x104 & n288 ;
  assign n13058 = ~n13056 & ~n13057 ;
  assign n13059 = ~n13055 & n13058 ;
  assign n13060 = n296 & n11648 ;
  assign n13061 = n13059 & ~n13060 ;
  assign n13062 = x5 & ~n13061 ;
  assign n13063 = x5 & ~n13062 ;
  assign n13064 = ~n13061 & ~n13062 ;
  assign n13065 = ~n13063 & ~n13064 ;
  assign n13066 = ~n12677 & ~n12679 ;
  assign n13067 = x96 & n1434 ;
  assign n13068 = x94 & n1646 ;
  assign n13069 = x95 & n1429 ;
  assign n13070 = ~n13068 & ~n13069 ;
  assign n13071 = ~n13067 & n13070 ;
  assign n13072 = n1437 & n7321 ;
  assign n13073 = n13071 & ~n13072 ;
  assign n13074 = x14 & ~n13073 ;
  assign n13075 = x14 & ~n13074 ;
  assign n13076 = ~n13073 & ~n13074 ;
  assign n13077 = ~n13075 & ~n13076 ;
  assign n13078 = ~n12657 & ~n12661 ;
  assign n13079 = x93 & n2093 ;
  assign n13080 = x91 & n2275 ;
  assign n13081 = x92 & n2088 ;
  assign n13082 = ~n13080 & ~n13081 ;
  assign n13083 = ~n13079 & n13082 ;
  assign n13084 = n2096 & n6094 ;
  assign n13085 = n13083 & ~n13084 ;
  assign n13086 = x17 & ~n13085 ;
  assign n13087 = x17 & ~n13086 ;
  assign n13088 = ~n13085 & ~n13086 ;
  assign n13089 = ~n13087 & ~n13088 ;
  assign n13090 = ~n12649 & ~n12654 ;
  assign n13091 = ~n12630 & ~n12636 ;
  assign n13092 = ~n12591 & ~n12598 ;
  assign n13093 = x81 & n5560 ;
  assign n13094 = x79 & n5943 ;
  assign n13095 = x80 & n5555 ;
  assign n13096 = ~n13094 & ~n13095 ;
  assign n13097 = ~n13093 & n13096 ;
  assign n13098 = n2348 & n5563 ;
  assign n13099 = n13097 & ~n13098 ;
  assign n13100 = x29 & ~n13099 ;
  assign n13101 = x29 & ~n13100 ;
  assign n13102 = ~n13099 & ~n13100 ;
  assign n13103 = ~n13101 & ~n13102 ;
  assign n13104 = ~n12575 & ~n12577 ;
  assign n13105 = x78 & n6725 ;
  assign n13106 = x76 & n7129 ;
  assign n13107 = x77 & n6720 ;
  assign n13108 = ~n13106 & ~n13107 ;
  assign n13109 = ~n13105 & n13108 ;
  assign n13110 = n1624 & n6728 ;
  assign n13111 = n13109 & ~n13110 ;
  assign n13112 = x32 & ~n13111 ;
  assign n13113 = x32 & ~n13112 ;
  assign n13114 = ~n13111 & ~n13112 ;
  assign n13115 = ~n13113 & ~n13114 ;
  assign n13116 = ~n12536 & ~n12542 ;
  assign n13117 = x72 & n9433 ;
  assign n13118 = x70 & n9915 ;
  assign n13119 = x71 & n9428 ;
  assign n13120 = ~n13118 & ~n13119 ;
  assign n13121 = ~n13117 & n13120 ;
  assign n13122 = n717 & n9436 ;
  assign n13123 = n13121 & ~n13122 ;
  assign n13124 = x38 & ~n13123 ;
  assign n13125 = x38 & ~n13124 ;
  assign n13126 = ~n13123 & ~n13124 ;
  assign n13127 = ~n13125 & ~n13126 ;
  assign n13128 = ~n12520 & ~n12522 ;
  assign n13129 = x66 & n12506 ;
  assign n13130 = n11958 & ~n12505 ;
  assign n13131 = n12500 & n13130 ;
  assign n13132 = x64 & n13131 ;
  assign n13133 = x65 & n12501 ;
  assign n13134 = ~n13132 & ~n13133 ;
  assign n13135 = ~n13129 & n13134 ;
  assign n13136 = n194 & n12509 ;
  assign n13137 = n13135 & ~n13136 ;
  assign n13138 = x44 & ~n13137 ;
  assign n13139 = x44 & ~n13138 ;
  assign n13140 = ~n13137 & ~n13138 ;
  assign n13141 = ~n13139 & ~n13140 ;
  assign n13142 = ~n12516 & n13141 ;
  assign n13143 = n12516 & ~n13141 ;
  assign n13144 = ~n13142 & ~n13143 ;
  assign n13145 = x69 & n10905 ;
  assign n13146 = x67 & n11466 ;
  assign n13147 = x68 & n10900 ;
  assign n13148 = ~n13146 & ~n13147 ;
  assign n13149 = ~n13145 & n13148 ;
  assign n13150 = n398 & n10908 ;
  assign n13151 = n13149 & ~n13150 ;
  assign n13152 = x41 & ~n13151 ;
  assign n13153 = x41 & ~n13152 ;
  assign n13154 = ~n13151 & ~n13152 ;
  assign n13155 = ~n13153 & ~n13154 ;
  assign n13156 = n13144 & ~n13155 ;
  assign n13157 = n13144 & ~n13156 ;
  assign n13158 = ~n13155 & ~n13156 ;
  assign n13159 = ~n13157 & ~n13158 ;
  assign n13160 = ~n13128 & ~n13159 ;
  assign n13161 = n13128 & n13159 ;
  assign n13162 = ~n13160 & ~n13161 ;
  assign n13163 = ~n13127 & n13162 ;
  assign n13164 = ~n13127 & ~n13163 ;
  assign n13165 = n13162 & ~n13163 ;
  assign n13166 = ~n13164 & ~n13165 ;
  assign n13167 = ~n13116 & ~n13166 ;
  assign n13168 = ~n13116 & ~n13167 ;
  assign n13169 = ~n13166 & ~n13167 ;
  assign n13170 = ~n13168 & ~n13169 ;
  assign n13171 = x75 & n8006 ;
  assign n13172 = x73 & n8474 ;
  assign n13173 = x74 & n8001 ;
  assign n13174 = ~n13172 & ~n13173 ;
  assign n13175 = ~n13171 & n13174 ;
  assign n13176 = n1150 & n8009 ;
  assign n13177 = n13175 & ~n13176 ;
  assign n13178 = x35 & ~n13177 ;
  assign n13179 = x35 & ~n13178 ;
  assign n13180 = ~n13177 & ~n13178 ;
  assign n13181 = ~n13179 & ~n13180 ;
  assign n13182 = n13170 & n13181 ;
  assign n13183 = ~n13170 & ~n13181 ;
  assign n13184 = ~n13182 & ~n13183 ;
  assign n13185 = ~n12560 & n13184 ;
  assign n13186 = n12560 & ~n13184 ;
  assign n13187 = ~n13185 & ~n13186 ;
  assign n13188 = n13115 & ~n13187 ;
  assign n13189 = ~n13115 & n13187 ;
  assign n13190 = ~n13188 & ~n13189 ;
  assign n13191 = ~n13104 & n13190 ;
  assign n13192 = n13104 & ~n13190 ;
  assign n13193 = ~n13191 & ~n13192 ;
  assign n13194 = n13103 & ~n13193 ;
  assign n13195 = ~n13103 & n13193 ;
  assign n13196 = ~n13194 & ~n13195 ;
  assign n13197 = ~n13092 & n13196 ;
  assign n13198 = n13092 & ~n13196 ;
  assign n13199 = ~n13197 & ~n13198 ;
  assign n13200 = x84 & n4531 ;
  assign n13201 = x82 & n4847 ;
  assign n13202 = x83 & n4526 ;
  assign n13203 = ~n13201 & ~n13202 ;
  assign n13204 = ~n13200 & n13203 ;
  assign n13205 = n3114 & n4534 ;
  assign n13206 = n13204 & ~n13205 ;
  assign n13207 = x26 & ~n13206 ;
  assign n13208 = x26 & ~n13207 ;
  assign n13209 = ~n13206 & ~n13207 ;
  assign n13210 = ~n13208 & ~n13209 ;
  assign n13211 = n13199 & ~n13210 ;
  assign n13212 = n13199 & ~n13211 ;
  assign n13213 = ~n13210 & ~n13211 ;
  assign n13214 = ~n13212 & ~n13213 ;
  assign n13215 = ~n12611 & ~n12617 ;
  assign n13216 = n13214 & n13215 ;
  assign n13217 = ~n13214 & ~n13215 ;
  assign n13218 = ~n13216 & ~n13217 ;
  assign n13219 = x87 & n3589 ;
  assign n13220 = x85 & n3878 ;
  assign n13221 = x86 & n3584 ;
  assign n13222 = ~n13220 & ~n13221 ;
  assign n13223 = ~n13219 & n13222 ;
  assign n13224 = n3592 & n3991 ;
  assign n13225 = n13223 & ~n13224 ;
  assign n13226 = x23 & ~n13225 ;
  assign n13227 = x23 & ~n13226 ;
  assign n13228 = ~n13225 & ~n13226 ;
  assign n13229 = ~n13227 & ~n13228 ;
  assign n13230 = n13218 & ~n13229 ;
  assign n13231 = ~n13218 & n13229 ;
  assign n13232 = ~n13091 & ~n13231 ;
  assign n13233 = ~n13230 & n13232 ;
  assign n13234 = ~n13091 & ~n13233 ;
  assign n13235 = ~n13230 & ~n13233 ;
  assign n13236 = ~n13231 & n13235 ;
  assign n13237 = ~n13234 & ~n13236 ;
  assign n13238 = x90 & n2751 ;
  assign n13239 = x88 & n3020 ;
  assign n13240 = x89 & n2746 ;
  assign n13241 = ~n13239 & ~n13240 ;
  assign n13242 = ~n13238 & n13241 ;
  assign n13243 = n2754 & n4986 ;
  assign n13244 = n13242 & ~n13243 ;
  assign n13245 = x20 & ~n13244 ;
  assign n13246 = x20 & ~n13245 ;
  assign n13247 = ~n13244 & ~n13245 ;
  assign n13248 = ~n13246 & ~n13247 ;
  assign n13249 = n13237 & n13248 ;
  assign n13250 = ~n13237 & ~n13248 ;
  assign n13251 = ~n13249 & ~n13250 ;
  assign n13252 = ~n13090 & n13251 ;
  assign n13253 = n13090 & ~n13251 ;
  assign n13254 = ~n13252 & ~n13253 ;
  assign n13255 = n13089 & ~n13254 ;
  assign n13256 = ~n13089 & n13254 ;
  assign n13257 = ~n13255 & ~n13256 ;
  assign n13258 = ~n13078 & n13257 ;
  assign n13259 = n13078 & ~n13257 ;
  assign n13260 = ~n13258 & ~n13259 ;
  assign n13261 = n13077 & ~n13260 ;
  assign n13262 = ~n13077 & n13260 ;
  assign n13263 = ~n13261 & ~n13262 ;
  assign n13264 = ~n13066 & n13263 ;
  assign n13265 = n13066 & ~n13263 ;
  assign n13266 = ~n13264 & ~n13265 ;
  assign n13267 = x99 & n945 ;
  assign n13268 = x97 & n1099 ;
  assign n13269 = x98 & n940 ;
  assign n13270 = ~n13268 & ~n13269 ;
  assign n13271 = ~n13267 & n13270 ;
  assign n13272 = n948 & n8660 ;
  assign n13273 = n13271 & ~n13272 ;
  assign n13274 = x11 & ~n13273 ;
  assign n13275 = x11 & ~n13274 ;
  assign n13276 = ~n13273 & ~n13274 ;
  assign n13277 = ~n13275 & ~n13276 ;
  assign n13278 = n13266 & ~n13277 ;
  assign n13279 = n13266 & ~n13278 ;
  assign n13280 = ~n13277 & ~n13278 ;
  assign n13281 = ~n13279 & ~n13280 ;
  assign n13282 = ~n12693 & ~n12700 ;
  assign n13283 = n13281 & n13282 ;
  assign n13284 = ~n13281 & ~n13282 ;
  assign n13285 = ~n13283 & ~n13284 ;
  assign n13286 = x102 & n574 ;
  assign n13287 = x100 & n673 ;
  assign n13288 = x101 & n569 ;
  assign n13289 = ~n13287 & ~n13288 ;
  assign n13290 = ~n13286 & n13289 ;
  assign n13291 = n577 & n10092 ;
  assign n13292 = n13290 & ~n13291 ;
  assign n13293 = x8 & ~n13292 ;
  assign n13294 = x8 & ~n13293 ;
  assign n13295 = ~n13292 & ~n13293 ;
  assign n13296 = ~n13294 & ~n13295 ;
  assign n13297 = n13285 & ~n13296 ;
  assign n13298 = n13285 & ~n13297 ;
  assign n13299 = ~n13296 & ~n13297 ;
  assign n13300 = ~n13298 & ~n13299 ;
  assign n13301 = ~n12718 & ~n13300 ;
  assign n13302 = n12718 & n13300 ;
  assign n13303 = ~n13301 & ~n13302 ;
  assign n13304 = ~n13065 & n13303 ;
  assign n13305 = ~n13065 & ~n13304 ;
  assign n13306 = n13303 & ~n13304 ;
  assign n13307 = ~n13305 & ~n13306 ;
  assign n13308 = ~n13054 & ~n13307 ;
  assign n13309 = ~n13054 & ~n13308 ;
  assign n13310 = ~n13307 & ~n13308 ;
  assign n13311 = ~n13309 & ~n13310 ;
  assign n13312 = x108 & n146 ;
  assign n13313 = x106 & n182 ;
  assign n13314 = x107 & n141 ;
  assign n13315 = ~n13313 & ~n13314 ;
  assign n13316 = ~n13312 & n13315 ;
  assign n13317 = ~n12745 & ~n12747 ;
  assign n13318 = ~x107 & ~x108 ;
  assign n13319 = x107 & x108 ;
  assign n13320 = ~n13318 & ~n13319 ;
  assign n13321 = ~n13317 & n13320 ;
  assign n13322 = n13317 & ~n13320 ;
  assign n13323 = ~n13321 & ~n13322 ;
  assign n13324 = n149 & n13323 ;
  assign n13325 = n13316 & ~n13324 ;
  assign n13326 = x2 & ~n13325 ;
  assign n13327 = x2 & ~n13326 ;
  assign n13328 = ~n13325 & ~n13326 ;
  assign n13329 = ~n13327 & ~n13328 ;
  assign n13330 = ~n13311 & n13329 ;
  assign n13331 = n13311 & ~n13329 ;
  assign n13332 = ~n13330 & ~n13331 ;
  assign n13333 = ~n13053 & ~n13332 ;
  assign n13334 = n13053 & n13332 ;
  assign n13335 = ~n13333 & ~n13334 ;
  assign n13615 = n13335 & x172 ;
  assign n13336 = ~n13041 & ~n13046 ;
  assign n13337 = ~n13021 & ~n13023 ;
  assign n13338 = ~x105 & n293 ;
  assign n13339 = ~x103 & n373 ;
  assign n13340 = ~x104 & n288 ;
  assign n13341 = ~n13339 & ~n13340 ;
  assign n13342 = ~n13338 & n13341 ;
  assign n13343 = n296 & n11907 ;
  assign n13344 = n13342 & ~n13343 ;
  assign n13345 = ~x5 & ~n13344 ;
  assign n13346 = ~x5 & ~n13345 ;
  assign n13347 = ~n13344 & ~n13345 ;
  assign n13348 = ~n13346 & ~n13347 ;
  assign n13349 = ~n12965 & ~n12967 ;
  assign n13350 = ~x96 & n1434 ;
  assign n13351 = ~x94 & n1646 ;
  assign n13352 = ~x95 & n1429 ;
  assign n13353 = ~n13351 & ~n13352 ;
  assign n13354 = ~n13350 & n13353 ;
  assign n13355 = n1437 & n7531 ;
  assign n13356 = n13354 & ~n13355 ;
  assign n13357 = ~x14 & ~n13356 ;
  assign n13358 = ~x14 & ~n13357 ;
  assign n13359 = ~n13356 & ~n13357 ;
  assign n13360 = ~n13358 & ~n13359 ;
  assign n13361 = ~n12945 & ~n12949 ;
  assign n13362 = ~x93 & n2093 ;
  assign n13363 = ~x91 & n2275 ;
  assign n13364 = ~x92 & n2088 ;
  assign n13365 = ~n13363 & ~n13364 ;
  assign n13366 = ~n13362 & n13365 ;
  assign n13367 = n2096 & n6285 ;
  assign n13368 = n13366 & ~n13367 ;
  assign n13369 = ~x17 & ~n13368 ;
  assign n13370 = ~x17 & ~n13369 ;
  assign n13371 = ~n13368 & ~n13369 ;
  assign n13372 = ~n13370 & ~n13371 ;
  assign n13373 = ~n12937 & ~n12942 ;
  assign n13374 = ~n12918 & ~n12924 ;
  assign n13375 = ~n12879 & ~n12886 ;
  assign n13376 = ~x81 & n5560 ;
  assign n13377 = ~x79 & n5943 ;
  assign n13378 = ~x80 & n5555 ;
  assign n13379 = ~n13377 & ~n13378 ;
  assign n13380 = ~n13376 & n13379 ;
  assign n13381 = n2460 & n5563 ;
  assign n13382 = n13380 & ~n13381 ;
  assign n13383 = ~x29 & ~n13382 ;
  assign n13384 = ~x29 & ~n13383 ;
  assign n13385 = ~n13382 & ~n13383 ;
  assign n13386 = ~n13384 & ~n13385 ;
  assign n13387 = ~n12863 & ~n12865 ;
  assign n13388 = ~x78 & n6725 ;
  assign n13389 = ~x76 & n7129 ;
  assign n13390 = ~x77 & n6720 ;
  assign n13391 = ~n13389 & ~n13390 ;
  assign n13392 = ~n13388 & n13391 ;
  assign n13393 = n1718 & n6728 ;
  assign n13394 = n13392 & ~n13393 ;
  assign n13395 = ~x32 & ~n13394 ;
  assign n13396 = ~x32 & ~n13395 ;
  assign n13397 = ~n13394 & ~n13395 ;
  assign n13398 = ~n13396 & ~n13397 ;
  assign n13399 = ~n12824 & ~n12830 ;
  assign n13400 = ~x72 & n9433 ;
  assign n13401 = ~x70 & n9915 ;
  assign n13402 = ~x71 & n9428 ;
  assign n13403 = ~n13401 & ~n13402 ;
  assign n13404 = ~n13400 & n13403 ;
  assign n13405 = n773 & n9436 ;
  assign n13406 = n13404 & ~n13405 ;
  assign n13407 = ~x38 & ~n13406 ;
  assign n13408 = ~x38 & ~n13407 ;
  assign n13409 = ~n13406 & ~n13407 ;
  assign n13410 = ~n13408 & ~n13409 ;
  assign n13411 = ~n12808 & ~n12810 ;
  assign n13412 = ~x66 & n12506 ;
  assign n13413 = ~x64 & n13131 ;
  assign n13414 = ~x65 & n12501 ;
  assign n13415 = ~n13413 & ~n13414 ;
  assign n13416 = ~n13412 & n13415 ;
  assign n13417 = n214 & n12509 ;
  assign n13418 = n13416 & ~n13417 ;
  assign n13419 = ~x44 & ~n13418 ;
  assign n13420 = ~x44 & ~n13419 ;
  assign n13421 = ~n13418 & ~n13419 ;
  assign n13422 = ~n13420 & ~n13421 ;
  assign n13423 = ~n12804 & n13422 ;
  assign n13424 = n12804 & ~n13422 ;
  assign n13425 = ~n13423 & ~n13424 ;
  assign n13426 = ~x69 & n10905 ;
  assign n13427 = ~x67 & n11466 ;
  assign n13428 = ~x68 & n10900 ;
  assign n13429 = ~n13427 & ~n13428 ;
  assign n13430 = ~n13426 & n13429 ;
  assign n13431 = n435 & n10908 ;
  assign n13432 = n13430 & ~n13431 ;
  assign n13433 = ~x41 & ~n13432 ;
  assign n13434 = ~x41 & ~n13433 ;
  assign n13435 = ~n13432 & ~n13433 ;
  assign n13436 = ~n13434 & ~n13435 ;
  assign n13437 = n13425 & ~n13436 ;
  assign n13438 = n13425 & ~n13437 ;
  assign n13439 = ~n13436 & ~n13437 ;
  assign n13440 = ~n13438 & ~n13439 ;
  assign n13441 = ~n13411 & ~n13440 ;
  assign n13442 = n13411 & n13440 ;
  assign n13443 = ~n13441 & ~n13442 ;
  assign n13444 = ~n13410 & n13443 ;
  assign n13445 = ~n13410 & ~n13444 ;
  assign n13446 = n13443 & ~n13444 ;
  assign n13447 = ~n13445 & ~n13446 ;
  assign n13448 = ~n13399 & ~n13447 ;
  assign n13449 = ~n13399 & ~n13448 ;
  assign n13450 = ~n13447 & ~n13448 ;
  assign n13451 = ~n13449 & ~n13450 ;
  assign n13452 = ~x75 & n8006 ;
  assign n13453 = ~x73 & n8474 ;
  assign n13454 = ~x74 & n8001 ;
  assign n13455 = ~n13453 & ~n13454 ;
  assign n13456 = ~n13452 & n13455 ;
  assign n13457 = n1225 & n8009 ;
  assign n13458 = n13456 & ~n13457 ;
  assign n13459 = ~x35 & ~n13458 ;
  assign n13460 = ~x35 & ~n13459 ;
  assign n13461 = ~n13458 & ~n13459 ;
  assign n13462 = ~n13460 & ~n13461 ;
  assign n13463 = n13451 & n13462 ;
  assign n13464 = ~n13451 & ~n13462 ;
  assign n13465 = ~n13463 & ~n13464 ;
  assign n13466 = ~n12848 & n13465 ;
  assign n13467 = n12848 & ~n13465 ;
  assign n13468 = ~n13466 & ~n13467 ;
  assign n13469 = n13398 & ~n13468 ;
  assign n13470 = ~n13398 & n13468 ;
  assign n13471 = ~n13469 & ~n13470 ;
  assign n13472 = ~n13387 & n13471 ;
  assign n13473 = n13387 & ~n13471 ;
  assign n13474 = ~n13472 & ~n13473 ;
  assign n13475 = n13386 & ~n13474 ;
  assign n13476 = ~n13386 & n13474 ;
  assign n13477 = ~n13475 & ~n13476 ;
  assign n13478 = ~n13375 & n13477 ;
  assign n13479 = n13375 & ~n13477 ;
  assign n13480 = ~n13478 & ~n13479 ;
  assign n13481 = ~x84 & n4531 ;
  assign n13482 = ~x82 & n4847 ;
  assign n13483 = ~x83 & n4526 ;
  assign n13484 = ~n13482 & ~n13483 ;
  assign n13485 = ~n13481 & n13484 ;
  assign n13486 = n3247 & n4534 ;
  assign n13487 = n13485 & ~n13486 ;
  assign n13488 = ~x26 & ~n13487 ;
  assign n13489 = ~x26 & ~n13488 ;
  assign n13490 = ~n13487 & ~n13488 ;
  assign n13491 = ~n13489 & ~n13490 ;
  assign n13492 = n13480 & ~n13491 ;
  assign n13493 = n13480 & ~n13492 ;
  assign n13494 = ~n13491 & ~n13492 ;
  assign n13495 = ~n13493 & ~n13494 ;
  assign n13496 = ~n12899 & ~n12905 ;
  assign n13497 = n13495 & n13496 ;
  assign n13498 = ~n13495 & ~n13496 ;
  assign n13499 = ~n13497 & ~n13498 ;
  assign n13500 = ~x87 & n3589 ;
  assign n13501 = ~x85 & n3878 ;
  assign n13502 = ~x86 & n3584 ;
  assign n13503 = ~n13501 & ~n13502 ;
  assign n13504 = ~n13500 & n13503 ;
  assign n13505 = n3592 & n4143 ;
  assign n13506 = n13504 & ~n13505 ;
  assign n13507 = ~x23 & ~n13506 ;
  assign n13508 = ~x23 & ~n13507 ;
  assign n13509 = ~n13506 & ~n13507 ;
  assign n13510 = ~n13508 & ~n13509 ;
  assign n13511 = n13499 & ~n13510 ;
  assign n13512 = ~n13499 & n13510 ;
  assign n13513 = ~n13374 & ~n13512 ;
  assign n13514 = ~n13511 & n13513 ;
  assign n13515 = ~n13374 & ~n13514 ;
  assign n13516 = ~n13511 & ~n13514 ;
  assign n13517 = ~n13512 & n13516 ;
  assign n13518 = ~n13515 & ~n13517 ;
  assign n13519 = ~x90 & n2751 ;
  assign n13520 = ~x88 & n3020 ;
  assign n13521 = ~x89 & n2746 ;
  assign n13522 = ~n13520 & ~n13521 ;
  assign n13523 = ~n13519 & n13522 ;
  assign n13524 = n2754 & n5155 ;
  assign n13525 = n13523 & ~n13524 ;
  assign n13526 = ~x20 & ~n13525 ;
  assign n13527 = ~x20 & ~n13526 ;
  assign n13528 = ~n13525 & ~n13526 ;
  assign n13529 = ~n13527 & ~n13528 ;
  assign n13530 = n13518 & n13529 ;
  assign n13531 = ~n13518 & ~n13529 ;
  assign n13532 = ~n13530 & ~n13531 ;
  assign n13533 = ~n13373 & n13532 ;
  assign n13534 = n13373 & ~n13532 ;
  assign n13535 = ~n13533 & ~n13534 ;
  assign n13536 = n13372 & ~n13535 ;
  assign n13537 = ~n13372 & n13535 ;
  assign n13538 = ~n13536 & ~n13537 ;
  assign n13539 = ~n13361 & n13538 ;
  assign n13540 = n13361 & ~n13538 ;
  assign n13541 = ~n13539 & ~n13540 ;
  assign n13542 = n13360 & ~n13541 ;
  assign n13543 = ~n13360 & n13541 ;
  assign n13544 = ~n13542 & ~n13543 ;
  assign n13545 = ~n13349 & n13544 ;
  assign n13546 = n13349 & ~n13544 ;
  assign n13547 = ~n13545 & ~n13546 ;
  assign n13548 = ~x99 & n945 ;
  assign n13549 = ~x97 & n1099 ;
  assign n13550 = ~x98 & n940 ;
  assign n13551 = ~n13549 & ~n13550 ;
  assign n13552 = ~n13548 & n13551 ;
  assign n13553 = n948 & n8885 ;
  assign n13554 = n13552 & ~n13553 ;
  assign n13555 = ~x11 & ~n13554 ;
  assign n13556 = ~x11 & ~n13555 ;
  assign n13557 = ~n13554 & ~n13555 ;
  assign n13558 = ~n13556 & ~n13557 ;
  assign n13559 = n13547 & ~n13558 ;
  assign n13560 = n13547 & ~n13559 ;
  assign n13561 = ~n13558 & ~n13559 ;
  assign n13562 = ~n13560 & ~n13561 ;
  assign n13563 = ~n12981 & ~n12988 ;
  assign n13564 = n13562 & n13563 ;
  assign n13565 = ~n13562 & ~n13563 ;
  assign n13566 = ~n13564 & ~n13565 ;
  assign n13567 = ~x102 & n574 ;
  assign n13568 = ~x100 & n673 ;
  assign n13569 = ~x101 & n569 ;
  assign n13570 = ~n13568 & ~n13569 ;
  assign n13571 = ~n13567 & n13570 ;
  assign n13572 = n577 & n10333 ;
  assign n13573 = n13571 & ~n13572 ;
  assign n13574 = ~x8 & ~n13573 ;
  assign n13575 = ~x8 & ~n13574 ;
  assign n13576 = ~n13573 & ~n13574 ;
  assign n13577 = ~n13575 & ~n13576 ;
  assign n13578 = n13566 & ~n13577 ;
  assign n13579 = n13566 & ~n13578 ;
  assign n13580 = ~n13577 & ~n13578 ;
  assign n13581 = ~n13579 & ~n13580 ;
  assign n13582 = ~n13006 & ~n13581 ;
  assign n13583 = n13006 & n13581 ;
  assign n13584 = ~n13582 & ~n13583 ;
  assign n13585 = ~n13348 & n13584 ;
  assign n13586 = ~n13348 & ~n13585 ;
  assign n13587 = n13584 & ~n13585 ;
  assign n13588 = ~n13586 & ~n13587 ;
  assign n13589 = ~n13337 & ~n13588 ;
  assign n13590 = ~n13337 & ~n13589 ;
  assign n13591 = ~n13588 & ~n13589 ;
  assign n13592 = ~n13590 & ~n13591 ;
  assign n13593 = ~x108 & n164 ;
  assign n13594 = ~x106 & n205 ;
  assign n13595 = ~x107 & n162 ;
  assign n13596 = ~n13594 & ~n13595 ;
  assign n13597 = ~n13593 & n13596 ;
  assign n13598 = ~n12744 & ~n13032 ;
  assign n13599 = n13320 & ~n13598 ;
  assign n13600 = ~n13320 & n13598 ;
  assign n13601 = ~n13599 & ~n13600 ;
  assign n13602 = n167 & n13601 ;
  assign n13603 = n13597 & ~n13602 ;
  assign n13604 = ~x2 & ~n13603 ;
  assign n13605 = ~x2 & ~n13604 ;
  assign n13606 = ~n13603 & ~n13604 ;
  assign n13607 = ~n13605 & ~n13606 ;
  assign n13608 = ~n13592 & n13607 ;
  assign n13609 = n13592 & ~n13607 ;
  assign n13610 = ~n13608 & ~n13609 ;
  assign n13611 = ~n13336 & ~n13610 ;
  assign n13612 = n13336 & n13610 ;
  assign n13613 = ~n13611 & ~n13612 ;
  assign n13616 = ~n13613 & ~x172 ;
  assign n13617 = ~n13615 & ~n13616 ;
  assign n13618 = ~n13311 & ~n13329 ;
  assign n13619 = ~n13333 & ~n13618 ;
  assign n13620 = ~n13278 & ~n13284 ;
  assign n13621 = ~n13262 & ~n13264 ;
  assign n13622 = ~n13256 & ~n13258 ;
  assign n13623 = ~n13250 & ~n13252 ;
  assign n13624 = ~n13195 & ~n13197 ;
  assign n13625 = ~n13189 & ~n13191 ;
  assign n13626 = ~n13183 & ~n13185 ;
  assign n13627 = x76 & n8006 ;
  assign n13628 = x74 & n8474 ;
  assign n13629 = x75 & n8001 ;
  assign n13630 = ~n13628 & ~n13629 ;
  assign n13631 = ~n13627 & n13630 ;
  assign n13632 = n1311 & n8009 ;
  assign n13633 = n13631 & ~n13632 ;
  assign n13634 = x35 & ~n13633 ;
  assign n13635 = x35 & ~n13634 ;
  assign n13636 = ~n13633 & ~n13634 ;
  assign n13637 = ~n13635 & ~n13636 ;
  assign n13638 = ~n13163 & ~n13167 ;
  assign n13639 = x44 & ~x45 ;
  assign n13640 = ~x44 & x45 ;
  assign n13641 = ~n13639 & ~n13640 ;
  assign n13642 = x64 & ~n13641 ;
  assign n13643 = ~n13143 & n13642 ;
  assign n13644 = n13143 & ~n13642 ;
  assign n13645 = ~n13643 & ~n13644 ;
  assign n13646 = x67 & n12506 ;
  assign n13647 = x65 & n13131 ;
  assign n13648 = x66 & n12501 ;
  assign n13649 = ~n13647 & ~n13648 ;
  assign n13650 = ~n13646 & n13649 ;
  assign n13651 = n240 & n12509 ;
  assign n13652 = n13650 & ~n13651 ;
  assign n13653 = x44 & ~n13652 ;
  assign n13654 = x44 & ~n13653 ;
  assign n13655 = ~n13652 & ~n13653 ;
  assign n13656 = ~n13654 & ~n13655 ;
  assign n13657 = ~n13645 & ~n13656 ;
  assign n13658 = n13645 & n13656 ;
  assign n13659 = ~n13657 & ~n13658 ;
  assign n13660 = x70 & n10905 ;
  assign n13661 = x68 & n11466 ;
  assign n13662 = x69 & n10900 ;
  assign n13663 = ~n13661 & ~n13662 ;
  assign n13664 = ~n13660 & n13663 ;
  assign n13665 = n488 & n10908 ;
  assign n13666 = n13664 & ~n13665 ;
  assign n13667 = x41 & ~n13666 ;
  assign n13668 = x41 & ~n13667 ;
  assign n13669 = ~n13666 & ~n13667 ;
  assign n13670 = ~n13668 & ~n13669 ;
  assign n13671 = n13659 & ~n13670 ;
  assign n13672 = n13659 & ~n13671 ;
  assign n13673 = ~n13670 & ~n13671 ;
  assign n13674 = ~n13672 & ~n13673 ;
  assign n13675 = ~n13156 & ~n13160 ;
  assign n13676 = n13674 & n13675 ;
  assign n13677 = ~n13674 & ~n13675 ;
  assign n13678 = ~n13676 & ~n13677 ;
  assign n13679 = x73 & n9433 ;
  assign n13680 = x71 & n9915 ;
  assign n13681 = x72 & n9428 ;
  assign n13682 = ~n13680 & ~n13681 ;
  assign n13683 = ~n13679 & n13682 ;
  assign n13684 = n843 & n9436 ;
  assign n13685 = n13683 & ~n13684 ;
  assign n13686 = x38 & ~n13685 ;
  assign n13687 = x38 & ~n13686 ;
  assign n13688 = ~n13685 & ~n13686 ;
  assign n13689 = ~n13687 & ~n13688 ;
  assign n13690 = ~n13678 & n13689 ;
  assign n13691 = n13678 & ~n13689 ;
  assign n13692 = ~n13690 & ~n13691 ;
  assign n13693 = ~n13638 & n13692 ;
  assign n13694 = n13638 & ~n13692 ;
  assign n13695 = ~n13693 & ~n13694 ;
  assign n13696 = ~n13637 & n13695 ;
  assign n13697 = ~n13637 & ~n13696 ;
  assign n13698 = n13695 & ~n13696 ;
  assign n13699 = ~n13697 & ~n13698 ;
  assign n13700 = ~n13626 & ~n13699 ;
  assign n13701 = ~n13626 & ~n13700 ;
  assign n13702 = ~n13699 & ~n13700 ;
  assign n13703 = ~n13701 & ~n13702 ;
  assign n13704 = x79 & n6725 ;
  assign n13705 = x77 & n7129 ;
  assign n13706 = x78 & n6720 ;
  assign n13707 = ~n13705 & ~n13706 ;
  assign n13708 = ~n13704 & n13707 ;
  assign n13709 = n1817 & n6728 ;
  assign n13710 = n13708 & ~n13709 ;
  assign n13711 = x32 & ~n13710 ;
  assign n13712 = x32 & ~n13711 ;
  assign n13713 = ~n13710 & ~n13711 ;
  assign n13714 = ~n13712 & ~n13713 ;
  assign n13715 = ~n13703 & ~n13714 ;
  assign n13716 = ~n13703 & ~n13715 ;
  assign n13717 = ~n13714 & ~n13715 ;
  assign n13718 = ~n13716 & ~n13717 ;
  assign n13719 = ~n13625 & n13718 ;
  assign n13720 = n13625 & ~n13718 ;
  assign n13721 = ~n13719 & ~n13720 ;
  assign n13722 = x82 & n5560 ;
  assign n13723 = x80 & n5943 ;
  assign n13724 = x81 & n5555 ;
  assign n13725 = ~n13723 & ~n13724 ;
  assign n13726 = ~n13722 & n13725 ;
  assign n13727 = n2584 & n5563 ;
  assign n13728 = n13726 & ~n13727 ;
  assign n13729 = x29 & ~n13728 ;
  assign n13730 = x29 & ~n13729 ;
  assign n13731 = ~n13728 & ~n13729 ;
  assign n13732 = ~n13730 & ~n13731 ;
  assign n13733 = ~n13721 & ~n13732 ;
  assign n13734 = n13721 & n13732 ;
  assign n13735 = ~n13733 & ~n13734 ;
  assign n13736 = ~n13624 & n13735 ;
  assign n13737 = n13624 & ~n13735 ;
  assign n13738 = ~n13736 & ~n13737 ;
  assign n13739 = x85 & n4531 ;
  assign n13740 = x83 & n4847 ;
  assign n13741 = x84 & n4526 ;
  assign n13742 = ~n13740 & ~n13741 ;
  assign n13743 = ~n13739 & n13742 ;
  assign n13744 = n3389 & n4534 ;
  assign n13745 = n13743 & ~n13744 ;
  assign n13746 = x26 & ~n13745 ;
  assign n13747 = x26 & ~n13746 ;
  assign n13748 = ~n13745 & ~n13746 ;
  assign n13749 = ~n13747 & ~n13748 ;
  assign n13750 = n13738 & ~n13749 ;
  assign n13751 = n13738 & ~n13750 ;
  assign n13752 = ~n13749 & ~n13750 ;
  assign n13753 = ~n13751 & ~n13752 ;
  assign n13754 = ~n13211 & ~n13217 ;
  assign n13755 = n13753 & n13754 ;
  assign n13756 = ~n13753 & ~n13754 ;
  assign n13757 = ~n13755 & ~n13756 ;
  assign n13758 = x88 & n3589 ;
  assign n13759 = x86 & n3878 ;
  assign n13760 = x87 & n3584 ;
  assign n13761 = ~n13759 & ~n13760 ;
  assign n13762 = ~n13758 & n13761 ;
  assign n13763 = n3592 & n4305 ;
  assign n13764 = n13762 & ~n13763 ;
  assign n13765 = x23 & ~n13764 ;
  assign n13766 = x23 & ~n13765 ;
  assign n13767 = ~n13764 & ~n13765 ;
  assign n13768 = ~n13766 & ~n13767 ;
  assign n13769 = ~n13757 & n13768 ;
  assign n13770 = n13757 & ~n13768 ;
  assign n13771 = ~n13769 & ~n13770 ;
  assign n13772 = ~n13235 & n13771 ;
  assign n13773 = n13235 & ~n13771 ;
  assign n13774 = ~n13772 & ~n13773 ;
  assign n13775 = x91 & n2751 ;
  assign n13776 = x89 & n3020 ;
  assign n13777 = x90 & n2746 ;
  assign n13778 = ~n13776 & ~n13777 ;
  assign n13779 = ~n13775 & n13778 ;
  assign n13780 = n2754 & n5336 ;
  assign n13781 = n13779 & ~n13780 ;
  assign n13782 = x20 & ~n13781 ;
  assign n13783 = x20 & ~n13782 ;
  assign n13784 = ~n13781 & ~n13782 ;
  assign n13785 = ~n13783 & ~n13784 ;
  assign n13786 = n13774 & ~n13785 ;
  assign n13787 = n13774 & ~n13786 ;
  assign n13788 = ~n13785 & ~n13786 ;
  assign n13789 = ~n13787 & ~n13788 ;
  assign n13790 = ~n13623 & n13789 ;
  assign n13791 = n13623 & ~n13789 ;
  assign n13792 = ~n13790 & ~n13791 ;
  assign n13793 = x94 & n2093 ;
  assign n13794 = x92 & n2275 ;
  assign n13795 = x93 & n2088 ;
  assign n13796 = ~n13794 & ~n13795 ;
  assign n13797 = ~n13793 & n13796 ;
  assign n13798 = n2096 & n6483 ;
  assign n13799 = n13797 & ~n13798 ;
  assign n13800 = x17 & ~n13799 ;
  assign n13801 = x17 & ~n13800 ;
  assign n13802 = ~n13799 & ~n13800 ;
  assign n13803 = ~n13801 & ~n13802 ;
  assign n13804 = ~n13792 & ~n13803 ;
  assign n13805 = n13792 & n13803 ;
  assign n13806 = ~n13804 & ~n13805 ;
  assign n13807 = ~n13622 & n13806 ;
  assign n13808 = n13622 & ~n13806 ;
  assign n13809 = ~n13807 & ~n13808 ;
  assign n13810 = x97 & n1434 ;
  assign n13811 = x95 & n1646 ;
  assign n13812 = x96 & n1429 ;
  assign n13813 = ~n13811 & ~n13812 ;
  assign n13814 = ~n13810 & n13813 ;
  assign n13815 = n1437 & n7745 ;
  assign n13816 = n13814 & ~n13815 ;
  assign n13817 = x14 & ~n13816 ;
  assign n13818 = x14 & ~n13817 ;
  assign n13819 = ~n13816 & ~n13817 ;
  assign n13820 = ~n13818 & ~n13819 ;
  assign n13821 = n13809 & ~n13820 ;
  assign n13822 = n13809 & ~n13821 ;
  assign n13823 = ~n13820 & ~n13821 ;
  assign n13824 = ~n13822 & ~n13823 ;
  assign n13825 = ~n13621 & n13824 ;
  assign n13826 = n13621 & ~n13824 ;
  assign n13827 = ~n13825 & ~n13826 ;
  assign n13828 = x100 & n945 ;
  assign n13829 = x98 & n1099 ;
  assign n13830 = x99 & n940 ;
  assign n13831 = ~n13829 & ~n13830 ;
  assign n13832 = ~n13828 & n13831 ;
  assign n13833 = n948 & n9115 ;
  assign n13834 = n13832 & ~n13833 ;
  assign n13835 = x11 & ~n13834 ;
  assign n13836 = x11 & ~n13835 ;
  assign n13837 = ~n13834 & ~n13835 ;
  assign n13838 = ~n13836 & ~n13837 ;
  assign n13839 = ~n13827 & ~n13838 ;
  assign n13840 = n13827 & n13838 ;
  assign n13841 = ~n13839 & ~n13840 ;
  assign n13842 = n13620 & ~n13841 ;
  assign n13843 = ~n13620 & n13841 ;
  assign n13844 = ~n13842 & ~n13843 ;
  assign n13845 = x103 & n574 ;
  assign n13846 = x101 & n673 ;
  assign n13847 = x102 & n569 ;
  assign n13848 = ~n13846 & ~n13847 ;
  assign n13849 = ~n13845 & n13848 ;
  assign n13850 = n577 & n10588 ;
  assign n13851 = n13849 & ~n13850 ;
  assign n13852 = x8 & ~n13851 ;
  assign n13853 = x8 & ~n13852 ;
  assign n13854 = ~n13851 & ~n13852 ;
  assign n13855 = ~n13853 & ~n13854 ;
  assign n13856 = n13844 & ~n13855 ;
  assign n13857 = n13844 & ~n13856 ;
  assign n13858 = ~n13855 & ~n13856 ;
  assign n13859 = ~n13857 & ~n13858 ;
  assign n13860 = ~n13297 & ~n13301 ;
  assign n13861 = n13859 & n13860 ;
  assign n13862 = ~n13859 & ~n13860 ;
  assign n13863 = ~n13861 & ~n13862 ;
  assign n13864 = x106 & n293 ;
  assign n13865 = x104 & n373 ;
  assign n13866 = x105 & n288 ;
  assign n13867 = ~n13865 & ~n13866 ;
  assign n13868 = ~n13864 & n13867 ;
  assign n13869 = n296 & n12181 ;
  assign n13870 = n13868 & ~n13869 ;
  assign n13871 = x5 & ~n13870 ;
  assign n13872 = x5 & ~n13871 ;
  assign n13873 = ~n13870 & ~n13871 ;
  assign n13874 = ~n13872 & ~n13873 ;
  assign n13875 = n13863 & ~n13874 ;
  assign n13876 = n13863 & ~n13875 ;
  assign n13877 = ~n13874 & ~n13875 ;
  assign n13878 = ~n13876 & ~n13877 ;
  assign n13879 = ~n13304 & ~n13308 ;
  assign n13880 = n13878 & n13879 ;
  assign n13881 = ~n13878 & ~n13879 ;
  assign n13882 = ~n13880 & ~n13881 ;
  assign n13883 = x109 & n146 ;
  assign n13884 = x107 & n182 ;
  assign n13885 = x108 & n141 ;
  assign n13886 = ~n13884 & ~n13885 ;
  assign n13887 = ~n13883 & n13886 ;
  assign n13888 = ~n13319 & ~n13321 ;
  assign n13889 = ~x108 & ~x109 ;
  assign n13890 = x108 & x109 ;
  assign n13891 = ~n13889 & ~n13890 ;
  assign n13892 = ~n13888 & n13891 ;
  assign n13893 = n13888 & ~n13891 ;
  assign n13894 = ~n13892 & ~n13893 ;
  assign n13895 = n149 & n13894 ;
  assign n13896 = n13887 & ~n13895 ;
  assign n13897 = x2 & ~n13896 ;
  assign n13898 = x2 & ~n13897 ;
  assign n13899 = ~n13896 & ~n13897 ;
  assign n13900 = ~n13898 & ~n13899 ;
  assign n13901 = ~n13882 & n13900 ;
  assign n13902 = n13882 & ~n13900 ;
  assign n13903 = ~n13901 & ~n13902 ;
  assign n13904 = ~n13619 & n13903 ;
  assign n13905 = n13619 & ~n13903 ;
  assign n13906 = ~n13904 & ~n13905 ;
  assign n14191 = n13906 & x173 ;
  assign n13907 = ~n13592 & ~n13607 ;
  assign n13908 = ~n13611 & ~n13907 ;
  assign n13909 = ~n13559 & ~n13565 ;
  assign n13910 = ~n13543 & ~n13545 ;
  assign n13911 = ~n13537 & ~n13539 ;
  assign n13912 = ~n13531 & ~n13533 ;
  assign n13913 = ~n13476 & ~n13478 ;
  assign n13914 = ~n13470 & ~n13472 ;
  assign n13915 = ~n13464 & ~n13466 ;
  assign n13916 = ~x76 & n8006 ;
  assign n13917 = ~x74 & n8474 ;
  assign n13918 = ~x75 & n8001 ;
  assign n13919 = ~n13917 & ~n13918 ;
  assign n13920 = ~n13916 & n13919 ;
  assign n13921 = n1390 & n8009 ;
  assign n13922 = n13920 & ~n13921 ;
  assign n13923 = ~x35 & ~n13922 ;
  assign n13924 = ~x35 & ~n13923 ;
  assign n13925 = ~n13922 & ~n13923 ;
  assign n13926 = ~n13924 & ~n13925 ;
  assign n13927 = ~n13444 & ~n13448 ;
  assign n13928 = ~x64 & ~n13641 ;
  assign n13929 = ~n13424 & n13928 ;
  assign n13930 = n13424 & ~n13928 ;
  assign n13931 = ~n13929 & ~n13930 ;
  assign n13932 = ~x67 & n12506 ;
  assign n13933 = ~x65 & n13131 ;
  assign n13934 = ~x66 & n12501 ;
  assign n13935 = ~n13933 & ~n13934 ;
  assign n13936 = ~n13932 & n13935 ;
  assign n13937 = n266 & n12509 ;
  assign n13938 = n13936 & ~n13937 ;
  assign n13939 = ~x44 & ~n13938 ;
  assign n13940 = ~x44 & ~n13939 ;
  assign n13941 = ~n13938 & ~n13939 ;
  assign n13942 = ~n13940 & ~n13941 ;
  assign n13943 = ~n13931 & ~n13942 ;
  assign n13944 = n13931 & n13942 ;
  assign n13945 = ~n13943 & ~n13944 ;
  assign n13946 = ~x70 & n10905 ;
  assign n13947 = ~x68 & n11466 ;
  assign n13948 = ~x69 & n10900 ;
  assign n13949 = ~n13947 & ~n13948 ;
  assign n13950 = ~n13946 & n13949 ;
  assign n13951 = n529 & n10908 ;
  assign n13952 = n13950 & ~n13951 ;
  assign n13953 = ~x41 & ~n13952 ;
  assign n13954 = ~x41 & ~n13953 ;
  assign n13955 = ~n13952 & ~n13953 ;
  assign n13956 = ~n13954 & ~n13955 ;
  assign n13957 = n13945 & ~n13956 ;
  assign n13958 = n13945 & ~n13957 ;
  assign n13959 = ~n13956 & ~n13957 ;
  assign n13960 = ~n13958 & ~n13959 ;
  assign n13961 = ~n13437 & ~n13441 ;
  assign n13962 = n13960 & n13961 ;
  assign n13963 = ~n13960 & ~n13961 ;
  assign n13964 = ~n13962 & ~n13963 ;
  assign n13965 = ~x73 & n9433 ;
  assign n13966 = ~x71 & n9915 ;
  assign n13967 = ~x72 & n9428 ;
  assign n13968 = ~n13966 & ~n13967 ;
  assign n13969 = ~n13965 & n13968 ;
  assign n13970 = n903 & n9436 ;
  assign n13971 = n13969 & ~n13970 ;
  assign n13972 = ~x38 & ~n13971 ;
  assign n13973 = ~x38 & ~n13972 ;
  assign n13974 = ~n13971 & ~n13972 ;
  assign n13975 = ~n13973 & ~n13974 ;
  assign n13976 = ~n13964 & n13975 ;
  assign n13977 = n13964 & ~n13975 ;
  assign n13978 = ~n13976 & ~n13977 ;
  assign n13979 = ~n13927 & n13978 ;
  assign n13980 = n13927 & ~n13978 ;
  assign n13981 = ~n13979 & ~n13980 ;
  assign n13982 = ~n13926 & n13981 ;
  assign n13983 = ~n13926 & ~n13982 ;
  assign n13984 = n13981 & ~n13982 ;
  assign n13985 = ~n13983 & ~n13984 ;
  assign n13986 = ~n13915 & ~n13985 ;
  assign n13987 = ~n13915 & ~n13986 ;
  assign n13988 = ~n13985 & ~n13986 ;
  assign n13989 = ~n13987 & ~n13988 ;
  assign n13990 = ~x79 & n6725 ;
  assign n13991 = ~x77 & n7129 ;
  assign n13992 = ~x78 & n6720 ;
  assign n13993 = ~n13991 & ~n13992 ;
  assign n13994 = ~n13990 & n13993 ;
  assign n13995 = n1921 & n6728 ;
  assign n13996 = n13994 & ~n13995 ;
  assign n13997 = ~x32 & ~n13996 ;
  assign n13998 = ~x32 & ~n13997 ;
  assign n13999 = ~n13996 & ~n13997 ;
  assign n14000 = ~n13998 & ~n13999 ;
  assign n14001 = ~n13989 & ~n14000 ;
  assign n14002 = ~n13989 & ~n14001 ;
  assign n14003 = ~n14000 & ~n14001 ;
  assign n14004 = ~n14002 & ~n14003 ;
  assign n14005 = ~n13914 & n14004 ;
  assign n14006 = n13914 & ~n14004 ;
  assign n14007 = ~n14005 & ~n14006 ;
  assign n14008 = ~x82 & n5560 ;
  assign n14009 = ~x80 & n5943 ;
  assign n14010 = ~x81 & n5555 ;
  assign n14011 = ~n14009 & ~n14010 ;
  assign n14012 = ~n14008 & n14011 ;
  assign n14013 = n2697 & n5563 ;
  assign n14014 = n14012 & ~n14013 ;
  assign n14015 = ~x29 & ~n14014 ;
  assign n14016 = ~x29 & ~n14015 ;
  assign n14017 = ~n14014 & ~n14015 ;
  assign n14018 = ~n14016 & ~n14017 ;
  assign n14019 = ~n14007 & ~n14018 ;
  assign n14020 = n14007 & n14018 ;
  assign n14021 = ~n14019 & ~n14020 ;
  assign n14022 = ~n13913 & n14021 ;
  assign n14023 = n13913 & ~n14021 ;
  assign n14024 = ~n14022 & ~n14023 ;
  assign n14025 = ~x85 & n4531 ;
  assign n14026 = ~x83 & n4847 ;
  assign n14027 = ~x84 & n4526 ;
  assign n14028 = ~n14026 & ~n14027 ;
  assign n14029 = ~n14025 & n14028 ;
  assign n14030 = n3521 & n4534 ;
  assign n14031 = n14029 & ~n14030 ;
  assign n14032 = ~x26 & ~n14031 ;
  assign n14033 = ~x26 & ~n14032 ;
  assign n14034 = ~n14031 & ~n14032 ;
  assign n14035 = ~n14033 & ~n14034 ;
  assign n14036 = n14024 & ~n14035 ;
  assign n14037 = n14024 & ~n14036 ;
  assign n14038 = ~n14035 & ~n14036 ;
  assign n14039 = ~n14037 & ~n14038 ;
  assign n14040 = ~n13492 & ~n13498 ;
  assign n14041 = n14039 & n14040 ;
  assign n14042 = ~n14039 & ~n14040 ;
  assign n14043 = ~n14041 & ~n14042 ;
  assign n14044 = ~x88 & n3589 ;
  assign n14045 = ~x86 & n3878 ;
  assign n14046 = ~x87 & n3584 ;
  assign n14047 = ~n14045 & ~n14046 ;
  assign n14048 = ~n14044 & n14047 ;
  assign n14049 = n3592 & n4457 ;
  assign n14050 = n14048 & ~n14049 ;
  assign n14051 = ~x23 & ~n14050 ;
  assign n14052 = ~x23 & ~n14051 ;
  assign n14053 = ~n14050 & ~n14051 ;
  assign n14054 = ~n14052 & ~n14053 ;
  assign n14055 = ~n14043 & n14054 ;
  assign n14056 = n14043 & ~n14054 ;
  assign n14057 = ~n14055 & ~n14056 ;
  assign n14058 = ~n13516 & n14057 ;
  assign n14059 = n13516 & ~n14057 ;
  assign n14060 = ~n14058 & ~n14059 ;
  assign n14061 = ~x91 & n2751 ;
  assign n14062 = ~x89 & n3020 ;
  assign n14063 = ~x90 & n2746 ;
  assign n14064 = ~n14062 & ~n14063 ;
  assign n14065 = ~n14061 & n14064 ;
  assign n14066 = n2754 & n5507 ;
  assign n14067 = n14065 & ~n14066 ;
  assign n14068 = ~x20 & ~n14067 ;
  assign n14069 = ~x20 & ~n14068 ;
  assign n14070 = ~n14067 & ~n14068 ;
  assign n14071 = ~n14069 & ~n14070 ;
  assign n14072 = n14060 & ~n14071 ;
  assign n14073 = n14060 & ~n14072 ;
  assign n14074 = ~n14071 & ~n14072 ;
  assign n14075 = ~n14073 & ~n14074 ;
  assign n14076 = ~n13912 & n14075 ;
  assign n14077 = n13912 & ~n14075 ;
  assign n14078 = ~n14076 & ~n14077 ;
  assign n14079 = ~x94 & n2093 ;
  assign n14080 = ~x92 & n2275 ;
  assign n14081 = ~x93 & n2088 ;
  assign n14082 = ~n14080 & ~n14081 ;
  assign n14083 = ~n14079 & n14082 ;
  assign n14084 = n2096 & n6671 ;
  assign n14085 = n14083 & ~n14084 ;
  assign n14086 = ~x17 & ~n14085 ;
  assign n14087 = ~x17 & ~n14086 ;
  assign n14088 = ~n14085 & ~n14086 ;
  assign n14089 = ~n14087 & ~n14088 ;
  assign n14090 = ~n14078 & ~n14089 ;
  assign n14091 = n14078 & n14089 ;
  assign n14092 = ~n14090 & ~n14091 ;
  assign n14093 = ~n13911 & n14092 ;
  assign n14094 = n13911 & ~n14092 ;
  assign n14095 = ~n14093 & ~n14094 ;
  assign n14096 = ~x97 & n1434 ;
  assign n14097 = ~x95 & n1646 ;
  assign n14098 = ~x96 & n1429 ;
  assign n14099 = ~n14097 & ~n14098 ;
  assign n14100 = ~n14096 & n14099 ;
  assign n14101 = n1437 & n7949 ;
  assign n14102 = n14100 & ~n14101 ;
  assign n14103 = ~x14 & ~n14102 ;
  assign n14104 = ~x14 & ~n14103 ;
  assign n14105 = ~n14102 & ~n14103 ;
  assign n14106 = ~n14104 & ~n14105 ;
  assign n14107 = n14095 & ~n14106 ;
  assign n14108 = n14095 & ~n14107 ;
  assign n14109 = ~n14106 & ~n14107 ;
  assign n14110 = ~n14108 & ~n14109 ;
  assign n14111 = ~n13910 & n14110 ;
  assign n14112 = n13910 & ~n14110 ;
  assign n14113 = ~n14111 & ~n14112 ;
  assign n14114 = ~x100 & n945 ;
  assign n14115 = ~x98 & n1099 ;
  assign n14116 = ~x99 & n940 ;
  assign n14117 = ~n14115 & ~n14116 ;
  assign n14118 = ~n14114 & n14117 ;
  assign n14119 = n948 & n9338 ;
  assign n14120 = n14118 & ~n14119 ;
  assign n14121 = ~x11 & ~n14120 ;
  assign n14122 = ~x11 & ~n14121 ;
  assign n14123 = ~n14120 & ~n14121 ;
  assign n14124 = ~n14122 & ~n14123 ;
  assign n14125 = ~n14113 & ~n14124 ;
  assign n14126 = n14113 & n14124 ;
  assign n14127 = ~n14125 & ~n14126 ;
  assign n14128 = n13909 & ~n14127 ;
  assign n14129 = ~n13909 & n14127 ;
  assign n14130 = ~n14128 & ~n14129 ;
  assign n14131 = ~x103 & n574 ;
  assign n14132 = ~x101 & n673 ;
  assign n14133 = ~x102 & n569 ;
  assign n14134 = ~n14132 & ~n14133 ;
  assign n14135 = ~n14131 & n14134 ;
  assign n14136 = n577 & n10833 ;
  assign n14137 = n14135 & ~n14136 ;
  assign n14138 = ~x8 & ~n14137 ;
  assign n14139 = ~x8 & ~n14138 ;
  assign n14140 = ~n14137 & ~n14138 ;
  assign n14141 = ~n14139 & ~n14140 ;
  assign n14142 = n14130 & ~n14141 ;
  assign n14143 = n14130 & ~n14142 ;
  assign n14144 = ~n14141 & ~n14142 ;
  assign n14145 = ~n14143 & ~n14144 ;
  assign n14146 = ~n13578 & ~n13582 ;
  assign n14147 = n14145 & n14146 ;
  assign n14148 = ~n14145 & ~n14146 ;
  assign n14149 = ~n14147 & ~n14148 ;
  assign n14150 = ~x106 & n293 ;
  assign n14151 = ~x104 & n373 ;
  assign n14152 = ~x105 & n288 ;
  assign n14153 = ~n14151 & ~n14152 ;
  assign n14154 = ~n14150 & n14153 ;
  assign n14155 = n296 & n12447 ;
  assign n14156 = n14154 & ~n14155 ;
  assign n14157 = ~x5 & ~n14156 ;
  assign n14158 = ~x5 & ~n14157 ;
  assign n14159 = ~n14156 & ~n14157 ;
  assign n14160 = ~n14158 & ~n14159 ;
  assign n14161 = n14149 & ~n14160 ;
  assign n14162 = n14149 & ~n14161 ;
  assign n14163 = ~n14160 & ~n14161 ;
  assign n14164 = ~n14162 & ~n14163 ;
  assign n14165 = ~n13585 & ~n13589 ;
  assign n14166 = n14164 & n14165 ;
  assign n14167 = ~n14164 & ~n14165 ;
  assign n14168 = ~n14166 & ~n14167 ;
  assign n14169 = ~x109 & n164 ;
  assign n14170 = ~x107 & n205 ;
  assign n14171 = ~x108 & n162 ;
  assign n14172 = ~n14170 & ~n14171 ;
  assign n14173 = ~n14169 & n14172 ;
  assign n14174 = ~n13318 & ~n13599 ;
  assign n14175 = n13891 & ~n14174 ;
  assign n14176 = ~n13891 & n14174 ;
  assign n14177 = ~n14175 & ~n14176 ;
  assign n14178 = n167 & n14177 ;
  assign n14179 = n14173 & ~n14178 ;
  assign n14180 = ~x2 & ~n14179 ;
  assign n14181 = ~x2 & ~n14180 ;
  assign n14182 = ~n14179 & ~n14180 ;
  assign n14183 = ~n14181 & ~n14182 ;
  assign n14184 = ~n14168 & n14183 ;
  assign n14185 = n14168 & ~n14183 ;
  assign n14186 = ~n14184 & ~n14185 ;
  assign n14187 = ~n13908 & n14186 ;
  assign n14188 = n13908 & ~n14186 ;
  assign n14189 = ~n14187 & ~n14188 ;
  assign n14192 = ~n14189 & ~x173 ;
  assign n14193 = ~n14191 & ~n14192 ;
  assign n14194 = ~n13856 & ~n13862 ;
  assign n14195 = ~n13804 & ~n13807 ;
  assign n14196 = ~n13623 & ~n13789 ;
  assign n14197 = ~n13786 & ~n14196 ;
  assign n14198 = x92 & n2751 ;
  assign n14199 = x90 & n3020 ;
  assign n14200 = x91 & n2746 ;
  assign n14201 = ~n14199 & ~n14200 ;
  assign n14202 = ~n14198 & n14201 ;
  assign n14203 = n2754 & n5710 ;
  assign n14204 = n14202 & ~n14203 ;
  assign n14205 = x20 & ~n14204 ;
  assign n14206 = x20 & ~n14205 ;
  assign n14207 = ~n14204 & ~n14205 ;
  assign n14208 = ~n14206 & ~n14207 ;
  assign n14209 = ~n13696 & ~n13700 ;
  assign n14210 = ~n13691 & ~n13693 ;
  assign n14211 = n13143 & n13642 ;
  assign n14212 = ~n13657 & ~n14211 ;
  assign n14213 = x68 & n12506 ;
  assign n14214 = x66 & n13131 ;
  assign n14215 = x67 & n12501 ;
  assign n14216 = ~n14214 & ~n14215 ;
  assign n14217 = ~n14213 & n14216 ;
  assign n14218 = n317 & n12509 ;
  assign n14219 = n14217 & ~n14218 ;
  assign n14220 = x44 & ~n14219 ;
  assign n14221 = x44 & ~n14220 ;
  assign n14222 = ~n14219 & ~n14220 ;
  assign n14223 = ~n14221 & ~n14222 ;
  assign n14224 = x47 & ~n13642 ;
  assign n14225 = ~x45 & x46 ;
  assign n14226 = x45 & ~x46 ;
  assign n14227 = ~n14225 & ~n14226 ;
  assign n14228 = n13641 & ~n14227 ;
  assign n14229 = x64 & n14228 ;
  assign n14230 = ~x46 & x47 ;
  assign n14231 = x46 & ~x47 ;
  assign n14232 = ~n14230 & ~n14231 ;
  assign n14233 = ~n13641 & n14232 ;
  assign n14234 = x65 & n14233 ;
  assign n14235 = ~n14229 & ~n14234 ;
  assign n14236 = ~n13641 & ~n14232 ;
  assign n14237 = ~n152 & n14236 ;
  assign n14238 = n14235 & ~n14237 ;
  assign n14239 = x47 & ~n14238 ;
  assign n14240 = x47 & ~n14239 ;
  assign n14241 = ~n14238 & ~n14239 ;
  assign n14242 = ~n14240 & ~n14241 ;
  assign n14243 = n14224 & ~n14242 ;
  assign n14244 = ~n14224 & n14242 ;
  assign n14245 = ~n14243 & ~n14244 ;
  assign n14246 = n14223 & ~n14245 ;
  assign n14247 = ~n14223 & n14245 ;
  assign n14248 = ~n14246 & ~n14247 ;
  assign n14249 = ~n14212 & n14248 ;
  assign n14250 = n14212 & ~n14248 ;
  assign n14251 = ~n14249 & ~n14250 ;
  assign n14252 = x71 & n10905 ;
  assign n14253 = x69 & n11466 ;
  assign n14254 = x70 & n10900 ;
  assign n14255 = ~n14253 & ~n14254 ;
  assign n14256 = ~n14252 & n14255 ;
  assign n14257 = n558 & n10908 ;
  assign n14258 = n14256 & ~n14257 ;
  assign n14259 = x41 & ~n14258 ;
  assign n14260 = x41 & ~n14259 ;
  assign n14261 = ~n14258 & ~n14259 ;
  assign n14262 = ~n14260 & ~n14261 ;
  assign n14263 = n14251 & ~n14262 ;
  assign n14264 = n14251 & ~n14263 ;
  assign n14265 = ~n14262 & ~n14263 ;
  assign n14266 = ~n14264 & ~n14265 ;
  assign n14267 = ~n13671 & ~n13677 ;
  assign n14268 = n14266 & n14267 ;
  assign n14269 = ~n14266 & ~n14267 ;
  assign n14270 = ~n14268 & ~n14269 ;
  assign n14271 = x74 & n9433 ;
  assign n14272 = x72 & n9915 ;
  assign n14273 = x73 & n9428 ;
  assign n14274 = ~n14272 & ~n14273 ;
  assign n14275 = ~n14271 & n14274 ;
  assign n14276 = n994 & n9436 ;
  assign n14277 = n14275 & ~n14276 ;
  assign n14278 = x38 & ~n14277 ;
  assign n14279 = x38 & ~n14278 ;
  assign n14280 = ~n14277 & ~n14278 ;
  assign n14281 = ~n14279 & ~n14280 ;
  assign n14282 = n14270 & ~n14281 ;
  assign n14283 = ~n14270 & n14281 ;
  assign n14284 = ~n14210 & ~n14283 ;
  assign n14285 = ~n14282 & n14284 ;
  assign n14286 = ~n14210 & ~n14285 ;
  assign n14287 = ~n14282 & ~n14285 ;
  assign n14288 = ~n14283 & n14287 ;
  assign n14289 = ~n14286 & ~n14288 ;
  assign n14290 = x77 & n8006 ;
  assign n14291 = x75 & n8474 ;
  assign n14292 = x76 & n8001 ;
  assign n14293 = ~n14291 & ~n14292 ;
  assign n14294 = ~n14290 & n14293 ;
  assign n14295 = n1502 & n8009 ;
  assign n14296 = n14294 & ~n14295 ;
  assign n14297 = x35 & ~n14296 ;
  assign n14298 = x35 & ~n14297 ;
  assign n14299 = ~n14296 & ~n14297 ;
  assign n14300 = ~n14298 & ~n14299 ;
  assign n14301 = n14289 & n14300 ;
  assign n14302 = ~n14289 & ~n14300 ;
  assign n14303 = ~n14301 & ~n14302 ;
  assign n14304 = ~n14209 & n14303 ;
  assign n14305 = n14209 & ~n14303 ;
  assign n14306 = ~n14304 & ~n14305 ;
  assign n14307 = x80 & n6725 ;
  assign n14308 = x78 & n7129 ;
  assign n14309 = x79 & n6720 ;
  assign n14310 = ~n14308 & ~n14309 ;
  assign n14311 = ~n14307 & n14310 ;
  assign n14312 = n2028 & n6728 ;
  assign n14313 = n14311 & ~n14312 ;
  assign n14314 = x32 & ~n14313 ;
  assign n14315 = x32 & ~n14314 ;
  assign n14316 = ~n14313 & ~n14314 ;
  assign n14317 = ~n14315 & ~n14316 ;
  assign n14318 = n14306 & ~n14317 ;
  assign n14319 = n14306 & ~n14318 ;
  assign n14320 = ~n14317 & ~n14318 ;
  assign n14321 = ~n14319 & ~n14320 ;
  assign n14322 = ~n13625 & ~n13718 ;
  assign n14323 = ~n13715 & ~n14322 ;
  assign n14324 = n14321 & n14323 ;
  assign n14325 = ~n14321 & ~n14323 ;
  assign n14326 = ~n14324 & ~n14325 ;
  assign n14327 = x83 & n5560 ;
  assign n14328 = x81 & n5943 ;
  assign n14329 = x82 & n5555 ;
  assign n14330 = ~n14328 & ~n14329 ;
  assign n14331 = ~n14327 & n14330 ;
  assign n14332 = n2843 & n5563 ;
  assign n14333 = n14331 & ~n14332 ;
  assign n14334 = x29 & ~n14333 ;
  assign n14335 = x29 & ~n14334 ;
  assign n14336 = ~n14333 & ~n14334 ;
  assign n14337 = ~n14335 & ~n14336 ;
  assign n14338 = n14326 & ~n14337 ;
  assign n14339 = n14326 & ~n14338 ;
  assign n14340 = ~n14337 & ~n14338 ;
  assign n14341 = ~n14339 & ~n14340 ;
  assign n14342 = ~n13733 & ~n13736 ;
  assign n14343 = n14341 & n14342 ;
  assign n14344 = ~n14341 & ~n14342 ;
  assign n14345 = ~n14343 & ~n14344 ;
  assign n14346 = x86 & n4531 ;
  assign n14347 = x84 & n4847 ;
  assign n14348 = x85 & n4526 ;
  assign n14349 = ~n14347 & ~n14348 ;
  assign n14350 = ~n14346 & n14349 ;
  assign n14351 = n3686 & n4534 ;
  assign n14352 = n14350 & ~n14351 ;
  assign n14353 = x26 & ~n14352 ;
  assign n14354 = x26 & ~n14353 ;
  assign n14355 = ~n14352 & ~n14353 ;
  assign n14356 = ~n14354 & ~n14355 ;
  assign n14357 = n14345 & ~n14356 ;
  assign n14358 = n14345 & ~n14357 ;
  assign n14359 = ~n14356 & ~n14357 ;
  assign n14360 = ~n14358 & ~n14359 ;
  assign n14361 = ~n13750 & ~n13756 ;
  assign n14362 = n14360 & n14361 ;
  assign n14363 = ~n14360 & ~n14361 ;
  assign n14364 = ~n14362 & ~n14363 ;
  assign n14365 = x89 & n3589 ;
  assign n14366 = x87 & n3878 ;
  assign n14367 = x88 & n3584 ;
  assign n14368 = ~n14366 & ~n14367 ;
  assign n14369 = ~n14365 & n14368 ;
  assign n14370 = n3592 & n4488 ;
  assign n14371 = n14369 & ~n14370 ;
  assign n14372 = x23 & ~n14371 ;
  assign n14373 = x23 & ~n14372 ;
  assign n14374 = ~n14371 & ~n14372 ;
  assign n14375 = ~n14373 & ~n14374 ;
  assign n14376 = n14364 & ~n14375 ;
  assign n14377 = n14364 & ~n14376 ;
  assign n14378 = ~n14375 & ~n14376 ;
  assign n14379 = ~n14377 & ~n14378 ;
  assign n14380 = ~n13770 & ~n13772 ;
  assign n14381 = ~n14379 & ~n14380 ;
  assign n14382 = n14379 & n14380 ;
  assign n14383 = ~n14381 & ~n14382 ;
  assign n14384 = ~n14208 & n14383 ;
  assign n14385 = ~n14208 & ~n14384 ;
  assign n14386 = n14383 & ~n14384 ;
  assign n14387 = ~n14385 & ~n14386 ;
  assign n14388 = ~n14197 & ~n14387 ;
  assign n14389 = ~n14197 & ~n14388 ;
  assign n14390 = ~n14387 & ~n14388 ;
  assign n14391 = ~n14389 & ~n14390 ;
  assign n14392 = x95 & n2093 ;
  assign n14393 = x93 & n2275 ;
  assign n14394 = x94 & n2088 ;
  assign n14395 = ~n14393 & ~n14394 ;
  assign n14396 = ~n14392 & n14395 ;
  assign n14397 = n2096 & n6894 ;
  assign n14398 = n14396 & ~n14397 ;
  assign n14399 = x17 & ~n14398 ;
  assign n14400 = x17 & ~n14399 ;
  assign n14401 = ~n14398 & ~n14399 ;
  assign n14402 = ~n14400 & ~n14401 ;
  assign n14403 = n14391 & n14402 ;
  assign n14404 = ~n14391 & ~n14402 ;
  assign n14405 = ~n14403 & ~n14404 ;
  assign n14406 = ~n14195 & n14405 ;
  assign n14407 = n14195 & ~n14405 ;
  assign n14408 = ~n14406 & ~n14407 ;
  assign n14409 = x98 & n1434 ;
  assign n14410 = x96 & n1646 ;
  assign n14411 = x97 & n1429 ;
  assign n14412 = ~n14410 & ~n14411 ;
  assign n14413 = ~n14409 & n14412 ;
  assign n14414 = n1437 & n8196 ;
  assign n14415 = n14413 & ~n14414 ;
  assign n14416 = x14 & ~n14415 ;
  assign n14417 = x14 & ~n14416 ;
  assign n14418 = ~n14415 & ~n14416 ;
  assign n14419 = ~n14417 & ~n14418 ;
  assign n14420 = n14408 & ~n14419 ;
  assign n14421 = n14408 & ~n14420 ;
  assign n14422 = ~n14419 & ~n14420 ;
  assign n14423 = ~n14421 & ~n14422 ;
  assign n14424 = ~n13621 & ~n13824 ;
  assign n14425 = ~n13821 & ~n14424 ;
  assign n14426 = n14423 & n14425 ;
  assign n14427 = ~n14423 & ~n14425 ;
  assign n14428 = ~n14426 & ~n14427 ;
  assign n14429 = x101 & n945 ;
  assign n14430 = x99 & n1099 ;
  assign n14431 = x100 & n940 ;
  assign n14432 = ~n14430 & ~n14431 ;
  assign n14433 = ~n14429 & n14432 ;
  assign n14434 = n948 & n9601 ;
  assign n14435 = n14433 & ~n14434 ;
  assign n14436 = x11 & ~n14435 ;
  assign n14437 = x11 & ~n14436 ;
  assign n14438 = ~n14435 & ~n14436 ;
  assign n14439 = ~n14437 & ~n14438 ;
  assign n14440 = n14428 & ~n14439 ;
  assign n14441 = n14428 & ~n14440 ;
  assign n14442 = ~n14439 & ~n14440 ;
  assign n14443 = ~n14441 & ~n14442 ;
  assign n14444 = ~n13839 & ~n13843 ;
  assign n14445 = n14443 & n14444 ;
  assign n14446 = ~n14443 & ~n14444 ;
  assign n14447 = ~n14445 & ~n14446 ;
  assign n14448 = x104 & n574 ;
  assign n14449 = x102 & n673 ;
  assign n14450 = x103 & n569 ;
  assign n14451 = ~n14449 & ~n14450 ;
  assign n14452 = ~n14448 & n14451 ;
  assign n14453 = n577 & n11116 ;
  assign n14454 = n14452 & ~n14453 ;
  assign n14455 = x8 & ~n14454 ;
  assign n14456 = x8 & ~n14455 ;
  assign n14457 = ~n14454 & ~n14455 ;
  assign n14458 = ~n14456 & ~n14457 ;
  assign n14459 = n14447 & ~n14458 ;
  assign n14460 = ~n14447 & n14458 ;
  assign n14461 = ~n14194 & ~n14460 ;
  assign n14462 = ~n14459 & n14461 ;
  assign n14463 = ~n14194 & ~n14462 ;
  assign n14464 = ~n14459 & ~n14462 ;
  assign n14465 = ~n14460 & n14464 ;
  assign n14466 = ~n14463 & ~n14465 ;
  assign n14467 = x107 & n293 ;
  assign n14468 = x105 & n373 ;
  assign n14469 = x106 & n288 ;
  assign n14470 = ~n14468 & ~n14469 ;
  assign n14471 = ~n14467 & n14470 ;
  assign n14472 = n296 & n12749 ;
  assign n14473 = n14471 & ~n14472 ;
  assign n14474 = x5 & ~n14473 ;
  assign n14475 = x5 & ~n14474 ;
  assign n14476 = ~n14473 & ~n14474 ;
  assign n14477 = ~n14475 & ~n14476 ;
  assign n14478 = ~n14466 & ~n14477 ;
  assign n14479 = ~n14466 & ~n14478 ;
  assign n14480 = ~n14477 & ~n14478 ;
  assign n14481 = ~n14479 & ~n14480 ;
  assign n14482 = ~n13875 & ~n13881 ;
  assign n14483 = n14481 & n14482 ;
  assign n14484 = ~n14481 & ~n14482 ;
  assign n14485 = ~n14483 & ~n14484 ;
  assign n14486 = x110 & n146 ;
  assign n14487 = x108 & n182 ;
  assign n14488 = x109 & n141 ;
  assign n14489 = ~n14487 & ~n14488 ;
  assign n14490 = ~n14486 & n14489 ;
  assign n14491 = ~n13890 & ~n13892 ;
  assign n14492 = ~x109 & ~x110 ;
  assign n14493 = x109 & x110 ;
  assign n14494 = ~n14492 & ~n14493 ;
  assign n14495 = ~n14491 & n14494 ;
  assign n14496 = n14491 & ~n14494 ;
  assign n14497 = ~n14495 & ~n14496 ;
  assign n14498 = n149 & n14497 ;
  assign n14499 = n14490 & ~n14498 ;
  assign n14500 = x2 & ~n14499 ;
  assign n14501 = x2 & ~n14500 ;
  assign n14502 = ~n14499 & ~n14500 ;
  assign n14503 = ~n14501 & ~n14502 ;
  assign n14504 = n14485 & ~n14503 ;
  assign n14505 = n14485 & ~n14504 ;
  assign n14506 = ~n14503 & ~n14504 ;
  assign n14507 = ~n14505 & ~n14506 ;
  assign n14508 = ~n13902 & ~n13904 ;
  assign n14509 = ~n14507 & ~n14508 ;
  assign n14510 = n14507 & n14508 ;
  assign n14511 = ~n14509 & ~n14510 ;
  assign n14818 = n14511 & x174 ;
  assign n14512 = ~n14142 & ~n14148 ;
  assign n14513 = ~n14090 & ~n14093 ;
  assign n14514 = ~n13912 & ~n14075 ;
  assign n14515 = ~n14072 & ~n14514 ;
  assign n14516 = ~x92 & n2751 ;
  assign n14517 = ~x90 & n3020 ;
  assign n14518 = ~x91 & n2746 ;
  assign n14519 = ~n14517 & ~n14518 ;
  assign n14520 = ~n14516 & n14519 ;
  assign n14521 = n2754 & n5896 ;
  assign n14522 = n14520 & ~n14521 ;
  assign n14523 = ~x20 & ~n14522 ;
  assign n14524 = ~x20 & ~n14523 ;
  assign n14525 = ~n14522 & ~n14523 ;
  assign n14526 = ~n14524 & ~n14525 ;
  assign n14527 = ~n13982 & ~n13986 ;
  assign n14528 = ~n13977 & ~n13979 ;
  assign n14529 = n13424 & n13928 ;
  assign n14530 = ~n13943 & ~n14529 ;
  assign n14531 = ~x68 & n12506 ;
  assign n14532 = ~x66 & n13131 ;
  assign n14533 = ~x67 & n12501 ;
  assign n14534 = ~n14532 & ~n14533 ;
  assign n14535 = ~n14531 & n14534 ;
  assign n14536 = n352 & n12509 ;
  assign n14537 = n14535 & ~n14536 ;
  assign n14538 = ~x44 & ~n14537 ;
  assign n14539 = ~x44 & ~n14538 ;
  assign n14540 = ~n14537 & ~n14538 ;
  assign n14541 = ~n14539 & ~n14540 ;
  assign n14542 = ~x47 & ~n13928 ;
  assign n14543 = ~x64 & n14228 ;
  assign n14544 = ~x65 & n14233 ;
  assign n14545 = ~n14543 & ~n14544 ;
  assign n14546 = ~n14237 & n14545 ;
  assign n14547 = ~x47 & ~n14546 ;
  assign n14548 = ~x47 & ~n14547 ;
  assign n14549 = ~n14546 & ~n14547 ;
  assign n14550 = ~n14548 & ~n14549 ;
  assign n14551 = n14542 & ~n14550 ;
  assign n14552 = ~n14542 & n14550 ;
  assign n14553 = ~n14551 & ~n14552 ;
  assign n14554 = n14541 & ~n14553 ;
  assign n14555 = ~n14541 & n14553 ;
  assign n14556 = ~n14554 & ~n14555 ;
  assign n14557 = ~n14530 & n14556 ;
  assign n14558 = n14530 & ~n14556 ;
  assign n14559 = ~n14557 & ~n14558 ;
  assign n14560 = ~x71 & n10905 ;
  assign n14561 = ~x69 & n11466 ;
  assign n14562 = ~x70 & n10900 ;
  assign n14563 = ~n14561 & ~n14562 ;
  assign n14564 = ~n14560 & n14563 ;
  assign n14565 = n622 & n10908 ;
  assign n14566 = n14564 & ~n14565 ;
  assign n14567 = ~x41 & ~n14566 ;
  assign n14568 = ~x41 & ~n14567 ;
  assign n14569 = ~n14566 & ~n14567 ;
  assign n14570 = ~n14568 & ~n14569 ;
  assign n14571 = n14559 & ~n14570 ;
  assign n14572 = n14559 & ~n14571 ;
  assign n14573 = ~n14570 & ~n14571 ;
  assign n14574 = ~n14572 & ~n14573 ;
  assign n14575 = ~n13957 & ~n13963 ;
  assign n14576 = n14574 & n14575 ;
  assign n14577 = ~n14574 & ~n14575 ;
  assign n14578 = ~n14576 & ~n14577 ;
  assign n14579 = ~x74 & n9433 ;
  assign n14580 = ~x72 & n9915 ;
  assign n14581 = ~x73 & n9428 ;
  assign n14582 = ~n14580 & ~n14581 ;
  assign n14583 = ~n14579 & n14582 ;
  assign n14584 = n1066 & n9436 ;
  assign n14585 = n14583 & ~n14584 ;
  assign n14586 = ~x38 & ~n14585 ;
  assign n14587 = ~x38 & ~n14586 ;
  assign n14588 = ~n14585 & ~n14586 ;
  assign n14589 = ~n14587 & ~n14588 ;
  assign n14590 = n14578 & ~n14589 ;
  assign n14591 = ~n14578 & n14589 ;
  assign n14592 = ~n14528 & ~n14591 ;
  assign n14593 = ~n14590 & n14592 ;
  assign n14594 = ~n14528 & ~n14593 ;
  assign n14595 = ~n14590 & ~n14593 ;
  assign n14596 = ~n14591 & n14595 ;
  assign n14597 = ~n14594 & ~n14596 ;
  assign n14598 = ~x77 & n8006 ;
  assign n14599 = ~x75 & n8474 ;
  assign n14600 = ~x76 & n8001 ;
  assign n14601 = ~n14599 & ~n14600 ;
  assign n14602 = ~n14598 & n14601 ;
  assign n14603 = n1594 & n8009 ;
  assign n14604 = n14602 & ~n14603 ;
  assign n14605 = ~x35 & ~n14604 ;
  assign n14606 = ~x35 & ~n14605 ;
  assign n14607 = ~n14604 & ~n14605 ;
  assign n14608 = ~n14606 & ~n14607 ;
  assign n14609 = n14597 & n14608 ;
  assign n14610 = ~n14597 & ~n14608 ;
  assign n14611 = ~n14609 & ~n14610 ;
  assign n14612 = ~n14527 & n14611 ;
  assign n14613 = n14527 & ~n14611 ;
  assign n14614 = ~n14612 & ~n14613 ;
  assign n14615 = ~x80 & n6725 ;
  assign n14616 = ~x78 & n7129 ;
  assign n14617 = ~x79 & n6720 ;
  assign n14618 = ~n14616 & ~n14617 ;
  assign n14619 = ~n14615 & n14618 ;
  assign n14620 = n2145 & n6728 ;
  assign n14621 = n14619 & ~n14620 ;
  assign n14622 = ~x32 & ~n14621 ;
  assign n14623 = ~x32 & ~n14622 ;
  assign n14624 = ~n14621 & ~n14622 ;
  assign n14625 = ~n14623 & ~n14624 ;
  assign n14626 = n14614 & ~n14625 ;
  assign n14627 = n14614 & ~n14626 ;
  assign n14628 = ~n14625 & ~n14626 ;
  assign n14629 = ~n14627 & ~n14628 ;
  assign n14630 = ~n13914 & ~n14004 ;
  assign n14631 = ~n14001 & ~n14630 ;
  assign n14632 = n14629 & n14631 ;
  assign n14633 = ~n14629 & ~n14631 ;
  assign n14634 = ~n14632 & ~n14633 ;
  assign n14635 = ~x83 & n5560 ;
  assign n14636 = ~x81 & n5943 ;
  assign n14637 = ~x82 & n5555 ;
  assign n14638 = ~n14636 & ~n14637 ;
  assign n14639 = ~n14635 & n14638 ;
  assign n14640 = n2972 & n5563 ;
  assign n14641 = n14639 & ~n14640 ;
  assign n14642 = ~x29 & ~n14641 ;
  assign n14643 = ~x29 & ~n14642 ;
  assign n14644 = ~n14641 & ~n14642 ;
  assign n14645 = ~n14643 & ~n14644 ;
  assign n14646 = n14634 & ~n14645 ;
  assign n14647 = n14634 & ~n14646 ;
  assign n14648 = ~n14645 & ~n14646 ;
  assign n14649 = ~n14647 & ~n14648 ;
  assign n14650 = ~n14019 & ~n14022 ;
  assign n14651 = n14649 & n14650 ;
  assign n14652 = ~n14649 & ~n14650 ;
  assign n14653 = ~n14651 & ~n14652 ;
  assign n14654 = ~x86 & n4531 ;
  assign n14655 = ~x84 & n4847 ;
  assign n14656 = ~x85 & n4526 ;
  assign n14657 = ~n14655 & ~n14656 ;
  assign n14658 = ~n14654 & n14657 ;
  assign n14659 = n3832 & n4534 ;
  assign n14660 = n14658 & ~n14659 ;
  assign n14661 = ~x26 & ~n14660 ;
  assign n14662 = ~x26 & ~n14661 ;
  assign n14663 = ~n14660 & ~n14661 ;
  assign n14664 = ~n14662 & ~n14663 ;
  assign n14665 = n14653 & ~n14664 ;
  assign n14666 = n14653 & ~n14665 ;
  assign n14667 = ~n14664 & ~n14665 ;
  assign n14668 = ~n14666 & ~n14667 ;
  assign n14669 = ~n14036 & ~n14042 ;
  assign n14670 = n14668 & n14669 ;
  assign n14671 = ~n14668 & ~n14669 ;
  assign n14672 = ~n14670 & ~n14671 ;
  assign n14673 = ~x89 & n3589 ;
  assign n14674 = ~x87 & n3878 ;
  assign n14675 = ~x88 & n3584 ;
  assign n14676 = ~n14674 & ~n14675 ;
  assign n14677 = ~n14673 & n14676 ;
  assign n14678 = n3592 & n4664 ;
  assign n14679 = n14677 & ~n14678 ;
  assign n14680 = ~x23 & ~n14679 ;
  assign n14681 = ~x23 & ~n14680 ;
  assign n14682 = ~n14679 & ~n14680 ;
  assign n14683 = ~n14681 & ~n14682 ;
  assign n14684 = n14672 & ~n14683 ;
  assign n14685 = n14672 & ~n14684 ;
  assign n14686 = ~n14683 & ~n14684 ;
  assign n14687 = ~n14685 & ~n14686 ;
  assign n14688 = ~n14056 & ~n14058 ;
  assign n14689 = ~n14687 & ~n14688 ;
  assign n14690 = n14687 & n14688 ;
  assign n14691 = ~n14689 & ~n14690 ;
  assign n14692 = ~n14526 & n14691 ;
  assign n14693 = ~n14526 & ~n14692 ;
  assign n14694 = n14691 & ~n14692 ;
  assign n14695 = ~n14693 & ~n14694 ;
  assign n14696 = ~n14515 & ~n14695 ;
  assign n14697 = ~n14515 & ~n14696 ;
  assign n14698 = ~n14695 & ~n14696 ;
  assign n14699 = ~n14697 & ~n14698 ;
  assign n14700 = ~x95 & n2093 ;
  assign n14701 = ~x93 & n2275 ;
  assign n14702 = ~x94 & n2088 ;
  assign n14703 = ~n14701 & ~n14702 ;
  assign n14704 = ~n14700 & n14703 ;
  assign n14705 = n2096 & n7100 ;
  assign n14706 = n14704 & ~n14705 ;
  assign n14707 = ~x17 & ~n14706 ;
  assign n14708 = ~x17 & ~n14707 ;
  assign n14709 = ~n14706 & ~n14707 ;
  assign n14710 = ~n14708 & ~n14709 ;
  assign n14711 = n14699 & n14710 ;
  assign n14712 = ~n14699 & ~n14710 ;
  assign n14713 = ~n14711 & ~n14712 ;
  assign n14714 = ~n14513 & n14713 ;
  assign n14715 = n14513 & ~n14713 ;
  assign n14716 = ~n14714 & ~n14715 ;
  assign n14717 = ~x98 & n1434 ;
  assign n14718 = ~x96 & n1646 ;
  assign n14719 = ~x97 & n1429 ;
  assign n14720 = ~n14718 & ~n14719 ;
  assign n14721 = ~n14717 & n14720 ;
  assign n14722 = n1437 & n8426 ;
  assign n14723 = n14721 & ~n14722 ;
  assign n14724 = ~x14 & ~n14723 ;
  assign n14725 = ~x14 & ~n14724 ;
  assign n14726 = ~n14723 & ~n14724 ;
  assign n14727 = ~n14725 & ~n14726 ;
  assign n14728 = n14716 & ~n14727 ;
  assign n14729 = n14716 & ~n14728 ;
  assign n14730 = ~n14727 & ~n14728 ;
  assign n14731 = ~n14729 & ~n14730 ;
  assign n14732 = ~n13910 & ~n14110 ;
  assign n14733 = ~n14107 & ~n14732 ;
  assign n14734 = n14731 & n14733 ;
  assign n14735 = ~n14731 & ~n14733 ;
  assign n14736 = ~n14734 & ~n14735 ;
  assign n14737 = ~x101 & n945 ;
  assign n14738 = ~x99 & n1099 ;
  assign n14739 = ~x100 & n940 ;
  assign n14740 = ~n14738 & ~n14739 ;
  assign n14741 = ~n14737 & n14740 ;
  assign n14742 = n948 & n9844 ;
  assign n14743 = n14741 & ~n14742 ;
  assign n14744 = ~x11 & ~n14743 ;
  assign n14745 = ~x11 & ~n14744 ;
  assign n14746 = ~n14743 & ~n14744 ;
  assign n14747 = ~n14745 & ~n14746 ;
  assign n14748 = n14736 & ~n14747 ;
  assign n14749 = n14736 & ~n14748 ;
  assign n14750 = ~n14747 & ~n14748 ;
  assign n14751 = ~n14749 & ~n14750 ;
  assign n14752 = ~n14125 & ~n14129 ;
  assign n14753 = n14751 & n14752 ;
  assign n14754 = ~n14751 & ~n14752 ;
  assign n14755 = ~n14753 & ~n14754 ;
  assign n14756 = ~x104 & n574 ;
  assign n14757 = ~x102 & n673 ;
  assign n14758 = ~x103 & n569 ;
  assign n14759 = ~n14757 & ~n14758 ;
  assign n14760 = ~n14756 & n14759 ;
  assign n14761 = n577 & n11380 ;
  assign n14762 = n14760 & ~n14761 ;
  assign n14763 = ~x8 & ~n14762 ;
  assign n14764 = ~x8 & ~n14763 ;
  assign n14765 = ~n14762 & ~n14763 ;
  assign n14766 = ~n14764 & ~n14765 ;
  assign n14767 = n14755 & ~n14766 ;
  assign n14768 = ~n14755 & n14766 ;
  assign n14769 = ~n14512 & ~n14768 ;
  assign n14770 = ~n14767 & n14769 ;
  assign n14771 = ~n14512 & ~n14770 ;
  assign n14772 = ~n14767 & ~n14770 ;
  assign n14773 = ~n14768 & n14772 ;
  assign n14774 = ~n14771 & ~n14773 ;
  assign n14775 = ~x107 & n293 ;
  assign n14776 = ~x105 & n373 ;
  assign n14777 = ~x106 & n288 ;
  assign n14778 = ~n14776 & ~n14777 ;
  assign n14779 = ~n14775 & n14778 ;
  assign n14780 = n296 & n13034 ;
  assign n14781 = n14779 & ~n14780 ;
  assign n14782 = ~x5 & ~n14781 ;
  assign n14783 = ~x5 & ~n14782 ;
  assign n14784 = ~n14781 & ~n14782 ;
  assign n14785 = ~n14783 & ~n14784 ;
  assign n14786 = ~n14774 & ~n14785 ;
  assign n14787 = ~n14774 & ~n14786 ;
  assign n14788 = ~n14785 & ~n14786 ;
  assign n14789 = ~n14787 & ~n14788 ;
  assign n14790 = ~n14161 & ~n14167 ;
  assign n14791 = n14789 & n14790 ;
  assign n14792 = ~n14789 & ~n14790 ;
  assign n14793 = ~n14791 & ~n14792 ;
  assign n14794 = ~x110 & n164 ;
  assign n14795 = ~x108 & n205 ;
  assign n14796 = ~x109 & n162 ;
  assign n14797 = ~n14795 & ~n14796 ;
  assign n14798 = ~n14794 & n14797 ;
  assign n14799 = ~n13889 & ~n14175 ;
  assign n14800 = n14494 & ~n14799 ;
  assign n14801 = ~n14494 & n14799 ;
  assign n14802 = ~n14800 & ~n14801 ;
  assign n14803 = n167 & n14802 ;
  assign n14804 = n14798 & ~n14803 ;
  assign n14805 = ~x2 & ~n14804 ;
  assign n14806 = ~x2 & ~n14805 ;
  assign n14807 = ~n14804 & ~n14805 ;
  assign n14808 = ~n14806 & ~n14807 ;
  assign n14809 = n14793 & ~n14808 ;
  assign n14810 = n14793 & ~n14809 ;
  assign n14811 = ~n14808 & ~n14809 ;
  assign n14812 = ~n14810 & ~n14811 ;
  assign n14813 = ~n14185 & ~n14187 ;
  assign n14814 = ~n14812 & ~n14813 ;
  assign n14815 = n14812 & n14813 ;
  assign n14816 = ~n14814 & ~n14815 ;
  assign n14819 = ~n14816 & ~x174 ;
  assign n14820 = ~n14818 & ~n14819 ;
  assign n14821 = ~n14478 & ~n14484 ;
  assign n14822 = ~n14404 & ~n14406 ;
  assign n14823 = x96 & n2093 ;
  assign n14824 = x94 & n2275 ;
  assign n14825 = x95 & n2088 ;
  assign n14826 = ~n14824 & ~n14825 ;
  assign n14827 = ~n14823 & n14826 ;
  assign n14828 = n2096 & n7321 ;
  assign n14829 = n14827 & ~n14828 ;
  assign n14830 = x17 & ~n14829 ;
  assign n14831 = x17 & ~n14830 ;
  assign n14832 = ~n14829 & ~n14830 ;
  assign n14833 = ~n14831 & ~n14832 ;
  assign n14834 = ~n14384 & ~n14388 ;
  assign n14835 = x93 & n2751 ;
  assign n14836 = x91 & n3020 ;
  assign n14837 = x92 & n2746 ;
  assign n14838 = ~n14836 & ~n14837 ;
  assign n14839 = ~n14835 & n14838 ;
  assign n14840 = n2754 & n6094 ;
  assign n14841 = n14839 & ~n14840 ;
  assign n14842 = x20 & ~n14841 ;
  assign n14843 = x20 & ~n14842 ;
  assign n14844 = ~n14841 & ~n14842 ;
  assign n14845 = ~n14843 & ~n14844 ;
  assign n14846 = ~n14376 & ~n14381 ;
  assign n14847 = ~n14357 & ~n14363 ;
  assign n14848 = ~n14318 & ~n14325 ;
  assign n14849 = x81 & n6725 ;
  assign n14850 = x79 & n7129 ;
  assign n14851 = x80 & n6720 ;
  assign n14852 = ~n14850 & ~n14851 ;
  assign n14853 = ~n14849 & n14852 ;
  assign n14854 = n2348 & n6728 ;
  assign n14855 = n14853 & ~n14854 ;
  assign n14856 = x32 & ~n14855 ;
  assign n14857 = x32 & ~n14856 ;
  assign n14858 = ~n14855 & ~n14856 ;
  assign n14859 = ~n14857 & ~n14858 ;
  assign n14860 = ~n14302 & ~n14304 ;
  assign n14861 = ~n14263 & ~n14269 ;
  assign n14862 = x72 & n10905 ;
  assign n14863 = x70 & n11466 ;
  assign n14864 = x71 & n10900 ;
  assign n14865 = ~n14863 & ~n14864 ;
  assign n14866 = ~n14862 & n14865 ;
  assign n14867 = n717 & n10908 ;
  assign n14868 = n14866 & ~n14867 ;
  assign n14869 = x41 & ~n14868 ;
  assign n14870 = x41 & ~n14869 ;
  assign n14871 = ~n14868 & ~n14869 ;
  assign n14872 = ~n14870 & ~n14871 ;
  assign n14873 = ~n14247 & ~n14249 ;
  assign n14874 = x66 & n14233 ;
  assign n14875 = n13641 & ~n14232 ;
  assign n14876 = n14227 & n14875 ;
  assign n14877 = x64 & n14876 ;
  assign n14878 = x65 & n14228 ;
  assign n14879 = ~n14877 & ~n14878 ;
  assign n14880 = ~n14874 & n14879 ;
  assign n14881 = n194 & n14236 ;
  assign n14882 = n14880 & ~n14881 ;
  assign n14883 = x47 & ~n14882 ;
  assign n14884 = x47 & ~n14883 ;
  assign n14885 = ~n14882 & ~n14883 ;
  assign n14886 = ~n14884 & ~n14885 ;
  assign n14887 = ~n14243 & n14886 ;
  assign n14888 = n14243 & ~n14886 ;
  assign n14889 = ~n14887 & ~n14888 ;
  assign n14890 = x69 & n12506 ;
  assign n14891 = x67 & n13131 ;
  assign n14892 = x68 & n12501 ;
  assign n14893 = ~n14891 & ~n14892 ;
  assign n14894 = ~n14890 & n14893 ;
  assign n14895 = n398 & n12509 ;
  assign n14896 = n14894 & ~n14895 ;
  assign n14897 = x44 & ~n14896 ;
  assign n14898 = x44 & ~n14897 ;
  assign n14899 = ~n14896 & ~n14897 ;
  assign n14900 = ~n14898 & ~n14899 ;
  assign n14901 = n14889 & ~n14900 ;
  assign n14902 = n14889 & ~n14901 ;
  assign n14903 = ~n14900 & ~n14901 ;
  assign n14904 = ~n14902 & ~n14903 ;
  assign n14905 = ~n14873 & ~n14904 ;
  assign n14906 = n14873 & n14904 ;
  assign n14907 = ~n14905 & ~n14906 ;
  assign n14908 = ~n14872 & n14907 ;
  assign n14909 = ~n14872 & ~n14908 ;
  assign n14910 = n14907 & ~n14908 ;
  assign n14911 = ~n14909 & ~n14910 ;
  assign n14912 = ~n14861 & ~n14911 ;
  assign n14913 = ~n14861 & ~n14912 ;
  assign n14914 = ~n14911 & ~n14912 ;
  assign n14915 = ~n14913 & ~n14914 ;
  assign n14916 = x75 & n9433 ;
  assign n14917 = x73 & n9915 ;
  assign n14918 = x74 & n9428 ;
  assign n14919 = ~n14917 & ~n14918 ;
  assign n14920 = ~n14916 & n14919 ;
  assign n14921 = n1150 & n9436 ;
  assign n14922 = n14920 & ~n14921 ;
  assign n14923 = x38 & ~n14922 ;
  assign n14924 = x38 & ~n14923 ;
  assign n14925 = ~n14922 & ~n14923 ;
  assign n14926 = ~n14924 & ~n14925 ;
  assign n14927 = n14915 & n14926 ;
  assign n14928 = ~n14915 & ~n14926 ;
  assign n14929 = ~n14927 & ~n14928 ;
  assign n14930 = ~n14287 & n14929 ;
  assign n14931 = n14287 & ~n14929 ;
  assign n14932 = ~n14930 & ~n14931 ;
  assign n14933 = x78 & n8006 ;
  assign n14934 = x76 & n8474 ;
  assign n14935 = x77 & n8001 ;
  assign n14936 = ~n14934 & ~n14935 ;
  assign n14937 = ~n14933 & n14936 ;
  assign n14938 = n1624 & n8009 ;
  assign n14939 = n14937 & ~n14938 ;
  assign n14940 = x35 & ~n14939 ;
  assign n14941 = x35 & ~n14940 ;
  assign n14942 = ~n14939 & ~n14940 ;
  assign n14943 = ~n14941 & ~n14942 ;
  assign n14944 = n14932 & ~n14943 ;
  assign n14945 = n14932 & ~n14944 ;
  assign n14946 = ~n14943 & ~n14944 ;
  assign n14947 = ~n14945 & ~n14946 ;
  assign n14948 = ~n14860 & ~n14947 ;
  assign n14949 = n14860 & n14947 ;
  assign n14950 = ~n14948 & ~n14949 ;
  assign n14951 = ~n14859 & n14950 ;
  assign n14952 = ~n14859 & ~n14951 ;
  assign n14953 = n14950 & ~n14951 ;
  assign n14954 = ~n14952 & ~n14953 ;
  assign n14955 = ~n14848 & ~n14954 ;
  assign n14956 = ~n14848 & ~n14955 ;
  assign n14957 = ~n14954 & ~n14955 ;
  assign n14958 = ~n14956 & ~n14957 ;
  assign n14959 = x84 & n5560 ;
  assign n14960 = x82 & n5943 ;
  assign n14961 = x83 & n5555 ;
  assign n14962 = ~n14960 & ~n14961 ;
  assign n14963 = ~n14959 & n14962 ;
  assign n14964 = n3114 & n5563 ;
  assign n14965 = n14963 & ~n14964 ;
  assign n14966 = x29 & ~n14965 ;
  assign n14967 = x29 & ~n14966 ;
  assign n14968 = ~n14965 & ~n14966 ;
  assign n14969 = ~n14967 & ~n14968 ;
  assign n14970 = ~n14958 & ~n14969 ;
  assign n14971 = ~n14958 & ~n14970 ;
  assign n14972 = ~n14969 & ~n14970 ;
  assign n14973 = ~n14971 & ~n14972 ;
  assign n14974 = ~n14338 & ~n14344 ;
  assign n14975 = n14973 & n14974 ;
  assign n14976 = ~n14973 & ~n14974 ;
  assign n14977 = ~n14975 & ~n14976 ;
  assign n14978 = x87 & n4531 ;
  assign n14979 = x85 & n4847 ;
  assign n14980 = x86 & n4526 ;
  assign n14981 = ~n14979 & ~n14980 ;
  assign n14982 = ~n14978 & n14981 ;
  assign n14983 = n3991 & n4534 ;
  assign n14984 = n14982 & ~n14983 ;
  assign n14985 = x26 & ~n14984 ;
  assign n14986 = x26 & ~n14985 ;
  assign n14987 = ~n14984 & ~n14985 ;
  assign n14988 = ~n14986 & ~n14987 ;
  assign n14989 = n14977 & ~n14988 ;
  assign n14990 = ~n14977 & n14988 ;
  assign n14991 = ~n14847 & ~n14990 ;
  assign n14992 = ~n14989 & n14991 ;
  assign n14993 = ~n14847 & ~n14992 ;
  assign n14994 = ~n14989 & ~n14992 ;
  assign n14995 = ~n14990 & n14994 ;
  assign n14996 = ~n14993 & ~n14995 ;
  assign n14997 = x90 & n3589 ;
  assign n14998 = x88 & n3878 ;
  assign n14999 = x89 & n3584 ;
  assign n15000 = ~n14998 & ~n14999 ;
  assign n15001 = ~n14997 & n15000 ;
  assign n15002 = n3592 & n4986 ;
  assign n15003 = n15001 & ~n15002 ;
  assign n15004 = x23 & ~n15003 ;
  assign n15005 = x23 & ~n15004 ;
  assign n15006 = ~n15003 & ~n15004 ;
  assign n15007 = ~n15005 & ~n15006 ;
  assign n15008 = n14996 & n15007 ;
  assign n15009 = ~n14996 & ~n15007 ;
  assign n15010 = ~n15008 & ~n15009 ;
  assign n15011 = ~n14846 & n15010 ;
  assign n15012 = n14846 & ~n15010 ;
  assign n15013 = ~n15011 & ~n15012 ;
  assign n15014 = n14845 & ~n15013 ;
  assign n15015 = ~n14845 & n15013 ;
  assign n15016 = ~n15014 & ~n15015 ;
  assign n15017 = ~n14834 & n15016 ;
  assign n15018 = n14834 & ~n15016 ;
  assign n15019 = ~n15017 & ~n15018 ;
  assign n15020 = n14833 & ~n15019 ;
  assign n15021 = ~n14833 & n15019 ;
  assign n15022 = ~n15020 & ~n15021 ;
  assign n15023 = ~n14822 & n15022 ;
  assign n15024 = n14822 & ~n15022 ;
  assign n15025 = ~n15023 & ~n15024 ;
  assign n15026 = x99 & n1434 ;
  assign n15027 = x97 & n1646 ;
  assign n15028 = x98 & n1429 ;
  assign n15029 = ~n15027 & ~n15028 ;
  assign n15030 = ~n15026 & n15029 ;
  assign n15031 = n1437 & n8660 ;
  assign n15032 = n15030 & ~n15031 ;
  assign n15033 = x14 & ~n15032 ;
  assign n15034 = x14 & ~n15033 ;
  assign n15035 = ~n15032 & ~n15033 ;
  assign n15036 = ~n15034 & ~n15035 ;
  assign n15037 = n15025 & ~n15036 ;
  assign n15038 = n15025 & ~n15037 ;
  assign n15039 = ~n15036 & ~n15037 ;
  assign n15040 = ~n15038 & ~n15039 ;
  assign n15041 = ~n14420 & ~n14427 ;
  assign n15042 = n15040 & n15041 ;
  assign n15043 = ~n15040 & ~n15041 ;
  assign n15044 = ~n15042 & ~n15043 ;
  assign n15045 = x102 & n945 ;
  assign n15046 = x100 & n1099 ;
  assign n15047 = x101 & n940 ;
  assign n15048 = ~n15046 & ~n15047 ;
  assign n15049 = ~n15045 & n15048 ;
  assign n15050 = n948 & n10092 ;
  assign n15051 = n15049 & ~n15050 ;
  assign n15052 = x11 & ~n15051 ;
  assign n15053 = x11 & ~n15052 ;
  assign n15054 = ~n15051 & ~n15052 ;
  assign n15055 = ~n15053 & ~n15054 ;
  assign n15056 = n15044 & ~n15055 ;
  assign n15057 = n15044 & ~n15056 ;
  assign n15058 = ~n15055 & ~n15056 ;
  assign n15059 = ~n15057 & ~n15058 ;
  assign n15060 = ~n14440 & ~n14446 ;
  assign n15061 = n15059 & n15060 ;
  assign n15062 = ~n15059 & ~n15060 ;
  assign n15063 = ~n15061 & ~n15062 ;
  assign n15064 = x105 & n574 ;
  assign n15065 = x103 & n673 ;
  assign n15066 = x104 & n569 ;
  assign n15067 = ~n15065 & ~n15066 ;
  assign n15068 = ~n15064 & n15067 ;
  assign n15069 = n577 & n11648 ;
  assign n15070 = n15068 & ~n15069 ;
  assign n15071 = x8 & ~n15070 ;
  assign n15072 = x8 & ~n15071 ;
  assign n15073 = ~n15070 & ~n15071 ;
  assign n15074 = ~n15072 & ~n15073 ;
  assign n15075 = n15063 & ~n15074 ;
  assign n15076 = ~n15063 & n15074 ;
  assign n15077 = ~n14464 & ~n15076 ;
  assign n15078 = ~n15075 & n15077 ;
  assign n15079 = ~n14464 & ~n15078 ;
  assign n15080 = ~n15075 & ~n15078 ;
  assign n15081 = ~n15076 & n15080 ;
  assign n15082 = ~n15079 & ~n15081 ;
  assign n15083 = x108 & n293 ;
  assign n15084 = x106 & n373 ;
  assign n15085 = x107 & n288 ;
  assign n15086 = ~n15084 & ~n15085 ;
  assign n15087 = ~n15083 & n15086 ;
  assign n15088 = n296 & n13323 ;
  assign n15089 = n15087 & ~n15088 ;
  assign n15090 = x5 & ~n15089 ;
  assign n15091 = x5 & ~n15090 ;
  assign n15092 = ~n15089 & ~n15090 ;
  assign n15093 = ~n15091 & ~n15092 ;
  assign n15094 = n15082 & n15093 ;
  assign n15095 = ~n15082 & ~n15093 ;
  assign n15096 = ~n15094 & ~n15095 ;
  assign n15097 = ~n14821 & n15096 ;
  assign n15098 = n14821 & ~n15096 ;
  assign n15099 = ~n15097 & ~n15098 ;
  assign n15100 = x111 & n146 ;
  assign n15101 = x109 & n182 ;
  assign n15102 = x110 & n141 ;
  assign n15103 = ~n15101 & ~n15102 ;
  assign n15104 = ~n15100 & n15103 ;
  assign n15105 = ~n14493 & ~n14495 ;
  assign n15106 = ~x110 & ~x111 ;
  assign n15107 = x110 & x111 ;
  assign n15108 = ~n15106 & ~n15107 ;
  assign n15109 = ~n15105 & n15108 ;
  assign n15110 = n15105 & ~n15108 ;
  assign n15111 = ~n15109 & ~n15110 ;
  assign n15112 = n149 & n15111 ;
  assign n15113 = n15104 & ~n15112 ;
  assign n15114 = x2 & ~n15113 ;
  assign n15115 = x2 & ~n15114 ;
  assign n15116 = ~n15113 & ~n15114 ;
  assign n15117 = ~n15115 & ~n15116 ;
  assign n15118 = n15099 & ~n15117 ;
  assign n15119 = n15099 & ~n15118 ;
  assign n15120 = ~n15117 & ~n15118 ;
  assign n15121 = ~n15119 & ~n15120 ;
  assign n15122 = ~n14504 & ~n14509 ;
  assign n15123 = ~n15121 & ~n15122 ;
  assign n15124 = n15121 & n15122 ;
  assign n15125 = ~n15123 & ~n15124 ;
  assign n15427 = n15125 & x175 ;
  assign n15126 = ~n14786 & ~n14792 ;
  assign n15127 = ~n14712 & ~n14714 ;
  assign n15128 = ~x96 & n2093 ;
  assign n15129 = ~x94 & n2275 ;
  assign n15130 = ~x95 & n2088 ;
  assign n15131 = ~n15129 & ~n15130 ;
  assign n15132 = ~n15128 & n15131 ;
  assign n15133 = n2096 & n7531 ;
  assign n15134 = n15132 & ~n15133 ;
  assign n15135 = ~x17 & ~n15134 ;
  assign n15136 = ~x17 & ~n15135 ;
  assign n15137 = ~n15134 & ~n15135 ;
  assign n15138 = ~n15136 & ~n15137 ;
  assign n15139 = ~n14692 & ~n14696 ;
  assign n15140 = ~x93 & n2751 ;
  assign n15141 = ~x91 & n3020 ;
  assign n15142 = ~x92 & n2746 ;
  assign n15143 = ~n15141 & ~n15142 ;
  assign n15144 = ~n15140 & n15143 ;
  assign n15145 = n2754 & n6285 ;
  assign n15146 = n15144 & ~n15145 ;
  assign n15147 = ~x20 & ~n15146 ;
  assign n15148 = ~x20 & ~n15147 ;
  assign n15149 = ~n15146 & ~n15147 ;
  assign n15150 = ~n15148 & ~n15149 ;
  assign n15151 = ~n14684 & ~n14689 ;
  assign n15152 = ~n14665 & ~n14671 ;
  assign n15153 = ~n14626 & ~n14633 ;
  assign n15154 = ~x81 & n6725 ;
  assign n15155 = ~x79 & n7129 ;
  assign n15156 = ~x80 & n6720 ;
  assign n15157 = ~n15155 & ~n15156 ;
  assign n15158 = ~n15154 & n15157 ;
  assign n15159 = n2460 & n6728 ;
  assign n15160 = n15158 & ~n15159 ;
  assign n15161 = ~x32 & ~n15160 ;
  assign n15162 = ~x32 & ~n15161 ;
  assign n15163 = ~n15160 & ~n15161 ;
  assign n15164 = ~n15162 & ~n15163 ;
  assign n15165 = ~n14610 & ~n14612 ;
  assign n15166 = ~n14571 & ~n14577 ;
  assign n15167 = ~x72 & n10905 ;
  assign n15168 = ~x70 & n11466 ;
  assign n15169 = ~x71 & n10900 ;
  assign n15170 = ~n15168 & ~n15169 ;
  assign n15171 = ~n15167 & n15170 ;
  assign n15172 = n773 & n10908 ;
  assign n15173 = n15171 & ~n15172 ;
  assign n15174 = ~x41 & ~n15173 ;
  assign n15175 = ~x41 & ~n15174 ;
  assign n15176 = ~n15173 & ~n15174 ;
  assign n15177 = ~n15175 & ~n15176 ;
  assign n15178 = ~n14555 & ~n14557 ;
  assign n15179 = ~x66 & n14233 ;
  assign n15180 = ~x64 & n14876 ;
  assign n15181 = ~x65 & n14228 ;
  assign n15182 = ~n15180 & ~n15181 ;
  assign n15183 = ~n15179 & n15182 ;
  assign n15184 = n214 & n14236 ;
  assign n15185 = n15183 & ~n15184 ;
  assign n15186 = ~x47 & ~n15185 ;
  assign n15187 = ~x47 & ~n15186 ;
  assign n15188 = ~n15185 & ~n15186 ;
  assign n15189 = ~n15187 & ~n15188 ;
  assign n15190 = ~n14551 & n15189 ;
  assign n15191 = n14551 & ~n15189 ;
  assign n15192 = ~n15190 & ~n15191 ;
  assign n15193 = ~x69 & n12506 ;
  assign n15194 = ~x67 & n13131 ;
  assign n15195 = ~x68 & n12501 ;
  assign n15196 = ~n15194 & ~n15195 ;
  assign n15197 = ~n15193 & n15196 ;
  assign n15198 = n435 & n12509 ;
  assign n15199 = n15197 & ~n15198 ;
  assign n15200 = ~x44 & ~n15199 ;
  assign n15201 = ~x44 & ~n15200 ;
  assign n15202 = ~n15199 & ~n15200 ;
  assign n15203 = ~n15201 & ~n15202 ;
  assign n15204 = n15192 & ~n15203 ;
  assign n15205 = n15192 & ~n15204 ;
  assign n15206 = ~n15203 & ~n15204 ;
  assign n15207 = ~n15205 & ~n15206 ;
  assign n15208 = ~n15178 & ~n15207 ;
  assign n15209 = n15178 & n15207 ;
  assign n15210 = ~n15208 & ~n15209 ;
  assign n15211 = ~n15177 & n15210 ;
  assign n15212 = ~n15177 & ~n15211 ;
  assign n15213 = n15210 & ~n15211 ;
  assign n15214 = ~n15212 & ~n15213 ;
  assign n15215 = ~n15166 & ~n15214 ;
  assign n15216 = ~n15166 & ~n15215 ;
  assign n15217 = ~n15214 & ~n15215 ;
  assign n15218 = ~n15216 & ~n15217 ;
  assign n15219 = ~x75 & n9433 ;
  assign n15220 = ~x73 & n9915 ;
  assign n15221 = ~x74 & n9428 ;
  assign n15222 = ~n15220 & ~n15221 ;
  assign n15223 = ~n15219 & n15222 ;
  assign n15224 = n1225 & n9436 ;
  assign n15225 = n15223 & ~n15224 ;
  assign n15226 = ~x38 & ~n15225 ;
  assign n15227 = ~x38 & ~n15226 ;
  assign n15228 = ~n15225 & ~n15226 ;
  assign n15229 = ~n15227 & ~n15228 ;
  assign n15230 = n15218 & n15229 ;
  assign n15231 = ~n15218 & ~n15229 ;
  assign n15232 = ~n15230 & ~n15231 ;
  assign n15233 = ~n14595 & n15232 ;
  assign n15234 = n14595 & ~n15232 ;
  assign n15235 = ~n15233 & ~n15234 ;
  assign n15236 = ~x78 & n8006 ;
  assign n15237 = ~x76 & n8474 ;
  assign n15238 = ~x77 & n8001 ;
  assign n15239 = ~n15237 & ~n15238 ;
  assign n15240 = ~n15236 & n15239 ;
  assign n15241 = n1718 & n8009 ;
  assign n15242 = n15240 & ~n15241 ;
  assign n15243 = ~x35 & ~n15242 ;
  assign n15244 = ~x35 & ~n15243 ;
  assign n15245 = ~n15242 & ~n15243 ;
  assign n15246 = ~n15244 & ~n15245 ;
  assign n15247 = n15235 & ~n15246 ;
  assign n15248 = n15235 & ~n15247 ;
  assign n15249 = ~n15246 & ~n15247 ;
  assign n15250 = ~n15248 & ~n15249 ;
  assign n15251 = ~n15165 & ~n15250 ;
  assign n15252 = n15165 & n15250 ;
  assign n15253 = ~n15251 & ~n15252 ;
  assign n15254 = ~n15164 & n15253 ;
  assign n15255 = ~n15164 & ~n15254 ;
  assign n15256 = n15253 & ~n15254 ;
  assign n15257 = ~n15255 & ~n15256 ;
  assign n15258 = ~n15153 & ~n15257 ;
  assign n15259 = ~n15153 & ~n15258 ;
  assign n15260 = ~n15257 & ~n15258 ;
  assign n15261 = ~n15259 & ~n15260 ;
  assign n15262 = ~x84 & n5560 ;
  assign n15263 = ~x82 & n5943 ;
  assign n15264 = ~x83 & n5555 ;
  assign n15265 = ~n15263 & ~n15264 ;
  assign n15266 = ~n15262 & n15265 ;
  assign n15267 = n3247 & n5563 ;
  assign n15268 = n15266 & ~n15267 ;
  assign n15269 = ~x29 & ~n15268 ;
  assign n15270 = ~x29 & ~n15269 ;
  assign n15271 = ~n15268 & ~n15269 ;
  assign n15272 = ~n15270 & ~n15271 ;
  assign n15273 = ~n15261 & ~n15272 ;
  assign n15274 = ~n15261 & ~n15273 ;
  assign n15275 = ~n15272 & ~n15273 ;
  assign n15276 = ~n15274 & ~n15275 ;
  assign n15277 = ~n14646 & ~n14652 ;
  assign n15278 = n15276 & n15277 ;
  assign n15279 = ~n15276 & ~n15277 ;
  assign n15280 = ~n15278 & ~n15279 ;
  assign n15281 = ~x87 & n4531 ;
  assign n15282 = ~x85 & n4847 ;
  assign n15283 = ~x86 & n4526 ;
  assign n15284 = ~n15282 & ~n15283 ;
  assign n15285 = ~n15281 & n15284 ;
  assign n15286 = n4143 & n4534 ;
  assign n15287 = n15285 & ~n15286 ;
  assign n15288 = ~x26 & ~n15287 ;
  assign n15289 = ~x26 & ~n15288 ;
  assign n15290 = ~n15287 & ~n15288 ;
  assign n15291 = ~n15289 & ~n15290 ;
  assign n15292 = n15280 & ~n15291 ;
  assign n15293 = ~n15280 & n15291 ;
  assign n15294 = ~n15152 & ~n15293 ;
  assign n15295 = ~n15292 & n15294 ;
  assign n15296 = ~n15152 & ~n15295 ;
  assign n15297 = ~n15292 & ~n15295 ;
  assign n15298 = ~n15293 & n15297 ;
  assign n15299 = ~n15296 & ~n15298 ;
  assign n15300 = ~x90 & n3589 ;
  assign n15301 = ~x88 & n3878 ;
  assign n15302 = ~x89 & n3584 ;
  assign n15303 = ~n15301 & ~n15302 ;
  assign n15304 = ~n15300 & n15303 ;
  assign n15305 = n3592 & n5155 ;
  assign n15306 = n15304 & ~n15305 ;
  assign n15307 = ~x23 & ~n15306 ;
  assign n15308 = ~x23 & ~n15307 ;
  assign n15309 = ~n15306 & ~n15307 ;
  assign n15310 = ~n15308 & ~n15309 ;
  assign n15311 = n15299 & n15310 ;
  assign n15312 = ~n15299 & ~n15310 ;
  assign n15313 = ~n15311 & ~n15312 ;
  assign n15314 = ~n15151 & n15313 ;
  assign n15315 = n15151 & ~n15313 ;
  assign n15316 = ~n15314 & ~n15315 ;
  assign n15317 = n15150 & ~n15316 ;
  assign n15318 = ~n15150 & n15316 ;
  assign n15319 = ~n15317 & ~n15318 ;
  assign n15320 = ~n15139 & n15319 ;
  assign n15321 = n15139 & ~n15319 ;
  assign n15322 = ~n15320 & ~n15321 ;
  assign n15323 = n15138 & ~n15322 ;
  assign n15324 = ~n15138 & n15322 ;
  assign n15325 = ~n15323 & ~n15324 ;
  assign n15326 = ~n15127 & n15325 ;
  assign n15327 = n15127 & ~n15325 ;
  assign n15328 = ~n15326 & ~n15327 ;
  assign n15329 = ~x99 & n1434 ;
  assign n15330 = ~x97 & n1646 ;
  assign n15331 = ~x98 & n1429 ;
  assign n15332 = ~n15330 & ~n15331 ;
  assign n15333 = ~n15329 & n15332 ;
  assign n15334 = n1437 & n8885 ;
  assign n15335 = n15333 & ~n15334 ;
  assign n15336 = ~x14 & ~n15335 ;
  assign n15337 = ~x14 & ~n15336 ;
  assign n15338 = ~n15335 & ~n15336 ;
  assign n15339 = ~n15337 & ~n15338 ;
  assign n15340 = n15328 & ~n15339 ;
  assign n15341 = n15328 & ~n15340 ;
  assign n15342 = ~n15339 & ~n15340 ;
  assign n15343 = ~n15341 & ~n15342 ;
  assign n15344 = ~n14728 & ~n14735 ;
  assign n15345 = n15343 & n15344 ;
  assign n15346 = ~n15343 & ~n15344 ;
  assign n15347 = ~n15345 & ~n15346 ;
  assign n15348 = ~x102 & n945 ;
  assign n15349 = ~x100 & n1099 ;
  assign n15350 = ~x101 & n940 ;
  assign n15351 = ~n15349 & ~n15350 ;
  assign n15352 = ~n15348 & n15351 ;
  assign n15353 = n948 & n10333 ;
  assign n15354 = n15352 & ~n15353 ;
  assign n15355 = ~x11 & ~n15354 ;
  assign n15356 = ~x11 & ~n15355 ;
  assign n15357 = ~n15354 & ~n15355 ;
  assign n15358 = ~n15356 & ~n15357 ;
  assign n15359 = n15347 & ~n15358 ;
  assign n15360 = n15347 & ~n15359 ;
  assign n15361 = ~n15358 & ~n15359 ;
  assign n15362 = ~n15360 & ~n15361 ;
  assign n15363 = ~n14748 & ~n14754 ;
  assign n15364 = n15362 & n15363 ;
  assign n15365 = ~n15362 & ~n15363 ;
  assign n15366 = ~n15364 & ~n15365 ;
  assign n15367 = ~x105 & n574 ;
  assign n15368 = ~x103 & n673 ;
  assign n15369 = ~x104 & n569 ;
  assign n15370 = ~n15368 & ~n15369 ;
  assign n15371 = ~n15367 & n15370 ;
  assign n15372 = n577 & n11907 ;
  assign n15373 = n15371 & ~n15372 ;
  assign n15374 = ~x8 & ~n15373 ;
  assign n15375 = ~x8 & ~n15374 ;
  assign n15376 = ~n15373 & ~n15374 ;
  assign n15377 = ~n15375 & ~n15376 ;
  assign n15378 = n15366 & ~n15377 ;
  assign n15379 = ~n15366 & n15377 ;
  assign n15380 = ~n14772 & ~n15379 ;
  assign n15381 = ~n15378 & n15380 ;
  assign n15382 = ~n14772 & ~n15381 ;
  assign n15383 = ~n15378 & ~n15381 ;
  assign n15384 = ~n15379 & n15383 ;
  assign n15385 = ~n15382 & ~n15384 ;
  assign n15386 = ~x108 & n293 ;
  assign n15387 = ~x106 & n373 ;
  assign n15388 = ~x107 & n288 ;
  assign n15389 = ~n15387 & ~n15388 ;
  assign n15390 = ~n15386 & n15389 ;
  assign n15391 = n296 & n13601 ;
  assign n15392 = n15390 & ~n15391 ;
  assign n15393 = ~x5 & ~n15392 ;
  assign n15394 = ~x5 & ~n15393 ;
  assign n15395 = ~n15392 & ~n15393 ;
  assign n15396 = ~n15394 & ~n15395 ;
  assign n15397 = n15385 & n15396 ;
  assign n15398 = ~n15385 & ~n15396 ;
  assign n15399 = ~n15397 & ~n15398 ;
  assign n15400 = ~n15126 & n15399 ;
  assign n15401 = n15126 & ~n15399 ;
  assign n15402 = ~n15400 & ~n15401 ;
  assign n15403 = ~x111 & n164 ;
  assign n15404 = ~x109 & n205 ;
  assign n15405 = ~x110 & n162 ;
  assign n15406 = ~n15404 & ~n15405 ;
  assign n15407 = ~n15403 & n15406 ;
  assign n15408 = ~n14492 & ~n14800 ;
  assign n15409 = n15108 & ~n15408 ;
  assign n15410 = ~n15108 & n15408 ;
  assign n15411 = ~n15409 & ~n15410 ;
  assign n15412 = n167 & n15411 ;
  assign n15413 = n15407 & ~n15412 ;
  assign n15414 = ~x2 & ~n15413 ;
  assign n15415 = ~x2 & ~n15414 ;
  assign n15416 = ~n15413 & ~n15414 ;
  assign n15417 = ~n15415 & ~n15416 ;
  assign n15418 = n15402 & ~n15417 ;
  assign n15419 = n15402 & ~n15418 ;
  assign n15420 = ~n15417 & ~n15418 ;
  assign n15421 = ~n15419 & ~n15420 ;
  assign n15422 = ~n14809 & ~n14814 ;
  assign n15423 = ~n15421 & ~n15422 ;
  assign n15424 = n15421 & n15422 ;
  assign n15425 = ~n15423 & ~n15424 ;
  assign n15428 = ~n15425 & ~x175 ;
  assign n15429 = ~n15427 & ~n15428 ;
  assign n15430 = ~n15118 & ~n15123 ;
  assign n15431 = x112 & n146 ;
  assign n15432 = x110 & n182 ;
  assign n15433 = x111 & n141 ;
  assign n15434 = ~n15432 & ~n15433 ;
  assign n15435 = ~n15431 & n15434 ;
  assign n15436 = ~n15107 & ~n15109 ;
  assign n15437 = ~x111 & ~x112 ;
  assign n15438 = x111 & x112 ;
  assign n15439 = ~n15437 & ~n15438 ;
  assign n15440 = ~n15436 & n15439 ;
  assign n15441 = n15436 & ~n15439 ;
  assign n15442 = ~n15440 & ~n15441 ;
  assign n15443 = n149 & n15442 ;
  assign n15444 = n15435 & ~n15443 ;
  assign n15445 = x2 & ~n15444 ;
  assign n15446 = x2 & ~n15445 ;
  assign n15447 = ~n15444 & ~n15445 ;
  assign n15448 = ~n15446 & ~n15447 ;
  assign n15449 = ~n15095 & ~n15097 ;
  assign n15450 = ~n15037 & ~n15043 ;
  assign n15451 = ~n15021 & ~n15023 ;
  assign n15452 = ~n15015 & ~n15017 ;
  assign n15453 = ~n15009 & ~n15011 ;
  assign n15454 = ~n14944 & ~n14948 ;
  assign n15455 = x79 & n8006 ;
  assign n15456 = x77 & n8474 ;
  assign n15457 = x78 & n8001 ;
  assign n15458 = ~n15456 & ~n15457 ;
  assign n15459 = ~n15455 & n15458 ;
  assign n15460 = n1817 & n8009 ;
  assign n15461 = n15459 & ~n15460 ;
  assign n15462 = x35 & ~n15461 ;
  assign n15463 = x35 & ~n15462 ;
  assign n15464 = ~n15461 & ~n15462 ;
  assign n15465 = ~n15463 & ~n15464 ;
  assign n15466 = ~n14928 & ~n14930 ;
  assign n15467 = x76 & n9433 ;
  assign n15468 = x74 & n9915 ;
  assign n15469 = x75 & n9428 ;
  assign n15470 = ~n15468 & ~n15469 ;
  assign n15471 = ~n15467 & n15470 ;
  assign n15472 = n1311 & n9436 ;
  assign n15473 = n15471 & ~n15472 ;
  assign n15474 = x38 & ~n15473 ;
  assign n15475 = x38 & ~n15474 ;
  assign n15476 = ~n15473 & ~n15474 ;
  assign n15477 = ~n15475 & ~n15476 ;
  assign n15478 = ~n14908 & ~n14912 ;
  assign n15479 = x47 & ~x48 ;
  assign n15480 = ~x47 & x48 ;
  assign n15481 = ~n15479 & ~n15480 ;
  assign n15482 = x64 & ~n15481 ;
  assign n15483 = ~n14888 & n15482 ;
  assign n15484 = n14888 & ~n15482 ;
  assign n15485 = ~n15483 & ~n15484 ;
  assign n15486 = x67 & n14233 ;
  assign n15487 = x65 & n14876 ;
  assign n15488 = x66 & n14228 ;
  assign n15489 = ~n15487 & ~n15488 ;
  assign n15490 = ~n15486 & n15489 ;
  assign n15491 = n240 & n14236 ;
  assign n15492 = n15490 & ~n15491 ;
  assign n15493 = x47 & ~n15492 ;
  assign n15494 = x47 & ~n15493 ;
  assign n15495 = ~n15492 & ~n15493 ;
  assign n15496 = ~n15494 & ~n15495 ;
  assign n15497 = ~n15485 & ~n15496 ;
  assign n15498 = n15485 & n15496 ;
  assign n15499 = ~n15497 & ~n15498 ;
  assign n15500 = x70 & n12506 ;
  assign n15501 = x68 & n13131 ;
  assign n15502 = x69 & n12501 ;
  assign n15503 = ~n15501 & ~n15502 ;
  assign n15504 = ~n15500 & n15503 ;
  assign n15505 = n488 & n12509 ;
  assign n15506 = n15504 & ~n15505 ;
  assign n15507 = x44 & ~n15506 ;
  assign n15508 = x44 & ~n15507 ;
  assign n15509 = ~n15506 & ~n15507 ;
  assign n15510 = ~n15508 & ~n15509 ;
  assign n15511 = n15499 & ~n15510 ;
  assign n15512 = n15499 & ~n15511 ;
  assign n15513 = ~n15510 & ~n15511 ;
  assign n15514 = ~n15512 & ~n15513 ;
  assign n15515 = ~n14901 & ~n14905 ;
  assign n15516 = n15514 & n15515 ;
  assign n15517 = ~n15514 & ~n15515 ;
  assign n15518 = ~n15516 & ~n15517 ;
  assign n15519 = x73 & n10905 ;
  assign n15520 = x71 & n11466 ;
  assign n15521 = x72 & n10900 ;
  assign n15522 = ~n15520 & ~n15521 ;
  assign n15523 = ~n15519 & n15522 ;
  assign n15524 = n843 & n10908 ;
  assign n15525 = n15523 & ~n15524 ;
  assign n15526 = x41 & ~n15525 ;
  assign n15527 = x41 & ~n15526 ;
  assign n15528 = ~n15525 & ~n15526 ;
  assign n15529 = ~n15527 & ~n15528 ;
  assign n15530 = ~n15518 & n15529 ;
  assign n15531 = n15518 & ~n15529 ;
  assign n15532 = ~n15530 & ~n15531 ;
  assign n15533 = ~n15478 & n15532 ;
  assign n15534 = n15478 & ~n15532 ;
  assign n15535 = ~n15533 & ~n15534 ;
  assign n15536 = ~n15477 & n15535 ;
  assign n15537 = ~n15477 & ~n15536 ;
  assign n15538 = n15535 & ~n15536 ;
  assign n15539 = ~n15537 & ~n15538 ;
  assign n15540 = ~n15466 & ~n15539 ;
  assign n15541 = n15466 & ~n15538 ;
  assign n15542 = ~n15537 & n15541 ;
  assign n15543 = ~n15540 & ~n15542 ;
  assign n15544 = ~n15465 & n15543 ;
  assign n15545 = n15465 & ~n15543 ;
  assign n15546 = ~n15544 & ~n15545 ;
  assign n15547 = ~n15454 & n15546 ;
  assign n15548 = n15454 & ~n15546 ;
  assign n15549 = ~n15547 & ~n15548 ;
  assign n15550 = x82 & n6725 ;
  assign n15551 = x80 & n7129 ;
  assign n15552 = x81 & n6720 ;
  assign n15553 = ~n15551 & ~n15552 ;
  assign n15554 = ~n15550 & n15553 ;
  assign n15555 = n2584 & n6728 ;
  assign n15556 = n15554 & ~n15555 ;
  assign n15557 = x32 & ~n15556 ;
  assign n15558 = x32 & ~n15557 ;
  assign n15559 = ~n15556 & ~n15557 ;
  assign n15560 = ~n15558 & ~n15559 ;
  assign n15561 = n15549 & ~n15560 ;
  assign n15562 = n15549 & ~n15561 ;
  assign n15563 = ~n15560 & ~n15561 ;
  assign n15564 = ~n15562 & ~n15563 ;
  assign n15565 = ~n14951 & ~n14955 ;
  assign n15566 = n15564 & n15565 ;
  assign n15567 = ~n15564 & ~n15565 ;
  assign n15568 = ~n15566 & ~n15567 ;
  assign n15569 = x85 & n5560 ;
  assign n15570 = x83 & n5943 ;
  assign n15571 = x84 & n5555 ;
  assign n15572 = ~n15570 & ~n15571 ;
  assign n15573 = ~n15569 & n15572 ;
  assign n15574 = n3389 & n5563 ;
  assign n15575 = n15573 & ~n15574 ;
  assign n15576 = x29 & ~n15575 ;
  assign n15577 = x29 & ~n15576 ;
  assign n15578 = ~n15575 & ~n15576 ;
  assign n15579 = ~n15577 & ~n15578 ;
  assign n15580 = n15568 & ~n15579 ;
  assign n15581 = n15568 & ~n15580 ;
  assign n15582 = ~n15579 & ~n15580 ;
  assign n15583 = ~n15581 & ~n15582 ;
  assign n15584 = ~n14970 & ~n14976 ;
  assign n15585 = n15583 & n15584 ;
  assign n15586 = ~n15583 & ~n15584 ;
  assign n15587 = ~n15585 & ~n15586 ;
  assign n15588 = x88 & n4531 ;
  assign n15589 = x86 & n4847 ;
  assign n15590 = x87 & n4526 ;
  assign n15591 = ~n15589 & ~n15590 ;
  assign n15592 = ~n15588 & n15591 ;
  assign n15593 = n4305 & n4534 ;
  assign n15594 = n15592 & ~n15593 ;
  assign n15595 = x26 & ~n15594 ;
  assign n15596 = x26 & ~n15595 ;
  assign n15597 = ~n15594 & ~n15595 ;
  assign n15598 = ~n15596 & ~n15597 ;
  assign n15599 = ~n15587 & n15598 ;
  assign n15600 = n15587 & ~n15598 ;
  assign n15601 = ~n15599 & ~n15600 ;
  assign n15602 = ~n14994 & n15601 ;
  assign n15603 = n14994 & ~n15601 ;
  assign n15604 = ~n15602 & ~n15603 ;
  assign n15605 = x91 & n3589 ;
  assign n15606 = x89 & n3878 ;
  assign n15607 = x90 & n3584 ;
  assign n15608 = ~n15606 & ~n15607 ;
  assign n15609 = ~n15605 & n15608 ;
  assign n15610 = n3592 & n5336 ;
  assign n15611 = n15609 & ~n15610 ;
  assign n15612 = x23 & ~n15611 ;
  assign n15613 = x23 & ~n15612 ;
  assign n15614 = ~n15611 & ~n15612 ;
  assign n15615 = ~n15613 & ~n15614 ;
  assign n15616 = n15604 & ~n15615 ;
  assign n15617 = n15604 & ~n15616 ;
  assign n15618 = ~n15615 & ~n15616 ;
  assign n15619 = ~n15617 & ~n15618 ;
  assign n15620 = ~n15453 & n15619 ;
  assign n15621 = n15453 & ~n15619 ;
  assign n15622 = ~n15620 & ~n15621 ;
  assign n15623 = x94 & n2751 ;
  assign n15624 = x92 & n3020 ;
  assign n15625 = x93 & n2746 ;
  assign n15626 = ~n15624 & ~n15625 ;
  assign n15627 = ~n15623 & n15626 ;
  assign n15628 = n2754 & n6483 ;
  assign n15629 = n15627 & ~n15628 ;
  assign n15630 = x20 & ~n15629 ;
  assign n15631 = x20 & ~n15630 ;
  assign n15632 = ~n15629 & ~n15630 ;
  assign n15633 = ~n15631 & ~n15632 ;
  assign n15634 = ~n15622 & ~n15633 ;
  assign n15635 = n15622 & n15633 ;
  assign n15636 = ~n15634 & ~n15635 ;
  assign n15637 = ~n15452 & n15636 ;
  assign n15638 = n15452 & ~n15636 ;
  assign n15639 = ~n15637 & ~n15638 ;
  assign n15640 = x97 & n2093 ;
  assign n15641 = x95 & n2275 ;
  assign n15642 = x96 & n2088 ;
  assign n15643 = ~n15641 & ~n15642 ;
  assign n15644 = ~n15640 & n15643 ;
  assign n15645 = n2096 & n7745 ;
  assign n15646 = n15644 & ~n15645 ;
  assign n15647 = x17 & ~n15646 ;
  assign n15648 = x17 & ~n15647 ;
  assign n15649 = ~n15646 & ~n15647 ;
  assign n15650 = ~n15648 & ~n15649 ;
  assign n15651 = n15639 & ~n15650 ;
  assign n15652 = n15639 & ~n15651 ;
  assign n15653 = ~n15650 & ~n15651 ;
  assign n15654 = ~n15652 & ~n15653 ;
  assign n15655 = ~n15451 & n15654 ;
  assign n15656 = n15451 & ~n15654 ;
  assign n15657 = ~n15655 & ~n15656 ;
  assign n15658 = x100 & n1434 ;
  assign n15659 = x98 & n1646 ;
  assign n15660 = x99 & n1429 ;
  assign n15661 = ~n15659 & ~n15660 ;
  assign n15662 = ~n15658 & n15661 ;
  assign n15663 = n1437 & n9115 ;
  assign n15664 = n15662 & ~n15663 ;
  assign n15665 = x14 & ~n15664 ;
  assign n15666 = x14 & ~n15665 ;
  assign n15667 = ~n15664 & ~n15665 ;
  assign n15668 = ~n15666 & ~n15667 ;
  assign n15669 = ~n15657 & ~n15668 ;
  assign n15670 = n15657 & n15668 ;
  assign n15671 = ~n15669 & ~n15670 ;
  assign n15672 = n15450 & ~n15671 ;
  assign n15673 = ~n15450 & n15671 ;
  assign n15674 = ~n15672 & ~n15673 ;
  assign n15675 = x103 & n945 ;
  assign n15676 = x101 & n1099 ;
  assign n15677 = x102 & n940 ;
  assign n15678 = ~n15676 & ~n15677 ;
  assign n15679 = ~n15675 & n15678 ;
  assign n15680 = n948 & n10588 ;
  assign n15681 = n15679 & ~n15680 ;
  assign n15682 = x11 & ~n15681 ;
  assign n15683 = x11 & ~n15682 ;
  assign n15684 = ~n15681 & ~n15682 ;
  assign n15685 = ~n15683 & ~n15684 ;
  assign n15686 = n15674 & ~n15685 ;
  assign n15687 = n15674 & ~n15686 ;
  assign n15688 = ~n15685 & ~n15686 ;
  assign n15689 = ~n15687 & ~n15688 ;
  assign n15690 = ~n15056 & ~n15062 ;
  assign n15691 = n15689 & n15690 ;
  assign n15692 = ~n15689 & ~n15690 ;
  assign n15693 = ~n15691 & ~n15692 ;
  assign n15694 = x106 & n574 ;
  assign n15695 = x104 & n673 ;
  assign n15696 = x105 & n569 ;
  assign n15697 = ~n15695 & ~n15696 ;
  assign n15698 = ~n15694 & n15697 ;
  assign n15699 = n577 & n12181 ;
  assign n15700 = n15698 & ~n15699 ;
  assign n15701 = x8 & ~n15700 ;
  assign n15702 = x8 & ~n15701 ;
  assign n15703 = ~n15700 & ~n15701 ;
  assign n15704 = ~n15702 & ~n15703 ;
  assign n15705 = n15693 & ~n15704 ;
  assign n15706 = n15693 & ~n15705 ;
  assign n15707 = ~n15704 & ~n15705 ;
  assign n15708 = ~n15706 & ~n15707 ;
  assign n15709 = ~n15080 & n15708 ;
  assign n15710 = n15080 & ~n15708 ;
  assign n15711 = ~n15709 & ~n15710 ;
  assign n15712 = x109 & n293 ;
  assign n15713 = x107 & n373 ;
  assign n15714 = x108 & n288 ;
  assign n15715 = ~n15713 & ~n15714 ;
  assign n15716 = ~n15712 & n15715 ;
  assign n15717 = n296 & n13894 ;
  assign n15718 = n15716 & ~n15717 ;
  assign n15719 = x5 & ~n15718 ;
  assign n15720 = x5 & ~n15719 ;
  assign n15721 = ~n15718 & ~n15719 ;
  assign n15722 = ~n15720 & ~n15721 ;
  assign n15723 = ~n15711 & ~n15722 ;
  assign n15724 = n15711 & n15722 ;
  assign n15725 = ~n15723 & ~n15724 ;
  assign n15726 = ~n15449 & n15725 ;
  assign n15727 = n15449 & ~n15725 ;
  assign n15728 = ~n15726 & ~n15727 ;
  assign n15729 = n15448 & ~n15728 ;
  assign n15730 = ~n15448 & n15728 ;
  assign n15731 = ~n15729 & ~n15730 ;
  assign n15732 = ~n15430 & n15731 ;
  assign n15733 = n15430 & ~n15731 ;
  assign n15734 = ~n15732 & ~n15733 ;
  assign n16035 = n15734 & x176 ;
  assign n15735 = ~n15418 & ~n15423 ;
  assign n15736 = ~x112 & n164 ;
  assign n15737 = ~x110 & n205 ;
  assign n15738 = ~x111 & n162 ;
  assign n15739 = ~n15737 & ~n15738 ;
  assign n15740 = ~n15736 & n15739 ;
  assign n15741 = ~n15106 & ~n15409 ;
  assign n15742 = n15439 & ~n15741 ;
  assign n15743 = ~n15439 & n15741 ;
  assign n15744 = ~n15742 & ~n15743 ;
  assign n15745 = n167 & n15744 ;
  assign n15746 = n15740 & ~n15745 ;
  assign n15747 = ~x2 & ~n15746 ;
  assign n15748 = ~x2 & ~n15747 ;
  assign n15749 = ~n15746 & ~n15747 ;
  assign n15750 = ~n15748 & ~n15749 ;
  assign n15751 = ~n15398 & ~n15400 ;
  assign n15752 = ~n15340 & ~n15346 ;
  assign n15753 = ~n15324 & ~n15326 ;
  assign n15754 = ~n15318 & ~n15320 ;
  assign n15755 = ~n15312 & ~n15314 ;
  assign n15756 = ~n15247 & ~n15251 ;
  assign n15757 = ~x79 & n8006 ;
  assign n15758 = ~x77 & n8474 ;
  assign n15759 = ~x78 & n8001 ;
  assign n15760 = ~n15758 & ~n15759 ;
  assign n15761 = ~n15757 & n15760 ;
  assign n15762 = n1921 & n8009 ;
  assign n15763 = n15761 & ~n15762 ;
  assign n15764 = ~x35 & ~n15763 ;
  assign n15765 = ~x35 & ~n15764 ;
  assign n15766 = ~n15763 & ~n15764 ;
  assign n15767 = ~n15765 & ~n15766 ;
  assign n15768 = ~n15231 & ~n15233 ;
  assign n15769 = ~x76 & n9433 ;
  assign n15770 = ~x74 & n9915 ;
  assign n15771 = ~x75 & n9428 ;
  assign n15772 = ~n15770 & ~n15771 ;
  assign n15773 = ~n15769 & n15772 ;
  assign n15774 = n1390 & n9436 ;
  assign n15775 = n15773 & ~n15774 ;
  assign n15776 = ~x38 & ~n15775 ;
  assign n15777 = ~x38 & ~n15776 ;
  assign n15778 = ~n15775 & ~n15776 ;
  assign n15779 = ~n15777 & ~n15778 ;
  assign n15780 = ~n15211 & ~n15215 ;
  assign n15781 = ~x64 & ~n15481 ;
  assign n15782 = ~n15191 & n15781 ;
  assign n15783 = n15191 & ~n15781 ;
  assign n15784 = ~n15782 & ~n15783 ;
  assign n15785 = ~x67 & n14233 ;
  assign n15786 = ~x65 & n14876 ;
  assign n15787 = ~x66 & n14228 ;
  assign n15788 = ~n15786 & ~n15787 ;
  assign n15789 = ~n15785 & n15788 ;
  assign n15790 = n266 & n14236 ;
  assign n15791 = n15789 & ~n15790 ;
  assign n15792 = ~x47 & ~n15791 ;
  assign n15793 = ~x47 & ~n15792 ;
  assign n15794 = ~n15791 & ~n15792 ;
  assign n15795 = ~n15793 & ~n15794 ;
  assign n15796 = ~n15784 & ~n15795 ;
  assign n15797 = n15784 & n15795 ;
  assign n15798 = ~n15796 & ~n15797 ;
  assign n15799 = ~x70 & n12506 ;
  assign n15800 = ~x68 & n13131 ;
  assign n15801 = ~x69 & n12501 ;
  assign n15802 = ~n15800 & ~n15801 ;
  assign n15803 = ~n15799 & n15802 ;
  assign n15804 = n529 & n12509 ;
  assign n15805 = n15803 & ~n15804 ;
  assign n15806 = ~x44 & ~n15805 ;
  assign n15807 = ~x44 & ~n15806 ;
  assign n15808 = ~n15805 & ~n15806 ;
  assign n15809 = ~n15807 & ~n15808 ;
  assign n15810 = n15798 & ~n15809 ;
  assign n15811 = n15798 & ~n15810 ;
  assign n15812 = ~n15809 & ~n15810 ;
  assign n15813 = ~n15811 & ~n15812 ;
  assign n15814 = ~n15204 & ~n15208 ;
  assign n15815 = n15813 & n15814 ;
  assign n15816 = ~n15813 & ~n15814 ;
  assign n15817 = ~n15815 & ~n15816 ;
  assign n15818 = ~x73 & n10905 ;
  assign n15819 = ~x71 & n11466 ;
  assign n15820 = ~x72 & n10900 ;
  assign n15821 = ~n15819 & ~n15820 ;
  assign n15822 = ~n15818 & n15821 ;
  assign n15823 = n903 & n10908 ;
  assign n15824 = n15822 & ~n15823 ;
  assign n15825 = ~x41 & ~n15824 ;
  assign n15826 = ~x41 & ~n15825 ;
  assign n15827 = ~n15824 & ~n15825 ;
  assign n15828 = ~n15826 & ~n15827 ;
  assign n15829 = ~n15817 & n15828 ;
  assign n15830 = n15817 & ~n15828 ;
  assign n15831 = ~n15829 & ~n15830 ;
  assign n15832 = ~n15780 & n15831 ;
  assign n15833 = n15780 & ~n15831 ;
  assign n15834 = ~n15832 & ~n15833 ;
  assign n15835 = ~n15779 & n15834 ;
  assign n15836 = ~n15779 & ~n15835 ;
  assign n15837 = n15834 & ~n15835 ;
  assign n15838 = ~n15836 & ~n15837 ;
  assign n15839 = ~n15768 & ~n15838 ;
  assign n15840 = n15768 & ~n15837 ;
  assign n15841 = ~n15836 & n15840 ;
  assign n15842 = ~n15839 & ~n15841 ;
  assign n15843 = ~n15767 & n15842 ;
  assign n15844 = n15767 & ~n15842 ;
  assign n15845 = ~n15843 & ~n15844 ;
  assign n15846 = ~n15756 & n15845 ;
  assign n15847 = n15756 & ~n15845 ;
  assign n15848 = ~n15846 & ~n15847 ;
  assign n15849 = ~x82 & n6725 ;
  assign n15850 = ~x80 & n7129 ;
  assign n15851 = ~x81 & n6720 ;
  assign n15852 = ~n15850 & ~n15851 ;
  assign n15853 = ~n15849 & n15852 ;
  assign n15854 = n2697 & n6728 ;
  assign n15855 = n15853 & ~n15854 ;
  assign n15856 = ~x32 & ~n15855 ;
  assign n15857 = ~x32 & ~n15856 ;
  assign n15858 = ~n15855 & ~n15856 ;
  assign n15859 = ~n15857 & ~n15858 ;
  assign n15860 = n15848 & ~n15859 ;
  assign n15861 = n15848 & ~n15860 ;
  assign n15862 = ~n15859 & ~n15860 ;
  assign n15863 = ~n15861 & ~n15862 ;
  assign n15864 = ~n15254 & ~n15258 ;
  assign n15865 = n15863 & n15864 ;
  assign n15866 = ~n15863 & ~n15864 ;
  assign n15867 = ~n15865 & ~n15866 ;
  assign n15868 = ~x85 & n5560 ;
  assign n15869 = ~x83 & n5943 ;
  assign n15870 = ~x84 & n5555 ;
  assign n15871 = ~n15869 & ~n15870 ;
  assign n15872 = ~n15868 & n15871 ;
  assign n15873 = n3521 & n5563 ;
  assign n15874 = n15872 & ~n15873 ;
  assign n15875 = ~x29 & ~n15874 ;
  assign n15876 = ~x29 & ~n15875 ;
  assign n15877 = ~n15874 & ~n15875 ;
  assign n15878 = ~n15876 & ~n15877 ;
  assign n15879 = n15867 & ~n15878 ;
  assign n15880 = n15867 & ~n15879 ;
  assign n15881 = ~n15878 & ~n15879 ;
  assign n15882 = ~n15880 & ~n15881 ;
  assign n15883 = ~n15273 & ~n15279 ;
  assign n15884 = n15882 & n15883 ;
  assign n15885 = ~n15882 & ~n15883 ;
  assign n15886 = ~n15884 & ~n15885 ;
  assign n15887 = ~x88 & n4531 ;
  assign n15888 = ~x86 & n4847 ;
  assign n15889 = ~x87 & n4526 ;
  assign n15890 = ~n15888 & ~n15889 ;
  assign n15891 = ~n15887 & n15890 ;
  assign n15892 = n4457 & n4534 ;
  assign n15893 = n15891 & ~n15892 ;
  assign n15894 = ~x26 & ~n15893 ;
  assign n15895 = ~x26 & ~n15894 ;
  assign n15896 = ~n15893 & ~n15894 ;
  assign n15897 = ~n15895 & ~n15896 ;
  assign n15898 = ~n15886 & n15897 ;
  assign n15899 = n15886 & ~n15897 ;
  assign n15900 = ~n15898 & ~n15899 ;
  assign n15901 = ~n15297 & n15900 ;
  assign n15902 = n15297 & ~n15900 ;
  assign n15903 = ~n15901 & ~n15902 ;
  assign n15904 = ~x91 & n3589 ;
  assign n15905 = ~x89 & n3878 ;
  assign n15906 = ~x90 & n3584 ;
  assign n15907 = ~n15905 & ~n15906 ;
  assign n15908 = ~n15904 & n15907 ;
  assign n15909 = n3592 & n5507 ;
  assign n15910 = n15908 & ~n15909 ;
  assign n15911 = ~x23 & ~n15910 ;
  assign n15912 = ~x23 & ~n15911 ;
  assign n15913 = ~n15910 & ~n15911 ;
  assign n15914 = ~n15912 & ~n15913 ;
  assign n15915 = n15903 & ~n15914 ;
  assign n15916 = n15903 & ~n15915 ;
  assign n15917 = ~n15914 & ~n15915 ;
  assign n15918 = ~n15916 & ~n15917 ;
  assign n15919 = ~n15755 & n15918 ;
  assign n15920 = n15755 & ~n15918 ;
  assign n15921 = ~n15919 & ~n15920 ;
  assign n15922 = ~x94 & n2751 ;
  assign n15923 = ~x92 & n3020 ;
  assign n15924 = ~x93 & n2746 ;
  assign n15925 = ~n15923 & ~n15924 ;
  assign n15926 = ~n15922 & n15925 ;
  assign n15927 = n2754 & n6671 ;
  assign n15928 = n15926 & ~n15927 ;
  assign n15929 = ~x20 & ~n15928 ;
  assign n15930 = ~x20 & ~n15929 ;
  assign n15931 = ~n15928 & ~n15929 ;
  assign n15932 = ~n15930 & ~n15931 ;
  assign n15933 = ~n15921 & ~n15932 ;
  assign n15934 = n15921 & n15932 ;
  assign n15935 = ~n15933 & ~n15934 ;
  assign n15936 = ~n15754 & n15935 ;
  assign n15937 = n15754 & ~n15935 ;
  assign n15938 = ~n15936 & ~n15937 ;
  assign n15939 = ~x97 & n2093 ;
  assign n15940 = ~x95 & n2275 ;
  assign n15941 = ~x96 & n2088 ;
  assign n15942 = ~n15940 & ~n15941 ;
  assign n15943 = ~n15939 & n15942 ;
  assign n15944 = n2096 & n7949 ;
  assign n15945 = n15943 & ~n15944 ;
  assign n15946 = ~x17 & ~n15945 ;
  assign n15947 = ~x17 & ~n15946 ;
  assign n15948 = ~n15945 & ~n15946 ;
  assign n15949 = ~n15947 & ~n15948 ;
  assign n15950 = n15938 & ~n15949 ;
  assign n15951 = n15938 & ~n15950 ;
  assign n15952 = ~n15949 & ~n15950 ;
  assign n15953 = ~n15951 & ~n15952 ;
  assign n15954 = ~n15753 & n15953 ;
  assign n15955 = n15753 & ~n15953 ;
  assign n15956 = ~n15954 & ~n15955 ;
  assign n15957 = ~x100 & n1434 ;
  assign n15958 = ~x98 & n1646 ;
  assign n15959 = ~x99 & n1429 ;
  assign n15960 = ~n15958 & ~n15959 ;
  assign n15961 = ~n15957 & n15960 ;
  assign n15962 = n1437 & n9338 ;
  assign n15963 = n15961 & ~n15962 ;
  assign n15964 = ~x14 & ~n15963 ;
  assign n15965 = ~x14 & ~n15964 ;
  assign n15966 = ~n15963 & ~n15964 ;
  assign n15967 = ~n15965 & ~n15966 ;
  assign n15968 = ~n15956 & ~n15967 ;
  assign n15969 = n15956 & n15967 ;
  assign n15970 = ~n15968 & ~n15969 ;
  assign n15971 = n15752 & ~n15970 ;
  assign n15972 = ~n15752 & n15970 ;
  assign n15973 = ~n15971 & ~n15972 ;
  assign n15974 = ~x103 & n945 ;
  assign n15975 = ~x101 & n1099 ;
  assign n15976 = ~x102 & n940 ;
  assign n15977 = ~n15975 & ~n15976 ;
  assign n15978 = ~n15974 & n15977 ;
  assign n15979 = n948 & n10833 ;
  assign n15980 = n15978 & ~n15979 ;
  assign n15981 = ~x11 & ~n15980 ;
  assign n15982 = ~x11 & ~n15981 ;
  assign n15983 = ~n15980 & ~n15981 ;
  assign n15984 = ~n15982 & ~n15983 ;
  assign n15985 = n15973 & ~n15984 ;
  assign n15986 = n15973 & ~n15985 ;
  assign n15987 = ~n15984 & ~n15985 ;
  assign n15988 = ~n15986 & ~n15987 ;
  assign n15989 = ~n15359 & ~n15365 ;
  assign n15990 = n15988 & n15989 ;
  assign n15991 = ~n15988 & ~n15989 ;
  assign n15992 = ~n15990 & ~n15991 ;
  assign n15993 = ~x106 & n574 ;
  assign n15994 = ~x104 & n673 ;
  assign n15995 = ~x105 & n569 ;
  assign n15996 = ~n15994 & ~n15995 ;
  assign n15997 = ~n15993 & n15996 ;
  assign n15998 = n577 & n12447 ;
  assign n15999 = n15997 & ~n15998 ;
  assign n16000 = ~x8 & ~n15999 ;
  assign n16001 = ~x8 & ~n16000 ;
  assign n16002 = ~n15999 & ~n16000 ;
  assign n16003 = ~n16001 & ~n16002 ;
  assign n16004 = n15992 & ~n16003 ;
  assign n16005 = n15992 & ~n16004 ;
  assign n16006 = ~n16003 & ~n16004 ;
  assign n16007 = ~n16005 & ~n16006 ;
  assign n16008 = ~n15383 & n16007 ;
  assign n16009 = n15383 & ~n16007 ;
  assign n16010 = ~n16008 & ~n16009 ;
  assign n16011 = ~x109 & n293 ;
  assign n16012 = ~x107 & n373 ;
  assign n16013 = ~x108 & n288 ;
  assign n16014 = ~n16012 & ~n16013 ;
  assign n16015 = ~n16011 & n16014 ;
  assign n16016 = n296 & n14177 ;
  assign n16017 = n16015 & ~n16016 ;
  assign n16018 = ~x5 & ~n16017 ;
  assign n16019 = ~x5 & ~n16018 ;
  assign n16020 = ~n16017 & ~n16018 ;
  assign n16021 = ~n16019 & ~n16020 ;
  assign n16022 = ~n16010 & ~n16021 ;
  assign n16023 = n16010 & n16021 ;
  assign n16024 = ~n16022 & ~n16023 ;
  assign n16025 = ~n15751 & n16024 ;
  assign n16026 = n15751 & ~n16024 ;
  assign n16027 = ~n16025 & ~n16026 ;
  assign n16028 = n15750 & ~n16027 ;
  assign n16029 = ~n15750 & n16027 ;
  assign n16030 = ~n16028 & ~n16029 ;
  assign n16031 = ~n15735 & n16030 ;
  assign n16032 = n15735 & ~n16030 ;
  assign n16033 = ~n16031 & ~n16032 ;
  assign n16036 = ~n16033 & ~x176 ;
  assign n16037 = ~n16035 & ~n16036 ;
  assign n16038 = ~n15730 & ~n15732 ;
  assign n16039 = ~n15453 & ~n15619 ;
  assign n16040 = ~n15616 & ~n16039 ;
  assign n16041 = x92 & n3589 ;
  assign n16042 = x90 & n3878 ;
  assign n16043 = x91 & n3584 ;
  assign n16044 = ~n16042 & ~n16043 ;
  assign n16045 = ~n16041 & n16044 ;
  assign n16046 = n3592 & n5710 ;
  assign n16047 = n16045 & ~n16046 ;
  assign n16048 = x23 & ~n16047 ;
  assign n16049 = x23 & ~n16048 ;
  assign n16050 = ~n16047 & ~n16048 ;
  assign n16051 = ~n16049 & ~n16050 ;
  assign n16052 = ~n15536 & ~n15540 ;
  assign n16053 = ~n15531 & ~n15533 ;
  assign n16054 = n14888 & n15482 ;
  assign n16055 = ~n15497 & ~n16054 ;
  assign n16056 = x68 & n14233 ;
  assign n16057 = x66 & n14876 ;
  assign n16058 = x67 & n14228 ;
  assign n16059 = ~n16057 & ~n16058 ;
  assign n16060 = ~n16056 & n16059 ;
  assign n16061 = n317 & n14236 ;
  assign n16062 = n16060 & ~n16061 ;
  assign n16063 = x47 & ~n16062 ;
  assign n16064 = x47 & ~n16063 ;
  assign n16065 = ~n16062 & ~n16063 ;
  assign n16066 = ~n16064 & ~n16065 ;
  assign n16067 = x50 & ~n15482 ;
  assign n16068 = ~x48 & x49 ;
  assign n16069 = x48 & ~x49 ;
  assign n16070 = ~n16068 & ~n16069 ;
  assign n16071 = n15481 & ~n16070 ;
  assign n16072 = x64 & n16071 ;
  assign n16073 = ~x49 & x50 ;
  assign n16074 = x49 & ~x50 ;
  assign n16075 = ~n16073 & ~n16074 ;
  assign n16076 = ~n15481 & n16075 ;
  assign n16077 = x65 & n16076 ;
  assign n16078 = ~n16072 & ~n16077 ;
  assign n16079 = ~n15481 & ~n16075 ;
  assign n16080 = ~n152 & n16079 ;
  assign n16081 = n16078 & ~n16080 ;
  assign n16082 = x50 & ~n16081 ;
  assign n16083 = x50 & ~n16082 ;
  assign n16084 = ~n16081 & ~n16082 ;
  assign n16085 = ~n16083 & ~n16084 ;
  assign n16086 = n16067 & ~n16085 ;
  assign n16087 = ~n16067 & n16085 ;
  assign n16088 = ~n16086 & ~n16087 ;
  assign n16089 = n16066 & ~n16088 ;
  assign n16090 = ~n16066 & n16088 ;
  assign n16091 = ~n16089 & ~n16090 ;
  assign n16092 = ~n16055 & n16091 ;
  assign n16093 = n16055 & ~n16091 ;
  assign n16094 = ~n16092 & ~n16093 ;
  assign n16095 = x71 & n12506 ;
  assign n16096 = x69 & n13131 ;
  assign n16097 = x70 & n12501 ;
  assign n16098 = ~n16096 & ~n16097 ;
  assign n16099 = ~n16095 & n16098 ;
  assign n16100 = n558 & n12509 ;
  assign n16101 = n16099 & ~n16100 ;
  assign n16102 = x44 & ~n16101 ;
  assign n16103 = x44 & ~n16102 ;
  assign n16104 = ~n16101 & ~n16102 ;
  assign n16105 = ~n16103 & ~n16104 ;
  assign n16106 = n16094 & ~n16105 ;
  assign n16107 = n16094 & ~n16106 ;
  assign n16108 = ~n16105 & ~n16106 ;
  assign n16109 = ~n16107 & ~n16108 ;
  assign n16110 = ~n15511 & ~n15517 ;
  assign n16111 = n16109 & n16110 ;
  assign n16112 = ~n16109 & ~n16110 ;
  assign n16113 = ~n16111 & ~n16112 ;
  assign n16114 = x74 & n10905 ;
  assign n16115 = x72 & n11466 ;
  assign n16116 = x73 & n10900 ;
  assign n16117 = ~n16115 & ~n16116 ;
  assign n16118 = ~n16114 & n16117 ;
  assign n16119 = n994 & n10908 ;
  assign n16120 = n16118 & ~n16119 ;
  assign n16121 = x41 & ~n16120 ;
  assign n16122 = x41 & ~n16121 ;
  assign n16123 = ~n16120 & ~n16121 ;
  assign n16124 = ~n16122 & ~n16123 ;
  assign n16125 = n16113 & ~n16124 ;
  assign n16126 = ~n16113 & n16124 ;
  assign n16127 = ~n16053 & ~n16126 ;
  assign n16128 = ~n16125 & n16127 ;
  assign n16129 = ~n16053 & ~n16128 ;
  assign n16130 = ~n16125 & ~n16128 ;
  assign n16131 = ~n16126 & n16130 ;
  assign n16132 = ~n16129 & ~n16131 ;
  assign n16133 = x77 & n9433 ;
  assign n16134 = x75 & n9915 ;
  assign n16135 = x76 & n9428 ;
  assign n16136 = ~n16134 & ~n16135 ;
  assign n16137 = ~n16133 & n16136 ;
  assign n16138 = n1502 & n9436 ;
  assign n16139 = n16137 & ~n16138 ;
  assign n16140 = x38 & ~n16139 ;
  assign n16141 = x38 & ~n16140 ;
  assign n16142 = ~n16139 & ~n16140 ;
  assign n16143 = ~n16141 & ~n16142 ;
  assign n16144 = n16132 & n16143 ;
  assign n16145 = ~n16132 & ~n16143 ;
  assign n16146 = ~n16144 & ~n16145 ;
  assign n16147 = ~n16052 & n16146 ;
  assign n16148 = n16052 & ~n16146 ;
  assign n16149 = ~n16147 & ~n16148 ;
  assign n16150 = x80 & n8006 ;
  assign n16151 = x78 & n8474 ;
  assign n16152 = x79 & n8001 ;
  assign n16153 = ~n16151 & ~n16152 ;
  assign n16154 = ~n16150 & n16153 ;
  assign n16155 = n2028 & n8009 ;
  assign n16156 = n16154 & ~n16155 ;
  assign n16157 = x35 & ~n16156 ;
  assign n16158 = x35 & ~n16157 ;
  assign n16159 = ~n16156 & ~n16157 ;
  assign n16160 = ~n16158 & ~n16159 ;
  assign n16161 = n16149 & ~n16160 ;
  assign n16162 = n16149 & ~n16161 ;
  assign n16163 = ~n16160 & ~n16161 ;
  assign n16164 = ~n16162 & ~n16163 ;
  assign n16165 = ~n15544 & ~n15547 ;
  assign n16166 = n16164 & n16165 ;
  assign n16167 = ~n16164 & ~n16165 ;
  assign n16168 = ~n16166 & ~n16167 ;
  assign n16169 = x83 & n6725 ;
  assign n16170 = x81 & n7129 ;
  assign n16171 = x82 & n6720 ;
  assign n16172 = ~n16170 & ~n16171 ;
  assign n16173 = ~n16169 & n16172 ;
  assign n16174 = n2843 & n6728 ;
  assign n16175 = n16173 & ~n16174 ;
  assign n16176 = x32 & ~n16175 ;
  assign n16177 = x32 & ~n16176 ;
  assign n16178 = ~n16175 & ~n16176 ;
  assign n16179 = ~n16177 & ~n16178 ;
  assign n16180 = n16168 & ~n16179 ;
  assign n16181 = n16168 & ~n16180 ;
  assign n16182 = ~n16179 & ~n16180 ;
  assign n16183 = ~n16181 & ~n16182 ;
  assign n16184 = ~n15561 & ~n15567 ;
  assign n16185 = n16183 & n16184 ;
  assign n16186 = ~n16183 & ~n16184 ;
  assign n16187 = ~n16185 & ~n16186 ;
  assign n16188 = x86 & n5560 ;
  assign n16189 = x84 & n5943 ;
  assign n16190 = x85 & n5555 ;
  assign n16191 = ~n16189 & ~n16190 ;
  assign n16192 = ~n16188 & n16191 ;
  assign n16193 = n3686 & n5563 ;
  assign n16194 = n16192 & ~n16193 ;
  assign n16195 = x29 & ~n16194 ;
  assign n16196 = x29 & ~n16195 ;
  assign n16197 = ~n16194 & ~n16195 ;
  assign n16198 = ~n16196 & ~n16197 ;
  assign n16199 = n16187 & ~n16198 ;
  assign n16200 = n16187 & ~n16199 ;
  assign n16201 = ~n16198 & ~n16199 ;
  assign n16202 = ~n16200 & ~n16201 ;
  assign n16203 = ~n15580 & ~n15586 ;
  assign n16204 = n16202 & n16203 ;
  assign n16205 = ~n16202 & ~n16203 ;
  assign n16206 = ~n16204 & ~n16205 ;
  assign n16207 = x89 & n4531 ;
  assign n16208 = x87 & n4847 ;
  assign n16209 = x88 & n4526 ;
  assign n16210 = ~n16208 & ~n16209 ;
  assign n16211 = ~n16207 & n16210 ;
  assign n16212 = n4488 & n4534 ;
  assign n16213 = n16211 & ~n16212 ;
  assign n16214 = x26 & ~n16213 ;
  assign n16215 = x26 & ~n16214 ;
  assign n16216 = ~n16213 & ~n16214 ;
  assign n16217 = ~n16215 & ~n16216 ;
  assign n16218 = n16206 & ~n16217 ;
  assign n16219 = n16206 & ~n16218 ;
  assign n16220 = ~n16217 & ~n16218 ;
  assign n16221 = ~n16219 & ~n16220 ;
  assign n16222 = ~n15600 & ~n15602 ;
  assign n16223 = ~n16221 & ~n16222 ;
  assign n16224 = n16221 & n16222 ;
  assign n16225 = ~n16223 & ~n16224 ;
  assign n16226 = ~n16051 & n16225 ;
  assign n16227 = ~n16051 & ~n16226 ;
  assign n16228 = n16225 & ~n16226 ;
  assign n16229 = ~n16227 & ~n16228 ;
  assign n16230 = ~n16040 & ~n16229 ;
  assign n16231 = ~n16040 & ~n16230 ;
  assign n16232 = ~n16229 & ~n16230 ;
  assign n16233 = ~n16231 & ~n16232 ;
  assign n16234 = x95 & n2751 ;
  assign n16235 = x93 & n3020 ;
  assign n16236 = x94 & n2746 ;
  assign n16237 = ~n16235 & ~n16236 ;
  assign n16238 = ~n16234 & n16237 ;
  assign n16239 = n2754 & n6894 ;
  assign n16240 = n16238 & ~n16239 ;
  assign n16241 = x20 & ~n16240 ;
  assign n16242 = x20 & ~n16241 ;
  assign n16243 = ~n16240 & ~n16241 ;
  assign n16244 = ~n16242 & ~n16243 ;
  assign n16245 = ~n16233 & ~n16244 ;
  assign n16246 = ~n16233 & ~n16245 ;
  assign n16247 = ~n16244 & ~n16245 ;
  assign n16248 = ~n16246 & ~n16247 ;
  assign n16249 = ~n15634 & ~n15637 ;
  assign n16250 = n16248 & n16249 ;
  assign n16251 = ~n16248 & ~n16249 ;
  assign n16252 = ~n16250 & ~n16251 ;
  assign n16253 = x98 & n2093 ;
  assign n16254 = x96 & n2275 ;
  assign n16255 = x97 & n2088 ;
  assign n16256 = ~n16254 & ~n16255 ;
  assign n16257 = ~n16253 & n16256 ;
  assign n16258 = n2096 & n8196 ;
  assign n16259 = n16257 & ~n16258 ;
  assign n16260 = x17 & ~n16259 ;
  assign n16261 = x17 & ~n16260 ;
  assign n16262 = ~n16259 & ~n16260 ;
  assign n16263 = ~n16261 & ~n16262 ;
  assign n16264 = n16252 & ~n16263 ;
  assign n16265 = n16252 & ~n16264 ;
  assign n16266 = ~n16263 & ~n16264 ;
  assign n16267 = ~n16265 & ~n16266 ;
  assign n16268 = ~n15451 & ~n15654 ;
  assign n16269 = ~n15651 & ~n16268 ;
  assign n16270 = n16267 & n16269 ;
  assign n16271 = ~n16267 & ~n16269 ;
  assign n16272 = ~n16270 & ~n16271 ;
  assign n16273 = x101 & n1434 ;
  assign n16274 = x99 & n1646 ;
  assign n16275 = x100 & n1429 ;
  assign n16276 = ~n16274 & ~n16275 ;
  assign n16277 = ~n16273 & n16276 ;
  assign n16278 = n1437 & n9601 ;
  assign n16279 = n16277 & ~n16278 ;
  assign n16280 = x14 & ~n16279 ;
  assign n16281 = x14 & ~n16280 ;
  assign n16282 = ~n16279 & ~n16280 ;
  assign n16283 = ~n16281 & ~n16282 ;
  assign n16284 = n16272 & ~n16283 ;
  assign n16285 = n16272 & ~n16284 ;
  assign n16286 = ~n16283 & ~n16284 ;
  assign n16287 = ~n16285 & ~n16286 ;
  assign n16288 = ~n15669 & ~n15673 ;
  assign n16289 = n16287 & n16288 ;
  assign n16290 = ~n16287 & ~n16288 ;
  assign n16291 = ~n16289 & ~n16290 ;
  assign n16292 = x104 & n945 ;
  assign n16293 = x102 & n1099 ;
  assign n16294 = x103 & n940 ;
  assign n16295 = ~n16293 & ~n16294 ;
  assign n16296 = ~n16292 & n16295 ;
  assign n16297 = n948 & n11116 ;
  assign n16298 = n16296 & ~n16297 ;
  assign n16299 = x11 & ~n16298 ;
  assign n16300 = x11 & ~n16299 ;
  assign n16301 = ~n16298 & ~n16299 ;
  assign n16302 = ~n16300 & ~n16301 ;
  assign n16303 = n16291 & ~n16302 ;
  assign n16304 = n16291 & ~n16303 ;
  assign n16305 = ~n16302 & ~n16303 ;
  assign n16306 = ~n16304 & ~n16305 ;
  assign n16307 = ~n15686 & ~n15692 ;
  assign n16308 = n16306 & n16307 ;
  assign n16309 = ~n16306 & ~n16307 ;
  assign n16310 = ~n16308 & ~n16309 ;
  assign n16311 = x107 & n574 ;
  assign n16312 = x105 & n673 ;
  assign n16313 = x106 & n569 ;
  assign n16314 = ~n16312 & ~n16313 ;
  assign n16315 = ~n16311 & n16314 ;
  assign n16316 = n577 & n12749 ;
  assign n16317 = n16315 & ~n16316 ;
  assign n16318 = x8 & ~n16317 ;
  assign n16319 = x8 & ~n16318 ;
  assign n16320 = ~n16317 & ~n16318 ;
  assign n16321 = ~n16319 & ~n16320 ;
  assign n16322 = n16310 & ~n16321 ;
  assign n16323 = n16310 & ~n16322 ;
  assign n16324 = ~n16321 & ~n16322 ;
  assign n16325 = ~n16323 & ~n16324 ;
  assign n16326 = ~n15080 & ~n15708 ;
  assign n16327 = ~n15705 & ~n16326 ;
  assign n16328 = n16325 & n16327 ;
  assign n16329 = ~n16325 & ~n16327 ;
  assign n16330 = ~n16328 & ~n16329 ;
  assign n16331 = x110 & n293 ;
  assign n16332 = x108 & n373 ;
  assign n16333 = x109 & n288 ;
  assign n16334 = ~n16332 & ~n16333 ;
  assign n16335 = ~n16331 & n16334 ;
  assign n16336 = n296 & n14497 ;
  assign n16337 = n16335 & ~n16336 ;
  assign n16338 = x5 & ~n16337 ;
  assign n16339 = x5 & ~n16338 ;
  assign n16340 = ~n16337 & ~n16338 ;
  assign n16341 = ~n16339 & ~n16340 ;
  assign n16342 = n16330 & ~n16341 ;
  assign n16343 = n16330 & ~n16342 ;
  assign n16344 = ~n16341 & ~n16342 ;
  assign n16345 = ~n16343 & ~n16344 ;
  assign n16346 = ~n15723 & ~n15726 ;
  assign n16347 = n16345 & n16346 ;
  assign n16348 = ~n16345 & ~n16346 ;
  assign n16349 = ~n16347 & ~n16348 ;
  assign n16350 = x113 & n146 ;
  assign n16351 = x111 & n182 ;
  assign n16352 = x112 & n141 ;
  assign n16353 = ~n16351 & ~n16352 ;
  assign n16354 = ~n16350 & n16353 ;
  assign n16355 = ~n15438 & ~n15440 ;
  assign n16356 = ~x112 & ~x113 ;
  assign n16357 = x112 & x113 ;
  assign n16358 = ~n16356 & ~n16357 ;
  assign n16359 = ~n16355 & n16358 ;
  assign n16360 = n16355 & ~n16358 ;
  assign n16361 = ~n16359 & ~n16360 ;
  assign n16362 = n149 & n16361 ;
  assign n16363 = n16354 & ~n16362 ;
  assign n16364 = x2 & ~n16363 ;
  assign n16365 = x2 & ~n16364 ;
  assign n16366 = ~n16363 & ~n16364 ;
  assign n16367 = ~n16365 & ~n16366 ;
  assign n16368 = ~n16349 & n16367 ;
  assign n16369 = n16349 & ~n16367 ;
  assign n16370 = ~n16368 & ~n16369 ;
  assign n16371 = ~n16038 & n16370 ;
  assign n16372 = n16038 & ~n16370 ;
  assign n16373 = ~n16371 & ~n16372 ;
  assign n16698 = n16373 & x177 ;
  assign n16374 = ~n16029 & ~n16031 ;
  assign n16375 = ~n15755 & ~n15918 ;
  assign n16376 = ~n15915 & ~n16375 ;
  assign n16377 = ~x92 & n3589 ;
  assign n16378 = ~x90 & n3878 ;
  assign n16379 = ~x91 & n3584 ;
  assign n16380 = ~n16378 & ~n16379 ;
  assign n16381 = ~n16377 & n16380 ;
  assign n16382 = n3592 & n5896 ;
  assign n16383 = n16381 & ~n16382 ;
  assign n16384 = ~x23 & ~n16383 ;
  assign n16385 = ~x23 & ~n16384 ;
  assign n16386 = ~n16383 & ~n16384 ;
  assign n16387 = ~n16385 & ~n16386 ;
  assign n16388 = ~n15835 & ~n15839 ;
  assign n16389 = ~n15830 & ~n15832 ;
  assign n16390 = n15191 & n15781 ;
  assign n16391 = ~n15796 & ~n16390 ;
  assign n16392 = ~x68 & n14233 ;
  assign n16393 = ~x66 & n14876 ;
  assign n16394 = ~x67 & n14228 ;
  assign n16395 = ~n16393 & ~n16394 ;
  assign n16396 = ~n16392 & n16395 ;
  assign n16397 = n352 & n14236 ;
  assign n16398 = n16396 & ~n16397 ;
  assign n16399 = ~x47 & ~n16398 ;
  assign n16400 = ~x47 & ~n16399 ;
  assign n16401 = ~n16398 & ~n16399 ;
  assign n16402 = ~n16400 & ~n16401 ;
  assign n16403 = ~x50 & ~n15781 ;
  assign n16404 = ~x64 & n16071 ;
  assign n16405 = ~x65 & n16076 ;
  assign n16406 = ~n16404 & ~n16405 ;
  assign n16407 = ~n16080 & n16406 ;
  assign n16408 = ~x50 & ~n16407 ;
  assign n16409 = ~x50 & ~n16408 ;
  assign n16410 = ~n16407 & ~n16408 ;
  assign n16411 = ~n16409 & ~n16410 ;
  assign n16412 = n16403 & ~n16411 ;
  assign n16413 = ~n16403 & n16411 ;
  assign n16414 = ~n16412 & ~n16413 ;
  assign n16415 = n16402 & ~n16414 ;
  assign n16416 = ~n16402 & n16414 ;
  assign n16417 = ~n16415 & ~n16416 ;
  assign n16418 = ~n16391 & n16417 ;
  assign n16419 = n16391 & ~n16417 ;
  assign n16420 = ~n16418 & ~n16419 ;
  assign n16421 = ~x71 & n12506 ;
  assign n16422 = ~x69 & n13131 ;
  assign n16423 = ~x70 & n12501 ;
  assign n16424 = ~n16422 & ~n16423 ;
  assign n16425 = ~n16421 & n16424 ;
  assign n16426 = n622 & n12509 ;
  assign n16427 = n16425 & ~n16426 ;
  assign n16428 = ~x44 & ~n16427 ;
  assign n16429 = ~x44 & ~n16428 ;
  assign n16430 = ~n16427 & ~n16428 ;
  assign n16431 = ~n16429 & ~n16430 ;
  assign n16432 = n16420 & ~n16431 ;
  assign n16433 = n16420 & ~n16432 ;
  assign n16434 = ~n16431 & ~n16432 ;
  assign n16435 = ~n16433 & ~n16434 ;
  assign n16436 = ~n15810 & ~n15816 ;
  assign n16437 = n16435 & n16436 ;
  assign n16438 = ~n16435 & ~n16436 ;
  assign n16439 = ~n16437 & ~n16438 ;
  assign n16440 = ~x74 & n10905 ;
  assign n16441 = ~x72 & n11466 ;
  assign n16442 = ~x73 & n10900 ;
  assign n16443 = ~n16441 & ~n16442 ;
  assign n16444 = ~n16440 & n16443 ;
  assign n16445 = n1066 & n10908 ;
  assign n16446 = n16444 & ~n16445 ;
  assign n16447 = ~x41 & ~n16446 ;
  assign n16448 = ~x41 & ~n16447 ;
  assign n16449 = ~n16446 & ~n16447 ;
  assign n16450 = ~n16448 & ~n16449 ;
  assign n16451 = n16439 & ~n16450 ;
  assign n16452 = ~n16439 & n16450 ;
  assign n16453 = ~n16389 & ~n16452 ;
  assign n16454 = ~n16451 & n16453 ;
  assign n16455 = ~n16389 & ~n16454 ;
  assign n16456 = ~n16451 & ~n16454 ;
  assign n16457 = ~n16452 & n16456 ;
  assign n16458 = ~n16455 & ~n16457 ;
  assign n16459 = ~x77 & n9433 ;
  assign n16460 = ~x75 & n9915 ;
  assign n16461 = ~x76 & n9428 ;
  assign n16462 = ~n16460 & ~n16461 ;
  assign n16463 = ~n16459 & n16462 ;
  assign n16464 = n1594 & n9436 ;
  assign n16465 = n16463 & ~n16464 ;
  assign n16466 = ~x38 & ~n16465 ;
  assign n16467 = ~x38 & ~n16466 ;
  assign n16468 = ~n16465 & ~n16466 ;
  assign n16469 = ~n16467 & ~n16468 ;
  assign n16470 = n16458 & n16469 ;
  assign n16471 = ~n16458 & ~n16469 ;
  assign n16472 = ~n16470 & ~n16471 ;
  assign n16473 = ~n16388 & n16472 ;
  assign n16474 = n16388 & ~n16472 ;
  assign n16475 = ~n16473 & ~n16474 ;
  assign n16476 = ~x80 & n8006 ;
  assign n16477 = ~x78 & n8474 ;
  assign n16478 = ~x79 & n8001 ;
  assign n16479 = ~n16477 & ~n16478 ;
  assign n16480 = ~n16476 & n16479 ;
  assign n16481 = n2145 & n8009 ;
  assign n16482 = n16480 & ~n16481 ;
  assign n16483 = ~x35 & ~n16482 ;
  assign n16484 = ~x35 & ~n16483 ;
  assign n16485 = ~n16482 & ~n16483 ;
  assign n16486 = ~n16484 & ~n16485 ;
  assign n16487 = n16475 & ~n16486 ;
  assign n16488 = n16475 & ~n16487 ;
  assign n16489 = ~n16486 & ~n16487 ;
  assign n16490 = ~n16488 & ~n16489 ;
  assign n16491 = ~n15843 & ~n15846 ;
  assign n16492 = n16490 & n16491 ;
  assign n16493 = ~n16490 & ~n16491 ;
  assign n16494 = ~n16492 & ~n16493 ;
  assign n16495 = ~x83 & n6725 ;
  assign n16496 = ~x81 & n7129 ;
  assign n16497 = ~x82 & n6720 ;
  assign n16498 = ~n16496 & ~n16497 ;
  assign n16499 = ~n16495 & n16498 ;
  assign n16500 = n2972 & n6728 ;
  assign n16501 = n16499 & ~n16500 ;
  assign n16502 = ~x32 & ~n16501 ;
  assign n16503 = ~x32 & ~n16502 ;
  assign n16504 = ~n16501 & ~n16502 ;
  assign n16505 = ~n16503 & ~n16504 ;
  assign n16506 = n16494 & ~n16505 ;
  assign n16507 = n16494 & ~n16506 ;
  assign n16508 = ~n16505 & ~n16506 ;
  assign n16509 = ~n16507 & ~n16508 ;
  assign n16510 = ~n15860 & ~n15866 ;
  assign n16511 = n16509 & n16510 ;
  assign n16512 = ~n16509 & ~n16510 ;
  assign n16513 = ~n16511 & ~n16512 ;
  assign n16514 = ~x86 & n5560 ;
  assign n16515 = ~x84 & n5943 ;
  assign n16516 = ~x85 & n5555 ;
  assign n16517 = ~n16515 & ~n16516 ;
  assign n16518 = ~n16514 & n16517 ;
  assign n16519 = n3832 & n5563 ;
  assign n16520 = n16518 & ~n16519 ;
  assign n16521 = ~x29 & ~n16520 ;
  assign n16522 = ~x29 & ~n16521 ;
  assign n16523 = ~n16520 & ~n16521 ;
  assign n16524 = ~n16522 & ~n16523 ;
  assign n16525 = n16513 & ~n16524 ;
  assign n16526 = n16513 & ~n16525 ;
  assign n16527 = ~n16524 & ~n16525 ;
  assign n16528 = ~n16526 & ~n16527 ;
  assign n16529 = ~n15879 & ~n15885 ;
  assign n16530 = n16528 & n16529 ;
  assign n16531 = ~n16528 & ~n16529 ;
  assign n16532 = ~n16530 & ~n16531 ;
  assign n16533 = ~x89 & n4531 ;
  assign n16534 = ~x87 & n4847 ;
  assign n16535 = ~x88 & n4526 ;
  assign n16536 = ~n16534 & ~n16535 ;
  assign n16537 = ~n16533 & n16536 ;
  assign n16538 = n4534 & n4664 ;
  assign n16539 = n16537 & ~n16538 ;
  assign n16540 = ~x26 & ~n16539 ;
  assign n16541 = ~x26 & ~n16540 ;
  assign n16542 = ~n16539 & ~n16540 ;
  assign n16543 = ~n16541 & ~n16542 ;
  assign n16544 = n16532 & ~n16543 ;
  assign n16545 = n16532 & ~n16544 ;
  assign n16546 = ~n16543 & ~n16544 ;
  assign n16547 = ~n16545 & ~n16546 ;
  assign n16548 = ~n15899 & ~n15901 ;
  assign n16549 = ~n16547 & ~n16548 ;
  assign n16550 = n16547 & n16548 ;
  assign n16551 = ~n16549 & ~n16550 ;
  assign n16552 = ~n16387 & n16551 ;
  assign n16553 = ~n16387 & ~n16552 ;
  assign n16554 = n16551 & ~n16552 ;
  assign n16555 = ~n16553 & ~n16554 ;
  assign n16556 = ~n16376 & ~n16555 ;
  assign n16557 = ~n16376 & ~n16556 ;
  assign n16558 = ~n16555 & ~n16556 ;
  assign n16559 = ~n16557 & ~n16558 ;
  assign n16560 = ~x95 & n2751 ;
  assign n16561 = ~x93 & n3020 ;
  assign n16562 = ~x94 & n2746 ;
  assign n16563 = ~n16561 & ~n16562 ;
  assign n16564 = ~n16560 & n16563 ;
  assign n16565 = n2754 & n7100 ;
  assign n16566 = n16564 & ~n16565 ;
  assign n16567 = ~x20 & ~n16566 ;
  assign n16568 = ~x20 & ~n16567 ;
  assign n16569 = ~n16566 & ~n16567 ;
  assign n16570 = ~n16568 & ~n16569 ;
  assign n16571 = ~n16559 & ~n16570 ;
  assign n16572 = ~n16559 & ~n16571 ;
  assign n16573 = ~n16570 & ~n16571 ;
  assign n16574 = ~n16572 & ~n16573 ;
  assign n16575 = ~n15933 & ~n15936 ;
  assign n16576 = n16574 & n16575 ;
  assign n16577 = ~n16574 & ~n16575 ;
  assign n16578 = ~n16576 & ~n16577 ;
  assign n16579 = ~x98 & n2093 ;
  assign n16580 = ~x96 & n2275 ;
  assign n16581 = ~x97 & n2088 ;
  assign n16582 = ~n16580 & ~n16581 ;
  assign n16583 = ~n16579 & n16582 ;
  assign n16584 = n2096 & n8426 ;
  assign n16585 = n16583 & ~n16584 ;
  assign n16586 = ~x17 & ~n16585 ;
  assign n16587 = ~x17 & ~n16586 ;
  assign n16588 = ~n16585 & ~n16586 ;
  assign n16589 = ~n16587 & ~n16588 ;
  assign n16590 = n16578 & ~n16589 ;
  assign n16591 = n16578 & ~n16590 ;
  assign n16592 = ~n16589 & ~n16590 ;
  assign n16593 = ~n16591 & ~n16592 ;
  assign n16594 = ~n15753 & ~n15953 ;
  assign n16595 = ~n15950 & ~n16594 ;
  assign n16596 = n16593 & n16595 ;
  assign n16597 = ~n16593 & ~n16595 ;
  assign n16598 = ~n16596 & ~n16597 ;
  assign n16599 = ~x101 & n1434 ;
  assign n16600 = ~x99 & n1646 ;
  assign n16601 = ~x100 & n1429 ;
  assign n16602 = ~n16600 & ~n16601 ;
  assign n16603 = ~n16599 & n16602 ;
  assign n16604 = n1437 & n9844 ;
  assign n16605 = n16603 & ~n16604 ;
  assign n16606 = ~x14 & ~n16605 ;
  assign n16607 = ~x14 & ~n16606 ;
  assign n16608 = ~n16605 & ~n16606 ;
  assign n16609 = ~n16607 & ~n16608 ;
  assign n16610 = n16598 & ~n16609 ;
  assign n16611 = n16598 & ~n16610 ;
  assign n16612 = ~n16609 & ~n16610 ;
  assign n16613 = ~n16611 & ~n16612 ;
  assign n16614 = ~n15968 & ~n15972 ;
  assign n16615 = n16613 & n16614 ;
  assign n16616 = ~n16613 & ~n16614 ;
  assign n16617 = ~n16615 & ~n16616 ;
  assign n16618 = ~x104 & n945 ;
  assign n16619 = ~x102 & n1099 ;
  assign n16620 = ~x103 & n940 ;
  assign n16621 = ~n16619 & ~n16620 ;
  assign n16622 = ~n16618 & n16621 ;
  assign n16623 = n948 & n11380 ;
  assign n16624 = n16622 & ~n16623 ;
  assign n16625 = ~x11 & ~n16624 ;
  assign n16626 = ~x11 & ~n16625 ;
  assign n16627 = ~n16624 & ~n16625 ;
  assign n16628 = ~n16626 & ~n16627 ;
  assign n16629 = n16617 & ~n16628 ;
  assign n16630 = n16617 & ~n16629 ;
  assign n16631 = ~n16628 & ~n16629 ;
  assign n16632 = ~n16630 & ~n16631 ;
  assign n16633 = ~n15985 & ~n15991 ;
  assign n16634 = n16632 & n16633 ;
  assign n16635 = ~n16632 & ~n16633 ;
  assign n16636 = ~n16634 & ~n16635 ;
  assign n16637 = ~x107 & n574 ;
  assign n16638 = ~x105 & n673 ;
  assign n16639 = ~x106 & n569 ;
  assign n16640 = ~n16638 & ~n16639 ;
  assign n16641 = ~n16637 & n16640 ;
  assign n16642 = n577 & n13034 ;
  assign n16643 = n16641 & ~n16642 ;
  assign n16644 = ~x8 & ~n16643 ;
  assign n16645 = ~x8 & ~n16644 ;
  assign n16646 = ~n16643 & ~n16644 ;
  assign n16647 = ~n16645 & ~n16646 ;
  assign n16648 = n16636 & ~n16647 ;
  assign n16649 = n16636 & ~n16648 ;
  assign n16650 = ~n16647 & ~n16648 ;
  assign n16651 = ~n16649 & ~n16650 ;
  assign n16652 = ~n15383 & ~n16007 ;
  assign n16653 = ~n16004 & ~n16652 ;
  assign n16654 = n16651 & n16653 ;
  assign n16655 = ~n16651 & ~n16653 ;
  assign n16656 = ~n16654 & ~n16655 ;
  assign n16657 = ~x110 & n293 ;
  assign n16658 = ~x108 & n373 ;
  assign n16659 = ~x109 & n288 ;
  assign n16660 = ~n16658 & ~n16659 ;
  assign n16661 = ~n16657 & n16660 ;
  assign n16662 = n296 & n14802 ;
  assign n16663 = n16661 & ~n16662 ;
  assign n16664 = ~x5 & ~n16663 ;
  assign n16665 = ~x5 & ~n16664 ;
  assign n16666 = ~n16663 & ~n16664 ;
  assign n16667 = ~n16665 & ~n16666 ;
  assign n16668 = n16656 & ~n16667 ;
  assign n16669 = n16656 & ~n16668 ;
  assign n16670 = ~n16667 & ~n16668 ;
  assign n16671 = ~n16669 & ~n16670 ;
  assign n16672 = ~n16022 & ~n16025 ;
  assign n16673 = n16671 & n16672 ;
  assign n16674 = ~n16671 & ~n16672 ;
  assign n16675 = ~n16673 & ~n16674 ;
  assign n16676 = ~x113 & n164 ;
  assign n16677 = ~x111 & n205 ;
  assign n16678 = ~x112 & n162 ;
  assign n16679 = ~n16677 & ~n16678 ;
  assign n16680 = ~n16676 & n16679 ;
  assign n16681 = ~n15437 & ~n15742 ;
  assign n16682 = n16358 & ~n16681 ;
  assign n16683 = ~n16358 & n16681 ;
  assign n16684 = ~n16682 & ~n16683 ;
  assign n16685 = n167 & n16684 ;
  assign n16686 = n16680 & ~n16685 ;
  assign n16687 = ~x2 & ~n16686 ;
  assign n16688 = ~x2 & ~n16687 ;
  assign n16689 = ~n16686 & ~n16687 ;
  assign n16690 = ~n16688 & ~n16689 ;
  assign n16691 = ~n16675 & n16690 ;
  assign n16692 = n16675 & ~n16690 ;
  assign n16693 = ~n16691 & ~n16692 ;
  assign n16694 = ~n16374 & n16693 ;
  assign n16695 = n16374 & ~n16693 ;
  assign n16696 = ~n16694 & ~n16695 ;
  assign n16699 = ~n16696 & ~x177 ;
  assign n16700 = ~n16698 & ~n16699 ;
  assign n16701 = ~n16322 & ~n16329 ;
  assign n16702 = ~n16245 & ~n16251 ;
  assign n16703 = x96 & n2751 ;
  assign n16704 = x94 & n3020 ;
  assign n16705 = x95 & n2746 ;
  assign n16706 = ~n16704 & ~n16705 ;
  assign n16707 = ~n16703 & n16706 ;
  assign n16708 = n2754 & n7321 ;
  assign n16709 = n16707 & ~n16708 ;
  assign n16710 = x20 & ~n16709 ;
  assign n16711 = x20 & ~n16710 ;
  assign n16712 = ~n16709 & ~n16710 ;
  assign n16713 = ~n16711 & ~n16712 ;
  assign n16714 = ~n16226 & ~n16230 ;
  assign n16715 = x93 & n3589 ;
  assign n16716 = x91 & n3878 ;
  assign n16717 = x92 & n3584 ;
  assign n16718 = ~n16716 & ~n16717 ;
  assign n16719 = ~n16715 & n16718 ;
  assign n16720 = n3592 & n6094 ;
  assign n16721 = n16719 & ~n16720 ;
  assign n16722 = x23 & ~n16721 ;
  assign n16723 = x23 & ~n16722 ;
  assign n16724 = ~n16721 & ~n16722 ;
  assign n16725 = ~n16723 & ~n16724 ;
  assign n16726 = ~n16218 & ~n16223 ;
  assign n16727 = ~n16199 & ~n16205 ;
  assign n16728 = ~n16161 & ~n16167 ;
  assign n16729 = x81 & n8006 ;
  assign n16730 = x79 & n8474 ;
  assign n16731 = x80 & n8001 ;
  assign n16732 = ~n16730 & ~n16731 ;
  assign n16733 = ~n16729 & n16732 ;
  assign n16734 = n2348 & n8009 ;
  assign n16735 = n16733 & ~n16734 ;
  assign n16736 = x35 & ~n16735 ;
  assign n16737 = x35 & ~n16736 ;
  assign n16738 = ~n16735 & ~n16736 ;
  assign n16739 = ~n16737 & ~n16738 ;
  assign n16740 = ~n16145 & ~n16147 ;
  assign n16741 = ~n16106 & ~n16112 ;
  assign n16742 = x72 & n12506 ;
  assign n16743 = x70 & n13131 ;
  assign n16744 = x71 & n12501 ;
  assign n16745 = ~n16743 & ~n16744 ;
  assign n16746 = ~n16742 & n16745 ;
  assign n16747 = n717 & n12509 ;
  assign n16748 = n16746 & ~n16747 ;
  assign n16749 = x44 & ~n16748 ;
  assign n16750 = x44 & ~n16749 ;
  assign n16751 = ~n16748 & ~n16749 ;
  assign n16752 = ~n16750 & ~n16751 ;
  assign n16753 = ~n16090 & ~n16092 ;
  assign n16754 = x66 & n16076 ;
  assign n16755 = n15481 & ~n16075 ;
  assign n16756 = n16070 & n16755 ;
  assign n16757 = x64 & n16756 ;
  assign n16758 = x65 & n16071 ;
  assign n16759 = ~n16757 & ~n16758 ;
  assign n16760 = ~n16754 & n16759 ;
  assign n16761 = n194 & n16079 ;
  assign n16762 = n16760 & ~n16761 ;
  assign n16763 = x50 & ~n16762 ;
  assign n16764 = x50 & ~n16763 ;
  assign n16765 = ~n16762 & ~n16763 ;
  assign n16766 = ~n16764 & ~n16765 ;
  assign n16767 = ~n16086 & n16766 ;
  assign n16768 = n16086 & ~n16766 ;
  assign n16769 = ~n16767 & ~n16768 ;
  assign n16770 = x69 & n14233 ;
  assign n16771 = x67 & n14876 ;
  assign n16772 = x68 & n14228 ;
  assign n16773 = ~n16771 & ~n16772 ;
  assign n16774 = ~n16770 & n16773 ;
  assign n16775 = n398 & n14236 ;
  assign n16776 = n16774 & ~n16775 ;
  assign n16777 = x47 & ~n16776 ;
  assign n16778 = x47 & ~n16777 ;
  assign n16779 = ~n16776 & ~n16777 ;
  assign n16780 = ~n16778 & ~n16779 ;
  assign n16781 = n16769 & ~n16780 ;
  assign n16782 = n16769 & ~n16781 ;
  assign n16783 = ~n16780 & ~n16781 ;
  assign n16784 = ~n16782 & ~n16783 ;
  assign n16785 = ~n16753 & ~n16784 ;
  assign n16786 = n16753 & n16784 ;
  assign n16787 = ~n16785 & ~n16786 ;
  assign n16788 = ~n16752 & n16787 ;
  assign n16789 = ~n16752 & ~n16788 ;
  assign n16790 = n16787 & ~n16788 ;
  assign n16791 = ~n16789 & ~n16790 ;
  assign n16792 = ~n16741 & ~n16791 ;
  assign n16793 = ~n16741 & ~n16792 ;
  assign n16794 = ~n16791 & ~n16792 ;
  assign n16795 = ~n16793 & ~n16794 ;
  assign n16796 = x75 & n10905 ;
  assign n16797 = x73 & n11466 ;
  assign n16798 = x74 & n10900 ;
  assign n16799 = ~n16797 & ~n16798 ;
  assign n16800 = ~n16796 & n16799 ;
  assign n16801 = n1150 & n10908 ;
  assign n16802 = n16800 & ~n16801 ;
  assign n16803 = x41 & ~n16802 ;
  assign n16804 = x41 & ~n16803 ;
  assign n16805 = ~n16802 & ~n16803 ;
  assign n16806 = ~n16804 & ~n16805 ;
  assign n16807 = n16795 & n16806 ;
  assign n16808 = ~n16795 & ~n16806 ;
  assign n16809 = ~n16807 & ~n16808 ;
  assign n16810 = ~n16130 & n16809 ;
  assign n16811 = n16130 & ~n16809 ;
  assign n16812 = ~n16810 & ~n16811 ;
  assign n16813 = x78 & n9433 ;
  assign n16814 = x76 & n9915 ;
  assign n16815 = x77 & n9428 ;
  assign n16816 = ~n16814 & ~n16815 ;
  assign n16817 = ~n16813 & n16816 ;
  assign n16818 = n1624 & n9436 ;
  assign n16819 = n16817 & ~n16818 ;
  assign n16820 = x38 & ~n16819 ;
  assign n16821 = x38 & ~n16820 ;
  assign n16822 = ~n16819 & ~n16820 ;
  assign n16823 = ~n16821 & ~n16822 ;
  assign n16824 = n16812 & ~n16823 ;
  assign n16825 = n16812 & ~n16824 ;
  assign n16826 = ~n16823 & ~n16824 ;
  assign n16827 = ~n16825 & ~n16826 ;
  assign n16828 = ~n16740 & ~n16827 ;
  assign n16829 = n16740 & n16827 ;
  assign n16830 = ~n16828 & ~n16829 ;
  assign n16831 = ~n16739 & n16830 ;
  assign n16832 = ~n16739 & ~n16831 ;
  assign n16833 = n16830 & ~n16831 ;
  assign n16834 = ~n16832 & ~n16833 ;
  assign n16835 = ~n16728 & ~n16834 ;
  assign n16836 = ~n16728 & ~n16835 ;
  assign n16837 = ~n16834 & ~n16835 ;
  assign n16838 = ~n16836 & ~n16837 ;
  assign n16839 = x84 & n6725 ;
  assign n16840 = x82 & n7129 ;
  assign n16841 = x83 & n6720 ;
  assign n16842 = ~n16840 & ~n16841 ;
  assign n16843 = ~n16839 & n16842 ;
  assign n16844 = n3114 & n6728 ;
  assign n16845 = n16843 & ~n16844 ;
  assign n16846 = x32 & ~n16845 ;
  assign n16847 = x32 & ~n16846 ;
  assign n16848 = ~n16845 & ~n16846 ;
  assign n16849 = ~n16847 & ~n16848 ;
  assign n16850 = ~n16838 & ~n16849 ;
  assign n16851 = ~n16838 & ~n16850 ;
  assign n16852 = ~n16849 & ~n16850 ;
  assign n16853 = ~n16851 & ~n16852 ;
  assign n16854 = ~n16180 & ~n16186 ;
  assign n16855 = n16853 & n16854 ;
  assign n16856 = ~n16853 & ~n16854 ;
  assign n16857 = ~n16855 & ~n16856 ;
  assign n16858 = x87 & n5560 ;
  assign n16859 = x85 & n5943 ;
  assign n16860 = x86 & n5555 ;
  assign n16861 = ~n16859 & ~n16860 ;
  assign n16862 = ~n16858 & n16861 ;
  assign n16863 = n3991 & n5563 ;
  assign n16864 = n16862 & ~n16863 ;
  assign n16865 = x29 & ~n16864 ;
  assign n16866 = x29 & ~n16865 ;
  assign n16867 = ~n16864 & ~n16865 ;
  assign n16868 = ~n16866 & ~n16867 ;
  assign n16869 = n16857 & ~n16868 ;
  assign n16870 = ~n16857 & n16868 ;
  assign n16871 = ~n16727 & ~n16870 ;
  assign n16872 = ~n16869 & n16871 ;
  assign n16873 = ~n16727 & ~n16872 ;
  assign n16874 = ~n16869 & ~n16872 ;
  assign n16875 = ~n16870 & n16874 ;
  assign n16876 = ~n16873 & ~n16875 ;
  assign n16877 = x90 & n4531 ;
  assign n16878 = x88 & n4847 ;
  assign n16879 = x89 & n4526 ;
  assign n16880 = ~n16878 & ~n16879 ;
  assign n16881 = ~n16877 & n16880 ;
  assign n16882 = n4534 & n4986 ;
  assign n16883 = n16881 & ~n16882 ;
  assign n16884 = x26 & ~n16883 ;
  assign n16885 = x26 & ~n16884 ;
  assign n16886 = ~n16883 & ~n16884 ;
  assign n16887 = ~n16885 & ~n16886 ;
  assign n16888 = n16876 & n16887 ;
  assign n16889 = ~n16876 & ~n16887 ;
  assign n16890 = ~n16888 & ~n16889 ;
  assign n16891 = ~n16726 & n16890 ;
  assign n16892 = n16726 & ~n16890 ;
  assign n16893 = ~n16891 & ~n16892 ;
  assign n16894 = n16725 & ~n16893 ;
  assign n16895 = ~n16725 & n16893 ;
  assign n16896 = ~n16894 & ~n16895 ;
  assign n16897 = ~n16714 & n16896 ;
  assign n16898 = n16714 & ~n16896 ;
  assign n16899 = ~n16897 & ~n16898 ;
  assign n16900 = n16713 & ~n16899 ;
  assign n16901 = ~n16713 & n16899 ;
  assign n16902 = ~n16900 & ~n16901 ;
  assign n16903 = ~n16702 & n16902 ;
  assign n16904 = n16702 & ~n16902 ;
  assign n16905 = ~n16903 & ~n16904 ;
  assign n16906 = x99 & n2093 ;
  assign n16907 = x97 & n2275 ;
  assign n16908 = x98 & n2088 ;
  assign n16909 = ~n16907 & ~n16908 ;
  assign n16910 = ~n16906 & n16909 ;
  assign n16911 = n2096 & n8660 ;
  assign n16912 = n16910 & ~n16911 ;
  assign n16913 = x17 & ~n16912 ;
  assign n16914 = x17 & ~n16913 ;
  assign n16915 = ~n16912 & ~n16913 ;
  assign n16916 = ~n16914 & ~n16915 ;
  assign n16917 = n16905 & ~n16916 ;
  assign n16918 = n16905 & ~n16917 ;
  assign n16919 = ~n16916 & ~n16917 ;
  assign n16920 = ~n16918 & ~n16919 ;
  assign n16921 = ~n16264 & ~n16271 ;
  assign n16922 = n16920 & n16921 ;
  assign n16923 = ~n16920 & ~n16921 ;
  assign n16924 = ~n16922 & ~n16923 ;
  assign n16925 = x102 & n1434 ;
  assign n16926 = x100 & n1646 ;
  assign n16927 = x101 & n1429 ;
  assign n16928 = ~n16926 & ~n16927 ;
  assign n16929 = ~n16925 & n16928 ;
  assign n16930 = n1437 & n10092 ;
  assign n16931 = n16929 & ~n16930 ;
  assign n16932 = x14 & ~n16931 ;
  assign n16933 = x14 & ~n16932 ;
  assign n16934 = ~n16931 & ~n16932 ;
  assign n16935 = ~n16933 & ~n16934 ;
  assign n16936 = n16924 & ~n16935 ;
  assign n16937 = n16924 & ~n16936 ;
  assign n16938 = ~n16935 & ~n16936 ;
  assign n16939 = ~n16937 & ~n16938 ;
  assign n16940 = ~n16284 & ~n16290 ;
  assign n16941 = n16939 & n16940 ;
  assign n16942 = ~n16939 & ~n16940 ;
  assign n16943 = ~n16941 & ~n16942 ;
  assign n16944 = x105 & n945 ;
  assign n16945 = x103 & n1099 ;
  assign n16946 = x104 & n940 ;
  assign n16947 = ~n16945 & ~n16946 ;
  assign n16948 = ~n16944 & n16947 ;
  assign n16949 = n948 & n11648 ;
  assign n16950 = n16948 & ~n16949 ;
  assign n16951 = x11 & ~n16950 ;
  assign n16952 = x11 & ~n16951 ;
  assign n16953 = ~n16950 & ~n16951 ;
  assign n16954 = ~n16952 & ~n16953 ;
  assign n16955 = n16943 & ~n16954 ;
  assign n16956 = n16943 & ~n16955 ;
  assign n16957 = ~n16954 & ~n16955 ;
  assign n16958 = ~n16956 & ~n16957 ;
  assign n16959 = ~n16303 & ~n16309 ;
  assign n16960 = n16958 & n16959 ;
  assign n16961 = ~n16958 & ~n16959 ;
  assign n16962 = ~n16960 & ~n16961 ;
  assign n16963 = x108 & n574 ;
  assign n16964 = x106 & n673 ;
  assign n16965 = x107 & n569 ;
  assign n16966 = ~n16964 & ~n16965 ;
  assign n16967 = ~n16963 & n16966 ;
  assign n16968 = n577 & n13323 ;
  assign n16969 = n16967 & ~n16968 ;
  assign n16970 = x8 & ~n16969 ;
  assign n16971 = x8 & ~n16970 ;
  assign n16972 = ~n16969 & ~n16970 ;
  assign n16973 = ~n16971 & ~n16972 ;
  assign n16974 = n16962 & ~n16973 ;
  assign n16975 = ~n16962 & n16973 ;
  assign n16976 = ~n16701 & ~n16975 ;
  assign n16977 = ~n16974 & n16976 ;
  assign n16978 = ~n16701 & ~n16977 ;
  assign n16979 = ~n16974 & ~n16977 ;
  assign n16980 = ~n16975 & n16979 ;
  assign n16981 = ~n16978 & ~n16980 ;
  assign n16982 = x111 & n293 ;
  assign n16983 = x109 & n373 ;
  assign n16984 = x110 & n288 ;
  assign n16985 = ~n16983 & ~n16984 ;
  assign n16986 = ~n16982 & n16985 ;
  assign n16987 = n296 & n15111 ;
  assign n16988 = n16986 & ~n16987 ;
  assign n16989 = x5 & ~n16988 ;
  assign n16990 = x5 & ~n16989 ;
  assign n16991 = ~n16988 & ~n16989 ;
  assign n16992 = ~n16990 & ~n16991 ;
  assign n16993 = ~n16981 & ~n16992 ;
  assign n16994 = ~n16981 & ~n16993 ;
  assign n16995 = ~n16992 & ~n16993 ;
  assign n16996 = ~n16994 & ~n16995 ;
  assign n16997 = ~n16342 & ~n16348 ;
  assign n16998 = n16996 & n16997 ;
  assign n16999 = ~n16996 & ~n16997 ;
  assign n17000 = ~n16998 & ~n16999 ;
  assign n17001 = x114 & n146 ;
  assign n17002 = x112 & n182 ;
  assign n17003 = x113 & n141 ;
  assign n17004 = ~n17002 & ~n17003 ;
  assign n17005 = ~n17001 & n17004 ;
  assign n17006 = ~n16357 & ~n16359 ;
  assign n17007 = ~x113 & ~x114 ;
  assign n17008 = x113 & x114 ;
  assign n17009 = ~n17007 & ~n17008 ;
  assign n17010 = ~n17006 & n17009 ;
  assign n17011 = n17006 & ~n17009 ;
  assign n17012 = ~n17010 & ~n17011 ;
  assign n17013 = n149 & n17012 ;
  assign n17014 = n17005 & ~n17013 ;
  assign n17015 = x2 & ~n17014 ;
  assign n17016 = x2 & ~n17015 ;
  assign n17017 = ~n17014 & ~n17015 ;
  assign n17018 = ~n17016 & ~n17017 ;
  assign n17019 = n17000 & ~n17018 ;
  assign n17020 = n17000 & ~n17019 ;
  assign n17021 = ~n17018 & ~n17019 ;
  assign n17022 = ~n17020 & ~n17021 ;
  assign n17023 = ~n16369 & ~n16371 ;
  assign n17024 = ~n17022 & ~n17023 ;
  assign n17025 = n17022 & n17023 ;
  assign n17026 = ~n17024 & ~n17025 ;
  assign n17349 = n17026 & x178 ;
  assign n17027 = ~n16648 & ~n16655 ;
  assign n17028 = ~n16571 & ~n16577 ;
  assign n17029 = ~x96 & n2751 ;
  assign n17030 = ~x94 & n3020 ;
  assign n17031 = ~x95 & n2746 ;
  assign n17032 = ~n17030 & ~n17031 ;
  assign n17033 = ~n17029 & n17032 ;
  assign n17034 = n2754 & n7531 ;
  assign n17035 = n17033 & ~n17034 ;
  assign n17036 = ~x20 & ~n17035 ;
  assign n17037 = ~x20 & ~n17036 ;
  assign n17038 = ~n17035 & ~n17036 ;
  assign n17039 = ~n17037 & ~n17038 ;
  assign n17040 = ~n16552 & ~n16556 ;
  assign n17041 = ~x93 & n3589 ;
  assign n17042 = ~x91 & n3878 ;
  assign n17043 = ~x92 & n3584 ;
  assign n17044 = ~n17042 & ~n17043 ;
  assign n17045 = ~n17041 & n17044 ;
  assign n17046 = n3592 & n6285 ;
  assign n17047 = n17045 & ~n17046 ;
  assign n17048 = ~x23 & ~n17047 ;
  assign n17049 = ~x23 & ~n17048 ;
  assign n17050 = ~n17047 & ~n17048 ;
  assign n17051 = ~n17049 & ~n17050 ;
  assign n17052 = ~n16544 & ~n16549 ;
  assign n17053 = ~n16525 & ~n16531 ;
  assign n17054 = ~n16487 & ~n16493 ;
  assign n17055 = ~x81 & n8006 ;
  assign n17056 = ~x79 & n8474 ;
  assign n17057 = ~x80 & n8001 ;
  assign n17058 = ~n17056 & ~n17057 ;
  assign n17059 = ~n17055 & n17058 ;
  assign n17060 = n2460 & n8009 ;
  assign n17061 = n17059 & ~n17060 ;
  assign n17062 = ~x35 & ~n17061 ;
  assign n17063 = ~x35 & ~n17062 ;
  assign n17064 = ~n17061 & ~n17062 ;
  assign n17065 = ~n17063 & ~n17064 ;
  assign n17066 = ~n16471 & ~n16473 ;
  assign n17067 = ~n16432 & ~n16438 ;
  assign n17068 = ~x72 & n12506 ;
  assign n17069 = ~x70 & n13131 ;
  assign n17070 = ~x71 & n12501 ;
  assign n17071 = ~n17069 & ~n17070 ;
  assign n17072 = ~n17068 & n17071 ;
  assign n17073 = n773 & n12509 ;
  assign n17074 = n17072 & ~n17073 ;
  assign n17075 = ~x44 & ~n17074 ;
  assign n17076 = ~x44 & ~n17075 ;
  assign n17077 = ~n17074 & ~n17075 ;
  assign n17078 = ~n17076 & ~n17077 ;
  assign n17079 = ~n16416 & ~n16418 ;
  assign n17080 = ~x66 & n16076 ;
  assign n17081 = ~x64 & n16756 ;
  assign n17082 = ~x65 & n16071 ;
  assign n17083 = ~n17081 & ~n17082 ;
  assign n17084 = ~n17080 & n17083 ;
  assign n17085 = n214 & n16079 ;
  assign n17086 = n17084 & ~n17085 ;
  assign n17087 = ~x50 & ~n17086 ;
  assign n17088 = ~x50 & ~n17087 ;
  assign n17089 = ~n17086 & ~n17087 ;
  assign n17090 = ~n17088 & ~n17089 ;
  assign n17091 = ~n16412 & n17090 ;
  assign n17092 = n16412 & ~n17090 ;
  assign n17093 = ~n17091 & ~n17092 ;
  assign n17094 = ~x69 & n14233 ;
  assign n17095 = ~x67 & n14876 ;
  assign n17096 = ~x68 & n14228 ;
  assign n17097 = ~n17095 & ~n17096 ;
  assign n17098 = ~n17094 & n17097 ;
  assign n17099 = n435 & n14236 ;
  assign n17100 = n17098 & ~n17099 ;
  assign n17101 = ~x47 & ~n17100 ;
  assign n17102 = ~x47 & ~n17101 ;
  assign n17103 = ~n17100 & ~n17101 ;
  assign n17104 = ~n17102 & ~n17103 ;
  assign n17105 = n17093 & ~n17104 ;
  assign n17106 = n17093 & ~n17105 ;
  assign n17107 = ~n17104 & ~n17105 ;
  assign n17108 = ~n17106 & ~n17107 ;
  assign n17109 = ~n17079 & ~n17108 ;
  assign n17110 = n17079 & n17108 ;
  assign n17111 = ~n17109 & ~n17110 ;
  assign n17112 = ~n17078 & n17111 ;
  assign n17113 = ~n17078 & ~n17112 ;
  assign n17114 = n17111 & ~n17112 ;
  assign n17115 = ~n17113 & ~n17114 ;
  assign n17116 = ~n17067 & ~n17115 ;
  assign n17117 = ~n17067 & ~n17116 ;
  assign n17118 = ~n17115 & ~n17116 ;
  assign n17119 = ~n17117 & ~n17118 ;
  assign n17120 = ~x75 & n10905 ;
  assign n17121 = ~x73 & n11466 ;
  assign n17122 = ~x74 & n10900 ;
  assign n17123 = ~n17121 & ~n17122 ;
  assign n17124 = ~n17120 & n17123 ;
  assign n17125 = n1225 & n10908 ;
  assign n17126 = n17124 & ~n17125 ;
  assign n17127 = ~x41 & ~n17126 ;
  assign n17128 = ~x41 & ~n17127 ;
  assign n17129 = ~n17126 & ~n17127 ;
  assign n17130 = ~n17128 & ~n17129 ;
  assign n17131 = n17119 & n17130 ;
  assign n17132 = ~n17119 & ~n17130 ;
  assign n17133 = ~n17131 & ~n17132 ;
  assign n17134 = ~n16456 & n17133 ;
  assign n17135 = n16456 & ~n17133 ;
  assign n17136 = ~n17134 & ~n17135 ;
  assign n17137 = ~x78 & n9433 ;
  assign n17138 = ~x76 & n9915 ;
  assign n17139 = ~x77 & n9428 ;
  assign n17140 = ~n17138 & ~n17139 ;
  assign n17141 = ~n17137 & n17140 ;
  assign n17142 = n1718 & n9436 ;
  assign n17143 = n17141 & ~n17142 ;
  assign n17144 = ~x38 & ~n17143 ;
  assign n17145 = ~x38 & ~n17144 ;
  assign n17146 = ~n17143 & ~n17144 ;
  assign n17147 = ~n17145 & ~n17146 ;
  assign n17148 = n17136 & ~n17147 ;
  assign n17149 = n17136 & ~n17148 ;
  assign n17150 = ~n17147 & ~n17148 ;
  assign n17151 = ~n17149 & ~n17150 ;
  assign n17152 = ~n17066 & ~n17151 ;
  assign n17153 = n17066 & n17151 ;
  assign n17154 = ~n17152 & ~n17153 ;
  assign n17155 = ~n17065 & n17154 ;
  assign n17156 = ~n17065 & ~n17155 ;
  assign n17157 = n17154 & ~n17155 ;
  assign n17158 = ~n17156 & ~n17157 ;
  assign n17159 = ~n17054 & ~n17158 ;
  assign n17160 = ~n17054 & ~n17159 ;
  assign n17161 = ~n17158 & ~n17159 ;
  assign n17162 = ~n17160 & ~n17161 ;
  assign n17163 = ~x84 & n6725 ;
  assign n17164 = ~x82 & n7129 ;
  assign n17165 = ~x83 & n6720 ;
  assign n17166 = ~n17164 & ~n17165 ;
  assign n17167 = ~n17163 & n17166 ;
  assign n17168 = n3247 & n6728 ;
  assign n17169 = n17167 & ~n17168 ;
  assign n17170 = ~x32 & ~n17169 ;
  assign n17171 = ~x32 & ~n17170 ;
  assign n17172 = ~n17169 & ~n17170 ;
  assign n17173 = ~n17171 & ~n17172 ;
  assign n17174 = ~n17162 & ~n17173 ;
  assign n17175 = ~n17162 & ~n17174 ;
  assign n17176 = ~n17173 & ~n17174 ;
  assign n17177 = ~n17175 & ~n17176 ;
  assign n17178 = ~n16506 & ~n16512 ;
  assign n17179 = n17177 & n17178 ;
  assign n17180 = ~n17177 & ~n17178 ;
  assign n17181 = ~n17179 & ~n17180 ;
  assign n17182 = ~x87 & n5560 ;
  assign n17183 = ~x85 & n5943 ;
  assign n17184 = ~x86 & n5555 ;
  assign n17185 = ~n17183 & ~n17184 ;
  assign n17186 = ~n17182 & n17185 ;
  assign n17187 = n4143 & n5563 ;
  assign n17188 = n17186 & ~n17187 ;
  assign n17189 = ~x29 & ~n17188 ;
  assign n17190 = ~x29 & ~n17189 ;
  assign n17191 = ~n17188 & ~n17189 ;
  assign n17192 = ~n17190 & ~n17191 ;
  assign n17193 = n17181 & ~n17192 ;
  assign n17194 = ~n17181 & n17192 ;
  assign n17195 = ~n17053 & ~n17194 ;
  assign n17196 = ~n17193 & n17195 ;
  assign n17197 = ~n17053 & ~n17196 ;
  assign n17198 = ~n17193 & ~n17196 ;
  assign n17199 = ~n17194 & n17198 ;
  assign n17200 = ~n17197 & ~n17199 ;
  assign n17201 = ~x90 & n4531 ;
  assign n17202 = ~x88 & n4847 ;
  assign n17203 = ~x89 & n4526 ;
  assign n17204 = ~n17202 & ~n17203 ;
  assign n17205 = ~n17201 & n17204 ;
  assign n17206 = n4534 & n5155 ;
  assign n17207 = n17205 & ~n17206 ;
  assign n17208 = ~x26 & ~n17207 ;
  assign n17209 = ~x26 & ~n17208 ;
  assign n17210 = ~n17207 & ~n17208 ;
  assign n17211 = ~n17209 & ~n17210 ;
  assign n17212 = n17200 & n17211 ;
  assign n17213 = ~n17200 & ~n17211 ;
  assign n17214 = ~n17212 & ~n17213 ;
  assign n17215 = ~n17052 & n17214 ;
  assign n17216 = n17052 & ~n17214 ;
  assign n17217 = ~n17215 & ~n17216 ;
  assign n17218 = n17051 & ~n17217 ;
  assign n17219 = ~n17051 & n17217 ;
  assign n17220 = ~n17218 & ~n17219 ;
  assign n17221 = ~n17040 & n17220 ;
  assign n17222 = n17040 & ~n17220 ;
  assign n17223 = ~n17221 & ~n17222 ;
  assign n17224 = n17039 & ~n17223 ;
  assign n17225 = ~n17039 & n17223 ;
  assign n17226 = ~n17224 & ~n17225 ;
  assign n17227 = ~n17028 & n17226 ;
  assign n17228 = n17028 & ~n17226 ;
  assign n17229 = ~n17227 & ~n17228 ;
  assign n17230 = ~x99 & n2093 ;
  assign n17231 = ~x97 & n2275 ;
  assign n17232 = ~x98 & n2088 ;
  assign n17233 = ~n17231 & ~n17232 ;
  assign n17234 = ~n17230 & n17233 ;
  assign n17235 = n2096 & n8885 ;
  assign n17236 = n17234 & ~n17235 ;
  assign n17237 = ~x17 & ~n17236 ;
  assign n17238 = ~x17 & ~n17237 ;
  assign n17239 = ~n17236 & ~n17237 ;
  assign n17240 = ~n17238 & ~n17239 ;
  assign n17241 = n17229 & ~n17240 ;
  assign n17242 = n17229 & ~n17241 ;
  assign n17243 = ~n17240 & ~n17241 ;
  assign n17244 = ~n17242 & ~n17243 ;
  assign n17245 = ~n16590 & ~n16597 ;
  assign n17246 = n17244 & n17245 ;
  assign n17247 = ~n17244 & ~n17245 ;
  assign n17248 = ~n17246 & ~n17247 ;
  assign n17249 = ~x102 & n1434 ;
  assign n17250 = ~x100 & n1646 ;
  assign n17251 = ~x101 & n1429 ;
  assign n17252 = ~n17250 & ~n17251 ;
  assign n17253 = ~n17249 & n17252 ;
  assign n17254 = n1437 & n10333 ;
  assign n17255 = n17253 & ~n17254 ;
  assign n17256 = ~x14 & ~n17255 ;
  assign n17257 = ~x14 & ~n17256 ;
  assign n17258 = ~n17255 & ~n17256 ;
  assign n17259 = ~n17257 & ~n17258 ;
  assign n17260 = n17248 & ~n17259 ;
  assign n17261 = n17248 & ~n17260 ;
  assign n17262 = ~n17259 & ~n17260 ;
  assign n17263 = ~n17261 & ~n17262 ;
  assign n17264 = ~n16610 & ~n16616 ;
  assign n17265 = n17263 & n17264 ;
  assign n17266 = ~n17263 & ~n17264 ;
  assign n17267 = ~n17265 & ~n17266 ;
  assign n17268 = ~x105 & n945 ;
  assign n17269 = ~x103 & n1099 ;
  assign n17270 = ~x104 & n940 ;
  assign n17271 = ~n17269 & ~n17270 ;
  assign n17272 = ~n17268 & n17271 ;
  assign n17273 = n948 & n11907 ;
  assign n17274 = n17272 & ~n17273 ;
  assign n17275 = ~x11 & ~n17274 ;
  assign n17276 = ~x11 & ~n17275 ;
  assign n17277 = ~n17274 & ~n17275 ;
  assign n17278 = ~n17276 & ~n17277 ;
  assign n17279 = n17267 & ~n17278 ;
  assign n17280 = n17267 & ~n17279 ;
  assign n17281 = ~n17278 & ~n17279 ;
  assign n17282 = ~n17280 & ~n17281 ;
  assign n17283 = ~n16629 & ~n16635 ;
  assign n17284 = n17282 & n17283 ;
  assign n17285 = ~n17282 & ~n17283 ;
  assign n17286 = ~n17284 & ~n17285 ;
  assign n17287 = ~x108 & n574 ;
  assign n17288 = ~x106 & n673 ;
  assign n17289 = ~x107 & n569 ;
  assign n17290 = ~n17288 & ~n17289 ;
  assign n17291 = ~n17287 & n17290 ;
  assign n17292 = n577 & n13601 ;
  assign n17293 = n17291 & ~n17292 ;
  assign n17294 = ~x8 & ~n17293 ;
  assign n17295 = ~x8 & ~n17294 ;
  assign n17296 = ~n17293 & ~n17294 ;
  assign n17297 = ~n17295 & ~n17296 ;
  assign n17298 = n17286 & ~n17297 ;
  assign n17299 = ~n17286 & n17297 ;
  assign n17300 = ~n17027 & ~n17299 ;
  assign n17301 = ~n17298 & n17300 ;
  assign n17302 = ~n17027 & ~n17301 ;
  assign n17303 = ~n17298 & ~n17301 ;
  assign n17304 = ~n17299 & n17303 ;
  assign n17305 = ~n17302 & ~n17304 ;
  assign n17306 = ~x111 & n293 ;
  assign n17307 = ~x109 & n373 ;
  assign n17308 = ~x110 & n288 ;
  assign n17309 = ~n17307 & ~n17308 ;
  assign n17310 = ~n17306 & n17309 ;
  assign n17311 = n296 & n15411 ;
  assign n17312 = n17310 & ~n17311 ;
  assign n17313 = ~x5 & ~n17312 ;
  assign n17314 = ~x5 & ~n17313 ;
  assign n17315 = ~n17312 & ~n17313 ;
  assign n17316 = ~n17314 & ~n17315 ;
  assign n17317 = ~n17305 & ~n17316 ;
  assign n17318 = ~n17305 & ~n17317 ;
  assign n17319 = ~n17316 & ~n17317 ;
  assign n17320 = ~n17318 & ~n17319 ;
  assign n17321 = ~n16668 & ~n16674 ;
  assign n17322 = n17320 & n17321 ;
  assign n17323 = ~n17320 & ~n17321 ;
  assign n17324 = ~n17322 & ~n17323 ;
  assign n17325 = ~x114 & n164 ;
  assign n17326 = ~x112 & n205 ;
  assign n17327 = ~x113 & n162 ;
  assign n17328 = ~n17326 & ~n17327 ;
  assign n17329 = ~n17325 & n17328 ;
  assign n17330 = ~n16356 & ~n16682 ;
  assign n17331 = n17009 & ~n17330 ;
  assign n17332 = ~n17009 & n17330 ;
  assign n17333 = ~n17331 & ~n17332 ;
  assign n17334 = n167 & n17333 ;
  assign n17335 = n17329 & ~n17334 ;
  assign n17336 = ~x2 & ~n17335 ;
  assign n17337 = ~x2 & ~n17336 ;
  assign n17338 = ~n17335 & ~n17336 ;
  assign n17339 = ~n17337 & ~n17338 ;
  assign n17340 = n17324 & ~n17339 ;
  assign n17341 = n17324 & ~n17340 ;
  assign n17342 = ~n17339 & ~n17340 ;
  assign n17343 = ~n17341 & ~n17342 ;
  assign n17344 = ~n16692 & ~n16694 ;
  assign n17345 = ~n17343 & ~n17344 ;
  assign n17346 = n17343 & n17344 ;
  assign n17347 = ~n17345 & ~n17346 ;
  assign n17350 = ~n17347 & ~x178 ;
  assign n17351 = ~n17349 & ~n17350 ;
  assign n17352 = ~n17019 & ~n17024 ;
  assign n17353 = x115 & n146 ;
  assign n17354 = x113 & n182 ;
  assign n17355 = x114 & n141 ;
  assign n17356 = ~n17354 & ~n17355 ;
  assign n17357 = ~n17353 & n17356 ;
  assign n17358 = ~n17008 & ~n17010 ;
  assign n17359 = ~x114 & ~x115 ;
  assign n17360 = x114 & x115 ;
  assign n17361 = ~n17359 & ~n17360 ;
  assign n17362 = ~n17358 & n17361 ;
  assign n17363 = n17358 & ~n17361 ;
  assign n17364 = ~n17362 & ~n17363 ;
  assign n17365 = n149 & n17364 ;
  assign n17366 = n17357 & ~n17365 ;
  assign n17367 = x2 & ~n17366 ;
  assign n17368 = x2 & ~n17367 ;
  assign n17369 = ~n17366 & ~n17367 ;
  assign n17370 = ~n17368 & ~n17369 ;
  assign n17371 = ~n16993 & ~n16999 ;
  assign n17372 = ~n16917 & ~n16923 ;
  assign n17373 = ~n16901 & ~n16903 ;
  assign n17374 = ~n16895 & ~n16897 ;
  assign n17375 = ~n16889 & ~n16891 ;
  assign n17376 = ~n16831 & ~n16835 ;
  assign n17377 = x82 & n8006 ;
  assign n17378 = x80 & n8474 ;
  assign n17379 = x81 & n8001 ;
  assign n17380 = ~n17378 & ~n17379 ;
  assign n17381 = ~n17377 & n17380 ;
  assign n17382 = n2584 & n8009 ;
  assign n17383 = n17381 & ~n17382 ;
  assign n17384 = x35 & ~n17383 ;
  assign n17385 = x35 & ~n17384 ;
  assign n17386 = ~n17383 & ~n17384 ;
  assign n17387 = ~n17385 & ~n17386 ;
  assign n17388 = ~n16824 & ~n16828 ;
  assign n17389 = x79 & n9433 ;
  assign n17390 = x77 & n9915 ;
  assign n17391 = x78 & n9428 ;
  assign n17392 = ~n17390 & ~n17391 ;
  assign n17393 = ~n17389 & n17392 ;
  assign n17394 = n1817 & n9436 ;
  assign n17395 = n17393 & ~n17394 ;
  assign n17396 = x38 & ~n17395 ;
  assign n17397 = x38 & ~n17396 ;
  assign n17398 = ~n17395 & ~n17396 ;
  assign n17399 = ~n17397 & ~n17398 ;
  assign n17400 = ~n16808 & ~n16810 ;
  assign n17401 = x76 & n10905 ;
  assign n17402 = x74 & n11466 ;
  assign n17403 = x75 & n10900 ;
  assign n17404 = ~n17402 & ~n17403 ;
  assign n17405 = ~n17401 & n17404 ;
  assign n17406 = n1311 & n10908 ;
  assign n17407 = n17405 & ~n17406 ;
  assign n17408 = x41 & ~n17407 ;
  assign n17409 = x41 & ~n17408 ;
  assign n17410 = ~n17407 & ~n17408 ;
  assign n17411 = ~n17409 & ~n17410 ;
  assign n17412 = ~n16788 & ~n16792 ;
  assign n17413 = x50 & ~x51 ;
  assign n17414 = ~x50 & x51 ;
  assign n17415 = ~n17413 & ~n17414 ;
  assign n17416 = x64 & ~n17415 ;
  assign n17417 = ~n16768 & n17416 ;
  assign n17418 = n16768 & ~n17416 ;
  assign n17419 = ~n17417 & ~n17418 ;
  assign n17420 = x67 & n16076 ;
  assign n17421 = x65 & n16756 ;
  assign n17422 = x66 & n16071 ;
  assign n17423 = ~n17421 & ~n17422 ;
  assign n17424 = ~n17420 & n17423 ;
  assign n17425 = n240 & n16079 ;
  assign n17426 = n17424 & ~n17425 ;
  assign n17427 = x50 & ~n17426 ;
  assign n17428 = x50 & ~n17427 ;
  assign n17429 = ~n17426 & ~n17427 ;
  assign n17430 = ~n17428 & ~n17429 ;
  assign n17431 = ~n17419 & ~n17430 ;
  assign n17432 = n17419 & n17430 ;
  assign n17433 = ~n17431 & ~n17432 ;
  assign n17434 = x70 & n14233 ;
  assign n17435 = x68 & n14876 ;
  assign n17436 = x69 & n14228 ;
  assign n17437 = ~n17435 & ~n17436 ;
  assign n17438 = ~n17434 & n17437 ;
  assign n17439 = n488 & n14236 ;
  assign n17440 = n17438 & ~n17439 ;
  assign n17441 = x47 & ~n17440 ;
  assign n17442 = x47 & ~n17441 ;
  assign n17443 = ~n17440 & ~n17441 ;
  assign n17444 = ~n17442 & ~n17443 ;
  assign n17445 = n17433 & ~n17444 ;
  assign n17446 = n17433 & ~n17445 ;
  assign n17447 = ~n17444 & ~n17445 ;
  assign n17448 = ~n17446 & ~n17447 ;
  assign n17449 = ~n16781 & ~n16785 ;
  assign n17450 = n17448 & n17449 ;
  assign n17451 = ~n17448 & ~n17449 ;
  assign n17452 = ~n17450 & ~n17451 ;
  assign n17453 = x73 & n12506 ;
  assign n17454 = x71 & n13131 ;
  assign n17455 = x72 & n12501 ;
  assign n17456 = ~n17454 & ~n17455 ;
  assign n17457 = ~n17453 & n17456 ;
  assign n17458 = n843 & n12509 ;
  assign n17459 = n17457 & ~n17458 ;
  assign n17460 = x44 & ~n17459 ;
  assign n17461 = x44 & ~n17460 ;
  assign n17462 = ~n17459 & ~n17460 ;
  assign n17463 = ~n17461 & ~n17462 ;
  assign n17464 = ~n17452 & n17463 ;
  assign n17465 = n17452 & ~n17463 ;
  assign n17466 = ~n17464 & ~n17465 ;
  assign n17467 = ~n17412 & n17466 ;
  assign n17468 = n17412 & ~n17466 ;
  assign n17469 = ~n17467 & ~n17468 ;
  assign n17470 = ~n17411 & n17469 ;
  assign n17471 = ~n17411 & ~n17470 ;
  assign n17472 = n17469 & ~n17470 ;
  assign n17473 = ~n17471 & ~n17472 ;
  assign n17474 = ~n17400 & ~n17473 ;
  assign n17475 = n17400 & ~n17472 ;
  assign n17476 = ~n17471 & n17475 ;
  assign n17477 = ~n17474 & ~n17476 ;
  assign n17478 = ~n17399 & n17477 ;
  assign n17479 = n17399 & ~n17477 ;
  assign n17480 = ~n17478 & ~n17479 ;
  assign n17481 = ~n17388 & n17480 ;
  assign n17482 = n17388 & ~n17480 ;
  assign n17483 = ~n17481 & ~n17482 ;
  assign n17484 = ~n17387 & n17483 ;
  assign n17485 = n17387 & ~n17483 ;
  assign n17486 = ~n17484 & ~n17485 ;
  assign n17487 = ~n17376 & n17486 ;
  assign n17488 = n17376 & ~n17486 ;
  assign n17489 = ~n17487 & ~n17488 ;
  assign n17490 = x85 & n6725 ;
  assign n17491 = x83 & n7129 ;
  assign n17492 = x84 & n6720 ;
  assign n17493 = ~n17491 & ~n17492 ;
  assign n17494 = ~n17490 & n17493 ;
  assign n17495 = n3389 & n6728 ;
  assign n17496 = n17494 & ~n17495 ;
  assign n17497 = x32 & ~n17496 ;
  assign n17498 = x32 & ~n17497 ;
  assign n17499 = ~n17496 & ~n17497 ;
  assign n17500 = ~n17498 & ~n17499 ;
  assign n17501 = n17489 & ~n17500 ;
  assign n17502 = n17489 & ~n17501 ;
  assign n17503 = ~n17500 & ~n17501 ;
  assign n17504 = ~n17502 & ~n17503 ;
  assign n17505 = ~n16850 & ~n16856 ;
  assign n17506 = n17504 & n17505 ;
  assign n17507 = ~n17504 & ~n17505 ;
  assign n17508 = ~n17506 & ~n17507 ;
  assign n17509 = x88 & n5560 ;
  assign n17510 = x86 & n5943 ;
  assign n17511 = x87 & n5555 ;
  assign n17512 = ~n17510 & ~n17511 ;
  assign n17513 = ~n17509 & n17512 ;
  assign n17514 = n4305 & n5563 ;
  assign n17515 = n17513 & ~n17514 ;
  assign n17516 = x29 & ~n17515 ;
  assign n17517 = x29 & ~n17516 ;
  assign n17518 = ~n17515 & ~n17516 ;
  assign n17519 = ~n17517 & ~n17518 ;
  assign n17520 = ~n17508 & n17519 ;
  assign n17521 = n17508 & ~n17519 ;
  assign n17522 = ~n17520 & ~n17521 ;
  assign n17523 = ~n16874 & n17522 ;
  assign n17524 = n16874 & ~n17522 ;
  assign n17525 = ~n17523 & ~n17524 ;
  assign n17526 = x91 & n4531 ;
  assign n17527 = x89 & n4847 ;
  assign n17528 = x90 & n4526 ;
  assign n17529 = ~n17527 & ~n17528 ;
  assign n17530 = ~n17526 & n17529 ;
  assign n17531 = n4534 & n5336 ;
  assign n17532 = n17530 & ~n17531 ;
  assign n17533 = x26 & ~n17532 ;
  assign n17534 = x26 & ~n17533 ;
  assign n17535 = ~n17532 & ~n17533 ;
  assign n17536 = ~n17534 & ~n17535 ;
  assign n17537 = n17525 & ~n17536 ;
  assign n17538 = n17525 & ~n17537 ;
  assign n17539 = ~n17536 & ~n17537 ;
  assign n17540 = ~n17538 & ~n17539 ;
  assign n17541 = ~n17375 & n17540 ;
  assign n17542 = n17375 & ~n17540 ;
  assign n17543 = ~n17541 & ~n17542 ;
  assign n17544 = x94 & n3589 ;
  assign n17545 = x92 & n3878 ;
  assign n17546 = x93 & n3584 ;
  assign n17547 = ~n17545 & ~n17546 ;
  assign n17548 = ~n17544 & n17547 ;
  assign n17549 = n3592 & n6483 ;
  assign n17550 = n17548 & ~n17549 ;
  assign n17551 = x23 & ~n17550 ;
  assign n17552 = x23 & ~n17551 ;
  assign n17553 = ~n17550 & ~n17551 ;
  assign n17554 = ~n17552 & ~n17553 ;
  assign n17555 = ~n17543 & ~n17554 ;
  assign n17556 = n17543 & n17554 ;
  assign n17557 = ~n17555 & ~n17556 ;
  assign n17558 = ~n17374 & n17557 ;
  assign n17559 = n17374 & ~n17557 ;
  assign n17560 = ~n17558 & ~n17559 ;
  assign n17561 = x97 & n2751 ;
  assign n17562 = x95 & n3020 ;
  assign n17563 = x96 & n2746 ;
  assign n17564 = ~n17562 & ~n17563 ;
  assign n17565 = ~n17561 & n17564 ;
  assign n17566 = n2754 & n7745 ;
  assign n17567 = n17565 & ~n17566 ;
  assign n17568 = x20 & ~n17567 ;
  assign n17569 = x20 & ~n17568 ;
  assign n17570 = ~n17567 & ~n17568 ;
  assign n17571 = ~n17569 & ~n17570 ;
  assign n17572 = n17560 & ~n17571 ;
  assign n17573 = n17560 & ~n17572 ;
  assign n17574 = ~n17571 & ~n17572 ;
  assign n17575 = ~n17573 & ~n17574 ;
  assign n17576 = ~n17373 & n17575 ;
  assign n17577 = n17373 & ~n17575 ;
  assign n17578 = ~n17576 & ~n17577 ;
  assign n17579 = x100 & n2093 ;
  assign n17580 = x98 & n2275 ;
  assign n17581 = x99 & n2088 ;
  assign n17582 = ~n17580 & ~n17581 ;
  assign n17583 = ~n17579 & n17582 ;
  assign n17584 = n2096 & n9115 ;
  assign n17585 = n17583 & ~n17584 ;
  assign n17586 = x17 & ~n17585 ;
  assign n17587 = x17 & ~n17586 ;
  assign n17588 = ~n17585 & ~n17586 ;
  assign n17589 = ~n17587 & ~n17588 ;
  assign n17590 = ~n17578 & ~n17589 ;
  assign n17591 = n17578 & n17589 ;
  assign n17592 = ~n17590 & ~n17591 ;
  assign n17593 = n17372 & ~n17592 ;
  assign n17594 = ~n17372 & n17592 ;
  assign n17595 = ~n17593 & ~n17594 ;
  assign n17596 = x103 & n1434 ;
  assign n17597 = x101 & n1646 ;
  assign n17598 = x102 & n1429 ;
  assign n17599 = ~n17597 & ~n17598 ;
  assign n17600 = ~n17596 & n17599 ;
  assign n17601 = n1437 & n10588 ;
  assign n17602 = n17600 & ~n17601 ;
  assign n17603 = x14 & ~n17602 ;
  assign n17604 = x14 & ~n17603 ;
  assign n17605 = ~n17602 & ~n17603 ;
  assign n17606 = ~n17604 & ~n17605 ;
  assign n17607 = n17595 & ~n17606 ;
  assign n17608 = n17595 & ~n17607 ;
  assign n17609 = ~n17606 & ~n17607 ;
  assign n17610 = ~n17608 & ~n17609 ;
  assign n17611 = ~n16936 & ~n16942 ;
  assign n17612 = n17610 & n17611 ;
  assign n17613 = ~n17610 & ~n17611 ;
  assign n17614 = ~n17612 & ~n17613 ;
  assign n17615 = x106 & n945 ;
  assign n17616 = x104 & n1099 ;
  assign n17617 = x105 & n940 ;
  assign n17618 = ~n17616 & ~n17617 ;
  assign n17619 = ~n17615 & n17618 ;
  assign n17620 = n948 & n12181 ;
  assign n17621 = n17619 & ~n17620 ;
  assign n17622 = x11 & ~n17621 ;
  assign n17623 = x11 & ~n17622 ;
  assign n17624 = ~n17621 & ~n17622 ;
  assign n17625 = ~n17623 & ~n17624 ;
  assign n17626 = ~n17614 & n17625 ;
  assign n17627 = n17614 & ~n17625 ;
  assign n17628 = ~n17626 & ~n17627 ;
  assign n17629 = ~n16955 & ~n16961 ;
  assign n17630 = n17628 & ~n17629 ;
  assign n17631 = ~n17628 & n17629 ;
  assign n17632 = ~n17630 & ~n17631 ;
  assign n17633 = x109 & n574 ;
  assign n17634 = x107 & n673 ;
  assign n17635 = x108 & n569 ;
  assign n17636 = ~n17634 & ~n17635 ;
  assign n17637 = ~n17633 & n17636 ;
  assign n17638 = n577 & n13894 ;
  assign n17639 = n17637 & ~n17638 ;
  assign n17640 = x8 & ~n17639 ;
  assign n17641 = x8 & ~n17640 ;
  assign n17642 = ~n17639 & ~n17640 ;
  assign n17643 = ~n17641 & ~n17642 ;
  assign n17644 = n17632 & ~n17643 ;
  assign n17645 = n17632 & ~n17644 ;
  assign n17646 = ~n17643 & ~n17644 ;
  assign n17647 = ~n17645 & ~n17646 ;
  assign n17648 = ~n16979 & n17647 ;
  assign n17649 = n16979 & ~n17647 ;
  assign n17650 = ~n17648 & ~n17649 ;
  assign n17651 = x112 & n293 ;
  assign n17652 = x110 & n373 ;
  assign n17653 = x111 & n288 ;
  assign n17654 = ~n17652 & ~n17653 ;
  assign n17655 = ~n17651 & n17654 ;
  assign n17656 = n296 & n15442 ;
  assign n17657 = n17655 & ~n17656 ;
  assign n17658 = x5 & ~n17657 ;
  assign n17659 = x5 & ~n17658 ;
  assign n17660 = ~n17657 & ~n17658 ;
  assign n17661 = ~n17659 & ~n17660 ;
  assign n17662 = n17650 & n17661 ;
  assign n17663 = ~n17650 & ~n17661 ;
  assign n17664 = ~n17662 & ~n17663 ;
  assign n17665 = ~n17371 & n17664 ;
  assign n17666 = n17371 & ~n17664 ;
  assign n17667 = ~n17665 & ~n17666 ;
  assign n17668 = ~n17370 & n17667 ;
  assign n17669 = n17370 & ~n17667 ;
  assign n17670 = ~n17668 & ~n17669 ;
  assign n17671 = ~n17352 & n17670 ;
  assign n17672 = n17352 & ~n17670 ;
  assign n17673 = ~n17671 & ~n17672 ;
  assign n17991 = n17673 & x179 ;
  assign n17674 = ~n17340 & ~n17345 ;
  assign n17675 = ~x115 & n164 ;
  assign n17676 = ~x113 & n205 ;
  assign n17677 = ~x114 & n162 ;
  assign n17678 = ~n17676 & ~n17677 ;
  assign n17679 = ~n17675 & n17678 ;
  assign n17680 = ~n17007 & ~n17331 ;
  assign n17681 = n17361 & ~n17680 ;
  assign n17682 = ~n17361 & n17680 ;
  assign n17683 = ~n17681 & ~n17682 ;
  assign n17684 = n167 & n17683 ;
  assign n17685 = n17679 & ~n17684 ;
  assign n17686 = ~x2 & ~n17685 ;
  assign n17687 = ~x2 & ~n17686 ;
  assign n17688 = ~n17685 & ~n17686 ;
  assign n17689 = ~n17687 & ~n17688 ;
  assign n17690 = ~n17317 & ~n17323 ;
  assign n17691 = ~n17241 & ~n17247 ;
  assign n17692 = ~n17225 & ~n17227 ;
  assign n17693 = ~n17219 & ~n17221 ;
  assign n17694 = ~n17213 & ~n17215 ;
  assign n17695 = ~n17155 & ~n17159 ;
  assign n17696 = ~x82 & n8006 ;
  assign n17697 = ~x80 & n8474 ;
  assign n17698 = ~x81 & n8001 ;
  assign n17699 = ~n17697 & ~n17698 ;
  assign n17700 = ~n17696 & n17699 ;
  assign n17701 = n2697 & n8009 ;
  assign n17702 = n17700 & ~n17701 ;
  assign n17703 = ~x35 & ~n17702 ;
  assign n17704 = ~x35 & ~n17703 ;
  assign n17705 = ~n17702 & ~n17703 ;
  assign n17706 = ~n17704 & ~n17705 ;
  assign n17707 = ~n17148 & ~n17152 ;
  assign n17708 = ~x79 & n9433 ;
  assign n17709 = ~x77 & n9915 ;
  assign n17710 = ~x78 & n9428 ;
  assign n17711 = ~n17709 & ~n17710 ;
  assign n17712 = ~n17708 & n17711 ;
  assign n17713 = n1921 & n9436 ;
  assign n17714 = n17712 & ~n17713 ;
  assign n17715 = ~x38 & ~n17714 ;
  assign n17716 = ~x38 & ~n17715 ;
  assign n17717 = ~n17714 & ~n17715 ;
  assign n17718 = ~n17716 & ~n17717 ;
  assign n17719 = ~n17132 & ~n17134 ;
  assign n17720 = ~x76 & n10905 ;
  assign n17721 = ~x74 & n11466 ;
  assign n17722 = ~x75 & n10900 ;
  assign n17723 = ~n17721 & ~n17722 ;
  assign n17724 = ~n17720 & n17723 ;
  assign n17725 = n1390 & n10908 ;
  assign n17726 = n17724 & ~n17725 ;
  assign n17727 = ~x41 & ~n17726 ;
  assign n17728 = ~x41 & ~n17727 ;
  assign n17729 = ~n17726 & ~n17727 ;
  assign n17730 = ~n17728 & ~n17729 ;
  assign n17731 = ~n17112 & ~n17116 ;
  assign n17732 = ~x64 & ~n17415 ;
  assign n17733 = ~n17092 & n17732 ;
  assign n17734 = n17092 & ~n17732 ;
  assign n17735 = ~n17733 & ~n17734 ;
  assign n17736 = ~x67 & n16076 ;
  assign n17737 = ~x65 & n16756 ;
  assign n17738 = ~x66 & n16071 ;
  assign n17739 = ~n17737 & ~n17738 ;
  assign n17740 = ~n17736 & n17739 ;
  assign n17741 = n266 & n16079 ;
  assign n17742 = n17740 & ~n17741 ;
  assign n17743 = ~x50 & ~n17742 ;
  assign n17744 = ~x50 & ~n17743 ;
  assign n17745 = ~n17742 & ~n17743 ;
  assign n17746 = ~n17744 & ~n17745 ;
  assign n17747 = ~n17735 & ~n17746 ;
  assign n17748 = n17735 & n17746 ;
  assign n17749 = ~n17747 & ~n17748 ;
  assign n17750 = ~x70 & n14233 ;
  assign n17751 = ~x68 & n14876 ;
  assign n17752 = ~x69 & n14228 ;
  assign n17753 = ~n17751 & ~n17752 ;
  assign n17754 = ~n17750 & n17753 ;
  assign n17755 = n529 & n14236 ;
  assign n17756 = n17754 & ~n17755 ;
  assign n17757 = ~x47 & ~n17756 ;
  assign n17758 = ~x47 & ~n17757 ;
  assign n17759 = ~n17756 & ~n17757 ;
  assign n17760 = ~n17758 & ~n17759 ;
  assign n17761 = n17749 & ~n17760 ;
  assign n17762 = n17749 & ~n17761 ;
  assign n17763 = ~n17760 & ~n17761 ;
  assign n17764 = ~n17762 & ~n17763 ;
  assign n17765 = ~n17105 & ~n17109 ;
  assign n17766 = n17764 & n17765 ;
  assign n17767 = ~n17764 & ~n17765 ;
  assign n17768 = ~n17766 & ~n17767 ;
  assign n17769 = ~x73 & n12506 ;
  assign n17770 = ~x71 & n13131 ;
  assign n17771 = ~x72 & n12501 ;
  assign n17772 = ~n17770 & ~n17771 ;
  assign n17773 = ~n17769 & n17772 ;
  assign n17774 = n903 & n12509 ;
  assign n17775 = n17773 & ~n17774 ;
  assign n17776 = ~x44 & ~n17775 ;
  assign n17777 = ~x44 & ~n17776 ;
  assign n17778 = ~n17775 & ~n17776 ;
  assign n17779 = ~n17777 & ~n17778 ;
  assign n17780 = ~n17768 & n17779 ;
  assign n17781 = n17768 & ~n17779 ;
  assign n17782 = ~n17780 & ~n17781 ;
  assign n17783 = ~n17731 & n17782 ;
  assign n17784 = n17731 & ~n17782 ;
  assign n17785 = ~n17783 & ~n17784 ;
  assign n17786 = ~n17730 & n17785 ;
  assign n17787 = ~n17730 & ~n17786 ;
  assign n17788 = n17785 & ~n17786 ;
  assign n17789 = ~n17787 & ~n17788 ;
  assign n17790 = ~n17719 & ~n17789 ;
  assign n17791 = n17719 & ~n17788 ;
  assign n17792 = ~n17787 & n17791 ;
  assign n17793 = ~n17790 & ~n17792 ;
  assign n17794 = ~n17718 & n17793 ;
  assign n17795 = n17718 & ~n17793 ;
  assign n17796 = ~n17794 & ~n17795 ;
  assign n17797 = ~n17707 & n17796 ;
  assign n17798 = n17707 & ~n17796 ;
  assign n17799 = ~n17797 & ~n17798 ;
  assign n17800 = ~n17706 & n17799 ;
  assign n17801 = n17706 & ~n17799 ;
  assign n17802 = ~n17800 & ~n17801 ;
  assign n17803 = ~n17695 & n17802 ;
  assign n17804 = n17695 & ~n17802 ;
  assign n17805 = ~n17803 & ~n17804 ;
  assign n17806 = ~x85 & n6725 ;
  assign n17807 = ~x83 & n7129 ;
  assign n17808 = ~x84 & n6720 ;
  assign n17809 = ~n17807 & ~n17808 ;
  assign n17810 = ~n17806 & n17809 ;
  assign n17811 = n3521 & n6728 ;
  assign n17812 = n17810 & ~n17811 ;
  assign n17813 = ~x32 & ~n17812 ;
  assign n17814 = ~x32 & ~n17813 ;
  assign n17815 = ~n17812 & ~n17813 ;
  assign n17816 = ~n17814 & ~n17815 ;
  assign n17817 = n17805 & ~n17816 ;
  assign n17818 = n17805 & ~n17817 ;
  assign n17819 = ~n17816 & ~n17817 ;
  assign n17820 = ~n17818 & ~n17819 ;
  assign n17821 = ~n17174 & ~n17180 ;
  assign n17822 = n17820 & n17821 ;
  assign n17823 = ~n17820 & ~n17821 ;
  assign n17824 = ~n17822 & ~n17823 ;
  assign n17825 = ~x88 & n5560 ;
  assign n17826 = ~x86 & n5943 ;
  assign n17827 = ~x87 & n5555 ;
  assign n17828 = ~n17826 & ~n17827 ;
  assign n17829 = ~n17825 & n17828 ;
  assign n17830 = n4457 & n5563 ;
  assign n17831 = n17829 & ~n17830 ;
  assign n17832 = ~x29 & ~n17831 ;
  assign n17833 = ~x29 & ~n17832 ;
  assign n17834 = ~n17831 & ~n17832 ;
  assign n17835 = ~n17833 & ~n17834 ;
  assign n17836 = ~n17824 & n17835 ;
  assign n17837 = n17824 & ~n17835 ;
  assign n17838 = ~n17836 & ~n17837 ;
  assign n17839 = ~n17198 & n17838 ;
  assign n17840 = n17198 & ~n17838 ;
  assign n17841 = ~n17839 & ~n17840 ;
  assign n17842 = ~x91 & n4531 ;
  assign n17843 = ~x89 & n4847 ;
  assign n17844 = ~x90 & n4526 ;
  assign n17845 = ~n17843 & ~n17844 ;
  assign n17846 = ~n17842 & n17845 ;
  assign n17847 = n4534 & n5507 ;
  assign n17848 = n17846 & ~n17847 ;
  assign n17849 = ~x26 & ~n17848 ;
  assign n17850 = ~x26 & ~n17849 ;
  assign n17851 = ~n17848 & ~n17849 ;
  assign n17852 = ~n17850 & ~n17851 ;
  assign n17853 = n17841 & ~n17852 ;
  assign n17854 = n17841 & ~n17853 ;
  assign n17855 = ~n17852 & ~n17853 ;
  assign n17856 = ~n17854 & ~n17855 ;
  assign n17857 = ~n17694 & n17856 ;
  assign n17858 = n17694 & ~n17856 ;
  assign n17859 = ~n17857 & ~n17858 ;
  assign n17860 = ~x94 & n3589 ;
  assign n17861 = ~x92 & n3878 ;
  assign n17862 = ~x93 & n3584 ;
  assign n17863 = ~n17861 & ~n17862 ;
  assign n17864 = ~n17860 & n17863 ;
  assign n17865 = n3592 & n6671 ;
  assign n17866 = n17864 & ~n17865 ;
  assign n17867 = ~x23 & ~n17866 ;
  assign n17868 = ~x23 & ~n17867 ;
  assign n17869 = ~n17866 & ~n17867 ;
  assign n17870 = ~n17868 & ~n17869 ;
  assign n17871 = ~n17859 & ~n17870 ;
  assign n17872 = n17859 & n17870 ;
  assign n17873 = ~n17871 & ~n17872 ;
  assign n17874 = ~n17693 & n17873 ;
  assign n17875 = n17693 & ~n17873 ;
  assign n17876 = ~n17874 & ~n17875 ;
  assign n17877 = ~x97 & n2751 ;
  assign n17878 = ~x95 & n3020 ;
  assign n17879 = ~x96 & n2746 ;
  assign n17880 = ~n17878 & ~n17879 ;
  assign n17881 = ~n17877 & n17880 ;
  assign n17882 = n2754 & n7949 ;
  assign n17883 = n17881 & ~n17882 ;
  assign n17884 = ~x20 & ~n17883 ;
  assign n17885 = ~x20 & ~n17884 ;
  assign n17886 = ~n17883 & ~n17884 ;
  assign n17887 = ~n17885 & ~n17886 ;
  assign n17888 = n17876 & ~n17887 ;
  assign n17889 = n17876 & ~n17888 ;
  assign n17890 = ~n17887 & ~n17888 ;
  assign n17891 = ~n17889 & ~n17890 ;
  assign n17892 = ~n17692 & n17891 ;
  assign n17893 = n17692 & ~n17891 ;
  assign n17894 = ~n17892 & ~n17893 ;
  assign n17895 = ~x100 & n2093 ;
  assign n17896 = ~x98 & n2275 ;
  assign n17897 = ~x99 & n2088 ;
  assign n17898 = ~n17896 & ~n17897 ;
  assign n17899 = ~n17895 & n17898 ;
  assign n17900 = n2096 & n9338 ;
  assign n17901 = n17899 & ~n17900 ;
  assign n17902 = ~x17 & ~n17901 ;
  assign n17903 = ~x17 & ~n17902 ;
  assign n17904 = ~n17901 & ~n17902 ;
  assign n17905 = ~n17903 & ~n17904 ;
  assign n17906 = ~n17894 & ~n17905 ;
  assign n17907 = n17894 & n17905 ;
  assign n17908 = ~n17906 & ~n17907 ;
  assign n17909 = n17691 & ~n17908 ;
  assign n17910 = ~n17691 & n17908 ;
  assign n17911 = ~n17909 & ~n17910 ;
  assign n17912 = ~x103 & n1434 ;
  assign n17913 = ~x101 & n1646 ;
  assign n17914 = ~x102 & n1429 ;
  assign n17915 = ~n17913 & ~n17914 ;
  assign n17916 = ~n17912 & n17915 ;
  assign n17917 = n1437 & n10833 ;
  assign n17918 = n17916 & ~n17917 ;
  assign n17919 = ~x14 & ~n17918 ;
  assign n17920 = ~x14 & ~n17919 ;
  assign n17921 = ~n17918 & ~n17919 ;
  assign n17922 = ~n17920 & ~n17921 ;
  assign n17923 = n17911 & ~n17922 ;
  assign n17924 = n17911 & ~n17923 ;
  assign n17925 = ~n17922 & ~n17923 ;
  assign n17926 = ~n17924 & ~n17925 ;
  assign n17927 = ~n17260 & ~n17266 ;
  assign n17928 = n17926 & n17927 ;
  assign n17929 = ~n17926 & ~n17927 ;
  assign n17930 = ~n17928 & ~n17929 ;
  assign n17931 = ~x106 & n945 ;
  assign n17932 = ~x104 & n1099 ;
  assign n17933 = ~x105 & n940 ;
  assign n17934 = ~n17932 & ~n17933 ;
  assign n17935 = ~n17931 & n17934 ;
  assign n17936 = n948 & n12447 ;
  assign n17937 = n17935 & ~n17936 ;
  assign n17938 = ~x11 & ~n17937 ;
  assign n17939 = ~x11 & ~n17938 ;
  assign n17940 = ~n17937 & ~n17938 ;
  assign n17941 = ~n17939 & ~n17940 ;
  assign n17942 = ~n17930 & n17941 ;
  assign n17943 = n17930 & ~n17941 ;
  assign n17944 = ~n17942 & ~n17943 ;
  assign n17945 = ~n17279 & ~n17285 ;
  assign n17946 = n17944 & ~n17945 ;
  assign n17947 = ~n17944 & n17945 ;
  assign n17948 = ~n17946 & ~n17947 ;
  assign n17949 = ~x109 & n574 ;
  assign n17950 = ~x107 & n673 ;
  assign n17951 = ~x108 & n569 ;
  assign n17952 = ~n17950 & ~n17951 ;
  assign n17953 = ~n17949 & n17952 ;
  assign n17954 = n577 & n14177 ;
  assign n17955 = n17953 & ~n17954 ;
  assign n17956 = ~x8 & ~n17955 ;
  assign n17957 = ~x8 & ~n17956 ;
  assign n17958 = ~n17955 & ~n17956 ;
  assign n17959 = ~n17957 & ~n17958 ;
  assign n17960 = n17948 & ~n17959 ;
  assign n17961 = n17948 & ~n17960 ;
  assign n17962 = ~n17959 & ~n17960 ;
  assign n17963 = ~n17961 & ~n17962 ;
  assign n17964 = ~n17303 & n17963 ;
  assign n17965 = n17303 & ~n17963 ;
  assign n17966 = ~n17964 & ~n17965 ;
  assign n17967 = ~x112 & n293 ;
  assign n17968 = ~x110 & n373 ;
  assign n17969 = ~x111 & n288 ;
  assign n17970 = ~n17968 & ~n17969 ;
  assign n17971 = ~n17967 & n17970 ;
  assign n17972 = n296 & n15744 ;
  assign n17973 = n17971 & ~n17972 ;
  assign n17974 = ~x5 & ~n17973 ;
  assign n17975 = ~x5 & ~n17974 ;
  assign n17976 = ~n17973 & ~n17974 ;
  assign n17977 = ~n17975 & ~n17976 ;
  assign n17978 = n17966 & n17977 ;
  assign n17979 = ~n17966 & ~n17977 ;
  assign n17980 = ~n17978 & ~n17979 ;
  assign n17981 = ~n17690 & n17980 ;
  assign n17982 = n17690 & ~n17980 ;
  assign n17983 = ~n17981 & ~n17982 ;
  assign n17984 = ~n17689 & n17983 ;
  assign n17985 = n17689 & ~n17983 ;
  assign n17986 = ~n17984 & ~n17985 ;
  assign n17987 = ~n17674 & n17986 ;
  assign n17988 = n17674 & ~n17986 ;
  assign n17989 = ~n17987 & ~n17988 ;
  assign n17992 = ~n17989 & ~x179 ;
  assign n17993 = ~n17991 & ~n17992 ;
  assign n17994 = ~n17668 & ~n17671 ;
  assign n17995 = ~n17663 & ~n17665 ;
  assign n17996 = ~n17627 & ~n17630 ;
  assign n17997 = ~n17375 & ~n17540 ;
  assign n17998 = ~n17537 & ~n17997 ;
  assign n17999 = ~n17521 & ~n17523 ;
  assign n18000 = ~n17484 & ~n17487 ;
  assign n18001 = ~n17470 & ~n17474 ;
  assign n18002 = ~n17465 & ~n17467 ;
  assign n18003 = n16768 & n17416 ;
  assign n18004 = ~n17431 & ~n18003 ;
  assign n18005 = x68 & n16076 ;
  assign n18006 = x66 & n16756 ;
  assign n18007 = x67 & n16071 ;
  assign n18008 = ~n18006 & ~n18007 ;
  assign n18009 = ~n18005 & n18008 ;
  assign n18010 = n317 & n16079 ;
  assign n18011 = n18009 & ~n18010 ;
  assign n18012 = x50 & ~n18011 ;
  assign n18013 = x50 & ~n18012 ;
  assign n18014 = ~n18011 & ~n18012 ;
  assign n18015 = ~n18013 & ~n18014 ;
  assign n18016 = x53 & ~n17416 ;
  assign n18017 = ~x51 & x52 ;
  assign n18018 = x51 & ~x52 ;
  assign n18019 = ~n18017 & ~n18018 ;
  assign n18020 = n17415 & ~n18019 ;
  assign n18021 = x64 & n18020 ;
  assign n18022 = ~x52 & x53 ;
  assign n18023 = x52 & ~x53 ;
  assign n18024 = ~n18022 & ~n18023 ;
  assign n18025 = ~n17415 & n18024 ;
  assign n18026 = x65 & n18025 ;
  assign n18027 = ~n18021 & ~n18026 ;
  assign n18028 = ~n17415 & ~n18024 ;
  assign n18029 = ~n152 & n18028 ;
  assign n18030 = n18027 & ~n18029 ;
  assign n18031 = x53 & ~n18030 ;
  assign n18032 = x53 & ~n18031 ;
  assign n18033 = ~n18030 & ~n18031 ;
  assign n18034 = ~n18032 & ~n18033 ;
  assign n18035 = n18016 & ~n18034 ;
  assign n18036 = ~n18016 & n18034 ;
  assign n18037 = ~n18035 & ~n18036 ;
  assign n18038 = n18015 & ~n18037 ;
  assign n18039 = ~n18015 & n18037 ;
  assign n18040 = ~n18038 & ~n18039 ;
  assign n18041 = ~n18004 & n18040 ;
  assign n18042 = n18004 & ~n18040 ;
  assign n18043 = ~n18041 & ~n18042 ;
  assign n18044 = x71 & n14233 ;
  assign n18045 = x69 & n14876 ;
  assign n18046 = x70 & n14228 ;
  assign n18047 = ~n18045 & ~n18046 ;
  assign n18048 = ~n18044 & n18047 ;
  assign n18049 = n558 & n14236 ;
  assign n18050 = n18048 & ~n18049 ;
  assign n18051 = x47 & ~n18050 ;
  assign n18052 = x47 & ~n18051 ;
  assign n18053 = ~n18050 & ~n18051 ;
  assign n18054 = ~n18052 & ~n18053 ;
  assign n18055 = n18043 & ~n18054 ;
  assign n18056 = n18043 & ~n18055 ;
  assign n18057 = ~n18054 & ~n18055 ;
  assign n18058 = ~n18056 & ~n18057 ;
  assign n18059 = ~n17445 & ~n17451 ;
  assign n18060 = n18058 & n18059 ;
  assign n18061 = ~n18058 & ~n18059 ;
  assign n18062 = ~n18060 & ~n18061 ;
  assign n18063 = x74 & n12506 ;
  assign n18064 = x72 & n13131 ;
  assign n18065 = x73 & n12501 ;
  assign n18066 = ~n18064 & ~n18065 ;
  assign n18067 = ~n18063 & n18066 ;
  assign n18068 = n994 & n12509 ;
  assign n18069 = n18067 & ~n18068 ;
  assign n18070 = x44 & ~n18069 ;
  assign n18071 = x44 & ~n18070 ;
  assign n18072 = ~n18069 & ~n18070 ;
  assign n18073 = ~n18071 & ~n18072 ;
  assign n18074 = n18062 & ~n18073 ;
  assign n18075 = ~n18062 & n18073 ;
  assign n18076 = ~n18002 & ~n18075 ;
  assign n18077 = ~n18074 & n18076 ;
  assign n18078 = ~n18002 & ~n18077 ;
  assign n18079 = ~n18074 & ~n18077 ;
  assign n18080 = ~n18075 & n18079 ;
  assign n18081 = ~n18078 & ~n18080 ;
  assign n18082 = x77 & n10905 ;
  assign n18083 = x75 & n11466 ;
  assign n18084 = x76 & n10900 ;
  assign n18085 = ~n18083 & ~n18084 ;
  assign n18086 = ~n18082 & n18085 ;
  assign n18087 = n1502 & n10908 ;
  assign n18088 = n18086 & ~n18087 ;
  assign n18089 = x41 & ~n18088 ;
  assign n18090 = x41 & ~n18089 ;
  assign n18091 = ~n18088 & ~n18089 ;
  assign n18092 = ~n18090 & ~n18091 ;
  assign n18093 = n18081 & n18092 ;
  assign n18094 = ~n18081 & ~n18092 ;
  assign n18095 = ~n18093 & ~n18094 ;
  assign n18096 = ~n18001 & n18095 ;
  assign n18097 = n18001 & ~n18095 ;
  assign n18098 = ~n18096 & ~n18097 ;
  assign n18099 = x80 & n9433 ;
  assign n18100 = x78 & n9915 ;
  assign n18101 = x79 & n9428 ;
  assign n18102 = ~n18100 & ~n18101 ;
  assign n18103 = ~n18099 & n18102 ;
  assign n18104 = n2028 & n9436 ;
  assign n18105 = n18103 & ~n18104 ;
  assign n18106 = x38 & ~n18105 ;
  assign n18107 = x38 & ~n18106 ;
  assign n18108 = ~n18105 & ~n18106 ;
  assign n18109 = ~n18107 & ~n18108 ;
  assign n18110 = n18098 & ~n18109 ;
  assign n18111 = n18098 & ~n18110 ;
  assign n18112 = ~n18109 & ~n18110 ;
  assign n18113 = ~n18111 & ~n18112 ;
  assign n18114 = ~n17478 & ~n17481 ;
  assign n18115 = n18113 & n18114 ;
  assign n18116 = ~n18113 & ~n18114 ;
  assign n18117 = ~n18115 & ~n18116 ;
  assign n18118 = x83 & n8006 ;
  assign n18119 = x81 & n8474 ;
  assign n18120 = x82 & n8001 ;
  assign n18121 = ~n18119 & ~n18120 ;
  assign n18122 = ~n18118 & n18121 ;
  assign n18123 = n2843 & n8009 ;
  assign n18124 = n18122 & ~n18123 ;
  assign n18125 = x35 & ~n18124 ;
  assign n18126 = x35 & ~n18125 ;
  assign n18127 = ~n18124 & ~n18125 ;
  assign n18128 = ~n18126 & ~n18127 ;
  assign n18129 = n18117 & ~n18128 ;
  assign n18130 = ~n18117 & n18128 ;
  assign n18131 = ~n18000 & ~n18130 ;
  assign n18132 = ~n18129 & n18131 ;
  assign n18133 = ~n18000 & ~n18132 ;
  assign n18134 = ~n18129 & ~n18132 ;
  assign n18135 = ~n18130 & n18134 ;
  assign n18136 = ~n18133 & ~n18135 ;
  assign n18137 = x86 & n6725 ;
  assign n18138 = x84 & n7129 ;
  assign n18139 = x85 & n6720 ;
  assign n18140 = ~n18138 & ~n18139 ;
  assign n18141 = ~n18137 & n18140 ;
  assign n18142 = n3686 & n6728 ;
  assign n18143 = n18141 & ~n18142 ;
  assign n18144 = x32 & ~n18143 ;
  assign n18145 = x32 & ~n18144 ;
  assign n18146 = ~n18143 & ~n18144 ;
  assign n18147 = ~n18145 & ~n18146 ;
  assign n18148 = ~n18136 & ~n18147 ;
  assign n18149 = ~n18136 & ~n18148 ;
  assign n18150 = ~n18147 & ~n18148 ;
  assign n18151 = ~n18149 & ~n18150 ;
  assign n18152 = ~n17501 & ~n17507 ;
  assign n18153 = n18151 & n18152 ;
  assign n18154 = ~n18151 & ~n18152 ;
  assign n18155 = ~n18153 & ~n18154 ;
  assign n18156 = x89 & n5560 ;
  assign n18157 = x87 & n5943 ;
  assign n18158 = x88 & n5555 ;
  assign n18159 = ~n18157 & ~n18158 ;
  assign n18160 = ~n18156 & n18159 ;
  assign n18161 = n4488 & n5563 ;
  assign n18162 = n18160 & ~n18161 ;
  assign n18163 = x29 & ~n18162 ;
  assign n18164 = x29 & ~n18163 ;
  assign n18165 = ~n18162 & ~n18163 ;
  assign n18166 = ~n18164 & ~n18165 ;
  assign n18167 = n18155 & ~n18166 ;
  assign n18168 = n18155 & ~n18167 ;
  assign n18169 = ~n18166 & ~n18167 ;
  assign n18170 = ~n18168 & ~n18169 ;
  assign n18171 = ~n17999 & n18170 ;
  assign n18172 = n17999 & ~n18170 ;
  assign n18173 = ~n18171 & ~n18172 ;
  assign n18174 = x92 & n4531 ;
  assign n18175 = x90 & n4847 ;
  assign n18176 = x91 & n4526 ;
  assign n18177 = ~n18175 & ~n18176 ;
  assign n18178 = ~n18174 & n18177 ;
  assign n18179 = n4534 & n5710 ;
  assign n18180 = n18178 & ~n18179 ;
  assign n18181 = x26 & ~n18180 ;
  assign n18182 = x26 & ~n18181 ;
  assign n18183 = ~n18180 & ~n18181 ;
  assign n18184 = ~n18182 & ~n18183 ;
  assign n18185 = ~n18173 & ~n18184 ;
  assign n18186 = n18173 & n18184 ;
  assign n18187 = ~n18185 & ~n18186 ;
  assign n18188 = n17998 & ~n18187 ;
  assign n18189 = ~n17998 & n18187 ;
  assign n18190 = ~n18188 & ~n18189 ;
  assign n18191 = x95 & n3589 ;
  assign n18192 = x93 & n3878 ;
  assign n18193 = x94 & n3584 ;
  assign n18194 = ~n18192 & ~n18193 ;
  assign n18195 = ~n18191 & n18194 ;
  assign n18196 = n3592 & n6894 ;
  assign n18197 = n18195 & ~n18196 ;
  assign n18198 = x23 & ~n18197 ;
  assign n18199 = x23 & ~n18198 ;
  assign n18200 = ~n18197 & ~n18198 ;
  assign n18201 = ~n18199 & ~n18200 ;
  assign n18202 = n18190 & ~n18201 ;
  assign n18203 = n18190 & ~n18202 ;
  assign n18204 = ~n18201 & ~n18202 ;
  assign n18205 = ~n18203 & ~n18204 ;
  assign n18206 = ~n17555 & ~n17558 ;
  assign n18207 = n18205 & n18206 ;
  assign n18208 = ~n18205 & ~n18206 ;
  assign n18209 = ~n18207 & ~n18208 ;
  assign n18210 = x98 & n2751 ;
  assign n18211 = x96 & n3020 ;
  assign n18212 = x97 & n2746 ;
  assign n18213 = ~n18211 & ~n18212 ;
  assign n18214 = ~n18210 & n18213 ;
  assign n18215 = n2754 & n8196 ;
  assign n18216 = n18214 & ~n18215 ;
  assign n18217 = x20 & ~n18216 ;
  assign n18218 = x20 & ~n18217 ;
  assign n18219 = ~n18216 & ~n18217 ;
  assign n18220 = ~n18218 & ~n18219 ;
  assign n18221 = n18209 & ~n18220 ;
  assign n18222 = n18209 & ~n18221 ;
  assign n18223 = ~n18220 & ~n18221 ;
  assign n18224 = ~n18222 & ~n18223 ;
  assign n18225 = ~n17373 & ~n17575 ;
  assign n18226 = ~n17572 & ~n18225 ;
  assign n18227 = n18224 & n18226 ;
  assign n18228 = ~n18224 & ~n18226 ;
  assign n18229 = ~n18227 & ~n18228 ;
  assign n18230 = x101 & n2093 ;
  assign n18231 = x99 & n2275 ;
  assign n18232 = x100 & n2088 ;
  assign n18233 = ~n18231 & ~n18232 ;
  assign n18234 = ~n18230 & n18233 ;
  assign n18235 = n2096 & n9601 ;
  assign n18236 = n18234 & ~n18235 ;
  assign n18237 = x17 & ~n18236 ;
  assign n18238 = x17 & ~n18237 ;
  assign n18239 = ~n18236 & ~n18237 ;
  assign n18240 = ~n18238 & ~n18239 ;
  assign n18241 = n18229 & ~n18240 ;
  assign n18242 = n18229 & ~n18241 ;
  assign n18243 = ~n18240 & ~n18241 ;
  assign n18244 = ~n18242 & ~n18243 ;
  assign n18245 = ~n17590 & ~n17594 ;
  assign n18246 = n18244 & n18245 ;
  assign n18247 = ~n18244 & ~n18245 ;
  assign n18248 = ~n18246 & ~n18247 ;
  assign n18249 = x104 & n1434 ;
  assign n18250 = x102 & n1646 ;
  assign n18251 = x103 & n1429 ;
  assign n18252 = ~n18250 & ~n18251 ;
  assign n18253 = ~n18249 & n18252 ;
  assign n18254 = n1437 & n11116 ;
  assign n18255 = n18253 & ~n18254 ;
  assign n18256 = x14 & ~n18255 ;
  assign n18257 = x14 & ~n18256 ;
  assign n18258 = ~n18255 & ~n18256 ;
  assign n18259 = ~n18257 & ~n18258 ;
  assign n18260 = n18248 & ~n18259 ;
  assign n18261 = n18248 & ~n18260 ;
  assign n18262 = ~n18259 & ~n18260 ;
  assign n18263 = ~n18261 & ~n18262 ;
  assign n18264 = ~n17607 & ~n17613 ;
  assign n18265 = n18263 & n18264 ;
  assign n18266 = ~n18263 & ~n18264 ;
  assign n18267 = ~n18265 & ~n18266 ;
  assign n18268 = x107 & n945 ;
  assign n18269 = x105 & n1099 ;
  assign n18270 = x106 & n940 ;
  assign n18271 = ~n18269 & ~n18270 ;
  assign n18272 = ~n18268 & n18271 ;
  assign n18273 = n948 & n12749 ;
  assign n18274 = n18272 & ~n18273 ;
  assign n18275 = x11 & ~n18274 ;
  assign n18276 = x11 & ~n18275 ;
  assign n18277 = ~n18274 & ~n18275 ;
  assign n18278 = ~n18276 & ~n18277 ;
  assign n18279 = n18267 & ~n18278 ;
  assign n18280 = ~n18267 & n18278 ;
  assign n18281 = ~n17996 & ~n18280 ;
  assign n18282 = ~n18279 & n18281 ;
  assign n18283 = ~n17996 & ~n18282 ;
  assign n18284 = ~n18279 & ~n18282 ;
  assign n18285 = ~n18280 & n18284 ;
  assign n18286 = ~n18283 & ~n18285 ;
  assign n18287 = x110 & n574 ;
  assign n18288 = x108 & n673 ;
  assign n18289 = x109 & n569 ;
  assign n18290 = ~n18288 & ~n18289 ;
  assign n18291 = ~n18287 & n18290 ;
  assign n18292 = n577 & n14497 ;
  assign n18293 = n18291 & ~n18292 ;
  assign n18294 = x8 & ~n18293 ;
  assign n18295 = x8 & ~n18294 ;
  assign n18296 = ~n18293 & ~n18294 ;
  assign n18297 = ~n18295 & ~n18296 ;
  assign n18298 = ~n18286 & ~n18297 ;
  assign n18299 = ~n18286 & ~n18298 ;
  assign n18300 = ~n18297 & ~n18298 ;
  assign n18301 = ~n18299 & ~n18300 ;
  assign n18302 = ~n16979 & ~n17647 ;
  assign n18303 = ~n17644 & ~n18302 ;
  assign n18304 = n18301 & n18303 ;
  assign n18305 = ~n18301 & ~n18303 ;
  assign n18306 = ~n18304 & ~n18305 ;
  assign n18307 = x113 & n293 ;
  assign n18308 = x111 & n373 ;
  assign n18309 = x112 & n288 ;
  assign n18310 = ~n18308 & ~n18309 ;
  assign n18311 = ~n18307 & n18310 ;
  assign n18312 = n296 & n16361 ;
  assign n18313 = n18311 & ~n18312 ;
  assign n18314 = x5 & ~n18313 ;
  assign n18315 = x5 & ~n18314 ;
  assign n18316 = ~n18313 & ~n18314 ;
  assign n18317 = ~n18315 & ~n18316 ;
  assign n18318 = n18306 & ~n18317 ;
  assign n18319 = n18306 & ~n18318 ;
  assign n18320 = ~n18317 & ~n18318 ;
  assign n18321 = ~n18319 & ~n18320 ;
  assign n18322 = ~n17995 & n18321 ;
  assign n18323 = n17995 & ~n18321 ;
  assign n18324 = ~n18322 & ~n18323 ;
  assign n18325 = x116 & n146 ;
  assign n18326 = x114 & n182 ;
  assign n18327 = x115 & n141 ;
  assign n18328 = ~n18326 & ~n18327 ;
  assign n18329 = ~n18325 & n18328 ;
  assign n18330 = ~n17360 & ~n17362 ;
  assign n18331 = ~x115 & ~x116 ;
  assign n18332 = x115 & x116 ;
  assign n18333 = ~n18331 & ~n18332 ;
  assign n18334 = ~n18330 & n18333 ;
  assign n18335 = n18330 & ~n18333 ;
  assign n18336 = ~n18334 & ~n18335 ;
  assign n18337 = n149 & n18336 ;
  assign n18338 = n18329 & ~n18337 ;
  assign n18339 = x2 & ~n18338 ;
  assign n18340 = x2 & ~n18339 ;
  assign n18341 = ~n18338 & ~n18339 ;
  assign n18342 = ~n18340 & ~n18341 ;
  assign n18343 = ~n18324 & ~n18342 ;
  assign n18344 = n18324 & n18342 ;
  assign n18345 = ~n18343 & ~n18344 ;
  assign n18346 = ~n17994 & n18345 ;
  assign n18347 = n17994 & ~n18345 ;
  assign n18348 = ~n18346 & ~n18347 ;
  assign n18692 = n18348 & x180 ;
  assign n18349 = ~n17984 & ~n17987 ;
  assign n18350 = ~n17979 & ~n17981 ;
  assign n18351 = ~n17943 & ~n17946 ;
  assign n18352 = ~n17694 & ~n17856 ;
  assign n18353 = ~n17853 & ~n18352 ;
  assign n18354 = ~n17837 & ~n17839 ;
  assign n18355 = ~n17800 & ~n17803 ;
  assign n18356 = ~n17786 & ~n17790 ;
  assign n18357 = ~n17781 & ~n17783 ;
  assign n18358 = n17092 & n17732 ;
  assign n18359 = ~n17747 & ~n18358 ;
  assign n18360 = ~x68 & n16076 ;
  assign n18361 = ~x66 & n16756 ;
  assign n18362 = ~x67 & n16071 ;
  assign n18363 = ~n18361 & ~n18362 ;
  assign n18364 = ~n18360 & n18363 ;
  assign n18365 = n352 & n16079 ;
  assign n18366 = n18364 & ~n18365 ;
  assign n18367 = ~x50 & ~n18366 ;
  assign n18368 = ~x50 & ~n18367 ;
  assign n18369 = ~n18366 & ~n18367 ;
  assign n18370 = ~n18368 & ~n18369 ;
  assign n18371 = ~x53 & ~n17732 ;
  assign n18372 = ~x64 & n18020 ;
  assign n18373 = ~x65 & n18025 ;
  assign n18374 = ~n18372 & ~n18373 ;
  assign n18375 = ~n18029 & n18374 ;
  assign n18376 = ~x53 & ~n18375 ;
  assign n18377 = ~x53 & ~n18376 ;
  assign n18378 = ~n18375 & ~n18376 ;
  assign n18379 = ~n18377 & ~n18378 ;
  assign n18380 = n18371 & ~n18379 ;
  assign n18381 = ~n18371 & n18379 ;
  assign n18382 = ~n18380 & ~n18381 ;
  assign n18383 = n18370 & ~n18382 ;
  assign n18384 = ~n18370 & n18382 ;
  assign n18385 = ~n18383 & ~n18384 ;
  assign n18386 = ~n18359 & n18385 ;
  assign n18387 = n18359 & ~n18385 ;
  assign n18388 = ~n18386 & ~n18387 ;
  assign n18389 = ~x71 & n14233 ;
  assign n18390 = ~x69 & n14876 ;
  assign n18391 = ~x70 & n14228 ;
  assign n18392 = ~n18390 & ~n18391 ;
  assign n18393 = ~n18389 & n18392 ;
  assign n18394 = n622 & n14236 ;
  assign n18395 = n18393 & ~n18394 ;
  assign n18396 = ~x47 & ~n18395 ;
  assign n18397 = ~x47 & ~n18396 ;
  assign n18398 = ~n18395 & ~n18396 ;
  assign n18399 = ~n18397 & ~n18398 ;
  assign n18400 = n18388 & ~n18399 ;
  assign n18401 = n18388 & ~n18400 ;
  assign n18402 = ~n18399 & ~n18400 ;
  assign n18403 = ~n18401 & ~n18402 ;
  assign n18404 = ~n17761 & ~n17767 ;
  assign n18405 = n18403 & n18404 ;
  assign n18406 = ~n18403 & ~n18404 ;
  assign n18407 = ~n18405 & ~n18406 ;
  assign n18408 = ~x74 & n12506 ;
  assign n18409 = ~x72 & n13131 ;
  assign n18410 = ~x73 & n12501 ;
  assign n18411 = ~n18409 & ~n18410 ;
  assign n18412 = ~n18408 & n18411 ;
  assign n18413 = n1066 & n12509 ;
  assign n18414 = n18412 & ~n18413 ;
  assign n18415 = ~x44 & ~n18414 ;
  assign n18416 = ~x44 & ~n18415 ;
  assign n18417 = ~n18414 & ~n18415 ;
  assign n18418 = ~n18416 & ~n18417 ;
  assign n18419 = n18407 & ~n18418 ;
  assign n18420 = ~n18407 & n18418 ;
  assign n18421 = ~n18357 & ~n18420 ;
  assign n18422 = ~n18419 & n18421 ;
  assign n18423 = ~n18357 & ~n18422 ;
  assign n18424 = ~n18419 & ~n18422 ;
  assign n18425 = ~n18420 & n18424 ;
  assign n18426 = ~n18423 & ~n18425 ;
  assign n18427 = ~x77 & n10905 ;
  assign n18428 = ~x75 & n11466 ;
  assign n18429 = ~x76 & n10900 ;
  assign n18430 = ~n18428 & ~n18429 ;
  assign n18431 = ~n18427 & n18430 ;
  assign n18432 = n1594 & n10908 ;
  assign n18433 = n18431 & ~n18432 ;
  assign n18434 = ~x41 & ~n18433 ;
  assign n18435 = ~x41 & ~n18434 ;
  assign n18436 = ~n18433 & ~n18434 ;
  assign n18437 = ~n18435 & ~n18436 ;
  assign n18438 = n18426 & n18437 ;
  assign n18439 = ~n18426 & ~n18437 ;
  assign n18440 = ~n18438 & ~n18439 ;
  assign n18441 = ~n18356 & n18440 ;
  assign n18442 = n18356 & ~n18440 ;
  assign n18443 = ~n18441 & ~n18442 ;
  assign n18444 = ~x80 & n9433 ;
  assign n18445 = ~x78 & n9915 ;
  assign n18446 = ~x79 & n9428 ;
  assign n18447 = ~n18445 & ~n18446 ;
  assign n18448 = ~n18444 & n18447 ;
  assign n18449 = n2145 & n9436 ;
  assign n18450 = n18448 & ~n18449 ;
  assign n18451 = ~x38 & ~n18450 ;
  assign n18452 = ~x38 & ~n18451 ;
  assign n18453 = ~n18450 & ~n18451 ;
  assign n18454 = ~n18452 & ~n18453 ;
  assign n18455 = n18443 & ~n18454 ;
  assign n18456 = n18443 & ~n18455 ;
  assign n18457 = ~n18454 & ~n18455 ;
  assign n18458 = ~n18456 & ~n18457 ;
  assign n18459 = ~n17794 & ~n17797 ;
  assign n18460 = n18458 & n18459 ;
  assign n18461 = ~n18458 & ~n18459 ;
  assign n18462 = ~n18460 & ~n18461 ;
  assign n18463 = ~x83 & n8006 ;
  assign n18464 = ~x81 & n8474 ;
  assign n18465 = ~x82 & n8001 ;
  assign n18466 = ~n18464 & ~n18465 ;
  assign n18467 = ~n18463 & n18466 ;
  assign n18468 = n2972 & n8009 ;
  assign n18469 = n18467 & ~n18468 ;
  assign n18470 = ~x35 & ~n18469 ;
  assign n18471 = ~x35 & ~n18470 ;
  assign n18472 = ~n18469 & ~n18470 ;
  assign n18473 = ~n18471 & ~n18472 ;
  assign n18474 = n18462 & ~n18473 ;
  assign n18475 = ~n18462 & n18473 ;
  assign n18476 = ~n18355 & ~n18475 ;
  assign n18477 = ~n18474 & n18476 ;
  assign n18478 = ~n18355 & ~n18477 ;
  assign n18479 = ~n18474 & ~n18477 ;
  assign n18480 = ~n18475 & n18479 ;
  assign n18481 = ~n18478 & ~n18480 ;
  assign n18482 = ~x86 & n6725 ;
  assign n18483 = ~x84 & n7129 ;
  assign n18484 = ~x85 & n6720 ;
  assign n18485 = ~n18483 & ~n18484 ;
  assign n18486 = ~n18482 & n18485 ;
  assign n18487 = n3832 & n6728 ;
  assign n18488 = n18486 & ~n18487 ;
  assign n18489 = ~x32 & ~n18488 ;
  assign n18490 = ~x32 & ~n18489 ;
  assign n18491 = ~n18488 & ~n18489 ;
  assign n18492 = ~n18490 & ~n18491 ;
  assign n18493 = ~n18481 & ~n18492 ;
  assign n18494 = ~n18481 & ~n18493 ;
  assign n18495 = ~n18492 & ~n18493 ;
  assign n18496 = ~n18494 & ~n18495 ;
  assign n18497 = ~n17817 & ~n17823 ;
  assign n18498 = n18496 & n18497 ;
  assign n18499 = ~n18496 & ~n18497 ;
  assign n18500 = ~n18498 & ~n18499 ;
  assign n18501 = ~x89 & n5560 ;
  assign n18502 = ~x87 & n5943 ;
  assign n18503 = ~x88 & n5555 ;
  assign n18504 = ~n18502 & ~n18503 ;
  assign n18505 = ~n18501 & n18504 ;
  assign n18506 = n4664 & n5563 ;
  assign n18507 = n18505 & ~n18506 ;
  assign n18508 = ~x29 & ~n18507 ;
  assign n18509 = ~x29 & ~n18508 ;
  assign n18510 = ~n18507 & ~n18508 ;
  assign n18511 = ~n18509 & ~n18510 ;
  assign n18512 = n18500 & ~n18511 ;
  assign n18513 = n18500 & ~n18512 ;
  assign n18514 = ~n18511 & ~n18512 ;
  assign n18515 = ~n18513 & ~n18514 ;
  assign n18516 = ~n18354 & n18515 ;
  assign n18517 = n18354 & ~n18515 ;
  assign n18518 = ~n18516 & ~n18517 ;
  assign n18519 = ~x92 & n4531 ;
  assign n18520 = ~x90 & n4847 ;
  assign n18521 = ~x91 & n4526 ;
  assign n18522 = ~n18520 & ~n18521 ;
  assign n18523 = ~n18519 & n18522 ;
  assign n18524 = n4534 & n5896 ;
  assign n18525 = n18523 & ~n18524 ;
  assign n18526 = ~x26 & ~n18525 ;
  assign n18527 = ~x26 & ~n18526 ;
  assign n18528 = ~n18525 & ~n18526 ;
  assign n18529 = ~n18527 & ~n18528 ;
  assign n18530 = ~n18518 & ~n18529 ;
  assign n18531 = n18518 & n18529 ;
  assign n18532 = ~n18530 & ~n18531 ;
  assign n18533 = n18353 & ~n18532 ;
  assign n18534 = ~n18353 & n18532 ;
  assign n18535 = ~n18533 & ~n18534 ;
  assign n18536 = ~x95 & n3589 ;
  assign n18537 = ~x93 & n3878 ;
  assign n18538 = ~x94 & n3584 ;
  assign n18539 = ~n18537 & ~n18538 ;
  assign n18540 = ~n18536 & n18539 ;
  assign n18541 = n3592 & n7100 ;
  assign n18542 = n18540 & ~n18541 ;
  assign n18543 = ~x23 & ~n18542 ;
  assign n18544 = ~x23 & ~n18543 ;
  assign n18545 = ~n18542 & ~n18543 ;
  assign n18546 = ~n18544 & ~n18545 ;
  assign n18547 = n18535 & ~n18546 ;
  assign n18548 = n18535 & ~n18547 ;
  assign n18549 = ~n18546 & ~n18547 ;
  assign n18550 = ~n18548 & ~n18549 ;
  assign n18551 = ~n17871 & ~n17874 ;
  assign n18552 = n18550 & n18551 ;
  assign n18553 = ~n18550 & ~n18551 ;
  assign n18554 = ~n18552 & ~n18553 ;
  assign n18555 = ~x98 & n2751 ;
  assign n18556 = ~x96 & n3020 ;
  assign n18557 = ~x97 & n2746 ;
  assign n18558 = ~n18556 & ~n18557 ;
  assign n18559 = ~n18555 & n18558 ;
  assign n18560 = n2754 & n8426 ;
  assign n18561 = n18559 & ~n18560 ;
  assign n18562 = ~x20 & ~n18561 ;
  assign n18563 = ~x20 & ~n18562 ;
  assign n18564 = ~n18561 & ~n18562 ;
  assign n18565 = ~n18563 & ~n18564 ;
  assign n18566 = n18554 & ~n18565 ;
  assign n18567 = n18554 & ~n18566 ;
  assign n18568 = ~n18565 & ~n18566 ;
  assign n18569 = ~n18567 & ~n18568 ;
  assign n18570 = ~n17692 & ~n17891 ;
  assign n18571 = ~n17888 & ~n18570 ;
  assign n18572 = n18569 & n18571 ;
  assign n18573 = ~n18569 & ~n18571 ;
  assign n18574 = ~n18572 & ~n18573 ;
  assign n18575 = ~x101 & n2093 ;
  assign n18576 = ~x99 & n2275 ;
  assign n18577 = ~x100 & n2088 ;
  assign n18578 = ~n18576 & ~n18577 ;
  assign n18579 = ~n18575 & n18578 ;
  assign n18580 = n2096 & n9844 ;
  assign n18581 = n18579 & ~n18580 ;
  assign n18582 = ~x17 & ~n18581 ;
  assign n18583 = ~x17 & ~n18582 ;
  assign n18584 = ~n18581 & ~n18582 ;
  assign n18585 = ~n18583 & ~n18584 ;
  assign n18586 = n18574 & ~n18585 ;
  assign n18587 = n18574 & ~n18586 ;
  assign n18588 = ~n18585 & ~n18586 ;
  assign n18589 = ~n18587 & ~n18588 ;
  assign n18590 = ~n17906 & ~n17910 ;
  assign n18591 = n18589 & n18590 ;
  assign n18592 = ~n18589 & ~n18590 ;
  assign n18593 = ~n18591 & ~n18592 ;
  assign n18594 = ~x104 & n1434 ;
  assign n18595 = ~x102 & n1646 ;
  assign n18596 = ~x103 & n1429 ;
  assign n18597 = ~n18595 & ~n18596 ;
  assign n18598 = ~n18594 & n18597 ;
  assign n18599 = n1437 & n11380 ;
  assign n18600 = n18598 & ~n18599 ;
  assign n18601 = ~x14 & ~n18600 ;
  assign n18602 = ~x14 & ~n18601 ;
  assign n18603 = ~n18600 & ~n18601 ;
  assign n18604 = ~n18602 & ~n18603 ;
  assign n18605 = n18593 & ~n18604 ;
  assign n18606 = n18593 & ~n18605 ;
  assign n18607 = ~n18604 & ~n18605 ;
  assign n18608 = ~n18606 & ~n18607 ;
  assign n18609 = ~n17923 & ~n17929 ;
  assign n18610 = n18608 & n18609 ;
  assign n18611 = ~n18608 & ~n18609 ;
  assign n18612 = ~n18610 & ~n18611 ;
  assign n18613 = ~x107 & n945 ;
  assign n18614 = ~x105 & n1099 ;
  assign n18615 = ~x106 & n940 ;
  assign n18616 = ~n18614 & ~n18615 ;
  assign n18617 = ~n18613 & n18616 ;
  assign n18618 = n948 & n13034 ;
  assign n18619 = n18617 & ~n18618 ;
  assign n18620 = ~x11 & ~n18619 ;
  assign n18621 = ~x11 & ~n18620 ;
  assign n18622 = ~n18619 & ~n18620 ;
  assign n18623 = ~n18621 & ~n18622 ;
  assign n18624 = n18612 & ~n18623 ;
  assign n18625 = ~n18612 & n18623 ;
  assign n18626 = ~n18351 & ~n18625 ;
  assign n18627 = ~n18624 & n18626 ;
  assign n18628 = ~n18351 & ~n18627 ;
  assign n18629 = ~n18624 & ~n18627 ;
  assign n18630 = ~n18625 & n18629 ;
  assign n18631 = ~n18628 & ~n18630 ;
  assign n18632 = ~x110 & n574 ;
  assign n18633 = ~x108 & n673 ;
  assign n18634 = ~x109 & n569 ;
  assign n18635 = ~n18633 & ~n18634 ;
  assign n18636 = ~n18632 & n18635 ;
  assign n18637 = n577 & n14802 ;
  assign n18638 = n18636 & ~n18637 ;
  assign n18639 = ~x8 & ~n18638 ;
  assign n18640 = ~x8 & ~n18639 ;
  assign n18641 = ~n18638 & ~n18639 ;
  assign n18642 = ~n18640 & ~n18641 ;
  assign n18643 = ~n18631 & ~n18642 ;
  assign n18644 = ~n18631 & ~n18643 ;
  assign n18645 = ~n18642 & ~n18643 ;
  assign n18646 = ~n18644 & ~n18645 ;
  assign n18647 = ~n17303 & ~n17963 ;
  assign n18648 = ~n17960 & ~n18647 ;
  assign n18649 = n18646 & n18648 ;
  assign n18650 = ~n18646 & ~n18648 ;
  assign n18651 = ~n18649 & ~n18650 ;
  assign n18652 = ~x113 & n293 ;
  assign n18653 = ~x111 & n373 ;
  assign n18654 = ~x112 & n288 ;
  assign n18655 = ~n18653 & ~n18654 ;
  assign n18656 = ~n18652 & n18655 ;
  assign n18657 = n296 & n16684 ;
  assign n18658 = n18656 & ~n18657 ;
  assign n18659 = ~x5 & ~n18658 ;
  assign n18660 = ~x5 & ~n18659 ;
  assign n18661 = ~n18658 & ~n18659 ;
  assign n18662 = ~n18660 & ~n18661 ;
  assign n18663 = n18651 & ~n18662 ;
  assign n18664 = n18651 & ~n18663 ;
  assign n18665 = ~n18662 & ~n18663 ;
  assign n18666 = ~n18664 & ~n18665 ;
  assign n18667 = ~n18350 & n18666 ;
  assign n18668 = n18350 & ~n18666 ;
  assign n18669 = ~n18667 & ~n18668 ;
  assign n18670 = ~x116 & n164 ;
  assign n18671 = ~x114 & n205 ;
  assign n18672 = ~x115 & n162 ;
  assign n18673 = ~n18671 & ~n18672 ;
  assign n18674 = ~n18670 & n18673 ;
  assign n18675 = ~n17359 & ~n17681 ;
  assign n18676 = n18333 & ~n18675 ;
  assign n18677 = ~n18333 & n18675 ;
  assign n18678 = ~n18676 & ~n18677 ;
  assign n18679 = n167 & n18678 ;
  assign n18680 = n18674 & ~n18679 ;
  assign n18681 = ~x2 & ~n18680 ;
  assign n18682 = ~x2 & ~n18681 ;
  assign n18683 = ~n18680 & ~n18681 ;
  assign n18684 = ~n18682 & ~n18683 ;
  assign n18685 = ~n18669 & ~n18684 ;
  assign n18686 = n18669 & n18684 ;
  assign n18687 = ~n18685 & ~n18686 ;
  assign n18688 = ~n18349 & n18687 ;
  assign n18689 = n18349 & ~n18687 ;
  assign n18690 = ~n18688 & ~n18689 ;
  assign n18693 = ~n18690 & ~x180 ;
  assign n18694 = ~n18692 & ~n18693 ;
  assign n18695 = ~n18343 & ~n18346 ;
  assign n18696 = ~n17995 & ~n18321 ;
  assign n18697 = ~n18318 & ~n18696 ;
  assign n18698 = ~n18202 & ~n18208 ;
  assign n18699 = x96 & n3589 ;
  assign n18700 = x94 & n3878 ;
  assign n18701 = x95 & n3584 ;
  assign n18702 = ~n18700 & ~n18701 ;
  assign n18703 = ~n18699 & n18702 ;
  assign n18704 = n3592 & n7321 ;
  assign n18705 = n18703 & ~n18704 ;
  assign n18706 = x23 & ~n18705 ;
  assign n18707 = x23 & ~n18706 ;
  assign n18708 = ~n18705 & ~n18706 ;
  assign n18709 = ~n18707 & ~n18708 ;
  assign n18710 = ~n18185 & ~n18189 ;
  assign n18711 = x93 & n4531 ;
  assign n18712 = x91 & n4847 ;
  assign n18713 = x92 & n4526 ;
  assign n18714 = ~n18712 & ~n18713 ;
  assign n18715 = ~n18711 & n18714 ;
  assign n18716 = n4534 & n6094 ;
  assign n18717 = n18715 & ~n18716 ;
  assign n18718 = x26 & ~n18717 ;
  assign n18719 = x26 & ~n18718 ;
  assign n18720 = ~n18717 & ~n18718 ;
  assign n18721 = ~n18719 & ~n18720 ;
  assign n18722 = ~n17999 & ~n18170 ;
  assign n18723 = ~n18167 & ~n18722 ;
  assign n18724 = ~n18148 & ~n18154 ;
  assign n18725 = x87 & n6725 ;
  assign n18726 = x85 & n7129 ;
  assign n18727 = x86 & n6720 ;
  assign n18728 = ~n18726 & ~n18727 ;
  assign n18729 = ~n18725 & n18728 ;
  assign n18730 = n3991 & n6728 ;
  assign n18731 = n18729 & ~n18730 ;
  assign n18732 = x32 & ~n18731 ;
  assign n18733 = x32 & ~n18732 ;
  assign n18734 = ~n18731 & ~n18732 ;
  assign n18735 = ~n18733 & ~n18734 ;
  assign n18736 = ~n18110 & ~n18116 ;
  assign n18737 = x81 & n9433 ;
  assign n18738 = x79 & n9915 ;
  assign n18739 = x80 & n9428 ;
  assign n18740 = ~n18738 & ~n18739 ;
  assign n18741 = ~n18737 & n18740 ;
  assign n18742 = n2348 & n9436 ;
  assign n18743 = n18741 & ~n18742 ;
  assign n18744 = x38 & ~n18743 ;
  assign n18745 = x38 & ~n18744 ;
  assign n18746 = ~n18743 & ~n18744 ;
  assign n18747 = ~n18745 & ~n18746 ;
  assign n18748 = ~n18094 & ~n18096 ;
  assign n18749 = x75 & n12506 ;
  assign n18750 = x73 & n13131 ;
  assign n18751 = x74 & n12501 ;
  assign n18752 = ~n18750 & ~n18751 ;
  assign n18753 = ~n18749 & n18752 ;
  assign n18754 = n1150 & n12509 ;
  assign n18755 = n18753 & ~n18754 ;
  assign n18756 = x44 & ~n18755 ;
  assign n18757 = x44 & ~n18756 ;
  assign n18758 = ~n18755 & ~n18756 ;
  assign n18759 = ~n18757 & ~n18758 ;
  assign n18760 = ~n18055 & ~n18061 ;
  assign n18761 = ~n18039 & ~n18041 ;
  assign n18762 = x66 & n18025 ;
  assign n18763 = n17415 & ~n18024 ;
  assign n18764 = n18019 & n18763 ;
  assign n18765 = x64 & n18764 ;
  assign n18766 = x65 & n18020 ;
  assign n18767 = ~n18765 & ~n18766 ;
  assign n18768 = ~n18762 & n18767 ;
  assign n18769 = n194 & n18028 ;
  assign n18770 = n18768 & ~n18769 ;
  assign n18771 = x53 & ~n18770 ;
  assign n18772 = x53 & ~n18771 ;
  assign n18773 = ~n18770 & ~n18771 ;
  assign n18774 = ~n18772 & ~n18773 ;
  assign n18775 = ~n18035 & n18774 ;
  assign n18776 = n18035 & ~n18774 ;
  assign n18777 = ~n18775 & ~n18776 ;
  assign n18778 = x69 & n16076 ;
  assign n18779 = x67 & n16756 ;
  assign n18780 = x68 & n16071 ;
  assign n18781 = ~n18779 & ~n18780 ;
  assign n18782 = ~n18778 & n18781 ;
  assign n18783 = n398 & n16079 ;
  assign n18784 = n18782 & ~n18783 ;
  assign n18785 = x50 & ~n18784 ;
  assign n18786 = x50 & ~n18785 ;
  assign n18787 = ~n18784 & ~n18785 ;
  assign n18788 = ~n18786 & ~n18787 ;
  assign n18789 = n18777 & ~n18788 ;
  assign n18790 = ~n18777 & n18788 ;
  assign n18791 = ~n18761 & ~n18790 ;
  assign n18792 = ~n18789 & n18791 ;
  assign n18793 = ~n18761 & ~n18792 ;
  assign n18794 = ~n18789 & ~n18792 ;
  assign n18795 = ~n18790 & n18794 ;
  assign n18796 = ~n18793 & ~n18795 ;
  assign n18797 = x72 & n14233 ;
  assign n18798 = x70 & n14876 ;
  assign n18799 = x71 & n14228 ;
  assign n18800 = ~n18798 & ~n18799 ;
  assign n18801 = ~n18797 & n18800 ;
  assign n18802 = n717 & n14236 ;
  assign n18803 = n18801 & ~n18802 ;
  assign n18804 = x47 & ~n18803 ;
  assign n18805 = x47 & ~n18804 ;
  assign n18806 = ~n18803 & ~n18804 ;
  assign n18807 = ~n18805 & ~n18806 ;
  assign n18808 = n18796 & n18807 ;
  assign n18809 = ~n18796 & ~n18807 ;
  assign n18810 = ~n18808 & ~n18809 ;
  assign n18811 = ~n18760 & n18810 ;
  assign n18812 = n18760 & ~n18810 ;
  assign n18813 = ~n18811 & ~n18812 ;
  assign n18814 = n18759 & ~n18813 ;
  assign n18815 = ~n18759 & n18813 ;
  assign n18816 = ~n18814 & ~n18815 ;
  assign n18817 = ~n18079 & n18816 ;
  assign n18818 = n18079 & ~n18816 ;
  assign n18819 = ~n18817 & ~n18818 ;
  assign n18820 = x78 & n10905 ;
  assign n18821 = x76 & n11466 ;
  assign n18822 = x77 & n10900 ;
  assign n18823 = ~n18821 & ~n18822 ;
  assign n18824 = ~n18820 & n18823 ;
  assign n18825 = n1624 & n10908 ;
  assign n18826 = n18824 & ~n18825 ;
  assign n18827 = x41 & ~n18826 ;
  assign n18828 = x41 & ~n18827 ;
  assign n18829 = ~n18826 & ~n18827 ;
  assign n18830 = ~n18828 & ~n18829 ;
  assign n18831 = n18819 & ~n18830 ;
  assign n18832 = n18819 & ~n18831 ;
  assign n18833 = ~n18830 & ~n18831 ;
  assign n18834 = ~n18832 & ~n18833 ;
  assign n18835 = ~n18748 & ~n18834 ;
  assign n18836 = n18748 & n18834 ;
  assign n18837 = ~n18835 & ~n18836 ;
  assign n18838 = ~n18747 & n18837 ;
  assign n18839 = ~n18747 & ~n18838 ;
  assign n18840 = n18837 & ~n18838 ;
  assign n18841 = ~n18839 & ~n18840 ;
  assign n18842 = ~n18736 & ~n18841 ;
  assign n18843 = ~n18736 & ~n18842 ;
  assign n18844 = ~n18841 & ~n18842 ;
  assign n18845 = ~n18843 & ~n18844 ;
  assign n18846 = x84 & n8006 ;
  assign n18847 = x82 & n8474 ;
  assign n18848 = x83 & n8001 ;
  assign n18849 = ~n18847 & ~n18848 ;
  assign n18850 = ~n18846 & n18849 ;
  assign n18851 = n3114 & n8009 ;
  assign n18852 = n18850 & ~n18851 ;
  assign n18853 = x35 & ~n18852 ;
  assign n18854 = x35 & ~n18853 ;
  assign n18855 = ~n18852 & ~n18853 ;
  assign n18856 = ~n18854 & ~n18855 ;
  assign n18857 = ~n18845 & ~n18856 ;
  assign n18858 = ~n18845 & ~n18857 ;
  assign n18859 = ~n18856 & ~n18857 ;
  assign n18860 = ~n18858 & ~n18859 ;
  assign n18861 = ~n18134 & ~n18860 ;
  assign n18862 = n18134 & n18860 ;
  assign n18863 = ~n18861 & ~n18862 ;
  assign n18864 = ~n18735 & n18863 ;
  assign n18865 = ~n18735 & ~n18864 ;
  assign n18866 = n18863 & ~n18864 ;
  assign n18867 = ~n18865 & ~n18866 ;
  assign n18868 = ~n18724 & ~n18867 ;
  assign n18869 = ~n18724 & ~n18868 ;
  assign n18870 = ~n18867 & ~n18868 ;
  assign n18871 = ~n18869 & ~n18870 ;
  assign n18872 = x90 & n5560 ;
  assign n18873 = x88 & n5943 ;
  assign n18874 = x89 & n5555 ;
  assign n18875 = ~n18873 & ~n18874 ;
  assign n18876 = ~n18872 & n18875 ;
  assign n18877 = n4986 & n5563 ;
  assign n18878 = n18876 & ~n18877 ;
  assign n18879 = x29 & ~n18878 ;
  assign n18880 = x29 & ~n18879 ;
  assign n18881 = ~n18878 & ~n18879 ;
  assign n18882 = ~n18880 & ~n18881 ;
  assign n18883 = n18871 & n18882 ;
  assign n18884 = ~n18871 & ~n18882 ;
  assign n18885 = ~n18883 & ~n18884 ;
  assign n18886 = ~n18723 & n18885 ;
  assign n18887 = n18723 & ~n18885 ;
  assign n18888 = ~n18886 & ~n18887 ;
  assign n18889 = n18721 & ~n18888 ;
  assign n18890 = ~n18721 & n18888 ;
  assign n18891 = ~n18889 & ~n18890 ;
  assign n18892 = ~n18710 & n18891 ;
  assign n18893 = n18710 & ~n18891 ;
  assign n18894 = ~n18892 & ~n18893 ;
  assign n18895 = n18709 & ~n18894 ;
  assign n18896 = ~n18709 & n18894 ;
  assign n18897 = ~n18895 & ~n18896 ;
  assign n18898 = ~n18698 & n18897 ;
  assign n18899 = n18698 & ~n18897 ;
  assign n18900 = ~n18898 & ~n18899 ;
  assign n18901 = x99 & n2751 ;
  assign n18902 = x97 & n3020 ;
  assign n18903 = x98 & n2746 ;
  assign n18904 = ~n18902 & ~n18903 ;
  assign n18905 = ~n18901 & n18904 ;
  assign n18906 = n2754 & n8660 ;
  assign n18907 = n18905 & ~n18906 ;
  assign n18908 = x20 & ~n18907 ;
  assign n18909 = x20 & ~n18908 ;
  assign n18910 = ~n18907 & ~n18908 ;
  assign n18911 = ~n18909 & ~n18910 ;
  assign n18912 = n18900 & ~n18911 ;
  assign n18913 = n18900 & ~n18912 ;
  assign n18914 = ~n18911 & ~n18912 ;
  assign n18915 = ~n18913 & ~n18914 ;
  assign n18916 = ~n18221 & ~n18228 ;
  assign n18917 = n18915 & n18916 ;
  assign n18918 = ~n18915 & ~n18916 ;
  assign n18919 = ~n18917 & ~n18918 ;
  assign n18920 = x102 & n2093 ;
  assign n18921 = x100 & n2275 ;
  assign n18922 = x101 & n2088 ;
  assign n18923 = ~n18921 & ~n18922 ;
  assign n18924 = ~n18920 & n18923 ;
  assign n18925 = n2096 & n10092 ;
  assign n18926 = n18924 & ~n18925 ;
  assign n18927 = x17 & ~n18926 ;
  assign n18928 = x17 & ~n18927 ;
  assign n18929 = ~n18926 & ~n18927 ;
  assign n18930 = ~n18928 & ~n18929 ;
  assign n18931 = n18919 & ~n18930 ;
  assign n18932 = n18919 & ~n18931 ;
  assign n18933 = ~n18930 & ~n18931 ;
  assign n18934 = ~n18932 & ~n18933 ;
  assign n18935 = ~n18241 & ~n18247 ;
  assign n18936 = n18934 & n18935 ;
  assign n18937 = ~n18934 & ~n18935 ;
  assign n18938 = ~n18936 & ~n18937 ;
  assign n18939 = x105 & n1434 ;
  assign n18940 = x103 & n1646 ;
  assign n18941 = x104 & n1429 ;
  assign n18942 = ~n18940 & ~n18941 ;
  assign n18943 = ~n18939 & n18942 ;
  assign n18944 = n1437 & n11648 ;
  assign n18945 = n18943 & ~n18944 ;
  assign n18946 = x14 & ~n18945 ;
  assign n18947 = x14 & ~n18946 ;
  assign n18948 = ~n18945 & ~n18946 ;
  assign n18949 = ~n18947 & ~n18948 ;
  assign n18950 = n18938 & ~n18949 ;
  assign n18951 = n18938 & ~n18950 ;
  assign n18952 = ~n18949 & ~n18950 ;
  assign n18953 = ~n18951 & ~n18952 ;
  assign n18954 = ~n18260 & ~n18266 ;
  assign n18955 = n18953 & n18954 ;
  assign n18956 = ~n18953 & ~n18954 ;
  assign n18957 = ~n18955 & ~n18956 ;
  assign n18958 = x108 & n945 ;
  assign n18959 = x106 & n1099 ;
  assign n18960 = x107 & n940 ;
  assign n18961 = ~n18959 & ~n18960 ;
  assign n18962 = ~n18958 & n18961 ;
  assign n18963 = n948 & n13323 ;
  assign n18964 = n18962 & ~n18963 ;
  assign n18965 = x11 & ~n18964 ;
  assign n18966 = x11 & ~n18965 ;
  assign n18967 = ~n18964 & ~n18965 ;
  assign n18968 = ~n18966 & ~n18967 ;
  assign n18969 = n18957 & ~n18968 ;
  assign n18970 = ~n18957 & n18968 ;
  assign n18971 = ~n18284 & ~n18970 ;
  assign n18972 = ~n18969 & n18971 ;
  assign n18973 = ~n18284 & ~n18972 ;
  assign n18974 = ~n18969 & ~n18972 ;
  assign n18975 = ~n18970 & n18974 ;
  assign n18976 = ~n18973 & ~n18975 ;
  assign n18977 = x111 & n574 ;
  assign n18978 = x109 & n673 ;
  assign n18979 = x110 & n569 ;
  assign n18980 = ~n18978 & ~n18979 ;
  assign n18981 = ~n18977 & n18980 ;
  assign n18982 = n577 & n15111 ;
  assign n18983 = n18981 & ~n18982 ;
  assign n18984 = x8 & ~n18983 ;
  assign n18985 = x8 & ~n18984 ;
  assign n18986 = ~n18983 & ~n18984 ;
  assign n18987 = ~n18985 & ~n18986 ;
  assign n18988 = ~n18976 & ~n18987 ;
  assign n18989 = ~n18976 & ~n18988 ;
  assign n18990 = ~n18987 & ~n18988 ;
  assign n18991 = ~n18989 & ~n18990 ;
  assign n18992 = ~n18298 & ~n18305 ;
  assign n18993 = n18991 & n18992 ;
  assign n18994 = ~n18991 & ~n18992 ;
  assign n18995 = ~n18993 & ~n18994 ;
  assign n18996 = x114 & n293 ;
  assign n18997 = x112 & n373 ;
  assign n18998 = x113 & n288 ;
  assign n18999 = ~n18997 & ~n18998 ;
  assign n19000 = ~n18996 & n18999 ;
  assign n19001 = n296 & n17012 ;
  assign n19002 = n19000 & ~n19001 ;
  assign n19003 = x5 & ~n19002 ;
  assign n19004 = x5 & ~n19003 ;
  assign n19005 = ~n19002 & ~n19003 ;
  assign n19006 = ~n19004 & ~n19005 ;
  assign n19007 = n18995 & ~n19006 ;
  assign n19008 = ~n18995 & n19006 ;
  assign n19009 = ~n18697 & ~n19008 ;
  assign n19010 = ~n19007 & n19009 ;
  assign n19011 = ~n18697 & ~n19010 ;
  assign n19012 = ~n19007 & ~n19010 ;
  assign n19013 = ~n19008 & n19012 ;
  assign n19014 = ~n19011 & ~n19013 ;
  assign n19015 = x117 & n146 ;
  assign n19016 = x115 & n182 ;
  assign n19017 = x116 & n141 ;
  assign n19018 = ~n19016 & ~n19017 ;
  assign n19019 = ~n19015 & n19018 ;
  assign n19020 = ~n18332 & ~n18334 ;
  assign n19021 = ~x116 & ~x117 ;
  assign n19022 = x116 & x117 ;
  assign n19023 = ~n19021 & ~n19022 ;
  assign n19024 = ~n19020 & n19023 ;
  assign n19025 = n19020 & ~n19023 ;
  assign n19026 = ~n19024 & ~n19025 ;
  assign n19027 = n149 & n19026 ;
  assign n19028 = n19019 & ~n19027 ;
  assign n19029 = x2 & ~n19028 ;
  assign n19030 = x2 & ~n19029 ;
  assign n19031 = ~n19028 & ~n19029 ;
  assign n19032 = ~n19030 & ~n19031 ;
  assign n19033 = ~n19014 & n19032 ;
  assign n19034 = n19014 & ~n19032 ;
  assign n19035 = ~n19033 & ~n19034 ;
  assign n19036 = ~n18695 & ~n19035 ;
  assign n19037 = n18695 & n19035 ;
  assign n19038 = ~n19036 & ~n19037 ;
  assign n19379 = n19038 & x181 ;
  assign n19039 = ~n18685 & ~n18688 ;
  assign n19040 = ~n18350 & ~n18666 ;
  assign n19041 = ~n18663 & ~n19040 ;
  assign n19042 = ~n18547 & ~n18553 ;
  assign n19043 = ~x96 & n3589 ;
  assign n19044 = ~x94 & n3878 ;
  assign n19045 = ~x95 & n3584 ;
  assign n19046 = ~n19044 & ~n19045 ;
  assign n19047 = ~n19043 & n19046 ;
  assign n19048 = n3592 & n7531 ;
  assign n19049 = n19047 & ~n19048 ;
  assign n19050 = ~x23 & ~n19049 ;
  assign n19051 = ~x23 & ~n19050 ;
  assign n19052 = ~n19049 & ~n19050 ;
  assign n19053 = ~n19051 & ~n19052 ;
  assign n19054 = ~n18530 & ~n18534 ;
  assign n19055 = ~x93 & n4531 ;
  assign n19056 = ~x91 & n4847 ;
  assign n19057 = ~x92 & n4526 ;
  assign n19058 = ~n19056 & ~n19057 ;
  assign n19059 = ~n19055 & n19058 ;
  assign n19060 = n4534 & n6285 ;
  assign n19061 = n19059 & ~n19060 ;
  assign n19062 = ~x26 & ~n19061 ;
  assign n19063 = ~x26 & ~n19062 ;
  assign n19064 = ~n19061 & ~n19062 ;
  assign n19065 = ~n19063 & ~n19064 ;
  assign n19066 = ~n18354 & ~n18515 ;
  assign n19067 = ~n18512 & ~n19066 ;
  assign n19068 = ~n18493 & ~n18499 ;
  assign n19069 = ~x87 & n6725 ;
  assign n19070 = ~x85 & n7129 ;
  assign n19071 = ~x86 & n6720 ;
  assign n19072 = ~n19070 & ~n19071 ;
  assign n19073 = ~n19069 & n19072 ;
  assign n19074 = n4143 & n6728 ;
  assign n19075 = n19073 & ~n19074 ;
  assign n19076 = ~x32 & ~n19075 ;
  assign n19077 = ~x32 & ~n19076 ;
  assign n19078 = ~n19075 & ~n19076 ;
  assign n19079 = ~n19077 & ~n19078 ;
  assign n19080 = ~n18455 & ~n18461 ;
  assign n19081 = ~x81 & n9433 ;
  assign n19082 = ~x79 & n9915 ;
  assign n19083 = ~x80 & n9428 ;
  assign n19084 = ~n19082 & ~n19083 ;
  assign n19085 = ~n19081 & n19084 ;
  assign n19086 = n2460 & n9436 ;
  assign n19087 = n19085 & ~n19086 ;
  assign n19088 = ~x38 & ~n19087 ;
  assign n19089 = ~x38 & ~n19088 ;
  assign n19090 = ~n19087 & ~n19088 ;
  assign n19091 = ~n19089 & ~n19090 ;
  assign n19092 = ~n18439 & ~n18441 ;
  assign n19093 = ~x75 & n12506 ;
  assign n19094 = ~x73 & n13131 ;
  assign n19095 = ~x74 & n12501 ;
  assign n19096 = ~n19094 & ~n19095 ;
  assign n19097 = ~n19093 & n19096 ;
  assign n19098 = n1225 & n12509 ;
  assign n19099 = n19097 & ~n19098 ;
  assign n19100 = ~x44 & ~n19099 ;
  assign n19101 = ~x44 & ~n19100 ;
  assign n19102 = ~n19099 & ~n19100 ;
  assign n19103 = ~n19101 & ~n19102 ;
  assign n19104 = ~n18400 & ~n18406 ;
  assign n19105 = ~n18384 & ~n18386 ;
  assign n19106 = ~x66 & n18025 ;
  assign n19107 = ~x64 & n18764 ;
  assign n19108 = ~x65 & n18020 ;
  assign n19109 = ~n19107 & ~n19108 ;
  assign n19110 = ~n19106 & n19109 ;
  assign n19111 = n214 & n18028 ;
  assign n19112 = n19110 & ~n19111 ;
  assign n19113 = ~x53 & ~n19112 ;
  assign n19114 = ~x53 & ~n19113 ;
  assign n19115 = ~n19112 & ~n19113 ;
  assign n19116 = ~n19114 & ~n19115 ;
  assign n19117 = ~n18380 & n19116 ;
  assign n19118 = n18380 & ~n19116 ;
  assign n19119 = ~n19117 & ~n19118 ;
  assign n19120 = ~x69 & n16076 ;
  assign n19121 = ~x67 & n16756 ;
  assign n19122 = ~x68 & n16071 ;
  assign n19123 = ~n19121 & ~n19122 ;
  assign n19124 = ~n19120 & n19123 ;
  assign n19125 = n435 & n16079 ;
  assign n19126 = n19124 & ~n19125 ;
  assign n19127 = ~x50 & ~n19126 ;
  assign n19128 = ~x50 & ~n19127 ;
  assign n19129 = ~n19126 & ~n19127 ;
  assign n19130 = ~n19128 & ~n19129 ;
  assign n19131 = n19119 & ~n19130 ;
  assign n19132 = ~n19119 & n19130 ;
  assign n19133 = ~n19105 & ~n19132 ;
  assign n19134 = ~n19131 & n19133 ;
  assign n19135 = ~n19105 & ~n19134 ;
  assign n19136 = ~n19131 & ~n19134 ;
  assign n19137 = ~n19132 & n19136 ;
  assign n19138 = ~n19135 & ~n19137 ;
  assign n19139 = ~x72 & n14233 ;
  assign n19140 = ~x70 & n14876 ;
  assign n19141 = ~x71 & n14228 ;
  assign n19142 = ~n19140 & ~n19141 ;
  assign n19143 = ~n19139 & n19142 ;
  assign n19144 = n773 & n14236 ;
  assign n19145 = n19143 & ~n19144 ;
  assign n19146 = ~x47 & ~n19145 ;
  assign n19147 = ~x47 & ~n19146 ;
  assign n19148 = ~n19145 & ~n19146 ;
  assign n19149 = ~n19147 & ~n19148 ;
  assign n19150 = n19138 & n19149 ;
  assign n19151 = ~n19138 & ~n19149 ;
  assign n19152 = ~n19150 & ~n19151 ;
  assign n19153 = ~n19104 & n19152 ;
  assign n19154 = n19104 & ~n19152 ;
  assign n19155 = ~n19153 & ~n19154 ;
  assign n19156 = n19103 & ~n19155 ;
  assign n19157 = ~n19103 & n19155 ;
  assign n19158 = ~n19156 & ~n19157 ;
  assign n19159 = ~n18424 & n19158 ;
  assign n19160 = n18424 & ~n19158 ;
  assign n19161 = ~n19159 & ~n19160 ;
  assign n19162 = ~x78 & n10905 ;
  assign n19163 = ~x76 & n11466 ;
  assign n19164 = ~x77 & n10900 ;
  assign n19165 = ~n19163 & ~n19164 ;
  assign n19166 = ~n19162 & n19165 ;
  assign n19167 = n1718 & n10908 ;
  assign n19168 = n19166 & ~n19167 ;
  assign n19169 = ~x41 & ~n19168 ;
  assign n19170 = ~x41 & ~n19169 ;
  assign n19171 = ~n19168 & ~n19169 ;
  assign n19172 = ~n19170 & ~n19171 ;
  assign n19173 = n19161 & ~n19172 ;
  assign n19174 = n19161 & ~n19173 ;
  assign n19175 = ~n19172 & ~n19173 ;
  assign n19176 = ~n19174 & ~n19175 ;
  assign n19177 = ~n19092 & ~n19176 ;
  assign n19178 = n19092 & n19176 ;
  assign n19179 = ~n19177 & ~n19178 ;
  assign n19180 = ~n19091 & n19179 ;
  assign n19181 = ~n19091 & ~n19180 ;
  assign n19182 = n19179 & ~n19180 ;
  assign n19183 = ~n19181 & ~n19182 ;
  assign n19184 = ~n19080 & ~n19183 ;
  assign n19185 = ~n19080 & ~n19184 ;
  assign n19186 = ~n19183 & ~n19184 ;
  assign n19187 = ~n19185 & ~n19186 ;
  assign n19188 = ~x84 & n8006 ;
  assign n19189 = ~x82 & n8474 ;
  assign n19190 = ~x83 & n8001 ;
  assign n19191 = ~n19189 & ~n19190 ;
  assign n19192 = ~n19188 & n19191 ;
  assign n19193 = n3247 & n8009 ;
  assign n19194 = n19192 & ~n19193 ;
  assign n19195 = ~x35 & ~n19194 ;
  assign n19196 = ~x35 & ~n19195 ;
  assign n19197 = ~n19194 & ~n19195 ;
  assign n19198 = ~n19196 & ~n19197 ;
  assign n19199 = ~n19187 & ~n19198 ;
  assign n19200 = ~n19187 & ~n19199 ;
  assign n19201 = ~n19198 & ~n19199 ;
  assign n19202 = ~n19200 & ~n19201 ;
  assign n19203 = ~n18479 & ~n19202 ;
  assign n19204 = n18479 & n19202 ;
  assign n19205 = ~n19203 & ~n19204 ;
  assign n19206 = ~n19079 & n19205 ;
  assign n19207 = ~n19079 & ~n19206 ;
  assign n19208 = n19205 & ~n19206 ;
  assign n19209 = ~n19207 & ~n19208 ;
  assign n19210 = ~n19068 & ~n19209 ;
  assign n19211 = ~n19068 & ~n19210 ;
  assign n19212 = ~n19209 & ~n19210 ;
  assign n19213 = ~n19211 & ~n19212 ;
  assign n19214 = ~x90 & n5560 ;
  assign n19215 = ~x88 & n5943 ;
  assign n19216 = ~x89 & n5555 ;
  assign n19217 = ~n19215 & ~n19216 ;
  assign n19218 = ~n19214 & n19217 ;
  assign n19219 = n5155 & n5563 ;
  assign n19220 = n19218 & ~n19219 ;
  assign n19221 = ~x29 & ~n19220 ;
  assign n19222 = ~x29 & ~n19221 ;
  assign n19223 = ~n19220 & ~n19221 ;
  assign n19224 = ~n19222 & ~n19223 ;
  assign n19225 = n19213 & n19224 ;
  assign n19226 = ~n19213 & ~n19224 ;
  assign n19227 = ~n19225 & ~n19226 ;
  assign n19228 = ~n19067 & n19227 ;
  assign n19229 = n19067 & ~n19227 ;
  assign n19230 = ~n19228 & ~n19229 ;
  assign n19231 = n19065 & ~n19230 ;
  assign n19232 = ~n19065 & n19230 ;
  assign n19233 = ~n19231 & ~n19232 ;
  assign n19234 = ~n19054 & n19233 ;
  assign n19235 = n19054 & ~n19233 ;
  assign n19236 = ~n19234 & ~n19235 ;
  assign n19237 = n19053 & ~n19236 ;
  assign n19238 = ~n19053 & n19236 ;
  assign n19239 = ~n19237 & ~n19238 ;
  assign n19240 = ~n19042 & n19239 ;
  assign n19241 = n19042 & ~n19239 ;
  assign n19242 = ~n19240 & ~n19241 ;
  assign n19243 = ~x99 & n2751 ;
  assign n19244 = ~x97 & n3020 ;
  assign n19245 = ~x98 & n2746 ;
  assign n19246 = ~n19244 & ~n19245 ;
  assign n19247 = ~n19243 & n19246 ;
  assign n19248 = n2754 & n8885 ;
  assign n19249 = n19247 & ~n19248 ;
  assign n19250 = ~x20 & ~n19249 ;
  assign n19251 = ~x20 & ~n19250 ;
  assign n19252 = ~n19249 & ~n19250 ;
  assign n19253 = ~n19251 & ~n19252 ;
  assign n19254 = n19242 & ~n19253 ;
  assign n19255 = n19242 & ~n19254 ;
  assign n19256 = ~n19253 & ~n19254 ;
  assign n19257 = ~n19255 & ~n19256 ;
  assign n19258 = ~n18566 & ~n18573 ;
  assign n19259 = n19257 & n19258 ;
  assign n19260 = ~n19257 & ~n19258 ;
  assign n19261 = ~n19259 & ~n19260 ;
  assign n19262 = ~x102 & n2093 ;
  assign n19263 = ~x100 & n2275 ;
  assign n19264 = ~x101 & n2088 ;
  assign n19265 = ~n19263 & ~n19264 ;
  assign n19266 = ~n19262 & n19265 ;
  assign n19267 = n2096 & n10333 ;
  assign n19268 = n19266 & ~n19267 ;
  assign n19269 = ~x17 & ~n19268 ;
  assign n19270 = ~x17 & ~n19269 ;
  assign n19271 = ~n19268 & ~n19269 ;
  assign n19272 = ~n19270 & ~n19271 ;
  assign n19273 = n19261 & ~n19272 ;
  assign n19274 = n19261 & ~n19273 ;
  assign n19275 = ~n19272 & ~n19273 ;
  assign n19276 = ~n19274 & ~n19275 ;
  assign n19277 = ~n18586 & ~n18592 ;
  assign n19278 = n19276 & n19277 ;
  assign n19279 = ~n19276 & ~n19277 ;
  assign n19280 = ~n19278 & ~n19279 ;
  assign n19281 = ~x105 & n1434 ;
  assign n19282 = ~x103 & n1646 ;
  assign n19283 = ~x104 & n1429 ;
  assign n19284 = ~n19282 & ~n19283 ;
  assign n19285 = ~n19281 & n19284 ;
  assign n19286 = n1437 & n11907 ;
  assign n19287 = n19285 & ~n19286 ;
  assign n19288 = ~x14 & ~n19287 ;
  assign n19289 = ~x14 & ~n19288 ;
  assign n19290 = ~n19287 & ~n19288 ;
  assign n19291 = ~n19289 & ~n19290 ;
  assign n19292 = n19280 & ~n19291 ;
  assign n19293 = n19280 & ~n19292 ;
  assign n19294 = ~n19291 & ~n19292 ;
  assign n19295 = ~n19293 & ~n19294 ;
  assign n19296 = ~n18605 & ~n18611 ;
  assign n19297 = n19295 & n19296 ;
  assign n19298 = ~n19295 & ~n19296 ;
  assign n19299 = ~n19297 & ~n19298 ;
  assign n19300 = ~x108 & n945 ;
  assign n19301 = ~x106 & n1099 ;
  assign n19302 = ~x107 & n940 ;
  assign n19303 = ~n19301 & ~n19302 ;
  assign n19304 = ~n19300 & n19303 ;
  assign n19305 = n948 & n13601 ;
  assign n19306 = n19304 & ~n19305 ;
  assign n19307 = ~x11 & ~n19306 ;
  assign n19308 = ~x11 & ~n19307 ;
  assign n19309 = ~n19306 & ~n19307 ;
  assign n19310 = ~n19308 & ~n19309 ;
  assign n19311 = n19299 & ~n19310 ;
  assign n19312 = ~n19299 & n19310 ;
  assign n19313 = ~n18629 & ~n19312 ;
  assign n19314 = ~n19311 & n19313 ;
  assign n19315 = ~n18629 & ~n19314 ;
  assign n19316 = ~n19311 & ~n19314 ;
  assign n19317 = ~n19312 & n19316 ;
  assign n19318 = ~n19315 & ~n19317 ;
  assign n19319 = ~x111 & n574 ;
  assign n19320 = ~x109 & n673 ;
  assign n19321 = ~x110 & n569 ;
  assign n19322 = ~n19320 & ~n19321 ;
  assign n19323 = ~n19319 & n19322 ;
  assign n19324 = n577 & n15411 ;
  assign n19325 = n19323 & ~n19324 ;
  assign n19326 = ~x8 & ~n19325 ;
  assign n19327 = ~x8 & ~n19326 ;
  assign n19328 = ~n19325 & ~n19326 ;
  assign n19329 = ~n19327 & ~n19328 ;
  assign n19330 = ~n19318 & ~n19329 ;
  assign n19331 = ~n19318 & ~n19330 ;
  assign n19332 = ~n19329 & ~n19330 ;
  assign n19333 = ~n19331 & ~n19332 ;
  assign n19334 = ~n18643 & ~n18650 ;
  assign n19335 = n19333 & n19334 ;
  assign n19336 = ~n19333 & ~n19334 ;
  assign n19337 = ~n19335 & ~n19336 ;
  assign n19338 = ~x114 & n293 ;
  assign n19339 = ~x112 & n373 ;
  assign n19340 = ~x113 & n288 ;
  assign n19341 = ~n19339 & ~n19340 ;
  assign n19342 = ~n19338 & n19341 ;
  assign n19343 = n296 & n17333 ;
  assign n19344 = n19342 & ~n19343 ;
  assign n19345 = ~x5 & ~n19344 ;
  assign n19346 = ~x5 & ~n19345 ;
  assign n19347 = ~n19344 & ~n19345 ;
  assign n19348 = ~n19346 & ~n19347 ;
  assign n19349 = n19337 & ~n19348 ;
  assign n19350 = ~n19337 & n19348 ;
  assign n19351 = ~n19041 & ~n19350 ;
  assign n19352 = ~n19349 & n19351 ;
  assign n19353 = ~n19041 & ~n19352 ;
  assign n19354 = ~n19349 & ~n19352 ;
  assign n19355 = ~n19350 & n19354 ;
  assign n19356 = ~n19353 & ~n19355 ;
  assign n19357 = ~x117 & n164 ;
  assign n19358 = ~x115 & n205 ;
  assign n19359 = ~x116 & n162 ;
  assign n19360 = ~n19358 & ~n19359 ;
  assign n19361 = ~n19357 & n19360 ;
  assign n19362 = ~n18331 & ~n18676 ;
  assign n19363 = n19023 & ~n19362 ;
  assign n19364 = ~n19023 & n19362 ;
  assign n19365 = ~n19363 & ~n19364 ;
  assign n19366 = n167 & n19365 ;
  assign n19367 = n19361 & ~n19366 ;
  assign n19368 = ~x2 & ~n19367 ;
  assign n19369 = ~x2 & ~n19368 ;
  assign n19370 = ~n19367 & ~n19368 ;
  assign n19371 = ~n19369 & ~n19370 ;
  assign n19372 = ~n19356 & n19371 ;
  assign n19373 = n19356 & ~n19371 ;
  assign n19374 = ~n19372 & ~n19373 ;
  assign n19375 = ~n19039 & ~n19374 ;
  assign n19376 = n19039 & n19374 ;
  assign n19377 = ~n19375 & ~n19376 ;
  assign n19380 = ~n19377 & ~x181 ;
  assign n19381 = ~n19379 & ~n19380 ;
  assign n19382 = ~n19014 & ~n19032 ;
  assign n19383 = ~n19036 & ~n19382 ;
  assign n19384 = x118 & n146 ;
  assign n19385 = x116 & n182 ;
  assign n19386 = x117 & n141 ;
  assign n19387 = ~n19385 & ~n19386 ;
  assign n19388 = ~n19384 & n19387 ;
  assign n19389 = ~n19022 & ~n19024 ;
  assign n19390 = ~x117 & ~x118 ;
  assign n19391 = x117 & x118 ;
  assign n19392 = ~n19390 & ~n19391 ;
  assign n19393 = ~n19389 & n19392 ;
  assign n19394 = n19389 & ~n19392 ;
  assign n19395 = ~n19393 & ~n19394 ;
  assign n19396 = n149 & n19395 ;
  assign n19397 = n19388 & ~n19396 ;
  assign n19398 = x2 & ~n19397 ;
  assign n19399 = x2 & ~n19398 ;
  assign n19400 = ~n19397 & ~n19398 ;
  assign n19401 = ~n19399 & ~n19400 ;
  assign n19402 = x109 & n945 ;
  assign n19403 = x107 & n1099 ;
  assign n19404 = x108 & n940 ;
  assign n19405 = ~n19403 & ~n19404 ;
  assign n19406 = ~n19402 & n19405 ;
  assign n19407 = n948 & n13894 ;
  assign n19408 = n19406 & ~n19407 ;
  assign n19409 = x11 & ~n19408 ;
  assign n19410 = x11 & ~n19409 ;
  assign n19411 = ~n19408 & ~n19409 ;
  assign n19412 = ~n19410 & ~n19411 ;
  assign n19413 = ~n18950 & ~n18956 ;
  assign n19414 = ~n18912 & ~n18918 ;
  assign n19415 = ~n18896 & ~n18898 ;
  assign n19416 = ~n18890 & ~n18892 ;
  assign n19417 = x94 & n4531 ;
  assign n19418 = x92 & n4847 ;
  assign n19419 = x93 & n4526 ;
  assign n19420 = ~n19418 & ~n19419 ;
  assign n19421 = ~n19417 & n19420 ;
  assign n19422 = n4534 & n6483 ;
  assign n19423 = n19421 & ~n19422 ;
  assign n19424 = x26 & ~n19423 ;
  assign n19425 = x26 & ~n19424 ;
  assign n19426 = ~n19423 & ~n19424 ;
  assign n19427 = ~n19425 & ~n19426 ;
  assign n19428 = ~n18884 & ~n18886 ;
  assign n19429 = x91 & n5560 ;
  assign n19430 = x89 & n5943 ;
  assign n19431 = x90 & n5555 ;
  assign n19432 = ~n19430 & ~n19431 ;
  assign n19433 = ~n19429 & n19432 ;
  assign n19434 = n5336 & n5563 ;
  assign n19435 = n19433 & ~n19434 ;
  assign n19436 = x29 & ~n19435 ;
  assign n19437 = x29 & ~n19436 ;
  assign n19438 = ~n19435 & ~n19436 ;
  assign n19439 = ~n19437 & ~n19438 ;
  assign n19440 = ~n18864 & ~n18868 ;
  assign n19441 = x88 & n6725 ;
  assign n19442 = x86 & n7129 ;
  assign n19443 = x87 & n6720 ;
  assign n19444 = ~n19442 & ~n19443 ;
  assign n19445 = ~n19441 & n19444 ;
  assign n19446 = n4305 & n6728 ;
  assign n19447 = n19445 & ~n19446 ;
  assign n19448 = x32 & ~n19447 ;
  assign n19449 = x32 & ~n19448 ;
  assign n19450 = ~n19447 & ~n19448 ;
  assign n19451 = ~n19449 & ~n19450 ;
  assign n19452 = ~n18857 & ~n18861 ;
  assign n19453 = x85 & n8006 ;
  assign n19454 = x83 & n8474 ;
  assign n19455 = x84 & n8001 ;
  assign n19456 = ~n19454 & ~n19455 ;
  assign n19457 = ~n19453 & n19456 ;
  assign n19458 = n3389 & n8009 ;
  assign n19459 = n19457 & ~n19458 ;
  assign n19460 = x35 & ~n19459 ;
  assign n19461 = x35 & ~n19460 ;
  assign n19462 = ~n19459 & ~n19460 ;
  assign n19463 = ~n19461 & ~n19462 ;
  assign n19464 = ~n18838 & ~n18842 ;
  assign n19465 = x82 & n9433 ;
  assign n19466 = x80 & n9915 ;
  assign n19467 = x81 & n9428 ;
  assign n19468 = ~n19466 & ~n19467 ;
  assign n19469 = ~n19465 & n19468 ;
  assign n19470 = n2584 & n9436 ;
  assign n19471 = n19469 & ~n19470 ;
  assign n19472 = x38 & ~n19471 ;
  assign n19473 = x38 & ~n19472 ;
  assign n19474 = ~n19471 & ~n19472 ;
  assign n19475 = ~n19473 & ~n19474 ;
  assign n19476 = ~n18831 & ~n18835 ;
  assign n19477 = x79 & n10905 ;
  assign n19478 = x77 & n11466 ;
  assign n19479 = x78 & n10900 ;
  assign n19480 = ~n19478 & ~n19479 ;
  assign n19481 = ~n19477 & n19480 ;
  assign n19482 = n1817 & n10908 ;
  assign n19483 = n19481 & ~n19482 ;
  assign n19484 = x41 & ~n19483 ;
  assign n19485 = x41 & ~n19484 ;
  assign n19486 = ~n19483 & ~n19484 ;
  assign n19487 = ~n19485 & ~n19486 ;
  assign n19488 = ~n18815 & ~n18817 ;
  assign n19489 = x76 & n12506 ;
  assign n19490 = x74 & n13131 ;
  assign n19491 = x75 & n12501 ;
  assign n19492 = ~n19490 & ~n19491 ;
  assign n19493 = ~n19489 & n19492 ;
  assign n19494 = n1311 & n12509 ;
  assign n19495 = n19493 & ~n19494 ;
  assign n19496 = x44 & ~n19495 ;
  assign n19497 = x44 & ~n19496 ;
  assign n19498 = ~n19495 & ~n19496 ;
  assign n19499 = ~n19497 & ~n19498 ;
  assign n19500 = ~n18809 & ~n18811 ;
  assign n19501 = x73 & n14233 ;
  assign n19502 = x71 & n14876 ;
  assign n19503 = x72 & n14228 ;
  assign n19504 = ~n19502 & ~n19503 ;
  assign n19505 = ~n19501 & n19504 ;
  assign n19506 = n843 & n14236 ;
  assign n19507 = n19505 & ~n19506 ;
  assign n19508 = x47 & ~n19507 ;
  assign n19509 = x47 & ~n19508 ;
  assign n19510 = ~n19507 & ~n19508 ;
  assign n19511 = ~n19509 & ~n19510 ;
  assign n19512 = x53 & ~x54 ;
  assign n19513 = ~x53 & x54 ;
  assign n19514 = ~n19512 & ~n19513 ;
  assign n19515 = x64 & ~n19514 ;
  assign n19516 = ~n18776 & n19515 ;
  assign n19517 = n18776 & ~n19515 ;
  assign n19518 = ~n19516 & ~n19517 ;
  assign n19519 = x67 & n18025 ;
  assign n19520 = x65 & n18764 ;
  assign n19521 = x66 & n18020 ;
  assign n19522 = ~n19520 & ~n19521 ;
  assign n19523 = ~n19519 & n19522 ;
  assign n19524 = n240 & n18028 ;
  assign n19525 = n19523 & ~n19524 ;
  assign n19526 = x53 & ~n19525 ;
  assign n19527 = x53 & ~n19526 ;
  assign n19528 = ~n19525 & ~n19526 ;
  assign n19529 = ~n19527 & ~n19528 ;
  assign n19530 = ~n19518 & ~n19529 ;
  assign n19531 = n19518 & n19529 ;
  assign n19532 = ~n19530 & ~n19531 ;
  assign n19533 = x70 & n16076 ;
  assign n19534 = x68 & n16756 ;
  assign n19535 = x69 & n16071 ;
  assign n19536 = ~n19534 & ~n19535 ;
  assign n19537 = ~n19533 & n19536 ;
  assign n19538 = n488 & n16079 ;
  assign n19539 = n19537 & ~n19538 ;
  assign n19540 = x50 & ~n19539 ;
  assign n19541 = x50 & ~n19540 ;
  assign n19542 = ~n19539 & ~n19540 ;
  assign n19543 = ~n19541 & ~n19542 ;
  assign n19544 = n19532 & ~n19543 ;
  assign n19545 = n19532 & ~n19544 ;
  assign n19546 = ~n19543 & ~n19544 ;
  assign n19547 = ~n19545 & ~n19546 ;
  assign n19548 = ~n18794 & ~n19547 ;
  assign n19549 = n18794 & n19547 ;
  assign n19550 = ~n19548 & ~n19549 ;
  assign n19551 = ~n19511 & n19550 ;
  assign n19552 = ~n19511 & ~n19551 ;
  assign n19553 = n19550 & ~n19551 ;
  assign n19554 = ~n19552 & ~n19553 ;
  assign n19555 = ~n19500 & ~n19554 ;
  assign n19556 = n19500 & ~n19553 ;
  assign n19557 = ~n19552 & n19556 ;
  assign n19558 = ~n19555 & ~n19557 ;
  assign n19559 = ~n19499 & n19558 ;
  assign n19560 = ~n19499 & ~n19559 ;
  assign n19561 = n19558 & ~n19559 ;
  assign n19562 = ~n19560 & ~n19561 ;
  assign n19563 = ~n19488 & ~n19562 ;
  assign n19564 = n19488 & ~n19561 ;
  assign n19565 = ~n19560 & n19564 ;
  assign n19566 = ~n19563 & ~n19565 ;
  assign n19567 = ~n19487 & n19566 ;
  assign n19568 = n19487 & ~n19566 ;
  assign n19569 = ~n19567 & ~n19568 ;
  assign n19570 = ~n19476 & n19569 ;
  assign n19571 = n19476 & ~n19569 ;
  assign n19572 = ~n19570 & ~n19571 ;
  assign n19573 = ~n19475 & n19572 ;
  assign n19574 = ~n19475 & ~n19573 ;
  assign n19575 = n19572 & ~n19573 ;
  assign n19576 = ~n19574 & ~n19575 ;
  assign n19577 = ~n19464 & ~n19576 ;
  assign n19578 = n19464 & ~n19575 ;
  assign n19579 = ~n19574 & n19578 ;
  assign n19580 = ~n19577 & ~n19579 ;
  assign n19581 = ~n19463 & n19580 ;
  assign n19582 = n19463 & ~n19580 ;
  assign n19583 = ~n19581 & ~n19582 ;
  assign n19584 = ~n19452 & n19583 ;
  assign n19585 = n19452 & ~n19583 ;
  assign n19586 = ~n19584 & ~n19585 ;
  assign n19587 = ~n19451 & n19586 ;
  assign n19588 = n19451 & ~n19586 ;
  assign n19589 = ~n19587 & ~n19588 ;
  assign n19590 = ~n19440 & n19589 ;
  assign n19591 = n19440 & ~n19589 ;
  assign n19592 = ~n19590 & ~n19591 ;
  assign n19593 = ~n19439 & n19592 ;
  assign n19594 = n19439 & ~n19592 ;
  assign n19595 = ~n19593 & ~n19594 ;
  assign n19596 = ~n19428 & n19595 ;
  assign n19597 = n19428 & ~n19595 ;
  assign n19598 = ~n19596 & ~n19597 ;
  assign n19599 = ~n19427 & n19598 ;
  assign n19600 = n19427 & ~n19598 ;
  assign n19601 = ~n19599 & ~n19600 ;
  assign n19602 = ~n19416 & n19601 ;
  assign n19603 = n19416 & ~n19601 ;
  assign n19604 = ~n19602 & ~n19603 ;
  assign n19605 = x97 & n3589 ;
  assign n19606 = x95 & n3878 ;
  assign n19607 = x96 & n3584 ;
  assign n19608 = ~n19606 & ~n19607 ;
  assign n19609 = ~n19605 & n19608 ;
  assign n19610 = n3592 & n7745 ;
  assign n19611 = n19609 & ~n19610 ;
  assign n19612 = x23 & ~n19611 ;
  assign n19613 = x23 & ~n19612 ;
  assign n19614 = ~n19611 & ~n19612 ;
  assign n19615 = ~n19613 & ~n19614 ;
  assign n19616 = n19604 & ~n19615 ;
  assign n19617 = n19604 & ~n19616 ;
  assign n19618 = ~n19615 & ~n19616 ;
  assign n19619 = ~n19617 & ~n19618 ;
  assign n19620 = ~n19415 & n19619 ;
  assign n19621 = n19415 & ~n19619 ;
  assign n19622 = ~n19620 & ~n19621 ;
  assign n19623 = x100 & n2751 ;
  assign n19624 = x98 & n3020 ;
  assign n19625 = x99 & n2746 ;
  assign n19626 = ~n19624 & ~n19625 ;
  assign n19627 = ~n19623 & n19626 ;
  assign n19628 = n2754 & n9115 ;
  assign n19629 = n19627 & ~n19628 ;
  assign n19630 = x20 & ~n19629 ;
  assign n19631 = x20 & ~n19630 ;
  assign n19632 = ~n19629 & ~n19630 ;
  assign n19633 = ~n19631 & ~n19632 ;
  assign n19634 = ~n19622 & ~n19633 ;
  assign n19635 = n19622 & n19633 ;
  assign n19636 = ~n19634 & ~n19635 ;
  assign n19637 = n19414 & ~n19636 ;
  assign n19638 = ~n19414 & n19636 ;
  assign n19639 = ~n19637 & ~n19638 ;
  assign n19640 = x103 & n2093 ;
  assign n19641 = x101 & n2275 ;
  assign n19642 = x102 & n2088 ;
  assign n19643 = ~n19641 & ~n19642 ;
  assign n19644 = ~n19640 & n19643 ;
  assign n19645 = n2096 & n10588 ;
  assign n19646 = n19644 & ~n19645 ;
  assign n19647 = x17 & ~n19646 ;
  assign n19648 = x17 & ~n19647 ;
  assign n19649 = ~n19646 & ~n19647 ;
  assign n19650 = ~n19648 & ~n19649 ;
  assign n19651 = n19639 & ~n19650 ;
  assign n19652 = n19639 & ~n19651 ;
  assign n19653 = ~n19650 & ~n19651 ;
  assign n19654 = ~n19652 & ~n19653 ;
  assign n19655 = ~n18931 & ~n18937 ;
  assign n19656 = n19654 & n19655 ;
  assign n19657 = ~n19654 & ~n19655 ;
  assign n19658 = ~n19656 & ~n19657 ;
  assign n19659 = x106 & n1434 ;
  assign n19660 = x104 & n1646 ;
  assign n19661 = x105 & n1429 ;
  assign n19662 = ~n19660 & ~n19661 ;
  assign n19663 = ~n19659 & n19662 ;
  assign n19664 = n1437 & n12181 ;
  assign n19665 = n19663 & ~n19664 ;
  assign n19666 = x14 & ~n19665 ;
  assign n19667 = x14 & ~n19666 ;
  assign n19668 = ~n19665 & ~n19666 ;
  assign n19669 = ~n19667 & ~n19668 ;
  assign n19670 = ~n19658 & n19669 ;
  assign n19671 = n19658 & ~n19669 ;
  assign n19672 = ~n19670 & ~n19671 ;
  assign n19673 = ~n19413 & n19672 ;
  assign n19674 = n19413 & ~n19672 ;
  assign n19675 = ~n19673 & ~n19674 ;
  assign n19676 = ~n19412 & n19675 ;
  assign n19677 = ~n19412 & ~n19676 ;
  assign n19678 = n19675 & ~n19676 ;
  assign n19679 = ~n19677 & ~n19678 ;
  assign n19680 = ~n18974 & ~n19679 ;
  assign n19681 = ~n18974 & ~n19680 ;
  assign n19682 = ~n19679 & ~n19680 ;
  assign n19683 = ~n19681 & ~n19682 ;
  assign n19684 = x112 & n574 ;
  assign n19685 = x110 & n673 ;
  assign n19686 = x111 & n569 ;
  assign n19687 = ~n19685 & ~n19686 ;
  assign n19688 = ~n19684 & n19687 ;
  assign n19689 = n577 & n15442 ;
  assign n19690 = n19688 & ~n19689 ;
  assign n19691 = x8 & ~n19690 ;
  assign n19692 = x8 & ~n19691 ;
  assign n19693 = ~n19690 & ~n19691 ;
  assign n19694 = ~n19692 & ~n19693 ;
  assign n19695 = ~n19683 & ~n19694 ;
  assign n19696 = ~n19683 & ~n19695 ;
  assign n19697 = ~n19694 & ~n19695 ;
  assign n19698 = ~n19696 & ~n19697 ;
  assign n19699 = ~n18988 & ~n18994 ;
  assign n19700 = n19698 & n19699 ;
  assign n19701 = ~n19698 & ~n19699 ;
  assign n19702 = ~n19700 & ~n19701 ;
  assign n19703 = x115 & n293 ;
  assign n19704 = x113 & n373 ;
  assign n19705 = x114 & n288 ;
  assign n19706 = ~n19704 & ~n19705 ;
  assign n19707 = ~n19703 & n19706 ;
  assign n19708 = n296 & n17364 ;
  assign n19709 = n19707 & ~n19708 ;
  assign n19710 = x5 & ~n19709 ;
  assign n19711 = x5 & ~n19710 ;
  assign n19712 = ~n19709 & ~n19710 ;
  assign n19713 = ~n19711 & ~n19712 ;
  assign n19714 = ~n19702 & n19713 ;
  assign n19715 = n19702 & ~n19713 ;
  assign n19716 = ~n19714 & ~n19715 ;
  assign n19717 = ~n19012 & n19716 ;
  assign n19718 = n19012 & ~n19716 ;
  assign n19719 = ~n19717 & ~n19718 ;
  assign n19720 = ~n19401 & n19719 ;
  assign n19721 = n19401 & ~n19719 ;
  assign n19722 = ~n19720 & ~n19721 ;
  assign n19723 = ~n19383 & n19722 ;
  assign n19724 = n19383 & ~n19722 ;
  assign n19725 = ~n19723 & ~n19724 ;
  assign n20065 = n19725 & x182 ;
  assign n19726 = ~n19356 & ~n19371 ;
  assign n19727 = ~n19375 & ~n19726 ;
  assign n19728 = ~x118 & n164 ;
  assign n19729 = ~x116 & n205 ;
  assign n19730 = ~x117 & n162 ;
  assign n19731 = ~n19729 & ~n19730 ;
  assign n19732 = ~n19728 & n19731 ;
  assign n19733 = ~n19021 & ~n19363 ;
  assign n19734 = n19392 & ~n19733 ;
  assign n19735 = ~n19392 & n19733 ;
  assign n19736 = ~n19734 & ~n19735 ;
  assign n19737 = n167 & n19736 ;
  assign n19738 = n19732 & ~n19737 ;
  assign n19739 = ~x2 & ~n19738 ;
  assign n19740 = ~x2 & ~n19739 ;
  assign n19741 = ~n19738 & ~n19739 ;
  assign n19742 = ~n19740 & ~n19741 ;
  assign n19743 = ~x109 & n945 ;
  assign n19744 = ~x107 & n1099 ;
  assign n19745 = ~x108 & n940 ;
  assign n19746 = ~n19744 & ~n19745 ;
  assign n19747 = ~n19743 & n19746 ;
  assign n19748 = n948 & n14177 ;
  assign n19749 = n19747 & ~n19748 ;
  assign n19750 = ~x11 & ~n19749 ;
  assign n19751 = ~x11 & ~n19750 ;
  assign n19752 = ~n19749 & ~n19750 ;
  assign n19753 = ~n19751 & ~n19752 ;
  assign n19754 = ~n19292 & ~n19298 ;
  assign n19755 = ~n19254 & ~n19260 ;
  assign n19756 = ~n19238 & ~n19240 ;
  assign n19757 = ~n19232 & ~n19234 ;
  assign n19758 = ~x94 & n4531 ;
  assign n19759 = ~x92 & n4847 ;
  assign n19760 = ~x93 & n4526 ;
  assign n19761 = ~n19759 & ~n19760 ;
  assign n19762 = ~n19758 & n19761 ;
  assign n19763 = n4534 & n6671 ;
  assign n19764 = n19762 & ~n19763 ;
  assign n19765 = ~x26 & ~n19764 ;
  assign n19766 = ~x26 & ~n19765 ;
  assign n19767 = ~n19764 & ~n19765 ;
  assign n19768 = ~n19766 & ~n19767 ;
  assign n19769 = ~n19226 & ~n19228 ;
  assign n19770 = ~x91 & n5560 ;
  assign n19771 = ~x89 & n5943 ;
  assign n19772 = ~x90 & n5555 ;
  assign n19773 = ~n19771 & ~n19772 ;
  assign n19774 = ~n19770 & n19773 ;
  assign n19775 = n5507 & n5563 ;
  assign n19776 = n19774 & ~n19775 ;
  assign n19777 = ~x29 & ~n19776 ;
  assign n19778 = ~x29 & ~n19777 ;
  assign n19779 = ~n19776 & ~n19777 ;
  assign n19780 = ~n19778 & ~n19779 ;
  assign n19781 = ~n19206 & ~n19210 ;
  assign n19782 = ~x88 & n6725 ;
  assign n19783 = ~x86 & n7129 ;
  assign n19784 = ~x87 & n6720 ;
  assign n19785 = ~n19783 & ~n19784 ;
  assign n19786 = ~n19782 & n19785 ;
  assign n19787 = n4457 & n6728 ;
  assign n19788 = n19786 & ~n19787 ;
  assign n19789 = ~x32 & ~n19788 ;
  assign n19790 = ~x32 & ~n19789 ;
  assign n19791 = ~n19788 & ~n19789 ;
  assign n19792 = ~n19790 & ~n19791 ;
  assign n19793 = ~n19199 & ~n19203 ;
  assign n19794 = ~x85 & n8006 ;
  assign n19795 = ~x83 & n8474 ;
  assign n19796 = ~x84 & n8001 ;
  assign n19797 = ~n19795 & ~n19796 ;
  assign n19798 = ~n19794 & n19797 ;
  assign n19799 = n3521 & n8009 ;
  assign n19800 = n19798 & ~n19799 ;
  assign n19801 = ~x35 & ~n19800 ;
  assign n19802 = ~x35 & ~n19801 ;
  assign n19803 = ~n19800 & ~n19801 ;
  assign n19804 = ~n19802 & ~n19803 ;
  assign n19805 = ~n19180 & ~n19184 ;
  assign n19806 = ~x82 & n9433 ;
  assign n19807 = ~x80 & n9915 ;
  assign n19808 = ~x81 & n9428 ;
  assign n19809 = ~n19807 & ~n19808 ;
  assign n19810 = ~n19806 & n19809 ;
  assign n19811 = n2697 & n9436 ;
  assign n19812 = n19810 & ~n19811 ;
  assign n19813 = ~x38 & ~n19812 ;
  assign n19814 = ~x38 & ~n19813 ;
  assign n19815 = ~n19812 & ~n19813 ;
  assign n19816 = ~n19814 & ~n19815 ;
  assign n19817 = ~n19173 & ~n19177 ;
  assign n19818 = ~x79 & n10905 ;
  assign n19819 = ~x77 & n11466 ;
  assign n19820 = ~x78 & n10900 ;
  assign n19821 = ~n19819 & ~n19820 ;
  assign n19822 = ~n19818 & n19821 ;
  assign n19823 = n1921 & n10908 ;
  assign n19824 = n19822 & ~n19823 ;
  assign n19825 = ~x41 & ~n19824 ;
  assign n19826 = ~x41 & ~n19825 ;
  assign n19827 = ~n19824 & ~n19825 ;
  assign n19828 = ~n19826 & ~n19827 ;
  assign n19829 = ~n19157 & ~n19159 ;
  assign n19830 = ~x76 & n12506 ;
  assign n19831 = ~x74 & n13131 ;
  assign n19832 = ~x75 & n12501 ;
  assign n19833 = ~n19831 & ~n19832 ;
  assign n19834 = ~n19830 & n19833 ;
  assign n19835 = n1390 & n12509 ;
  assign n19836 = n19834 & ~n19835 ;
  assign n19837 = ~x44 & ~n19836 ;
  assign n19838 = ~x44 & ~n19837 ;
  assign n19839 = ~n19836 & ~n19837 ;
  assign n19840 = ~n19838 & ~n19839 ;
  assign n19841 = ~n19151 & ~n19153 ;
  assign n19842 = ~x73 & n14233 ;
  assign n19843 = ~x71 & n14876 ;
  assign n19844 = ~x72 & n14228 ;
  assign n19845 = ~n19843 & ~n19844 ;
  assign n19846 = ~n19842 & n19845 ;
  assign n19847 = n903 & n14236 ;
  assign n19848 = n19846 & ~n19847 ;
  assign n19849 = ~x47 & ~n19848 ;
  assign n19850 = ~x47 & ~n19849 ;
  assign n19851 = ~n19848 & ~n19849 ;
  assign n19852 = ~n19850 & ~n19851 ;
  assign n19853 = ~x64 & ~n19514 ;
  assign n19854 = ~n19118 & n19853 ;
  assign n19855 = n19118 & ~n19853 ;
  assign n19856 = ~n19854 & ~n19855 ;
  assign n19857 = ~x67 & n18025 ;
  assign n19858 = ~x65 & n18764 ;
  assign n19859 = ~x66 & n18020 ;
  assign n19860 = ~n19858 & ~n19859 ;
  assign n19861 = ~n19857 & n19860 ;
  assign n19862 = n266 & n18028 ;
  assign n19863 = n19861 & ~n19862 ;
  assign n19864 = ~x53 & ~n19863 ;
  assign n19865 = ~x53 & ~n19864 ;
  assign n19866 = ~n19863 & ~n19864 ;
  assign n19867 = ~n19865 & ~n19866 ;
  assign n19868 = ~n19856 & ~n19867 ;
  assign n19869 = n19856 & n19867 ;
  assign n19870 = ~n19868 & ~n19869 ;
  assign n19871 = ~x70 & n16076 ;
  assign n19872 = ~x68 & n16756 ;
  assign n19873 = ~x69 & n16071 ;
  assign n19874 = ~n19872 & ~n19873 ;
  assign n19875 = ~n19871 & n19874 ;
  assign n19876 = n529 & n16079 ;
  assign n19877 = n19875 & ~n19876 ;
  assign n19878 = ~x50 & ~n19877 ;
  assign n19879 = ~x50 & ~n19878 ;
  assign n19880 = ~n19877 & ~n19878 ;
  assign n19881 = ~n19879 & ~n19880 ;
  assign n19882 = n19870 & ~n19881 ;
  assign n19883 = n19870 & ~n19882 ;
  assign n19884 = ~n19881 & ~n19882 ;
  assign n19885 = ~n19883 & ~n19884 ;
  assign n19886 = ~n19136 & ~n19885 ;
  assign n19887 = n19136 & n19885 ;
  assign n19888 = ~n19886 & ~n19887 ;
  assign n19889 = ~n19852 & n19888 ;
  assign n19890 = ~n19852 & ~n19889 ;
  assign n19891 = n19888 & ~n19889 ;
  assign n19892 = ~n19890 & ~n19891 ;
  assign n19893 = ~n19841 & ~n19892 ;
  assign n19894 = n19841 & ~n19891 ;
  assign n19895 = ~n19890 & n19894 ;
  assign n19896 = ~n19893 & ~n19895 ;
  assign n19897 = ~n19840 & n19896 ;
  assign n19898 = ~n19840 & ~n19897 ;
  assign n19899 = n19896 & ~n19897 ;
  assign n19900 = ~n19898 & ~n19899 ;
  assign n19901 = ~n19829 & ~n19900 ;
  assign n19902 = n19829 & ~n19899 ;
  assign n19903 = ~n19898 & n19902 ;
  assign n19904 = ~n19901 & ~n19903 ;
  assign n19905 = ~n19828 & n19904 ;
  assign n19906 = n19828 & ~n19904 ;
  assign n19907 = ~n19905 & ~n19906 ;
  assign n19908 = ~n19817 & n19907 ;
  assign n19909 = n19817 & ~n19907 ;
  assign n19910 = ~n19908 & ~n19909 ;
  assign n19911 = ~n19816 & n19910 ;
  assign n19912 = ~n19816 & ~n19911 ;
  assign n19913 = n19910 & ~n19911 ;
  assign n19914 = ~n19912 & ~n19913 ;
  assign n19915 = ~n19805 & ~n19914 ;
  assign n19916 = n19805 & ~n19913 ;
  assign n19917 = ~n19912 & n19916 ;
  assign n19918 = ~n19915 & ~n19917 ;
  assign n19919 = ~n19804 & n19918 ;
  assign n19920 = n19804 & ~n19918 ;
  assign n19921 = ~n19919 & ~n19920 ;
  assign n19922 = ~n19793 & n19921 ;
  assign n19923 = n19793 & ~n19921 ;
  assign n19924 = ~n19922 & ~n19923 ;
  assign n19925 = ~n19792 & n19924 ;
  assign n19926 = n19792 & ~n19924 ;
  assign n19927 = ~n19925 & ~n19926 ;
  assign n19928 = ~n19781 & n19927 ;
  assign n19929 = n19781 & ~n19927 ;
  assign n19930 = ~n19928 & ~n19929 ;
  assign n19931 = ~n19780 & n19930 ;
  assign n19932 = n19780 & ~n19930 ;
  assign n19933 = ~n19931 & ~n19932 ;
  assign n19934 = ~n19769 & n19933 ;
  assign n19935 = n19769 & ~n19933 ;
  assign n19936 = ~n19934 & ~n19935 ;
  assign n19937 = ~n19768 & n19936 ;
  assign n19938 = n19768 & ~n19936 ;
  assign n19939 = ~n19937 & ~n19938 ;
  assign n19940 = ~n19757 & n19939 ;
  assign n19941 = n19757 & ~n19939 ;
  assign n19942 = ~n19940 & ~n19941 ;
  assign n19943 = ~x97 & n3589 ;
  assign n19944 = ~x95 & n3878 ;
  assign n19945 = ~x96 & n3584 ;
  assign n19946 = ~n19944 & ~n19945 ;
  assign n19947 = ~n19943 & n19946 ;
  assign n19948 = n3592 & n7949 ;
  assign n19949 = n19947 & ~n19948 ;
  assign n19950 = ~x23 & ~n19949 ;
  assign n19951 = ~x23 & ~n19950 ;
  assign n19952 = ~n19949 & ~n19950 ;
  assign n19953 = ~n19951 & ~n19952 ;
  assign n19954 = n19942 & ~n19953 ;
  assign n19955 = n19942 & ~n19954 ;
  assign n19956 = ~n19953 & ~n19954 ;
  assign n19957 = ~n19955 & ~n19956 ;
  assign n19958 = ~n19756 & n19957 ;
  assign n19959 = n19756 & ~n19957 ;
  assign n19960 = ~n19958 & ~n19959 ;
  assign n19961 = ~x100 & n2751 ;
  assign n19962 = ~x98 & n3020 ;
  assign n19963 = ~x99 & n2746 ;
  assign n19964 = ~n19962 & ~n19963 ;
  assign n19965 = ~n19961 & n19964 ;
  assign n19966 = n2754 & n9338 ;
  assign n19967 = n19965 & ~n19966 ;
  assign n19968 = ~x20 & ~n19967 ;
  assign n19969 = ~x20 & ~n19968 ;
  assign n19970 = ~n19967 & ~n19968 ;
  assign n19971 = ~n19969 & ~n19970 ;
  assign n19972 = ~n19960 & ~n19971 ;
  assign n19973 = n19960 & n19971 ;
  assign n19974 = ~n19972 & ~n19973 ;
  assign n19975 = n19755 & ~n19974 ;
  assign n19976 = ~n19755 & n19974 ;
  assign n19977 = ~n19975 & ~n19976 ;
  assign n19978 = ~x103 & n2093 ;
  assign n19979 = ~x101 & n2275 ;
  assign n19980 = ~x102 & n2088 ;
  assign n19981 = ~n19979 & ~n19980 ;
  assign n19982 = ~n19978 & n19981 ;
  assign n19983 = n2096 & n10833 ;
  assign n19984 = n19982 & ~n19983 ;
  assign n19985 = ~x17 & ~n19984 ;
  assign n19986 = ~x17 & ~n19985 ;
  assign n19987 = ~n19984 & ~n19985 ;
  assign n19988 = ~n19986 & ~n19987 ;
  assign n19989 = n19977 & ~n19988 ;
  assign n19990 = n19977 & ~n19989 ;
  assign n19991 = ~n19988 & ~n19989 ;
  assign n19992 = ~n19990 & ~n19991 ;
  assign n19993 = ~n19273 & ~n19279 ;
  assign n19994 = n19992 & n19993 ;
  assign n19995 = ~n19992 & ~n19993 ;
  assign n19996 = ~n19994 & ~n19995 ;
  assign n19997 = ~x106 & n1434 ;
  assign n19998 = ~x104 & n1646 ;
  assign n19999 = ~x105 & n1429 ;
  assign n20000 = ~n19998 & ~n19999 ;
  assign n20001 = ~n19997 & n20000 ;
  assign n20002 = n1437 & n12447 ;
  assign n20003 = n20001 & ~n20002 ;
  assign n20004 = ~x14 & ~n20003 ;
  assign n20005 = ~x14 & ~n20004 ;
  assign n20006 = ~n20003 & ~n20004 ;
  assign n20007 = ~n20005 & ~n20006 ;
  assign n20008 = ~n19996 & n20007 ;
  assign n20009 = n19996 & ~n20007 ;
  assign n20010 = ~n20008 & ~n20009 ;
  assign n20011 = ~n19754 & n20010 ;
  assign n20012 = n19754 & ~n20010 ;
  assign n20013 = ~n20011 & ~n20012 ;
  assign n20014 = ~n19753 & n20013 ;
  assign n20015 = ~n19753 & ~n20014 ;
  assign n20016 = n20013 & ~n20014 ;
  assign n20017 = ~n20015 & ~n20016 ;
  assign n20018 = ~n19316 & ~n20017 ;
  assign n20019 = ~n19316 & ~n20018 ;
  assign n20020 = ~n20017 & ~n20018 ;
  assign n20021 = ~n20019 & ~n20020 ;
  assign n20022 = ~x112 & n574 ;
  assign n20023 = ~x110 & n673 ;
  assign n20024 = ~x111 & n569 ;
  assign n20025 = ~n20023 & ~n20024 ;
  assign n20026 = ~n20022 & n20025 ;
  assign n20027 = n577 & n15744 ;
  assign n20028 = n20026 & ~n20027 ;
  assign n20029 = ~x8 & ~n20028 ;
  assign n20030 = ~x8 & ~n20029 ;
  assign n20031 = ~n20028 & ~n20029 ;
  assign n20032 = ~n20030 & ~n20031 ;
  assign n20033 = ~n20021 & ~n20032 ;
  assign n20034 = ~n20021 & ~n20033 ;
  assign n20035 = ~n20032 & ~n20033 ;
  assign n20036 = ~n20034 & ~n20035 ;
  assign n20037 = ~n19330 & ~n19336 ;
  assign n20038 = n20036 & n20037 ;
  assign n20039 = ~n20036 & ~n20037 ;
  assign n20040 = ~n20038 & ~n20039 ;
  assign n20041 = ~x115 & n293 ;
  assign n20042 = ~x113 & n373 ;
  assign n20043 = ~x114 & n288 ;
  assign n20044 = ~n20042 & ~n20043 ;
  assign n20045 = ~n20041 & n20044 ;
  assign n20046 = n296 & n17683 ;
  assign n20047 = n20045 & ~n20046 ;
  assign n20048 = ~x5 & ~n20047 ;
  assign n20049 = ~x5 & ~n20048 ;
  assign n20050 = ~n20047 & ~n20048 ;
  assign n20051 = ~n20049 & ~n20050 ;
  assign n20052 = ~n20040 & n20051 ;
  assign n20053 = n20040 & ~n20051 ;
  assign n20054 = ~n20052 & ~n20053 ;
  assign n20055 = ~n19354 & n20054 ;
  assign n20056 = n19354 & ~n20054 ;
  assign n20057 = ~n20055 & ~n20056 ;
  assign n20058 = ~n19742 & n20057 ;
  assign n20059 = n19742 & ~n20057 ;
  assign n20060 = ~n20058 & ~n20059 ;
  assign n20061 = ~n19727 & n20060 ;
  assign n20062 = n19727 & ~n20060 ;
  assign n20063 = ~n20061 & ~n20062 ;
  assign n20066 = ~n20063 & ~x182 ;
  assign n20067 = ~n20065 & ~n20066 ;
  assign n20068 = ~n19720 & ~n19723 ;
  assign n20069 = ~n19715 & ~n19717 ;
  assign n20070 = ~n19695 & ~n19701 ;
  assign n20071 = x113 & n574 ;
  assign n20072 = x111 & n673 ;
  assign n20073 = x112 & n569 ;
  assign n20074 = ~n20072 & ~n20073 ;
  assign n20075 = ~n20071 & n20074 ;
  assign n20076 = n577 & n16361 ;
  assign n20077 = n20075 & ~n20076 ;
  assign n20078 = x8 & ~n20077 ;
  assign n20079 = x8 & ~n20078 ;
  assign n20080 = ~n20077 & ~n20078 ;
  assign n20081 = ~n20079 & ~n20080 ;
  assign n20082 = ~n19676 & ~n19680 ;
  assign n20083 = ~n19671 & ~n19673 ;
  assign n20084 = ~n19573 & ~n19577 ;
  assign n20085 = ~n19559 & ~n19563 ;
  assign n20086 = x77 & n12506 ;
  assign n20087 = x75 & n13131 ;
  assign n20088 = x76 & n12501 ;
  assign n20089 = ~n20087 & ~n20088 ;
  assign n20090 = ~n20086 & n20089 ;
  assign n20091 = n1502 & n12509 ;
  assign n20092 = n20090 & ~n20091 ;
  assign n20093 = x44 & ~n20092 ;
  assign n20094 = x44 & ~n20093 ;
  assign n20095 = ~n20092 & ~n20093 ;
  assign n20096 = ~n20094 & ~n20095 ;
  assign n20097 = ~n19551 & ~n19555 ;
  assign n20098 = x74 & n14233 ;
  assign n20099 = x72 & n14876 ;
  assign n20100 = x73 & n14228 ;
  assign n20101 = ~n20099 & ~n20100 ;
  assign n20102 = ~n20098 & n20101 ;
  assign n20103 = n994 & n14236 ;
  assign n20104 = n20102 & ~n20103 ;
  assign n20105 = x47 & ~n20104 ;
  assign n20106 = x47 & ~n20105 ;
  assign n20107 = ~n20104 & ~n20105 ;
  assign n20108 = ~n20106 & ~n20107 ;
  assign n20109 = ~n19544 & ~n19548 ;
  assign n20110 = x71 & n16076 ;
  assign n20111 = x69 & n16756 ;
  assign n20112 = x70 & n16071 ;
  assign n20113 = ~n20111 & ~n20112 ;
  assign n20114 = ~n20110 & n20113 ;
  assign n20115 = n558 & n16079 ;
  assign n20116 = n20114 & ~n20115 ;
  assign n20117 = x50 & ~n20116 ;
  assign n20118 = x50 & ~n20117 ;
  assign n20119 = ~n20116 & ~n20117 ;
  assign n20120 = ~n20118 & ~n20119 ;
  assign n20121 = n18776 & n19515 ;
  assign n20122 = ~n19530 & ~n20121 ;
  assign n20123 = x68 & n18025 ;
  assign n20124 = x66 & n18764 ;
  assign n20125 = x67 & n18020 ;
  assign n20126 = ~n20124 & ~n20125 ;
  assign n20127 = ~n20123 & n20126 ;
  assign n20128 = n317 & n18028 ;
  assign n20129 = n20127 & ~n20128 ;
  assign n20130 = x53 & ~n20129 ;
  assign n20131 = x53 & ~n20130 ;
  assign n20132 = ~n20129 & ~n20130 ;
  assign n20133 = ~n20131 & ~n20132 ;
  assign n20134 = x56 & ~n19515 ;
  assign n20135 = ~x54 & x55 ;
  assign n20136 = x54 & ~x55 ;
  assign n20137 = ~n20135 & ~n20136 ;
  assign n20138 = n19514 & ~n20137 ;
  assign n20139 = x64 & n20138 ;
  assign n20140 = ~x55 & x56 ;
  assign n20141 = x55 & ~x56 ;
  assign n20142 = ~n20140 & ~n20141 ;
  assign n20143 = ~n19514 & n20142 ;
  assign n20144 = x65 & n20143 ;
  assign n20145 = ~n20139 & ~n20144 ;
  assign n20146 = ~n19514 & ~n20142 ;
  assign n20147 = ~n152 & n20146 ;
  assign n20148 = n20145 & ~n20147 ;
  assign n20149 = x56 & ~n20148 ;
  assign n20150 = x56 & ~n20149 ;
  assign n20151 = ~n20148 & ~n20149 ;
  assign n20152 = ~n20150 & ~n20151 ;
  assign n20153 = n20134 & ~n20152 ;
  assign n20154 = ~n20134 & n20152 ;
  assign n20155 = ~n20153 & ~n20154 ;
  assign n20156 = n20133 & ~n20155 ;
  assign n20157 = ~n20133 & n20155 ;
  assign n20158 = ~n20156 & ~n20157 ;
  assign n20159 = ~n20122 & n20158 ;
  assign n20160 = n20122 & ~n20158 ;
  assign n20161 = ~n20159 & ~n20160 ;
  assign n20162 = n20120 & ~n20161 ;
  assign n20163 = ~n20120 & n20161 ;
  assign n20164 = ~n20162 & ~n20163 ;
  assign n20165 = ~n20109 & n20164 ;
  assign n20166 = n20109 & ~n20164 ;
  assign n20167 = ~n20165 & ~n20166 ;
  assign n20168 = n20108 & ~n20167 ;
  assign n20169 = ~n20108 & n20167 ;
  assign n20170 = ~n20168 & ~n20169 ;
  assign n20171 = ~n20097 & n20170 ;
  assign n20172 = n20097 & ~n20170 ;
  assign n20173 = ~n20171 & ~n20172 ;
  assign n20174 = n20096 & ~n20173 ;
  assign n20175 = ~n20096 & n20173 ;
  assign n20176 = ~n20174 & ~n20175 ;
  assign n20177 = ~n20085 & n20176 ;
  assign n20178 = n20085 & ~n20176 ;
  assign n20179 = ~n20177 & ~n20178 ;
  assign n20180 = x80 & n10905 ;
  assign n20181 = x78 & n11466 ;
  assign n20182 = x79 & n10900 ;
  assign n20183 = ~n20181 & ~n20182 ;
  assign n20184 = ~n20180 & n20183 ;
  assign n20185 = n2028 & n10908 ;
  assign n20186 = n20184 & ~n20185 ;
  assign n20187 = x41 & ~n20186 ;
  assign n20188 = x41 & ~n20187 ;
  assign n20189 = ~n20186 & ~n20187 ;
  assign n20190 = ~n20188 & ~n20189 ;
  assign n20191 = n20179 & ~n20190 ;
  assign n20192 = n20179 & ~n20191 ;
  assign n20193 = ~n20190 & ~n20191 ;
  assign n20194 = ~n20192 & ~n20193 ;
  assign n20195 = ~n19567 & ~n19570 ;
  assign n20196 = n20194 & n20195 ;
  assign n20197 = ~n20194 & ~n20195 ;
  assign n20198 = ~n20196 & ~n20197 ;
  assign n20199 = x83 & n9433 ;
  assign n20200 = x81 & n9915 ;
  assign n20201 = x82 & n9428 ;
  assign n20202 = ~n20200 & ~n20201 ;
  assign n20203 = ~n20199 & n20202 ;
  assign n20204 = n2843 & n9436 ;
  assign n20205 = n20203 & ~n20204 ;
  assign n20206 = x38 & ~n20205 ;
  assign n20207 = x38 & ~n20206 ;
  assign n20208 = ~n20205 & ~n20206 ;
  assign n20209 = ~n20207 & ~n20208 ;
  assign n20210 = n20198 & ~n20209 ;
  assign n20211 = ~n20198 & n20209 ;
  assign n20212 = ~n20084 & ~n20211 ;
  assign n20213 = ~n20210 & n20212 ;
  assign n20214 = ~n20084 & ~n20213 ;
  assign n20215 = ~n20210 & ~n20213 ;
  assign n20216 = ~n20211 & n20215 ;
  assign n20217 = ~n20214 & ~n20216 ;
  assign n20218 = x86 & n8006 ;
  assign n20219 = x84 & n8474 ;
  assign n20220 = x85 & n8001 ;
  assign n20221 = ~n20219 & ~n20220 ;
  assign n20222 = ~n20218 & n20221 ;
  assign n20223 = n3686 & n8009 ;
  assign n20224 = n20222 & ~n20223 ;
  assign n20225 = x35 & ~n20224 ;
  assign n20226 = x35 & ~n20225 ;
  assign n20227 = ~n20224 & ~n20225 ;
  assign n20228 = ~n20226 & ~n20227 ;
  assign n20229 = ~n20217 & ~n20228 ;
  assign n20230 = ~n20217 & ~n20229 ;
  assign n20231 = ~n20228 & ~n20229 ;
  assign n20232 = ~n20230 & ~n20231 ;
  assign n20233 = ~n19581 & ~n19584 ;
  assign n20234 = n20232 & n20233 ;
  assign n20235 = ~n20232 & ~n20233 ;
  assign n20236 = ~n20234 & ~n20235 ;
  assign n20237 = x89 & n6725 ;
  assign n20238 = x87 & n7129 ;
  assign n20239 = x88 & n6720 ;
  assign n20240 = ~n20238 & ~n20239 ;
  assign n20241 = ~n20237 & n20240 ;
  assign n20242 = n4488 & n6728 ;
  assign n20243 = n20241 & ~n20242 ;
  assign n20244 = x32 & ~n20243 ;
  assign n20245 = x32 & ~n20244 ;
  assign n20246 = ~n20243 & ~n20244 ;
  assign n20247 = ~n20245 & ~n20246 ;
  assign n20248 = n20236 & ~n20247 ;
  assign n20249 = n20236 & ~n20248 ;
  assign n20250 = ~n20247 & ~n20248 ;
  assign n20251 = ~n20249 & ~n20250 ;
  assign n20252 = ~n19587 & ~n19590 ;
  assign n20253 = n20251 & n20252 ;
  assign n20254 = ~n20251 & ~n20252 ;
  assign n20255 = ~n20253 & ~n20254 ;
  assign n20256 = x92 & n5560 ;
  assign n20257 = x90 & n5943 ;
  assign n20258 = x91 & n5555 ;
  assign n20259 = ~n20257 & ~n20258 ;
  assign n20260 = ~n20256 & n20259 ;
  assign n20261 = n5563 & n5710 ;
  assign n20262 = n20260 & ~n20261 ;
  assign n20263 = x29 & ~n20262 ;
  assign n20264 = x29 & ~n20263 ;
  assign n20265 = ~n20262 & ~n20263 ;
  assign n20266 = ~n20264 & ~n20265 ;
  assign n20267 = n20255 & ~n20266 ;
  assign n20268 = n20255 & ~n20267 ;
  assign n20269 = ~n20266 & ~n20267 ;
  assign n20270 = ~n20268 & ~n20269 ;
  assign n20271 = ~n19593 & ~n19596 ;
  assign n20272 = n20270 & n20271 ;
  assign n20273 = ~n20270 & ~n20271 ;
  assign n20274 = ~n20272 & ~n20273 ;
  assign n20275 = x95 & n4531 ;
  assign n20276 = x93 & n4847 ;
  assign n20277 = x94 & n4526 ;
  assign n20278 = ~n20276 & ~n20277 ;
  assign n20279 = ~n20275 & n20278 ;
  assign n20280 = n4534 & n6894 ;
  assign n20281 = n20279 & ~n20280 ;
  assign n20282 = x26 & ~n20281 ;
  assign n20283 = x26 & ~n20282 ;
  assign n20284 = ~n20281 & ~n20282 ;
  assign n20285 = ~n20283 & ~n20284 ;
  assign n20286 = n20274 & ~n20285 ;
  assign n20287 = n20274 & ~n20286 ;
  assign n20288 = ~n20285 & ~n20286 ;
  assign n20289 = ~n20287 & ~n20288 ;
  assign n20290 = ~n19599 & ~n19602 ;
  assign n20291 = n20289 & n20290 ;
  assign n20292 = ~n20289 & ~n20290 ;
  assign n20293 = ~n20291 & ~n20292 ;
  assign n20294 = x98 & n3589 ;
  assign n20295 = x96 & n3878 ;
  assign n20296 = x97 & n3584 ;
  assign n20297 = ~n20295 & ~n20296 ;
  assign n20298 = ~n20294 & n20297 ;
  assign n20299 = n3592 & n8196 ;
  assign n20300 = n20298 & ~n20299 ;
  assign n20301 = x23 & ~n20300 ;
  assign n20302 = x23 & ~n20301 ;
  assign n20303 = ~n20300 & ~n20301 ;
  assign n20304 = ~n20302 & ~n20303 ;
  assign n20305 = n20293 & ~n20304 ;
  assign n20306 = n20293 & ~n20305 ;
  assign n20307 = ~n20304 & ~n20305 ;
  assign n20308 = ~n20306 & ~n20307 ;
  assign n20309 = ~n19415 & ~n19619 ;
  assign n20310 = ~n19616 & ~n20309 ;
  assign n20311 = n20308 & n20310 ;
  assign n20312 = ~n20308 & ~n20310 ;
  assign n20313 = ~n20311 & ~n20312 ;
  assign n20314 = x101 & n2751 ;
  assign n20315 = x99 & n3020 ;
  assign n20316 = x100 & n2746 ;
  assign n20317 = ~n20315 & ~n20316 ;
  assign n20318 = ~n20314 & n20317 ;
  assign n20319 = n2754 & n9601 ;
  assign n20320 = n20318 & ~n20319 ;
  assign n20321 = x20 & ~n20320 ;
  assign n20322 = x20 & ~n20321 ;
  assign n20323 = ~n20320 & ~n20321 ;
  assign n20324 = ~n20322 & ~n20323 ;
  assign n20325 = n20313 & ~n20324 ;
  assign n20326 = n20313 & ~n20325 ;
  assign n20327 = ~n20324 & ~n20325 ;
  assign n20328 = ~n20326 & ~n20327 ;
  assign n20329 = ~n19634 & ~n19638 ;
  assign n20330 = n20328 & n20329 ;
  assign n20331 = ~n20328 & ~n20329 ;
  assign n20332 = ~n20330 & ~n20331 ;
  assign n20333 = x104 & n2093 ;
  assign n20334 = x102 & n2275 ;
  assign n20335 = x103 & n2088 ;
  assign n20336 = ~n20334 & ~n20335 ;
  assign n20337 = ~n20333 & n20336 ;
  assign n20338 = n2096 & n11116 ;
  assign n20339 = n20337 & ~n20338 ;
  assign n20340 = x17 & ~n20339 ;
  assign n20341 = x17 & ~n20340 ;
  assign n20342 = ~n20339 & ~n20340 ;
  assign n20343 = ~n20341 & ~n20342 ;
  assign n20344 = n20332 & ~n20343 ;
  assign n20345 = n20332 & ~n20344 ;
  assign n20346 = ~n20343 & ~n20344 ;
  assign n20347 = ~n20345 & ~n20346 ;
  assign n20348 = ~n19651 & ~n19657 ;
  assign n20349 = n20347 & n20348 ;
  assign n20350 = ~n20347 & ~n20348 ;
  assign n20351 = ~n20349 & ~n20350 ;
  assign n20352 = x107 & n1434 ;
  assign n20353 = x105 & n1646 ;
  assign n20354 = x106 & n1429 ;
  assign n20355 = ~n20353 & ~n20354 ;
  assign n20356 = ~n20352 & n20355 ;
  assign n20357 = n1437 & n12749 ;
  assign n20358 = n20356 & ~n20357 ;
  assign n20359 = x14 & ~n20358 ;
  assign n20360 = x14 & ~n20359 ;
  assign n20361 = ~n20358 & ~n20359 ;
  assign n20362 = ~n20360 & ~n20361 ;
  assign n20363 = n20351 & ~n20362 ;
  assign n20364 = ~n20351 & n20362 ;
  assign n20365 = ~n20083 & ~n20364 ;
  assign n20366 = ~n20363 & n20365 ;
  assign n20367 = ~n20083 & ~n20366 ;
  assign n20368 = ~n20363 & ~n20366 ;
  assign n20369 = ~n20364 & n20368 ;
  assign n20370 = ~n20367 & ~n20369 ;
  assign n20371 = x110 & n945 ;
  assign n20372 = x108 & n1099 ;
  assign n20373 = x109 & n940 ;
  assign n20374 = ~n20372 & ~n20373 ;
  assign n20375 = ~n20371 & n20374 ;
  assign n20376 = n948 & n14497 ;
  assign n20377 = n20375 & ~n20376 ;
  assign n20378 = x11 & ~n20377 ;
  assign n20379 = x11 & ~n20378 ;
  assign n20380 = ~n20377 & ~n20378 ;
  assign n20381 = ~n20379 & ~n20380 ;
  assign n20382 = n20370 & n20381 ;
  assign n20383 = ~n20370 & ~n20381 ;
  assign n20384 = ~n20382 & ~n20383 ;
  assign n20385 = ~n20082 & n20384 ;
  assign n20386 = n20082 & ~n20384 ;
  assign n20387 = ~n20385 & ~n20386 ;
  assign n20388 = n20081 & ~n20387 ;
  assign n20389 = ~n20081 & n20387 ;
  assign n20390 = ~n20388 & ~n20389 ;
  assign n20391 = ~n20070 & n20390 ;
  assign n20392 = n20070 & ~n20390 ;
  assign n20393 = ~n20391 & ~n20392 ;
  assign n20394 = x116 & n293 ;
  assign n20395 = x114 & n373 ;
  assign n20396 = x115 & n288 ;
  assign n20397 = ~n20395 & ~n20396 ;
  assign n20398 = ~n20394 & n20397 ;
  assign n20399 = n296 & n18336 ;
  assign n20400 = n20398 & ~n20399 ;
  assign n20401 = x5 & ~n20400 ;
  assign n20402 = x5 & ~n20401 ;
  assign n20403 = ~n20400 & ~n20401 ;
  assign n20404 = ~n20402 & ~n20403 ;
  assign n20405 = n20393 & ~n20404 ;
  assign n20406 = n20393 & ~n20405 ;
  assign n20407 = ~n20404 & ~n20405 ;
  assign n20408 = ~n20406 & ~n20407 ;
  assign n20409 = ~n20069 & n20408 ;
  assign n20410 = n20069 & ~n20408 ;
  assign n20411 = ~n20409 & ~n20410 ;
  assign n20412 = x119 & n146 ;
  assign n20413 = x117 & n182 ;
  assign n20414 = x118 & n141 ;
  assign n20415 = ~n20413 & ~n20414 ;
  assign n20416 = ~n20412 & n20415 ;
  assign n20417 = ~n19391 & ~n19393 ;
  assign n20418 = ~x118 & ~x119 ;
  assign n20419 = x118 & x119 ;
  assign n20420 = ~n20418 & ~n20419 ;
  assign n20421 = ~n20417 & n20420 ;
  assign n20422 = n20417 & ~n20420 ;
  assign n20423 = ~n20421 & ~n20422 ;
  assign n20424 = n149 & n20423 ;
  assign n20425 = n20416 & ~n20424 ;
  assign n20426 = x2 & ~n20425 ;
  assign n20427 = x2 & ~n20426 ;
  assign n20428 = ~n20425 & ~n20426 ;
  assign n20429 = ~n20427 & ~n20428 ;
  assign n20430 = ~n20411 & ~n20429 ;
  assign n20431 = n20411 & n20429 ;
  assign n20432 = ~n20430 & ~n20431 ;
  assign n20433 = ~n20068 & n20432 ;
  assign n20434 = n20068 & ~n20432 ;
  assign n20435 = ~n20433 & ~n20434 ;
  assign n20792 = n20435 & x183 ;
  assign n20436 = ~n20058 & ~n20061 ;
  assign n20437 = ~n20053 & ~n20055 ;
  assign n20438 = ~n20033 & ~n20039 ;
  assign n20439 = ~x113 & n574 ;
  assign n20440 = ~x111 & n673 ;
  assign n20441 = ~x112 & n569 ;
  assign n20442 = ~n20440 & ~n20441 ;
  assign n20443 = ~n20439 & n20442 ;
  assign n20444 = n577 & n16684 ;
  assign n20445 = n20443 & ~n20444 ;
  assign n20446 = ~x8 & ~n20445 ;
  assign n20447 = ~x8 & ~n20446 ;
  assign n20448 = ~n20445 & ~n20446 ;
  assign n20449 = ~n20447 & ~n20448 ;
  assign n20450 = ~n20014 & ~n20018 ;
  assign n20451 = ~n20009 & ~n20011 ;
  assign n20452 = ~n19911 & ~n19915 ;
  assign n20453 = ~n19897 & ~n19901 ;
  assign n20454 = ~x77 & n12506 ;
  assign n20455 = ~x75 & n13131 ;
  assign n20456 = ~x76 & n12501 ;
  assign n20457 = ~n20455 & ~n20456 ;
  assign n20458 = ~n20454 & n20457 ;
  assign n20459 = n1594 & n12509 ;
  assign n20460 = n20458 & ~n20459 ;
  assign n20461 = ~x44 & ~n20460 ;
  assign n20462 = ~x44 & ~n20461 ;
  assign n20463 = ~n20460 & ~n20461 ;
  assign n20464 = ~n20462 & ~n20463 ;
  assign n20465 = ~n19889 & ~n19893 ;
  assign n20466 = ~x74 & n14233 ;
  assign n20467 = ~x72 & n14876 ;
  assign n20468 = ~x73 & n14228 ;
  assign n20469 = ~n20467 & ~n20468 ;
  assign n20470 = ~n20466 & n20469 ;
  assign n20471 = n1066 & n14236 ;
  assign n20472 = n20470 & ~n20471 ;
  assign n20473 = ~x47 & ~n20472 ;
  assign n20474 = ~x47 & ~n20473 ;
  assign n20475 = ~n20472 & ~n20473 ;
  assign n20476 = ~n20474 & ~n20475 ;
  assign n20477 = ~n19882 & ~n19886 ;
  assign n20478 = ~x71 & n16076 ;
  assign n20479 = ~x69 & n16756 ;
  assign n20480 = ~x70 & n16071 ;
  assign n20481 = ~n20479 & ~n20480 ;
  assign n20482 = ~n20478 & n20481 ;
  assign n20483 = n622 & n16079 ;
  assign n20484 = n20482 & ~n20483 ;
  assign n20485 = ~x50 & ~n20484 ;
  assign n20486 = ~x50 & ~n20485 ;
  assign n20487 = ~n20484 & ~n20485 ;
  assign n20488 = ~n20486 & ~n20487 ;
  assign n20489 = n19118 & n19853 ;
  assign n20490 = ~n19868 & ~n20489 ;
  assign n20491 = ~x68 & n18025 ;
  assign n20492 = ~x66 & n18764 ;
  assign n20493 = ~x67 & n18020 ;
  assign n20494 = ~n20492 & ~n20493 ;
  assign n20495 = ~n20491 & n20494 ;
  assign n20496 = n352 & n18028 ;
  assign n20497 = n20495 & ~n20496 ;
  assign n20498 = ~x53 & ~n20497 ;
  assign n20499 = ~x53 & ~n20498 ;
  assign n20500 = ~n20497 & ~n20498 ;
  assign n20501 = ~n20499 & ~n20500 ;
  assign n20502 = ~x56 & ~n19853 ;
  assign n20503 = ~x64 & n20138 ;
  assign n20504 = ~x65 & n20143 ;
  assign n20505 = ~n20503 & ~n20504 ;
  assign n20506 = ~n20147 & n20505 ;
  assign n20507 = ~x56 & ~n20506 ;
  assign n20508 = ~x56 & ~n20507 ;
  assign n20509 = ~n20506 & ~n20507 ;
  assign n20510 = ~n20508 & ~n20509 ;
  assign n20511 = n20502 & ~n20510 ;
  assign n20512 = ~n20502 & n20510 ;
  assign n20513 = ~n20511 & ~n20512 ;
  assign n20514 = n20501 & ~n20513 ;
  assign n20515 = ~n20501 & n20513 ;
  assign n20516 = ~n20514 & ~n20515 ;
  assign n20517 = ~n20490 & n20516 ;
  assign n20518 = n20490 & ~n20516 ;
  assign n20519 = ~n20517 & ~n20518 ;
  assign n20520 = n20488 & ~n20519 ;
  assign n20521 = ~n20488 & n20519 ;
  assign n20522 = ~n20520 & ~n20521 ;
  assign n20523 = ~n20477 & n20522 ;
  assign n20524 = n20477 & ~n20522 ;
  assign n20525 = ~n20523 & ~n20524 ;
  assign n20526 = n20476 & ~n20525 ;
  assign n20527 = ~n20476 & n20525 ;
  assign n20528 = ~n20526 & ~n20527 ;
  assign n20529 = ~n20465 & n20528 ;
  assign n20530 = n20465 & ~n20528 ;
  assign n20531 = ~n20529 & ~n20530 ;
  assign n20532 = n20464 & ~n20531 ;
  assign n20533 = ~n20464 & n20531 ;
  assign n20534 = ~n20532 & ~n20533 ;
  assign n20535 = ~n20453 & n20534 ;
  assign n20536 = n20453 & ~n20534 ;
  assign n20537 = ~n20535 & ~n20536 ;
  assign n20538 = ~x80 & n10905 ;
  assign n20539 = ~x78 & n11466 ;
  assign n20540 = ~x79 & n10900 ;
  assign n20541 = ~n20539 & ~n20540 ;
  assign n20542 = ~n20538 & n20541 ;
  assign n20543 = n2145 & n10908 ;
  assign n20544 = n20542 & ~n20543 ;
  assign n20545 = ~x41 & ~n20544 ;
  assign n20546 = ~x41 & ~n20545 ;
  assign n20547 = ~n20544 & ~n20545 ;
  assign n20548 = ~n20546 & ~n20547 ;
  assign n20549 = n20537 & ~n20548 ;
  assign n20550 = n20537 & ~n20549 ;
  assign n20551 = ~n20548 & ~n20549 ;
  assign n20552 = ~n20550 & ~n20551 ;
  assign n20553 = ~n19905 & ~n19908 ;
  assign n20554 = n20552 & n20553 ;
  assign n20555 = ~n20552 & ~n20553 ;
  assign n20556 = ~n20554 & ~n20555 ;
  assign n20557 = ~x83 & n9433 ;
  assign n20558 = ~x81 & n9915 ;
  assign n20559 = ~x82 & n9428 ;
  assign n20560 = ~n20558 & ~n20559 ;
  assign n20561 = ~n20557 & n20560 ;
  assign n20562 = n2972 & n9436 ;
  assign n20563 = n20561 & ~n20562 ;
  assign n20564 = ~x38 & ~n20563 ;
  assign n20565 = ~x38 & ~n20564 ;
  assign n20566 = ~n20563 & ~n20564 ;
  assign n20567 = ~n20565 & ~n20566 ;
  assign n20568 = n20556 & ~n20567 ;
  assign n20569 = ~n20556 & n20567 ;
  assign n20570 = ~n20452 & ~n20569 ;
  assign n20571 = ~n20568 & n20570 ;
  assign n20572 = ~n20452 & ~n20571 ;
  assign n20573 = ~n20568 & ~n20571 ;
  assign n20574 = ~n20569 & n20573 ;
  assign n20575 = ~n20572 & ~n20574 ;
  assign n20576 = ~x86 & n8006 ;
  assign n20577 = ~x84 & n8474 ;
  assign n20578 = ~x85 & n8001 ;
  assign n20579 = ~n20577 & ~n20578 ;
  assign n20580 = ~n20576 & n20579 ;
  assign n20581 = n3832 & n8009 ;
  assign n20582 = n20580 & ~n20581 ;
  assign n20583 = ~x35 & ~n20582 ;
  assign n20584 = ~x35 & ~n20583 ;
  assign n20585 = ~n20582 & ~n20583 ;
  assign n20586 = ~n20584 & ~n20585 ;
  assign n20587 = ~n20575 & ~n20586 ;
  assign n20588 = ~n20575 & ~n20587 ;
  assign n20589 = ~n20586 & ~n20587 ;
  assign n20590 = ~n20588 & ~n20589 ;
  assign n20591 = ~n19919 & ~n19922 ;
  assign n20592 = n20590 & n20591 ;
  assign n20593 = ~n20590 & ~n20591 ;
  assign n20594 = ~n20592 & ~n20593 ;
  assign n20595 = ~x89 & n6725 ;
  assign n20596 = ~x87 & n7129 ;
  assign n20597 = ~x88 & n6720 ;
  assign n20598 = ~n20596 & ~n20597 ;
  assign n20599 = ~n20595 & n20598 ;
  assign n20600 = n4664 & n6728 ;
  assign n20601 = n20599 & ~n20600 ;
  assign n20602 = ~x32 & ~n20601 ;
  assign n20603 = ~x32 & ~n20602 ;
  assign n20604 = ~n20601 & ~n20602 ;
  assign n20605 = ~n20603 & ~n20604 ;
  assign n20606 = n20594 & ~n20605 ;
  assign n20607 = n20594 & ~n20606 ;
  assign n20608 = ~n20605 & ~n20606 ;
  assign n20609 = ~n20607 & ~n20608 ;
  assign n20610 = ~n19925 & ~n19928 ;
  assign n20611 = n20609 & n20610 ;
  assign n20612 = ~n20609 & ~n20610 ;
  assign n20613 = ~n20611 & ~n20612 ;
  assign n20614 = ~x92 & n5560 ;
  assign n20615 = ~x90 & n5943 ;
  assign n20616 = ~x91 & n5555 ;
  assign n20617 = ~n20615 & ~n20616 ;
  assign n20618 = ~n20614 & n20617 ;
  assign n20619 = n5563 & n5896 ;
  assign n20620 = n20618 & ~n20619 ;
  assign n20621 = ~x29 & ~n20620 ;
  assign n20622 = ~x29 & ~n20621 ;
  assign n20623 = ~n20620 & ~n20621 ;
  assign n20624 = ~n20622 & ~n20623 ;
  assign n20625 = n20613 & ~n20624 ;
  assign n20626 = n20613 & ~n20625 ;
  assign n20627 = ~n20624 & ~n20625 ;
  assign n20628 = ~n20626 & ~n20627 ;
  assign n20629 = ~n19931 & ~n19934 ;
  assign n20630 = n20628 & n20629 ;
  assign n20631 = ~n20628 & ~n20629 ;
  assign n20632 = ~n20630 & ~n20631 ;
  assign n20633 = ~x95 & n4531 ;
  assign n20634 = ~x93 & n4847 ;
  assign n20635 = ~x94 & n4526 ;
  assign n20636 = ~n20634 & ~n20635 ;
  assign n20637 = ~n20633 & n20636 ;
  assign n20638 = n4534 & n7100 ;
  assign n20639 = n20637 & ~n20638 ;
  assign n20640 = ~x26 & ~n20639 ;
  assign n20641 = ~x26 & ~n20640 ;
  assign n20642 = ~n20639 & ~n20640 ;
  assign n20643 = ~n20641 & ~n20642 ;
  assign n20644 = n20632 & ~n20643 ;
  assign n20645 = n20632 & ~n20644 ;
  assign n20646 = ~n20643 & ~n20644 ;
  assign n20647 = ~n20645 & ~n20646 ;
  assign n20648 = ~n19937 & ~n19940 ;
  assign n20649 = n20647 & n20648 ;
  assign n20650 = ~n20647 & ~n20648 ;
  assign n20651 = ~n20649 & ~n20650 ;
  assign n20652 = ~x98 & n3589 ;
  assign n20653 = ~x96 & n3878 ;
  assign n20654 = ~x97 & n3584 ;
  assign n20655 = ~n20653 & ~n20654 ;
  assign n20656 = ~n20652 & n20655 ;
  assign n20657 = n3592 & n8426 ;
  assign n20658 = n20656 & ~n20657 ;
  assign n20659 = ~x23 & ~n20658 ;
  assign n20660 = ~x23 & ~n20659 ;
  assign n20661 = ~n20658 & ~n20659 ;
  assign n20662 = ~n20660 & ~n20661 ;
  assign n20663 = n20651 & ~n20662 ;
  assign n20664 = n20651 & ~n20663 ;
  assign n20665 = ~n20662 & ~n20663 ;
  assign n20666 = ~n20664 & ~n20665 ;
  assign n20667 = ~n19756 & ~n19957 ;
  assign n20668 = ~n19954 & ~n20667 ;
  assign n20669 = n20666 & n20668 ;
  assign n20670 = ~n20666 & ~n20668 ;
  assign n20671 = ~n20669 & ~n20670 ;
  assign n20672 = ~x101 & n2751 ;
  assign n20673 = ~x99 & n3020 ;
  assign n20674 = ~x100 & n2746 ;
  assign n20675 = ~n20673 & ~n20674 ;
  assign n20676 = ~n20672 & n20675 ;
  assign n20677 = n2754 & n9844 ;
  assign n20678 = n20676 & ~n20677 ;
  assign n20679 = ~x20 & ~n20678 ;
  assign n20680 = ~x20 & ~n20679 ;
  assign n20681 = ~n20678 & ~n20679 ;
  assign n20682 = ~n20680 & ~n20681 ;
  assign n20683 = n20671 & ~n20682 ;
  assign n20684 = n20671 & ~n20683 ;
  assign n20685 = ~n20682 & ~n20683 ;
  assign n20686 = ~n20684 & ~n20685 ;
  assign n20687 = ~n19972 & ~n19976 ;
  assign n20688 = n20686 & n20687 ;
  assign n20689 = ~n20686 & ~n20687 ;
  assign n20690 = ~n20688 & ~n20689 ;
  assign n20691 = ~x104 & n2093 ;
  assign n20692 = ~x102 & n2275 ;
  assign n20693 = ~x103 & n2088 ;
  assign n20694 = ~n20692 & ~n20693 ;
  assign n20695 = ~n20691 & n20694 ;
  assign n20696 = n2096 & n11380 ;
  assign n20697 = n20695 & ~n20696 ;
  assign n20698 = ~x17 & ~n20697 ;
  assign n20699 = ~x17 & ~n20698 ;
  assign n20700 = ~n20697 & ~n20698 ;
  assign n20701 = ~n20699 & ~n20700 ;
  assign n20702 = n20690 & ~n20701 ;
  assign n20703 = n20690 & ~n20702 ;
  assign n20704 = ~n20701 & ~n20702 ;
  assign n20705 = ~n20703 & ~n20704 ;
  assign n20706 = ~n19989 & ~n19995 ;
  assign n20707 = n20705 & n20706 ;
  assign n20708 = ~n20705 & ~n20706 ;
  assign n20709 = ~n20707 & ~n20708 ;
  assign n20710 = ~x107 & n1434 ;
  assign n20711 = ~x105 & n1646 ;
  assign n20712 = ~x106 & n1429 ;
  assign n20713 = ~n20711 & ~n20712 ;
  assign n20714 = ~n20710 & n20713 ;
  assign n20715 = n1437 & n13034 ;
  assign n20716 = n20714 & ~n20715 ;
  assign n20717 = ~x14 & ~n20716 ;
  assign n20718 = ~x14 & ~n20717 ;
  assign n20719 = ~n20716 & ~n20717 ;
  assign n20720 = ~n20718 & ~n20719 ;
  assign n20721 = n20709 & ~n20720 ;
  assign n20722 = ~n20709 & n20720 ;
  assign n20723 = ~n20451 & ~n20722 ;
  assign n20724 = ~n20721 & n20723 ;
  assign n20725 = ~n20451 & ~n20724 ;
  assign n20726 = ~n20721 & ~n20724 ;
  assign n20727 = ~n20722 & n20726 ;
  assign n20728 = ~n20725 & ~n20727 ;
  assign n20729 = ~x110 & n945 ;
  assign n20730 = ~x108 & n1099 ;
  assign n20731 = ~x109 & n940 ;
  assign n20732 = ~n20730 & ~n20731 ;
  assign n20733 = ~n20729 & n20732 ;
  assign n20734 = n948 & n14802 ;
  assign n20735 = n20733 & ~n20734 ;
  assign n20736 = ~x11 & ~n20735 ;
  assign n20737 = ~x11 & ~n20736 ;
  assign n20738 = ~n20735 & ~n20736 ;
  assign n20739 = ~n20737 & ~n20738 ;
  assign n20740 = n20728 & n20739 ;
  assign n20741 = ~n20728 & ~n20739 ;
  assign n20742 = ~n20740 & ~n20741 ;
  assign n20743 = ~n20450 & n20742 ;
  assign n20744 = n20450 & ~n20742 ;
  assign n20745 = ~n20743 & ~n20744 ;
  assign n20746 = n20449 & ~n20745 ;
  assign n20747 = ~n20449 & n20745 ;
  assign n20748 = ~n20746 & ~n20747 ;
  assign n20749 = ~n20438 & n20748 ;
  assign n20750 = n20438 & ~n20748 ;
  assign n20751 = ~n20749 & ~n20750 ;
  assign n20752 = ~x116 & n293 ;
  assign n20753 = ~x114 & n373 ;
  assign n20754 = ~x115 & n288 ;
  assign n20755 = ~n20753 & ~n20754 ;
  assign n20756 = ~n20752 & n20755 ;
  assign n20757 = n296 & n18678 ;
  assign n20758 = n20756 & ~n20757 ;
  assign n20759 = ~x5 & ~n20758 ;
  assign n20760 = ~x5 & ~n20759 ;
  assign n20761 = ~n20758 & ~n20759 ;
  assign n20762 = ~n20760 & ~n20761 ;
  assign n20763 = n20751 & ~n20762 ;
  assign n20764 = n20751 & ~n20763 ;
  assign n20765 = ~n20762 & ~n20763 ;
  assign n20766 = ~n20764 & ~n20765 ;
  assign n20767 = ~n20437 & n20766 ;
  assign n20768 = n20437 & ~n20766 ;
  assign n20769 = ~n20767 & ~n20768 ;
  assign n20770 = ~x119 & n164 ;
  assign n20771 = ~x117 & n205 ;
  assign n20772 = ~x118 & n162 ;
  assign n20773 = ~n20771 & ~n20772 ;
  assign n20774 = ~n20770 & n20773 ;
  assign n20775 = ~n19390 & ~n19734 ;
  assign n20776 = n20420 & ~n20775 ;
  assign n20777 = ~n20420 & n20775 ;
  assign n20778 = ~n20776 & ~n20777 ;
  assign n20779 = n167 & n20778 ;
  assign n20780 = n20774 & ~n20779 ;
  assign n20781 = ~x2 & ~n20780 ;
  assign n20782 = ~x2 & ~n20781 ;
  assign n20783 = ~n20780 & ~n20781 ;
  assign n20784 = ~n20782 & ~n20783 ;
  assign n20785 = ~n20769 & ~n20784 ;
  assign n20786 = n20769 & n20784 ;
  assign n20787 = ~n20785 & ~n20786 ;
  assign n20788 = ~n20436 & n20787 ;
  assign n20789 = n20436 & ~n20787 ;
  assign n20790 = ~n20788 & ~n20789 ;
  assign n20793 = ~n20790 & ~x183 ;
  assign n20794 = ~n20792 & ~n20793 ;
  assign n20795 = ~n20069 & ~n20408 ;
  assign n20796 = ~n20405 & ~n20795 ;
  assign n20797 = ~n20389 & ~n20391 ;
  assign n20798 = x114 & n574 ;
  assign n20799 = x112 & n673 ;
  assign n20800 = x113 & n569 ;
  assign n20801 = ~n20799 & ~n20800 ;
  assign n20802 = ~n20798 & n20801 ;
  assign n20803 = n577 & n17012 ;
  assign n20804 = n20802 & ~n20803 ;
  assign n20805 = x8 & ~n20804 ;
  assign n20806 = x8 & ~n20805 ;
  assign n20807 = ~n20804 & ~n20805 ;
  assign n20808 = ~n20806 & ~n20807 ;
  assign n20809 = ~n20383 & ~n20385 ;
  assign n20810 = ~n20286 & ~n20292 ;
  assign n20811 = x96 & n4531 ;
  assign n20812 = x94 & n4847 ;
  assign n20813 = x95 & n4526 ;
  assign n20814 = ~n20812 & ~n20813 ;
  assign n20815 = ~n20811 & n20814 ;
  assign n20816 = n4534 & n7321 ;
  assign n20817 = n20815 & ~n20816 ;
  assign n20818 = x26 & ~n20817 ;
  assign n20819 = x26 & ~n20818 ;
  assign n20820 = ~n20817 & ~n20818 ;
  assign n20821 = ~n20819 & ~n20820 ;
  assign n20822 = ~n20267 & ~n20273 ;
  assign n20823 = ~n20248 & ~n20254 ;
  assign n20824 = ~n20229 & ~n20235 ;
  assign n20825 = ~n20191 & ~n20197 ;
  assign n20826 = x81 & n10905 ;
  assign n20827 = x79 & n11466 ;
  assign n20828 = x80 & n10900 ;
  assign n20829 = ~n20827 & ~n20828 ;
  assign n20830 = ~n20826 & n20829 ;
  assign n20831 = n2348 & n10908 ;
  assign n20832 = n20830 & ~n20831 ;
  assign n20833 = x41 & ~n20832 ;
  assign n20834 = x41 & ~n20833 ;
  assign n20835 = ~n20832 & ~n20833 ;
  assign n20836 = ~n20834 & ~n20835 ;
  assign n20837 = ~n20175 & ~n20177 ;
  assign n20838 = ~n20169 & ~n20171 ;
  assign n20839 = x75 & n14233 ;
  assign n20840 = x73 & n14876 ;
  assign n20841 = x74 & n14228 ;
  assign n20842 = ~n20840 & ~n20841 ;
  assign n20843 = ~n20839 & n20842 ;
  assign n20844 = n1150 & n14236 ;
  assign n20845 = n20843 & ~n20844 ;
  assign n20846 = x47 & ~n20845 ;
  assign n20847 = x47 & ~n20846 ;
  assign n20848 = ~n20845 & ~n20846 ;
  assign n20849 = ~n20847 & ~n20848 ;
  assign n20850 = ~n20163 & ~n20165 ;
  assign n20851 = ~n20157 & ~n20159 ;
  assign n20852 = x66 & n20143 ;
  assign n20853 = n19514 & ~n20142 ;
  assign n20854 = n20137 & n20853 ;
  assign n20855 = x64 & n20854 ;
  assign n20856 = x65 & n20138 ;
  assign n20857 = ~n20855 & ~n20856 ;
  assign n20858 = ~n20852 & n20857 ;
  assign n20859 = n194 & n20146 ;
  assign n20860 = n20858 & ~n20859 ;
  assign n20861 = x56 & ~n20860 ;
  assign n20862 = x56 & ~n20861 ;
  assign n20863 = ~n20860 & ~n20861 ;
  assign n20864 = ~n20862 & ~n20863 ;
  assign n20865 = ~n20153 & n20864 ;
  assign n20866 = n20153 & ~n20864 ;
  assign n20867 = ~n20865 & ~n20866 ;
  assign n20868 = x69 & n18025 ;
  assign n20869 = x67 & n18764 ;
  assign n20870 = x68 & n18020 ;
  assign n20871 = ~n20869 & ~n20870 ;
  assign n20872 = ~n20868 & n20871 ;
  assign n20873 = n398 & n18028 ;
  assign n20874 = n20872 & ~n20873 ;
  assign n20875 = x53 & ~n20874 ;
  assign n20876 = x53 & ~n20875 ;
  assign n20877 = ~n20874 & ~n20875 ;
  assign n20878 = ~n20876 & ~n20877 ;
  assign n20879 = n20867 & ~n20878 ;
  assign n20880 = ~n20867 & n20878 ;
  assign n20881 = ~n20851 & ~n20880 ;
  assign n20882 = ~n20879 & n20881 ;
  assign n20883 = ~n20851 & ~n20882 ;
  assign n20884 = ~n20879 & ~n20882 ;
  assign n20885 = ~n20880 & n20884 ;
  assign n20886 = ~n20883 & ~n20885 ;
  assign n20887 = x72 & n16076 ;
  assign n20888 = x70 & n16756 ;
  assign n20889 = x71 & n16071 ;
  assign n20890 = ~n20888 & ~n20889 ;
  assign n20891 = ~n20887 & n20890 ;
  assign n20892 = n717 & n16079 ;
  assign n20893 = n20891 & ~n20892 ;
  assign n20894 = x50 & ~n20893 ;
  assign n20895 = x50 & ~n20894 ;
  assign n20896 = ~n20893 & ~n20894 ;
  assign n20897 = ~n20895 & ~n20896 ;
  assign n20898 = n20886 & n20897 ;
  assign n20899 = ~n20886 & ~n20897 ;
  assign n20900 = ~n20898 & ~n20899 ;
  assign n20901 = ~n20850 & n20900 ;
  assign n20902 = n20850 & ~n20900 ;
  assign n20903 = ~n20901 & ~n20902 ;
  assign n20904 = n20849 & ~n20903 ;
  assign n20905 = ~n20849 & n20903 ;
  assign n20906 = ~n20904 & ~n20905 ;
  assign n20907 = ~n20838 & n20906 ;
  assign n20908 = n20838 & ~n20906 ;
  assign n20909 = ~n20907 & ~n20908 ;
  assign n20910 = x78 & n12506 ;
  assign n20911 = x76 & n13131 ;
  assign n20912 = x77 & n12501 ;
  assign n20913 = ~n20911 & ~n20912 ;
  assign n20914 = ~n20910 & n20913 ;
  assign n20915 = n1624 & n12509 ;
  assign n20916 = n20914 & ~n20915 ;
  assign n20917 = x44 & ~n20916 ;
  assign n20918 = x44 & ~n20917 ;
  assign n20919 = ~n20916 & ~n20917 ;
  assign n20920 = ~n20918 & ~n20919 ;
  assign n20921 = n20909 & ~n20920 ;
  assign n20922 = n20909 & ~n20921 ;
  assign n20923 = ~n20920 & ~n20921 ;
  assign n20924 = ~n20922 & ~n20923 ;
  assign n20925 = ~n20837 & ~n20924 ;
  assign n20926 = n20837 & n20924 ;
  assign n20927 = ~n20925 & ~n20926 ;
  assign n20928 = ~n20836 & n20927 ;
  assign n20929 = ~n20836 & ~n20928 ;
  assign n20930 = n20927 & ~n20928 ;
  assign n20931 = ~n20929 & ~n20930 ;
  assign n20932 = ~n20825 & ~n20931 ;
  assign n20933 = ~n20825 & ~n20932 ;
  assign n20934 = ~n20931 & ~n20932 ;
  assign n20935 = ~n20933 & ~n20934 ;
  assign n20936 = x84 & n9433 ;
  assign n20937 = x82 & n9915 ;
  assign n20938 = x83 & n9428 ;
  assign n20939 = ~n20937 & ~n20938 ;
  assign n20940 = ~n20936 & n20939 ;
  assign n20941 = n3114 & n9436 ;
  assign n20942 = n20940 & ~n20941 ;
  assign n20943 = x38 & ~n20942 ;
  assign n20944 = x38 & ~n20943 ;
  assign n20945 = ~n20942 & ~n20943 ;
  assign n20946 = ~n20944 & ~n20945 ;
  assign n20947 = ~n20935 & ~n20946 ;
  assign n20948 = ~n20935 & ~n20947 ;
  assign n20949 = ~n20946 & ~n20947 ;
  assign n20950 = ~n20948 & ~n20949 ;
  assign n20951 = ~n20215 & n20950 ;
  assign n20952 = n20215 & ~n20950 ;
  assign n20953 = ~n20951 & ~n20952 ;
  assign n20954 = x87 & n8006 ;
  assign n20955 = x85 & n8474 ;
  assign n20956 = x86 & n8001 ;
  assign n20957 = ~n20955 & ~n20956 ;
  assign n20958 = ~n20954 & n20957 ;
  assign n20959 = n3991 & n8009 ;
  assign n20960 = n20958 & ~n20959 ;
  assign n20961 = x35 & ~n20960 ;
  assign n20962 = x35 & ~n20961 ;
  assign n20963 = ~n20960 & ~n20961 ;
  assign n20964 = ~n20962 & ~n20963 ;
  assign n20965 = ~n20953 & ~n20964 ;
  assign n20966 = n20953 & n20964 ;
  assign n20967 = ~n20965 & ~n20966 ;
  assign n20968 = n20824 & ~n20967 ;
  assign n20969 = ~n20824 & n20967 ;
  assign n20970 = ~n20968 & ~n20969 ;
  assign n20971 = x90 & n6725 ;
  assign n20972 = x88 & n7129 ;
  assign n20973 = x89 & n6720 ;
  assign n20974 = ~n20972 & ~n20973 ;
  assign n20975 = ~n20971 & n20974 ;
  assign n20976 = n4986 & n6728 ;
  assign n20977 = n20975 & ~n20976 ;
  assign n20978 = x32 & ~n20977 ;
  assign n20979 = x32 & ~n20978 ;
  assign n20980 = ~n20977 & ~n20978 ;
  assign n20981 = ~n20979 & ~n20980 ;
  assign n20982 = n20970 & ~n20981 ;
  assign n20983 = ~n20970 & n20981 ;
  assign n20984 = ~n20823 & ~n20983 ;
  assign n20985 = ~n20982 & n20984 ;
  assign n20986 = ~n20823 & ~n20985 ;
  assign n20987 = ~n20982 & ~n20985 ;
  assign n20988 = ~n20983 & n20987 ;
  assign n20989 = ~n20986 & ~n20988 ;
  assign n20990 = x93 & n5560 ;
  assign n20991 = x91 & n5943 ;
  assign n20992 = x92 & n5555 ;
  assign n20993 = ~n20991 & ~n20992 ;
  assign n20994 = ~n20990 & n20993 ;
  assign n20995 = n5563 & n6094 ;
  assign n20996 = n20994 & ~n20995 ;
  assign n20997 = x29 & ~n20996 ;
  assign n20998 = x29 & ~n20997 ;
  assign n20999 = ~n20996 & ~n20997 ;
  assign n21000 = ~n20998 & ~n20999 ;
  assign n21001 = n20989 & n21000 ;
  assign n21002 = ~n20989 & ~n21000 ;
  assign n21003 = ~n21001 & ~n21002 ;
  assign n21004 = ~n20822 & n21003 ;
  assign n21005 = n20822 & ~n21003 ;
  assign n21006 = ~n21004 & ~n21005 ;
  assign n21007 = n20821 & ~n21006 ;
  assign n21008 = ~n20821 & n21006 ;
  assign n21009 = ~n21007 & ~n21008 ;
  assign n21010 = ~n20810 & n21009 ;
  assign n21011 = n20810 & ~n21009 ;
  assign n21012 = ~n21010 & ~n21011 ;
  assign n21013 = x99 & n3589 ;
  assign n21014 = x97 & n3878 ;
  assign n21015 = x98 & n3584 ;
  assign n21016 = ~n21014 & ~n21015 ;
  assign n21017 = ~n21013 & n21016 ;
  assign n21018 = n3592 & n8660 ;
  assign n21019 = n21017 & ~n21018 ;
  assign n21020 = x23 & ~n21019 ;
  assign n21021 = x23 & ~n21020 ;
  assign n21022 = ~n21019 & ~n21020 ;
  assign n21023 = ~n21021 & ~n21022 ;
  assign n21024 = n21012 & ~n21023 ;
  assign n21025 = n21012 & ~n21024 ;
  assign n21026 = ~n21023 & ~n21024 ;
  assign n21027 = ~n21025 & ~n21026 ;
  assign n21028 = ~n20305 & ~n20312 ;
  assign n21029 = n21027 & n21028 ;
  assign n21030 = ~n21027 & ~n21028 ;
  assign n21031 = ~n21029 & ~n21030 ;
  assign n21032 = x102 & n2751 ;
  assign n21033 = x100 & n3020 ;
  assign n21034 = x101 & n2746 ;
  assign n21035 = ~n21033 & ~n21034 ;
  assign n21036 = ~n21032 & n21035 ;
  assign n21037 = n2754 & n10092 ;
  assign n21038 = n21036 & ~n21037 ;
  assign n21039 = x20 & ~n21038 ;
  assign n21040 = x20 & ~n21039 ;
  assign n21041 = ~n21038 & ~n21039 ;
  assign n21042 = ~n21040 & ~n21041 ;
  assign n21043 = n21031 & ~n21042 ;
  assign n21044 = n21031 & ~n21043 ;
  assign n21045 = ~n21042 & ~n21043 ;
  assign n21046 = ~n21044 & ~n21045 ;
  assign n21047 = ~n20325 & ~n20331 ;
  assign n21048 = n21046 & n21047 ;
  assign n21049 = ~n21046 & ~n21047 ;
  assign n21050 = ~n21048 & ~n21049 ;
  assign n21051 = x105 & n2093 ;
  assign n21052 = x103 & n2275 ;
  assign n21053 = x104 & n2088 ;
  assign n21054 = ~n21052 & ~n21053 ;
  assign n21055 = ~n21051 & n21054 ;
  assign n21056 = n2096 & n11648 ;
  assign n21057 = n21055 & ~n21056 ;
  assign n21058 = x17 & ~n21057 ;
  assign n21059 = x17 & ~n21058 ;
  assign n21060 = ~n21057 & ~n21058 ;
  assign n21061 = ~n21059 & ~n21060 ;
  assign n21062 = n21050 & ~n21061 ;
  assign n21063 = n21050 & ~n21062 ;
  assign n21064 = ~n21061 & ~n21062 ;
  assign n21065 = ~n21063 & ~n21064 ;
  assign n21066 = ~n20344 & ~n20350 ;
  assign n21067 = n21065 & n21066 ;
  assign n21068 = ~n21065 & ~n21066 ;
  assign n21069 = ~n21067 & ~n21068 ;
  assign n21070 = x108 & n1434 ;
  assign n21071 = x106 & n1646 ;
  assign n21072 = x107 & n1429 ;
  assign n21073 = ~n21071 & ~n21072 ;
  assign n21074 = ~n21070 & n21073 ;
  assign n21075 = n1437 & n13323 ;
  assign n21076 = n21074 & ~n21075 ;
  assign n21077 = x14 & ~n21076 ;
  assign n21078 = x14 & ~n21077 ;
  assign n21079 = ~n21076 & ~n21077 ;
  assign n21080 = ~n21078 & ~n21079 ;
  assign n21081 = n21069 & ~n21080 ;
  assign n21082 = ~n21069 & n21080 ;
  assign n21083 = ~n20368 & ~n21082 ;
  assign n21084 = ~n21081 & n21083 ;
  assign n21085 = ~n20368 & ~n21084 ;
  assign n21086 = ~n21081 & ~n21084 ;
  assign n21087 = ~n21082 & n21086 ;
  assign n21088 = ~n21085 & ~n21087 ;
  assign n21089 = x111 & n945 ;
  assign n21090 = x109 & n1099 ;
  assign n21091 = x110 & n940 ;
  assign n21092 = ~n21090 & ~n21091 ;
  assign n21093 = ~n21089 & n21092 ;
  assign n21094 = n948 & n15111 ;
  assign n21095 = n21093 & ~n21094 ;
  assign n21096 = x11 & ~n21095 ;
  assign n21097 = x11 & ~n21096 ;
  assign n21098 = ~n21095 & ~n21096 ;
  assign n21099 = ~n21097 & ~n21098 ;
  assign n21100 = ~n21088 & ~n21099 ;
  assign n21101 = ~n21088 & ~n21100 ;
  assign n21102 = ~n21099 & ~n21100 ;
  assign n21103 = ~n21101 & ~n21102 ;
  assign n21104 = ~n20809 & ~n21103 ;
  assign n21105 = n20809 & n21103 ;
  assign n21106 = ~n21104 & ~n21105 ;
  assign n21107 = ~n20808 & n21106 ;
  assign n21108 = ~n20808 & ~n21107 ;
  assign n21109 = n21106 & ~n21107 ;
  assign n21110 = ~n21108 & ~n21109 ;
  assign n21111 = ~n20797 & ~n21110 ;
  assign n21112 = ~n20797 & ~n21111 ;
  assign n21113 = ~n21110 & ~n21111 ;
  assign n21114 = ~n21112 & ~n21113 ;
  assign n21115 = x117 & n293 ;
  assign n21116 = x115 & n373 ;
  assign n21117 = x116 & n288 ;
  assign n21118 = ~n21116 & ~n21117 ;
  assign n21119 = ~n21115 & n21118 ;
  assign n21120 = n296 & n19026 ;
  assign n21121 = n21119 & ~n21120 ;
  assign n21122 = x5 & ~n21121 ;
  assign n21123 = x5 & ~n21122 ;
  assign n21124 = ~n21121 & ~n21122 ;
  assign n21125 = ~n21123 & ~n21124 ;
  assign n21126 = n21114 & n21125 ;
  assign n21127 = ~n21114 & ~n21125 ;
  assign n21128 = ~n21126 & ~n21127 ;
  assign n21129 = ~n20796 & n21128 ;
  assign n21130 = n20796 & ~n21128 ;
  assign n21131 = ~n21129 & ~n21130 ;
  assign n21132 = x120 & n146 ;
  assign n21133 = x118 & n182 ;
  assign n21134 = x119 & n141 ;
  assign n21135 = ~n21133 & ~n21134 ;
  assign n21136 = ~n21132 & n21135 ;
  assign n21137 = ~n20419 & ~n20421 ;
  assign n21138 = ~x119 & ~x120 ;
  assign n21139 = x119 & x120 ;
  assign n21140 = ~n21138 & ~n21139 ;
  assign n21141 = ~n21137 & n21140 ;
  assign n21142 = n21137 & ~n21140 ;
  assign n21143 = ~n21141 & ~n21142 ;
  assign n21144 = n149 & n21143 ;
  assign n21145 = n21136 & ~n21144 ;
  assign n21146 = x2 & ~n21145 ;
  assign n21147 = x2 & ~n21146 ;
  assign n21148 = ~n21145 & ~n21146 ;
  assign n21149 = ~n21147 & ~n21148 ;
  assign n21150 = n21131 & ~n21149 ;
  assign n21151 = n21131 & ~n21150 ;
  assign n21152 = ~n21149 & ~n21150 ;
  assign n21153 = ~n21151 & ~n21152 ;
  assign n21154 = ~n20430 & ~n20433 ;
  assign n21155 = ~n21153 & ~n21154 ;
  assign n21156 = n21153 & n21154 ;
  assign n21157 = ~n21155 & ~n21156 ;
  assign n21517 = n21157 & x184 ;
  assign n21158 = ~n20437 & ~n20766 ;
  assign n21159 = ~n20763 & ~n21158 ;
  assign n21160 = ~n20747 & ~n20749 ;
  assign n21161 = ~x114 & n574 ;
  assign n21162 = ~x112 & n673 ;
  assign n21163 = ~x113 & n569 ;
  assign n21164 = ~n21162 & ~n21163 ;
  assign n21165 = ~n21161 & n21164 ;
  assign n21166 = n577 & n17333 ;
  assign n21167 = n21165 & ~n21166 ;
  assign n21168 = ~x8 & ~n21167 ;
  assign n21169 = ~x8 & ~n21168 ;
  assign n21170 = ~n21167 & ~n21168 ;
  assign n21171 = ~n21169 & ~n21170 ;
  assign n21172 = ~n20741 & ~n20743 ;
  assign n21173 = ~n20644 & ~n20650 ;
  assign n21174 = ~x96 & n4531 ;
  assign n21175 = ~x94 & n4847 ;
  assign n21176 = ~x95 & n4526 ;
  assign n21177 = ~n21175 & ~n21176 ;
  assign n21178 = ~n21174 & n21177 ;
  assign n21179 = n4534 & n7531 ;
  assign n21180 = n21178 & ~n21179 ;
  assign n21181 = ~x26 & ~n21180 ;
  assign n21182 = ~x26 & ~n21181 ;
  assign n21183 = ~n21180 & ~n21181 ;
  assign n21184 = ~n21182 & ~n21183 ;
  assign n21185 = ~n20625 & ~n20631 ;
  assign n21186 = ~n20606 & ~n20612 ;
  assign n21187 = ~n20587 & ~n20593 ;
  assign n21188 = ~n20549 & ~n20555 ;
  assign n21189 = ~x81 & n10905 ;
  assign n21190 = ~x79 & n11466 ;
  assign n21191 = ~x80 & n10900 ;
  assign n21192 = ~n21190 & ~n21191 ;
  assign n21193 = ~n21189 & n21192 ;
  assign n21194 = n2460 & n10908 ;
  assign n21195 = n21193 & ~n21194 ;
  assign n21196 = ~x41 & ~n21195 ;
  assign n21197 = ~x41 & ~n21196 ;
  assign n21198 = ~n21195 & ~n21196 ;
  assign n21199 = ~n21197 & ~n21198 ;
  assign n21200 = ~n20533 & ~n20535 ;
  assign n21201 = ~n20527 & ~n20529 ;
  assign n21202 = ~x75 & n14233 ;
  assign n21203 = ~x73 & n14876 ;
  assign n21204 = ~x74 & n14228 ;
  assign n21205 = ~n21203 & ~n21204 ;
  assign n21206 = ~n21202 & n21205 ;
  assign n21207 = n1225 & n14236 ;
  assign n21208 = n21206 & ~n21207 ;
  assign n21209 = ~x47 & ~n21208 ;
  assign n21210 = ~x47 & ~n21209 ;
  assign n21211 = ~n21208 & ~n21209 ;
  assign n21212 = ~n21210 & ~n21211 ;
  assign n21213 = ~n20521 & ~n20523 ;
  assign n21214 = ~n20515 & ~n20517 ;
  assign n21215 = ~x66 & n20143 ;
  assign n21216 = ~x64 & n20854 ;
  assign n21217 = ~x65 & n20138 ;
  assign n21218 = ~n21216 & ~n21217 ;
  assign n21219 = ~n21215 & n21218 ;
  assign n21220 = n214 & n20146 ;
  assign n21221 = n21219 & ~n21220 ;
  assign n21222 = ~x56 & ~n21221 ;
  assign n21223 = ~x56 & ~n21222 ;
  assign n21224 = ~n21221 & ~n21222 ;
  assign n21225 = ~n21223 & ~n21224 ;
  assign n21226 = ~n20511 & n21225 ;
  assign n21227 = n20511 & ~n21225 ;
  assign n21228 = ~n21226 & ~n21227 ;
  assign n21229 = ~x69 & n18025 ;
  assign n21230 = ~x67 & n18764 ;
  assign n21231 = ~x68 & n18020 ;
  assign n21232 = ~n21230 & ~n21231 ;
  assign n21233 = ~n21229 & n21232 ;
  assign n21234 = n435 & n18028 ;
  assign n21235 = n21233 & ~n21234 ;
  assign n21236 = ~x53 & ~n21235 ;
  assign n21237 = ~x53 & ~n21236 ;
  assign n21238 = ~n21235 & ~n21236 ;
  assign n21239 = ~n21237 & ~n21238 ;
  assign n21240 = n21228 & ~n21239 ;
  assign n21241 = ~n21228 & n21239 ;
  assign n21242 = ~n21214 & ~n21241 ;
  assign n21243 = ~n21240 & n21242 ;
  assign n21244 = ~n21214 & ~n21243 ;
  assign n21245 = ~n21240 & ~n21243 ;
  assign n21246 = ~n21241 & n21245 ;
  assign n21247 = ~n21244 & ~n21246 ;
  assign n21248 = ~x72 & n16076 ;
  assign n21249 = ~x70 & n16756 ;
  assign n21250 = ~x71 & n16071 ;
  assign n21251 = ~n21249 & ~n21250 ;
  assign n21252 = ~n21248 & n21251 ;
  assign n21253 = n773 & n16079 ;
  assign n21254 = n21252 & ~n21253 ;
  assign n21255 = ~x50 & ~n21254 ;
  assign n21256 = ~x50 & ~n21255 ;
  assign n21257 = ~n21254 & ~n21255 ;
  assign n21258 = ~n21256 & ~n21257 ;
  assign n21259 = n21247 & n21258 ;
  assign n21260 = ~n21247 & ~n21258 ;
  assign n21261 = ~n21259 & ~n21260 ;
  assign n21262 = ~n21213 & n21261 ;
  assign n21263 = n21213 & ~n21261 ;
  assign n21264 = ~n21262 & ~n21263 ;
  assign n21265 = n21212 & ~n21264 ;
  assign n21266 = ~n21212 & n21264 ;
  assign n21267 = ~n21265 & ~n21266 ;
  assign n21268 = ~n21201 & n21267 ;
  assign n21269 = n21201 & ~n21267 ;
  assign n21270 = ~n21268 & ~n21269 ;
  assign n21271 = ~x78 & n12506 ;
  assign n21272 = ~x76 & n13131 ;
  assign n21273 = ~x77 & n12501 ;
  assign n21274 = ~n21272 & ~n21273 ;
  assign n21275 = ~n21271 & n21274 ;
  assign n21276 = n1718 & n12509 ;
  assign n21277 = n21275 & ~n21276 ;
  assign n21278 = ~x44 & ~n21277 ;
  assign n21279 = ~x44 & ~n21278 ;
  assign n21280 = ~n21277 & ~n21278 ;
  assign n21281 = ~n21279 & ~n21280 ;
  assign n21282 = n21270 & ~n21281 ;
  assign n21283 = n21270 & ~n21282 ;
  assign n21284 = ~n21281 & ~n21282 ;
  assign n21285 = ~n21283 & ~n21284 ;
  assign n21286 = ~n21200 & ~n21285 ;
  assign n21287 = n21200 & n21285 ;
  assign n21288 = ~n21286 & ~n21287 ;
  assign n21289 = ~n21199 & n21288 ;
  assign n21290 = ~n21199 & ~n21289 ;
  assign n21291 = n21288 & ~n21289 ;
  assign n21292 = ~n21290 & ~n21291 ;
  assign n21293 = ~n21188 & ~n21292 ;
  assign n21294 = ~n21188 & ~n21293 ;
  assign n21295 = ~n21292 & ~n21293 ;
  assign n21296 = ~n21294 & ~n21295 ;
  assign n21297 = ~x84 & n9433 ;
  assign n21298 = ~x82 & n9915 ;
  assign n21299 = ~x83 & n9428 ;
  assign n21300 = ~n21298 & ~n21299 ;
  assign n21301 = ~n21297 & n21300 ;
  assign n21302 = n3247 & n9436 ;
  assign n21303 = n21301 & ~n21302 ;
  assign n21304 = ~x38 & ~n21303 ;
  assign n21305 = ~x38 & ~n21304 ;
  assign n21306 = ~n21303 & ~n21304 ;
  assign n21307 = ~n21305 & ~n21306 ;
  assign n21308 = ~n21296 & ~n21307 ;
  assign n21309 = ~n21296 & ~n21308 ;
  assign n21310 = ~n21307 & ~n21308 ;
  assign n21311 = ~n21309 & ~n21310 ;
  assign n21312 = ~n20573 & n21311 ;
  assign n21313 = n20573 & ~n21311 ;
  assign n21314 = ~n21312 & ~n21313 ;
  assign n21315 = ~x87 & n8006 ;
  assign n21316 = ~x85 & n8474 ;
  assign n21317 = ~x86 & n8001 ;
  assign n21318 = ~n21316 & ~n21317 ;
  assign n21319 = ~n21315 & n21318 ;
  assign n21320 = n4143 & n8009 ;
  assign n21321 = n21319 & ~n21320 ;
  assign n21322 = ~x35 & ~n21321 ;
  assign n21323 = ~x35 & ~n21322 ;
  assign n21324 = ~n21321 & ~n21322 ;
  assign n21325 = ~n21323 & ~n21324 ;
  assign n21326 = ~n21314 & ~n21325 ;
  assign n21327 = n21314 & n21325 ;
  assign n21328 = ~n21326 & ~n21327 ;
  assign n21329 = n21187 & ~n21328 ;
  assign n21330 = ~n21187 & n21328 ;
  assign n21331 = ~n21329 & ~n21330 ;
  assign n21332 = ~x90 & n6725 ;
  assign n21333 = ~x88 & n7129 ;
  assign n21334 = ~x89 & n6720 ;
  assign n21335 = ~n21333 & ~n21334 ;
  assign n21336 = ~n21332 & n21335 ;
  assign n21337 = n5155 & n6728 ;
  assign n21338 = n21336 & ~n21337 ;
  assign n21339 = ~x32 & ~n21338 ;
  assign n21340 = ~x32 & ~n21339 ;
  assign n21341 = ~n21338 & ~n21339 ;
  assign n21342 = ~n21340 & ~n21341 ;
  assign n21343 = n21331 & ~n21342 ;
  assign n21344 = ~n21331 & n21342 ;
  assign n21345 = ~n21186 & ~n21344 ;
  assign n21346 = ~n21343 & n21345 ;
  assign n21347 = ~n21186 & ~n21346 ;
  assign n21348 = ~n21343 & ~n21346 ;
  assign n21349 = ~n21344 & n21348 ;
  assign n21350 = ~n21347 & ~n21349 ;
  assign n21351 = ~x93 & n5560 ;
  assign n21352 = ~x91 & n5943 ;
  assign n21353 = ~x92 & n5555 ;
  assign n21354 = ~n21352 & ~n21353 ;
  assign n21355 = ~n21351 & n21354 ;
  assign n21356 = n5563 & n6285 ;
  assign n21357 = n21355 & ~n21356 ;
  assign n21358 = ~x29 & ~n21357 ;
  assign n21359 = ~x29 & ~n21358 ;
  assign n21360 = ~n21357 & ~n21358 ;
  assign n21361 = ~n21359 & ~n21360 ;
  assign n21362 = n21350 & n21361 ;
  assign n21363 = ~n21350 & ~n21361 ;
  assign n21364 = ~n21362 & ~n21363 ;
  assign n21365 = ~n21185 & n21364 ;
  assign n21366 = n21185 & ~n21364 ;
  assign n21367 = ~n21365 & ~n21366 ;
  assign n21368 = n21184 & ~n21367 ;
  assign n21369 = ~n21184 & n21367 ;
  assign n21370 = ~n21368 & ~n21369 ;
  assign n21371 = ~n21173 & n21370 ;
  assign n21372 = n21173 & ~n21370 ;
  assign n21373 = ~n21371 & ~n21372 ;
  assign n21374 = ~x99 & n3589 ;
  assign n21375 = ~x97 & n3878 ;
  assign n21376 = ~x98 & n3584 ;
  assign n21377 = ~n21375 & ~n21376 ;
  assign n21378 = ~n21374 & n21377 ;
  assign n21379 = n3592 & n8885 ;
  assign n21380 = n21378 & ~n21379 ;
  assign n21381 = ~x23 & ~n21380 ;
  assign n21382 = ~x23 & ~n21381 ;
  assign n21383 = ~n21380 & ~n21381 ;
  assign n21384 = ~n21382 & ~n21383 ;
  assign n21385 = n21373 & ~n21384 ;
  assign n21386 = n21373 & ~n21385 ;
  assign n21387 = ~n21384 & ~n21385 ;
  assign n21388 = ~n21386 & ~n21387 ;
  assign n21389 = ~n20663 & ~n20670 ;
  assign n21390 = n21388 & n21389 ;
  assign n21391 = ~n21388 & ~n21389 ;
  assign n21392 = ~n21390 & ~n21391 ;
  assign n21393 = ~x102 & n2751 ;
  assign n21394 = ~x100 & n3020 ;
  assign n21395 = ~x101 & n2746 ;
  assign n21396 = ~n21394 & ~n21395 ;
  assign n21397 = ~n21393 & n21396 ;
  assign n21398 = n2754 & n10333 ;
  assign n21399 = n21397 & ~n21398 ;
  assign n21400 = ~x20 & ~n21399 ;
  assign n21401 = ~x20 & ~n21400 ;
  assign n21402 = ~n21399 & ~n21400 ;
  assign n21403 = ~n21401 & ~n21402 ;
  assign n21404 = n21392 & ~n21403 ;
  assign n21405 = n21392 & ~n21404 ;
  assign n21406 = ~n21403 & ~n21404 ;
  assign n21407 = ~n21405 & ~n21406 ;
  assign n21408 = ~n20683 & ~n20689 ;
  assign n21409 = n21407 & n21408 ;
  assign n21410 = ~n21407 & ~n21408 ;
  assign n21411 = ~n21409 & ~n21410 ;
  assign n21412 = ~x105 & n2093 ;
  assign n21413 = ~x103 & n2275 ;
  assign n21414 = ~x104 & n2088 ;
  assign n21415 = ~n21413 & ~n21414 ;
  assign n21416 = ~n21412 & n21415 ;
  assign n21417 = n2096 & n11907 ;
  assign n21418 = n21416 & ~n21417 ;
  assign n21419 = ~x17 & ~n21418 ;
  assign n21420 = ~x17 & ~n21419 ;
  assign n21421 = ~n21418 & ~n21419 ;
  assign n21422 = ~n21420 & ~n21421 ;
  assign n21423 = n21411 & ~n21422 ;
  assign n21424 = n21411 & ~n21423 ;
  assign n21425 = ~n21422 & ~n21423 ;
  assign n21426 = ~n21424 & ~n21425 ;
  assign n21427 = ~n20702 & ~n20708 ;
  assign n21428 = n21426 & n21427 ;
  assign n21429 = ~n21426 & ~n21427 ;
  assign n21430 = ~n21428 & ~n21429 ;
  assign n21431 = ~x108 & n1434 ;
  assign n21432 = ~x106 & n1646 ;
  assign n21433 = ~x107 & n1429 ;
  assign n21434 = ~n21432 & ~n21433 ;
  assign n21435 = ~n21431 & n21434 ;
  assign n21436 = n1437 & n13601 ;
  assign n21437 = n21435 & ~n21436 ;
  assign n21438 = ~x14 & ~n21437 ;
  assign n21439 = ~x14 & ~n21438 ;
  assign n21440 = ~n21437 & ~n21438 ;
  assign n21441 = ~n21439 & ~n21440 ;
  assign n21442 = n21430 & ~n21441 ;
  assign n21443 = ~n21430 & n21441 ;
  assign n21444 = ~n20726 & ~n21443 ;
  assign n21445 = ~n21442 & n21444 ;
  assign n21446 = ~n20726 & ~n21445 ;
  assign n21447 = ~n21442 & ~n21445 ;
  assign n21448 = ~n21443 & n21447 ;
  assign n21449 = ~n21446 & ~n21448 ;
  assign n21450 = ~x111 & n945 ;
  assign n21451 = ~x109 & n1099 ;
  assign n21452 = ~x110 & n940 ;
  assign n21453 = ~n21451 & ~n21452 ;
  assign n21454 = ~n21450 & n21453 ;
  assign n21455 = n948 & n15411 ;
  assign n21456 = n21454 & ~n21455 ;
  assign n21457 = ~x11 & ~n21456 ;
  assign n21458 = ~x11 & ~n21457 ;
  assign n21459 = ~n21456 & ~n21457 ;
  assign n21460 = ~n21458 & ~n21459 ;
  assign n21461 = ~n21449 & ~n21460 ;
  assign n21462 = ~n21449 & ~n21461 ;
  assign n21463 = ~n21460 & ~n21461 ;
  assign n21464 = ~n21462 & ~n21463 ;
  assign n21465 = ~n21172 & ~n21464 ;
  assign n21466 = n21172 & n21464 ;
  assign n21467 = ~n21465 & ~n21466 ;
  assign n21468 = ~n21171 & n21467 ;
  assign n21469 = ~n21171 & ~n21468 ;
  assign n21470 = n21467 & ~n21468 ;
  assign n21471 = ~n21469 & ~n21470 ;
  assign n21472 = ~n21160 & ~n21471 ;
  assign n21473 = ~n21160 & ~n21472 ;
  assign n21474 = ~n21471 & ~n21472 ;
  assign n21475 = ~n21473 & ~n21474 ;
  assign n21476 = ~x117 & n293 ;
  assign n21477 = ~x115 & n373 ;
  assign n21478 = ~x116 & n288 ;
  assign n21479 = ~n21477 & ~n21478 ;
  assign n21480 = ~n21476 & n21479 ;
  assign n21481 = n296 & n19365 ;
  assign n21482 = n21480 & ~n21481 ;
  assign n21483 = ~x5 & ~n21482 ;
  assign n21484 = ~x5 & ~n21483 ;
  assign n21485 = ~n21482 & ~n21483 ;
  assign n21486 = ~n21484 & ~n21485 ;
  assign n21487 = n21475 & n21486 ;
  assign n21488 = ~n21475 & ~n21486 ;
  assign n21489 = ~n21487 & ~n21488 ;
  assign n21490 = ~n21159 & n21489 ;
  assign n21491 = n21159 & ~n21489 ;
  assign n21492 = ~n21490 & ~n21491 ;
  assign n21493 = ~x120 & n164 ;
  assign n21494 = ~x118 & n205 ;
  assign n21495 = ~x119 & n162 ;
  assign n21496 = ~n21494 & ~n21495 ;
  assign n21497 = ~n21493 & n21496 ;
  assign n21498 = ~n20418 & ~n20776 ;
  assign n21499 = n21140 & ~n21498 ;
  assign n21500 = ~n21140 & n21498 ;
  assign n21501 = ~n21499 & ~n21500 ;
  assign n21502 = n167 & n21501 ;
  assign n21503 = n21497 & ~n21502 ;
  assign n21504 = ~x2 & ~n21503 ;
  assign n21505 = ~x2 & ~n21504 ;
  assign n21506 = ~n21503 & ~n21504 ;
  assign n21507 = ~n21505 & ~n21506 ;
  assign n21508 = n21492 & ~n21507 ;
  assign n21509 = n21492 & ~n21508 ;
  assign n21510 = ~n21507 & ~n21508 ;
  assign n21511 = ~n21509 & ~n21510 ;
  assign n21512 = ~n20785 & ~n20788 ;
  assign n21513 = ~n21511 & ~n21512 ;
  assign n21514 = n21511 & n21512 ;
  assign n21515 = ~n21513 & ~n21514 ;
  assign n21518 = ~n21515 & ~x184 ;
  assign n21519 = ~n21517 & ~n21518 ;
  assign n21520 = ~n21127 & ~n21129 ;
  assign n21521 = x118 & n293 ;
  assign n21522 = x116 & n373 ;
  assign n21523 = x117 & n288 ;
  assign n21524 = ~n21522 & ~n21523 ;
  assign n21525 = ~n21521 & n21524 ;
  assign n21526 = n296 & n19395 ;
  assign n21527 = n21525 & ~n21526 ;
  assign n21528 = x5 & ~n21527 ;
  assign n21529 = x5 & ~n21528 ;
  assign n21530 = ~n21527 & ~n21528 ;
  assign n21531 = ~n21529 & ~n21530 ;
  assign n21532 = ~n21107 & ~n21111 ;
  assign n21533 = x115 & n574 ;
  assign n21534 = x113 & n673 ;
  assign n21535 = x114 & n569 ;
  assign n21536 = ~n21534 & ~n21535 ;
  assign n21537 = ~n21533 & n21536 ;
  assign n21538 = n577 & n17364 ;
  assign n21539 = n21537 & ~n21538 ;
  assign n21540 = x8 & ~n21539 ;
  assign n21541 = x8 & ~n21540 ;
  assign n21542 = ~n21539 & ~n21540 ;
  assign n21543 = ~n21541 & ~n21542 ;
  assign n21544 = ~n21100 & ~n21104 ;
  assign n21545 = x112 & n945 ;
  assign n21546 = x110 & n1099 ;
  assign n21547 = x111 & n940 ;
  assign n21548 = ~n21546 & ~n21547 ;
  assign n21549 = ~n21545 & n21548 ;
  assign n21550 = n948 & n15442 ;
  assign n21551 = n21549 & ~n21550 ;
  assign n21552 = x11 & ~n21551 ;
  assign n21553 = x11 & ~n21552 ;
  assign n21554 = ~n21551 & ~n21552 ;
  assign n21555 = ~n21553 & ~n21554 ;
  assign n21556 = x109 & n1434 ;
  assign n21557 = x107 & n1646 ;
  assign n21558 = x108 & n1429 ;
  assign n21559 = ~n21557 & ~n21558 ;
  assign n21560 = ~n21556 & n21559 ;
  assign n21561 = n1437 & n13894 ;
  assign n21562 = n21560 & ~n21561 ;
  assign n21563 = x14 & ~n21562 ;
  assign n21564 = x14 & ~n21563 ;
  assign n21565 = ~n21562 & ~n21563 ;
  assign n21566 = ~n21564 & ~n21565 ;
  assign n21567 = ~n21062 & ~n21068 ;
  assign n21568 = ~n21024 & ~n21030 ;
  assign n21569 = ~n21008 & ~n21010 ;
  assign n21570 = ~n21002 & ~n21004 ;
  assign n21571 = x94 & n5560 ;
  assign n21572 = x92 & n5943 ;
  assign n21573 = x93 & n5555 ;
  assign n21574 = ~n21572 & ~n21573 ;
  assign n21575 = ~n21571 & n21574 ;
  assign n21576 = n5563 & n6483 ;
  assign n21577 = n21575 & ~n21576 ;
  assign n21578 = x29 & ~n21577 ;
  assign n21579 = x29 & ~n21578 ;
  assign n21580 = ~n21577 & ~n21578 ;
  assign n21581 = ~n21579 & ~n21580 ;
  assign n21582 = ~n20215 & ~n20950 ;
  assign n21583 = ~n20947 & ~n21582 ;
  assign n21584 = x85 & n9433 ;
  assign n21585 = x83 & n9915 ;
  assign n21586 = x84 & n9428 ;
  assign n21587 = ~n21585 & ~n21586 ;
  assign n21588 = ~n21584 & n21587 ;
  assign n21589 = n3389 & n9436 ;
  assign n21590 = n21588 & ~n21589 ;
  assign n21591 = x38 & ~n21590 ;
  assign n21592 = x38 & ~n21591 ;
  assign n21593 = ~n21590 & ~n21591 ;
  assign n21594 = ~n21592 & ~n21593 ;
  assign n21595 = ~n20928 & ~n20932 ;
  assign n21596 = x82 & n10905 ;
  assign n21597 = x80 & n11466 ;
  assign n21598 = x81 & n10900 ;
  assign n21599 = ~n21597 & ~n21598 ;
  assign n21600 = ~n21596 & n21599 ;
  assign n21601 = n2584 & n10908 ;
  assign n21602 = n21600 & ~n21601 ;
  assign n21603 = x41 & ~n21602 ;
  assign n21604 = x41 & ~n21603 ;
  assign n21605 = ~n21602 & ~n21603 ;
  assign n21606 = ~n21604 & ~n21605 ;
  assign n21607 = ~n20921 & ~n20925 ;
  assign n21608 = x79 & n12506 ;
  assign n21609 = x77 & n13131 ;
  assign n21610 = x78 & n12501 ;
  assign n21611 = ~n21609 & ~n21610 ;
  assign n21612 = ~n21608 & n21611 ;
  assign n21613 = n1817 & n12509 ;
  assign n21614 = n21612 & ~n21613 ;
  assign n21615 = x44 & ~n21614 ;
  assign n21616 = x44 & ~n21615 ;
  assign n21617 = ~n21614 & ~n21615 ;
  assign n21618 = ~n21616 & ~n21617 ;
  assign n21619 = ~n20905 & ~n20907 ;
  assign n21620 = x76 & n14233 ;
  assign n21621 = x74 & n14876 ;
  assign n21622 = x75 & n14228 ;
  assign n21623 = ~n21621 & ~n21622 ;
  assign n21624 = ~n21620 & n21623 ;
  assign n21625 = n1311 & n14236 ;
  assign n21626 = n21624 & ~n21625 ;
  assign n21627 = x47 & ~n21626 ;
  assign n21628 = x47 & ~n21627 ;
  assign n21629 = ~n21626 & ~n21627 ;
  assign n21630 = ~n21628 & ~n21629 ;
  assign n21631 = ~n20899 & ~n20901 ;
  assign n21632 = x56 & ~x57 ;
  assign n21633 = ~x56 & x57 ;
  assign n21634 = ~n21632 & ~n21633 ;
  assign n21635 = x64 & ~n21634 ;
  assign n21636 = ~n20866 & n21635 ;
  assign n21637 = n20866 & ~n21635 ;
  assign n21638 = ~n21636 & ~n21637 ;
  assign n21639 = x67 & n20143 ;
  assign n21640 = x65 & n20854 ;
  assign n21641 = x66 & n20138 ;
  assign n21642 = ~n21640 & ~n21641 ;
  assign n21643 = ~n21639 & n21642 ;
  assign n21644 = n240 & n20146 ;
  assign n21645 = n21643 & ~n21644 ;
  assign n21646 = x56 & ~n21645 ;
  assign n21647 = x56 & ~n21646 ;
  assign n21648 = ~n21645 & ~n21646 ;
  assign n21649 = ~n21647 & ~n21648 ;
  assign n21650 = ~n21638 & ~n21649 ;
  assign n21651 = n21638 & n21649 ;
  assign n21652 = ~n21650 & ~n21651 ;
  assign n21653 = x70 & n18025 ;
  assign n21654 = x68 & n18764 ;
  assign n21655 = x69 & n18020 ;
  assign n21656 = ~n21654 & ~n21655 ;
  assign n21657 = ~n21653 & n21656 ;
  assign n21658 = n488 & n18028 ;
  assign n21659 = n21657 & ~n21658 ;
  assign n21660 = x53 & ~n21659 ;
  assign n21661 = x53 & ~n21660 ;
  assign n21662 = ~n21659 & ~n21660 ;
  assign n21663 = ~n21661 & ~n21662 ;
  assign n21664 = n21652 & ~n21663 ;
  assign n21665 = n21652 & ~n21664 ;
  assign n21666 = ~n21663 & ~n21664 ;
  assign n21667 = ~n21665 & ~n21666 ;
  assign n21668 = ~n20884 & n21667 ;
  assign n21669 = n20884 & ~n21667 ;
  assign n21670 = ~n21668 & ~n21669 ;
  assign n21671 = x73 & n16076 ;
  assign n21672 = x71 & n16756 ;
  assign n21673 = x72 & n16071 ;
  assign n21674 = ~n21672 & ~n21673 ;
  assign n21675 = ~n21671 & n21674 ;
  assign n21676 = n843 & n16079 ;
  assign n21677 = n21675 & ~n21676 ;
  assign n21678 = x50 & ~n21677 ;
  assign n21679 = x50 & ~n21678 ;
  assign n21680 = ~n21677 & ~n21678 ;
  assign n21681 = ~n21679 & ~n21680 ;
  assign n21682 = ~n21670 & ~n21681 ;
  assign n21683 = n21670 & n21681 ;
  assign n21684 = ~n21682 & ~n21683 ;
  assign n21685 = ~n21631 & n21684 ;
  assign n21686 = n21631 & ~n21684 ;
  assign n21687 = ~n21685 & ~n21686 ;
  assign n21688 = n21630 & ~n21687 ;
  assign n21689 = ~n21630 & n21687 ;
  assign n21690 = ~n21688 & ~n21689 ;
  assign n21691 = ~n21619 & n21690 ;
  assign n21692 = n21619 & ~n21690 ;
  assign n21693 = ~n21691 & ~n21692 ;
  assign n21694 = ~n21618 & n21693 ;
  assign n21695 = n21618 & ~n21693 ;
  assign n21696 = ~n21694 & ~n21695 ;
  assign n21697 = ~n21607 & n21696 ;
  assign n21698 = n21607 & ~n21696 ;
  assign n21699 = ~n21697 & ~n21698 ;
  assign n21700 = ~n21606 & n21699 ;
  assign n21701 = ~n21606 & ~n21700 ;
  assign n21702 = n21699 & ~n21700 ;
  assign n21703 = ~n21701 & ~n21702 ;
  assign n21704 = ~n21595 & ~n21703 ;
  assign n21705 = n21595 & ~n21702 ;
  assign n21706 = ~n21701 & n21705 ;
  assign n21707 = ~n21704 & ~n21706 ;
  assign n21708 = ~n21594 & n21707 ;
  assign n21709 = n21594 & ~n21707 ;
  assign n21710 = ~n21708 & ~n21709 ;
  assign n21711 = ~n21583 & n21710 ;
  assign n21712 = n21583 & ~n21710 ;
  assign n21713 = ~n21711 & ~n21712 ;
  assign n21714 = x88 & n8006 ;
  assign n21715 = x86 & n8474 ;
  assign n21716 = x87 & n8001 ;
  assign n21717 = ~n21715 & ~n21716 ;
  assign n21718 = ~n21714 & n21717 ;
  assign n21719 = n4305 & n8009 ;
  assign n21720 = n21718 & ~n21719 ;
  assign n21721 = x35 & ~n21720 ;
  assign n21722 = x35 & ~n21721 ;
  assign n21723 = ~n21720 & ~n21721 ;
  assign n21724 = ~n21722 & ~n21723 ;
  assign n21725 = n21713 & ~n21724 ;
  assign n21726 = n21713 & ~n21725 ;
  assign n21727 = ~n21724 & ~n21725 ;
  assign n21728 = ~n21726 & ~n21727 ;
  assign n21729 = ~n20965 & ~n20969 ;
  assign n21730 = n21728 & n21729 ;
  assign n21731 = ~n21728 & ~n21729 ;
  assign n21732 = ~n21730 & ~n21731 ;
  assign n21733 = x91 & n6725 ;
  assign n21734 = x89 & n7129 ;
  assign n21735 = x90 & n6720 ;
  assign n21736 = ~n21734 & ~n21735 ;
  assign n21737 = ~n21733 & n21736 ;
  assign n21738 = n5336 & n6728 ;
  assign n21739 = n21737 & ~n21738 ;
  assign n21740 = x32 & ~n21739 ;
  assign n21741 = x32 & ~n21740 ;
  assign n21742 = ~n21739 & ~n21740 ;
  assign n21743 = ~n21741 & ~n21742 ;
  assign n21744 = ~n21732 & n21743 ;
  assign n21745 = n21732 & ~n21743 ;
  assign n21746 = ~n21744 & ~n21745 ;
  assign n21747 = ~n20987 & n21746 ;
  assign n21748 = n20987 & ~n21746 ;
  assign n21749 = ~n21747 & ~n21748 ;
  assign n21750 = ~n21581 & n21749 ;
  assign n21751 = n21581 & ~n21749 ;
  assign n21752 = ~n21750 & ~n21751 ;
  assign n21753 = ~n21570 & n21752 ;
  assign n21754 = n21570 & ~n21752 ;
  assign n21755 = ~n21753 & ~n21754 ;
  assign n21756 = x97 & n4531 ;
  assign n21757 = x95 & n4847 ;
  assign n21758 = x96 & n4526 ;
  assign n21759 = ~n21757 & ~n21758 ;
  assign n21760 = ~n21756 & n21759 ;
  assign n21761 = n4534 & n7745 ;
  assign n21762 = n21760 & ~n21761 ;
  assign n21763 = x26 & ~n21762 ;
  assign n21764 = x26 & ~n21763 ;
  assign n21765 = ~n21762 & ~n21763 ;
  assign n21766 = ~n21764 & ~n21765 ;
  assign n21767 = n21755 & ~n21766 ;
  assign n21768 = n21755 & ~n21767 ;
  assign n21769 = ~n21766 & ~n21767 ;
  assign n21770 = ~n21768 & ~n21769 ;
  assign n21771 = ~n21569 & n21770 ;
  assign n21772 = n21569 & ~n21770 ;
  assign n21773 = ~n21771 & ~n21772 ;
  assign n21774 = x100 & n3589 ;
  assign n21775 = x98 & n3878 ;
  assign n21776 = x99 & n3584 ;
  assign n21777 = ~n21775 & ~n21776 ;
  assign n21778 = ~n21774 & n21777 ;
  assign n21779 = n3592 & n9115 ;
  assign n21780 = n21778 & ~n21779 ;
  assign n21781 = x23 & ~n21780 ;
  assign n21782 = x23 & ~n21781 ;
  assign n21783 = ~n21780 & ~n21781 ;
  assign n21784 = ~n21782 & ~n21783 ;
  assign n21785 = ~n21773 & ~n21784 ;
  assign n21786 = n21773 & n21784 ;
  assign n21787 = ~n21785 & ~n21786 ;
  assign n21788 = n21568 & ~n21787 ;
  assign n21789 = ~n21568 & n21787 ;
  assign n21790 = ~n21788 & ~n21789 ;
  assign n21791 = x103 & n2751 ;
  assign n21792 = x101 & n3020 ;
  assign n21793 = x102 & n2746 ;
  assign n21794 = ~n21792 & ~n21793 ;
  assign n21795 = ~n21791 & n21794 ;
  assign n21796 = n2754 & n10588 ;
  assign n21797 = n21795 & ~n21796 ;
  assign n21798 = x20 & ~n21797 ;
  assign n21799 = x20 & ~n21798 ;
  assign n21800 = ~n21797 & ~n21798 ;
  assign n21801 = ~n21799 & ~n21800 ;
  assign n21802 = n21790 & ~n21801 ;
  assign n21803 = n21790 & ~n21802 ;
  assign n21804 = ~n21801 & ~n21802 ;
  assign n21805 = ~n21803 & ~n21804 ;
  assign n21806 = ~n21043 & ~n21049 ;
  assign n21807 = n21805 & n21806 ;
  assign n21808 = ~n21805 & ~n21806 ;
  assign n21809 = ~n21807 & ~n21808 ;
  assign n21810 = x106 & n2093 ;
  assign n21811 = x104 & n2275 ;
  assign n21812 = x105 & n2088 ;
  assign n21813 = ~n21811 & ~n21812 ;
  assign n21814 = ~n21810 & n21813 ;
  assign n21815 = n2096 & n12181 ;
  assign n21816 = n21814 & ~n21815 ;
  assign n21817 = x17 & ~n21816 ;
  assign n21818 = x17 & ~n21817 ;
  assign n21819 = ~n21816 & ~n21817 ;
  assign n21820 = ~n21818 & ~n21819 ;
  assign n21821 = ~n21809 & n21820 ;
  assign n21822 = n21809 & ~n21820 ;
  assign n21823 = ~n21821 & ~n21822 ;
  assign n21824 = ~n21567 & n21823 ;
  assign n21825 = n21567 & ~n21823 ;
  assign n21826 = ~n21824 & ~n21825 ;
  assign n21827 = ~n21566 & n21826 ;
  assign n21828 = ~n21566 & ~n21827 ;
  assign n21829 = n21826 & ~n21827 ;
  assign n21830 = ~n21828 & ~n21829 ;
  assign n21831 = ~n21086 & ~n21830 ;
  assign n21832 = n21086 & ~n21829 ;
  assign n21833 = ~n21828 & n21832 ;
  assign n21834 = ~n21831 & ~n21833 ;
  assign n21835 = ~n21555 & n21834 ;
  assign n21836 = ~n21555 & ~n21835 ;
  assign n21837 = n21834 & ~n21835 ;
  assign n21838 = ~n21836 & ~n21837 ;
  assign n21839 = ~n21544 & ~n21838 ;
  assign n21840 = n21544 & ~n21837 ;
  assign n21841 = ~n21836 & n21840 ;
  assign n21842 = ~n21839 & ~n21841 ;
  assign n21843 = ~n21543 & n21842 ;
  assign n21844 = ~n21543 & ~n21843 ;
  assign n21845 = n21842 & ~n21843 ;
  assign n21846 = ~n21844 & ~n21845 ;
  assign n21847 = ~n21532 & ~n21846 ;
  assign n21848 = n21532 & ~n21845 ;
  assign n21849 = ~n21844 & n21848 ;
  assign n21850 = ~n21847 & ~n21849 ;
  assign n21851 = ~n21531 & n21850 ;
  assign n21852 = ~n21531 & ~n21851 ;
  assign n21853 = n21850 & ~n21851 ;
  assign n21854 = ~n21852 & ~n21853 ;
  assign n21855 = ~n21520 & ~n21854 ;
  assign n21856 = ~n21520 & ~n21855 ;
  assign n21857 = ~n21854 & ~n21855 ;
  assign n21858 = ~n21856 & ~n21857 ;
  assign n21859 = x121 & n146 ;
  assign n21860 = x119 & n182 ;
  assign n21861 = x120 & n141 ;
  assign n21862 = ~n21860 & ~n21861 ;
  assign n21863 = ~n21859 & n21862 ;
  assign n21864 = ~n21139 & ~n21141 ;
  assign n21865 = ~x120 & ~x121 ;
  assign n21866 = x120 & x121 ;
  assign n21867 = ~n21865 & ~n21866 ;
  assign n21868 = ~n21864 & n21867 ;
  assign n21869 = n21864 & ~n21867 ;
  assign n21870 = ~n21868 & ~n21869 ;
  assign n21871 = n149 & n21870 ;
  assign n21872 = n21863 & ~n21871 ;
  assign n21873 = x2 & ~n21872 ;
  assign n21874 = x2 & ~n21873 ;
  assign n21875 = ~n21872 & ~n21873 ;
  assign n21876 = ~n21874 & ~n21875 ;
  assign n21877 = ~n21858 & ~n21876 ;
  assign n21878 = ~n21858 & ~n21877 ;
  assign n21879 = ~n21876 & ~n21877 ;
  assign n21880 = ~n21878 & ~n21879 ;
  assign n21881 = ~n21150 & ~n21155 ;
  assign n21882 = ~n21880 & ~n21881 ;
  assign n21883 = n21880 & n21881 ;
  assign n21884 = ~n21882 & ~n21883 ;
  assign n22245 = n21884 & x185 ;
  assign n21885 = ~n21488 & ~n21490 ;
  assign n21886 = ~x118 & n293 ;
  assign n21887 = ~x116 & n373 ;
  assign n21888 = ~x117 & n288 ;
  assign n21889 = ~n21887 & ~n21888 ;
  assign n21890 = ~n21886 & n21889 ;
  assign n21891 = n296 & n19736 ;
  assign n21892 = n21890 & ~n21891 ;
  assign n21893 = ~x5 & ~n21892 ;
  assign n21894 = ~x5 & ~n21893 ;
  assign n21895 = ~n21892 & ~n21893 ;
  assign n21896 = ~n21894 & ~n21895 ;
  assign n21897 = ~n21468 & ~n21472 ;
  assign n21898 = ~x115 & n574 ;
  assign n21899 = ~x113 & n673 ;
  assign n21900 = ~x114 & n569 ;
  assign n21901 = ~n21899 & ~n21900 ;
  assign n21902 = ~n21898 & n21901 ;
  assign n21903 = n577 & n17683 ;
  assign n21904 = n21902 & ~n21903 ;
  assign n21905 = ~x8 & ~n21904 ;
  assign n21906 = ~x8 & ~n21905 ;
  assign n21907 = ~n21904 & ~n21905 ;
  assign n21908 = ~n21906 & ~n21907 ;
  assign n21909 = ~n21461 & ~n21465 ;
  assign n21910 = ~x112 & n945 ;
  assign n21911 = ~x110 & n1099 ;
  assign n21912 = ~x111 & n940 ;
  assign n21913 = ~n21911 & ~n21912 ;
  assign n21914 = ~n21910 & n21913 ;
  assign n21915 = n948 & n15744 ;
  assign n21916 = n21914 & ~n21915 ;
  assign n21917 = ~x11 & ~n21916 ;
  assign n21918 = ~x11 & ~n21917 ;
  assign n21919 = ~n21916 & ~n21917 ;
  assign n21920 = ~n21918 & ~n21919 ;
  assign n21921 = ~x109 & n1434 ;
  assign n21922 = ~x107 & n1646 ;
  assign n21923 = ~x108 & n1429 ;
  assign n21924 = ~n21922 & ~n21923 ;
  assign n21925 = ~n21921 & n21924 ;
  assign n21926 = n1437 & n14177 ;
  assign n21927 = n21925 & ~n21926 ;
  assign n21928 = ~x14 & ~n21927 ;
  assign n21929 = ~x14 & ~n21928 ;
  assign n21930 = ~n21927 & ~n21928 ;
  assign n21931 = ~n21929 & ~n21930 ;
  assign n21932 = ~n21423 & ~n21429 ;
  assign n21933 = ~n21385 & ~n21391 ;
  assign n21934 = ~n21369 & ~n21371 ;
  assign n21935 = ~n21363 & ~n21365 ;
  assign n21936 = ~x94 & n5560 ;
  assign n21937 = ~x92 & n5943 ;
  assign n21938 = ~x93 & n5555 ;
  assign n21939 = ~n21937 & ~n21938 ;
  assign n21940 = ~n21936 & n21939 ;
  assign n21941 = n5563 & n6671 ;
  assign n21942 = n21940 & ~n21941 ;
  assign n21943 = ~x29 & ~n21942 ;
  assign n21944 = ~x29 & ~n21943 ;
  assign n21945 = ~n21942 & ~n21943 ;
  assign n21946 = ~n21944 & ~n21945 ;
  assign n21947 = ~n20573 & ~n21311 ;
  assign n21948 = ~n21308 & ~n21947 ;
  assign n21949 = ~x85 & n9433 ;
  assign n21950 = ~x83 & n9915 ;
  assign n21951 = ~x84 & n9428 ;
  assign n21952 = ~n21950 & ~n21951 ;
  assign n21953 = ~n21949 & n21952 ;
  assign n21954 = n3521 & n9436 ;
  assign n21955 = n21953 & ~n21954 ;
  assign n21956 = ~x38 & ~n21955 ;
  assign n21957 = ~x38 & ~n21956 ;
  assign n21958 = ~n21955 & ~n21956 ;
  assign n21959 = ~n21957 & ~n21958 ;
  assign n21960 = ~n21289 & ~n21293 ;
  assign n21961 = ~x82 & n10905 ;
  assign n21962 = ~x80 & n11466 ;
  assign n21963 = ~x81 & n10900 ;
  assign n21964 = ~n21962 & ~n21963 ;
  assign n21965 = ~n21961 & n21964 ;
  assign n21966 = n2697 & n10908 ;
  assign n21967 = n21965 & ~n21966 ;
  assign n21968 = ~x41 & ~n21967 ;
  assign n21969 = ~x41 & ~n21968 ;
  assign n21970 = ~n21967 & ~n21968 ;
  assign n21971 = ~n21969 & ~n21970 ;
  assign n21972 = ~n21282 & ~n21286 ;
  assign n21973 = ~x79 & n12506 ;
  assign n21974 = ~x77 & n13131 ;
  assign n21975 = ~x78 & n12501 ;
  assign n21976 = ~n21974 & ~n21975 ;
  assign n21977 = ~n21973 & n21976 ;
  assign n21978 = n1921 & n12509 ;
  assign n21979 = n21977 & ~n21978 ;
  assign n21980 = ~x44 & ~n21979 ;
  assign n21981 = ~x44 & ~n21980 ;
  assign n21982 = ~n21979 & ~n21980 ;
  assign n21983 = ~n21981 & ~n21982 ;
  assign n21984 = ~n21266 & ~n21268 ;
  assign n21985 = ~x76 & n14233 ;
  assign n21986 = ~x74 & n14876 ;
  assign n21987 = ~x75 & n14228 ;
  assign n21988 = ~n21986 & ~n21987 ;
  assign n21989 = ~n21985 & n21988 ;
  assign n21990 = n1390 & n14236 ;
  assign n21991 = n21989 & ~n21990 ;
  assign n21992 = ~x47 & ~n21991 ;
  assign n21993 = ~x47 & ~n21992 ;
  assign n21994 = ~n21991 & ~n21992 ;
  assign n21995 = ~n21993 & ~n21994 ;
  assign n21996 = ~n21260 & ~n21262 ;
  assign n21997 = ~x64 & ~n21634 ;
  assign n21998 = ~n21227 & n21997 ;
  assign n21999 = n21227 & ~n21997 ;
  assign n22000 = ~n21998 & ~n21999 ;
  assign n22001 = ~x67 & n20143 ;
  assign n22002 = ~x65 & n20854 ;
  assign n22003 = ~x66 & n20138 ;
  assign n22004 = ~n22002 & ~n22003 ;
  assign n22005 = ~n22001 & n22004 ;
  assign n22006 = n266 & n20146 ;
  assign n22007 = n22005 & ~n22006 ;
  assign n22008 = ~x56 & ~n22007 ;
  assign n22009 = ~x56 & ~n22008 ;
  assign n22010 = ~n22007 & ~n22008 ;
  assign n22011 = ~n22009 & ~n22010 ;
  assign n22012 = ~n22000 & ~n22011 ;
  assign n22013 = n22000 & n22011 ;
  assign n22014 = ~n22012 & ~n22013 ;
  assign n22015 = ~x70 & n18025 ;
  assign n22016 = ~x68 & n18764 ;
  assign n22017 = ~x69 & n18020 ;
  assign n22018 = ~n22016 & ~n22017 ;
  assign n22019 = ~n22015 & n22018 ;
  assign n22020 = n529 & n18028 ;
  assign n22021 = n22019 & ~n22020 ;
  assign n22022 = ~x53 & ~n22021 ;
  assign n22023 = ~x53 & ~n22022 ;
  assign n22024 = ~n22021 & ~n22022 ;
  assign n22025 = ~n22023 & ~n22024 ;
  assign n22026 = n22014 & ~n22025 ;
  assign n22027 = n22014 & ~n22026 ;
  assign n22028 = ~n22025 & ~n22026 ;
  assign n22029 = ~n22027 & ~n22028 ;
  assign n22030 = ~n21245 & n22029 ;
  assign n22031 = n21245 & ~n22029 ;
  assign n22032 = ~n22030 & ~n22031 ;
  assign n22033 = ~x73 & n16076 ;
  assign n22034 = ~x71 & n16756 ;
  assign n22035 = ~x72 & n16071 ;
  assign n22036 = ~n22034 & ~n22035 ;
  assign n22037 = ~n22033 & n22036 ;
  assign n22038 = n903 & n16079 ;
  assign n22039 = n22037 & ~n22038 ;
  assign n22040 = ~x50 & ~n22039 ;
  assign n22041 = ~x50 & ~n22040 ;
  assign n22042 = ~n22039 & ~n22040 ;
  assign n22043 = ~n22041 & ~n22042 ;
  assign n22044 = ~n22032 & ~n22043 ;
  assign n22045 = n22032 & n22043 ;
  assign n22046 = ~n22044 & ~n22045 ;
  assign n22047 = ~n21996 & n22046 ;
  assign n22048 = n21996 & ~n22046 ;
  assign n22049 = ~n22047 & ~n22048 ;
  assign n22050 = n21995 & ~n22049 ;
  assign n22051 = ~n21995 & n22049 ;
  assign n22052 = ~n22050 & ~n22051 ;
  assign n22053 = ~n21984 & n22052 ;
  assign n22054 = n21984 & ~n22052 ;
  assign n22055 = ~n22053 & ~n22054 ;
  assign n22056 = ~n21983 & n22055 ;
  assign n22057 = n21983 & ~n22055 ;
  assign n22058 = ~n22056 & ~n22057 ;
  assign n22059 = ~n21972 & n22058 ;
  assign n22060 = n21972 & ~n22058 ;
  assign n22061 = ~n22059 & ~n22060 ;
  assign n22062 = ~n21971 & n22061 ;
  assign n22063 = ~n21971 & ~n22062 ;
  assign n22064 = n22061 & ~n22062 ;
  assign n22065 = ~n22063 & ~n22064 ;
  assign n22066 = ~n21960 & ~n22065 ;
  assign n22067 = n21960 & ~n22064 ;
  assign n22068 = ~n22063 & n22067 ;
  assign n22069 = ~n22066 & ~n22068 ;
  assign n22070 = ~n21959 & n22069 ;
  assign n22071 = n21959 & ~n22069 ;
  assign n22072 = ~n22070 & ~n22071 ;
  assign n22073 = ~n21948 & n22072 ;
  assign n22074 = n21948 & ~n22072 ;
  assign n22075 = ~n22073 & ~n22074 ;
  assign n22076 = ~x88 & n8006 ;
  assign n22077 = ~x86 & n8474 ;
  assign n22078 = ~x87 & n8001 ;
  assign n22079 = ~n22077 & ~n22078 ;
  assign n22080 = ~n22076 & n22079 ;
  assign n22081 = n4457 & n8009 ;
  assign n22082 = n22080 & ~n22081 ;
  assign n22083 = ~x35 & ~n22082 ;
  assign n22084 = ~x35 & ~n22083 ;
  assign n22085 = ~n22082 & ~n22083 ;
  assign n22086 = ~n22084 & ~n22085 ;
  assign n22087 = n22075 & ~n22086 ;
  assign n22088 = n22075 & ~n22087 ;
  assign n22089 = ~n22086 & ~n22087 ;
  assign n22090 = ~n22088 & ~n22089 ;
  assign n22091 = ~n21326 & ~n21330 ;
  assign n22092 = n22090 & n22091 ;
  assign n22093 = ~n22090 & ~n22091 ;
  assign n22094 = ~n22092 & ~n22093 ;
  assign n22095 = ~x91 & n6725 ;
  assign n22096 = ~x89 & n7129 ;
  assign n22097 = ~x90 & n6720 ;
  assign n22098 = ~n22096 & ~n22097 ;
  assign n22099 = ~n22095 & n22098 ;
  assign n22100 = n5507 & n6728 ;
  assign n22101 = n22099 & ~n22100 ;
  assign n22102 = ~x32 & ~n22101 ;
  assign n22103 = ~x32 & ~n22102 ;
  assign n22104 = ~n22101 & ~n22102 ;
  assign n22105 = ~n22103 & ~n22104 ;
  assign n22106 = ~n22094 & n22105 ;
  assign n22107 = n22094 & ~n22105 ;
  assign n22108 = ~n22106 & ~n22107 ;
  assign n22109 = ~n21348 & n22108 ;
  assign n22110 = n21348 & ~n22108 ;
  assign n22111 = ~n22109 & ~n22110 ;
  assign n22112 = ~n21946 & n22111 ;
  assign n22113 = n21946 & ~n22111 ;
  assign n22114 = ~n22112 & ~n22113 ;
  assign n22115 = ~n21935 & n22114 ;
  assign n22116 = n21935 & ~n22114 ;
  assign n22117 = ~n22115 & ~n22116 ;
  assign n22118 = ~x97 & n4531 ;
  assign n22119 = ~x95 & n4847 ;
  assign n22120 = ~x96 & n4526 ;
  assign n22121 = ~n22119 & ~n22120 ;
  assign n22122 = ~n22118 & n22121 ;
  assign n22123 = n4534 & n7949 ;
  assign n22124 = n22122 & ~n22123 ;
  assign n22125 = ~x26 & ~n22124 ;
  assign n22126 = ~x26 & ~n22125 ;
  assign n22127 = ~n22124 & ~n22125 ;
  assign n22128 = ~n22126 & ~n22127 ;
  assign n22129 = n22117 & ~n22128 ;
  assign n22130 = n22117 & ~n22129 ;
  assign n22131 = ~n22128 & ~n22129 ;
  assign n22132 = ~n22130 & ~n22131 ;
  assign n22133 = ~n21934 & n22132 ;
  assign n22134 = n21934 & ~n22132 ;
  assign n22135 = ~n22133 & ~n22134 ;
  assign n22136 = ~x100 & n3589 ;
  assign n22137 = ~x98 & n3878 ;
  assign n22138 = ~x99 & n3584 ;
  assign n22139 = ~n22137 & ~n22138 ;
  assign n22140 = ~n22136 & n22139 ;
  assign n22141 = n3592 & n9338 ;
  assign n22142 = n22140 & ~n22141 ;
  assign n22143 = ~x23 & ~n22142 ;
  assign n22144 = ~x23 & ~n22143 ;
  assign n22145 = ~n22142 & ~n22143 ;
  assign n22146 = ~n22144 & ~n22145 ;
  assign n22147 = ~n22135 & ~n22146 ;
  assign n22148 = n22135 & n22146 ;
  assign n22149 = ~n22147 & ~n22148 ;
  assign n22150 = n21933 & ~n22149 ;
  assign n22151 = ~n21933 & n22149 ;
  assign n22152 = ~n22150 & ~n22151 ;
  assign n22153 = ~x103 & n2751 ;
  assign n22154 = ~x101 & n3020 ;
  assign n22155 = ~x102 & n2746 ;
  assign n22156 = ~n22154 & ~n22155 ;
  assign n22157 = ~n22153 & n22156 ;
  assign n22158 = n2754 & n10833 ;
  assign n22159 = n22157 & ~n22158 ;
  assign n22160 = ~x20 & ~n22159 ;
  assign n22161 = ~x20 & ~n22160 ;
  assign n22162 = ~n22159 & ~n22160 ;
  assign n22163 = ~n22161 & ~n22162 ;
  assign n22164 = n22152 & ~n22163 ;
  assign n22165 = n22152 & ~n22164 ;
  assign n22166 = ~n22163 & ~n22164 ;
  assign n22167 = ~n22165 & ~n22166 ;
  assign n22168 = ~n21404 & ~n21410 ;
  assign n22169 = n22167 & n22168 ;
  assign n22170 = ~n22167 & ~n22168 ;
  assign n22171 = ~n22169 & ~n22170 ;
  assign n22172 = ~x106 & n2093 ;
  assign n22173 = ~x104 & n2275 ;
  assign n22174 = ~x105 & n2088 ;
  assign n22175 = ~n22173 & ~n22174 ;
  assign n22176 = ~n22172 & n22175 ;
  assign n22177 = n2096 & n12447 ;
  assign n22178 = n22176 & ~n22177 ;
  assign n22179 = ~x17 & ~n22178 ;
  assign n22180 = ~x17 & ~n22179 ;
  assign n22181 = ~n22178 & ~n22179 ;
  assign n22182 = ~n22180 & ~n22181 ;
  assign n22183 = ~n22171 & n22182 ;
  assign n22184 = n22171 & ~n22182 ;
  assign n22185 = ~n22183 & ~n22184 ;
  assign n22186 = ~n21932 & n22185 ;
  assign n22187 = n21932 & ~n22185 ;
  assign n22188 = ~n22186 & ~n22187 ;
  assign n22189 = ~n21931 & n22188 ;
  assign n22190 = ~n21931 & ~n22189 ;
  assign n22191 = n22188 & ~n22189 ;
  assign n22192 = ~n22190 & ~n22191 ;
  assign n22193 = ~n21447 & ~n22192 ;
  assign n22194 = n21447 & ~n22191 ;
  assign n22195 = ~n22190 & n22194 ;
  assign n22196 = ~n22193 & ~n22195 ;
  assign n22197 = ~n21920 & n22196 ;
  assign n22198 = ~n21920 & ~n22197 ;
  assign n22199 = n22196 & ~n22197 ;
  assign n22200 = ~n22198 & ~n22199 ;
  assign n22201 = ~n21909 & ~n22200 ;
  assign n22202 = n21909 & ~n22199 ;
  assign n22203 = ~n22198 & n22202 ;
  assign n22204 = ~n22201 & ~n22203 ;
  assign n22205 = ~n21908 & n22204 ;
  assign n22206 = ~n21908 & ~n22205 ;
  assign n22207 = n22204 & ~n22205 ;
  assign n22208 = ~n22206 & ~n22207 ;
  assign n22209 = ~n21897 & ~n22208 ;
  assign n22210 = n21897 & ~n22207 ;
  assign n22211 = ~n22206 & n22210 ;
  assign n22212 = ~n22209 & ~n22211 ;
  assign n22213 = ~n21896 & n22212 ;
  assign n22214 = ~n21896 & ~n22213 ;
  assign n22215 = n22212 & ~n22213 ;
  assign n22216 = ~n22214 & ~n22215 ;
  assign n22217 = ~n21885 & ~n22216 ;
  assign n22218 = ~n21885 & ~n22217 ;
  assign n22219 = ~n22216 & ~n22217 ;
  assign n22220 = ~n22218 & ~n22219 ;
  assign n22221 = ~x121 & n164 ;
  assign n22222 = ~x119 & n205 ;
  assign n22223 = ~x120 & n162 ;
  assign n22224 = ~n22222 & ~n22223 ;
  assign n22225 = ~n22221 & n22224 ;
  assign n22226 = ~n21138 & ~n21499 ;
  assign n22227 = n21867 & ~n22226 ;
  assign n22228 = ~n21867 & n22226 ;
  assign n22229 = ~n22227 & ~n22228 ;
  assign n22230 = n167 & n22229 ;
  assign n22231 = n22225 & ~n22230 ;
  assign n22232 = ~x2 & ~n22231 ;
  assign n22233 = ~x2 & ~n22232 ;
  assign n22234 = ~n22231 & ~n22232 ;
  assign n22235 = ~n22233 & ~n22234 ;
  assign n22236 = ~n22220 & ~n22235 ;
  assign n22237 = ~n22220 & ~n22236 ;
  assign n22238 = ~n22235 & ~n22236 ;
  assign n22239 = ~n22237 & ~n22238 ;
  assign n22240 = ~n21508 & ~n21513 ;
  assign n22241 = ~n22239 & ~n22240 ;
  assign n22242 = n22239 & n22240 ;
  assign n22243 = ~n22241 & ~n22242 ;
  assign n22246 = ~n22243 & ~x185 ;
  assign n22247 = ~n22245 & ~n22246 ;
  assign n22248 = ~n21851 & ~n21855 ;
  assign n22249 = x119 & n293 ;
  assign n22250 = x117 & n373 ;
  assign n22251 = x118 & n288 ;
  assign n22252 = ~n22250 & ~n22251 ;
  assign n22253 = ~n22249 & n22252 ;
  assign n22254 = n296 & n20423 ;
  assign n22255 = n22253 & ~n22254 ;
  assign n22256 = x5 & ~n22255 ;
  assign n22257 = x5 & ~n22256 ;
  assign n22258 = ~n22255 & ~n22256 ;
  assign n22259 = ~n22257 & ~n22258 ;
  assign n22260 = ~n21843 & ~n21847 ;
  assign n22261 = x116 & n574 ;
  assign n22262 = x114 & n673 ;
  assign n22263 = x115 & n569 ;
  assign n22264 = ~n22262 & ~n22263 ;
  assign n22265 = ~n22261 & n22264 ;
  assign n22266 = n577 & n18336 ;
  assign n22267 = n22265 & ~n22266 ;
  assign n22268 = x8 & ~n22267 ;
  assign n22269 = x8 & ~n22268 ;
  assign n22270 = ~n22267 & ~n22268 ;
  assign n22271 = ~n22269 & ~n22270 ;
  assign n22272 = ~n21835 & ~n21839 ;
  assign n22273 = x113 & n945 ;
  assign n22274 = x111 & n1099 ;
  assign n22275 = x112 & n940 ;
  assign n22276 = ~n22274 & ~n22275 ;
  assign n22277 = ~n22273 & n22276 ;
  assign n22278 = n948 & n16361 ;
  assign n22279 = n22277 & ~n22278 ;
  assign n22280 = x11 & ~n22279 ;
  assign n22281 = x11 & ~n22280 ;
  assign n22282 = ~n22279 & ~n22280 ;
  assign n22283 = ~n22281 & ~n22282 ;
  assign n22284 = ~n21827 & ~n21831 ;
  assign n22285 = ~n21822 & ~n21824 ;
  assign n22286 = ~n21750 & ~n21753 ;
  assign n22287 = ~n21745 & ~n21747 ;
  assign n22288 = ~n21700 & ~n21704 ;
  assign n22289 = ~n21689 & ~n21691 ;
  assign n22290 = ~n20884 & ~n21667 ;
  assign n22291 = ~n21664 & ~n22290 ;
  assign n22292 = x71 & n18025 ;
  assign n22293 = x69 & n18764 ;
  assign n22294 = x70 & n18020 ;
  assign n22295 = ~n22293 & ~n22294 ;
  assign n22296 = ~n22292 & n22295 ;
  assign n22297 = n558 & n18028 ;
  assign n22298 = n22296 & ~n22297 ;
  assign n22299 = x53 & ~n22298 ;
  assign n22300 = x53 & ~n22299 ;
  assign n22301 = ~n22298 & ~n22299 ;
  assign n22302 = ~n22300 & ~n22301 ;
  assign n22303 = n20866 & n21635 ;
  assign n22304 = ~n21650 & ~n22303 ;
  assign n22305 = x68 & n20143 ;
  assign n22306 = x66 & n20854 ;
  assign n22307 = x67 & n20138 ;
  assign n22308 = ~n22306 & ~n22307 ;
  assign n22309 = ~n22305 & n22308 ;
  assign n22310 = n317 & n20146 ;
  assign n22311 = n22309 & ~n22310 ;
  assign n22312 = x56 & ~n22311 ;
  assign n22313 = x56 & ~n22312 ;
  assign n22314 = ~n22311 & ~n22312 ;
  assign n22315 = ~n22313 & ~n22314 ;
  assign n22316 = x59 & ~n21635 ;
  assign n22317 = ~x57 & x58 ;
  assign n22318 = x57 & ~x58 ;
  assign n22319 = ~n22317 & ~n22318 ;
  assign n22320 = n21634 & ~n22319 ;
  assign n22321 = x64 & n22320 ;
  assign n22322 = ~x58 & x59 ;
  assign n22323 = x58 & ~x59 ;
  assign n22324 = ~n22322 & ~n22323 ;
  assign n22325 = ~n21634 & n22324 ;
  assign n22326 = x65 & n22325 ;
  assign n22327 = ~n22321 & ~n22326 ;
  assign n22328 = ~n21634 & ~n22324 ;
  assign n22329 = ~n152 & n22328 ;
  assign n22330 = n22327 & ~n22329 ;
  assign n22331 = x59 & ~n22330 ;
  assign n22332 = x59 & ~n22331 ;
  assign n22333 = ~n22330 & ~n22331 ;
  assign n22334 = ~n22332 & ~n22333 ;
  assign n22335 = n22316 & ~n22334 ;
  assign n22336 = ~n22316 & n22334 ;
  assign n22337 = ~n22335 & ~n22336 ;
  assign n22338 = n22315 & ~n22337 ;
  assign n22339 = ~n22315 & n22337 ;
  assign n22340 = ~n22338 & ~n22339 ;
  assign n22341 = ~n22304 & n22340 ;
  assign n22342 = n22304 & ~n22340 ;
  assign n22343 = ~n22341 & ~n22342 ;
  assign n22344 = n22302 & ~n22343 ;
  assign n22345 = ~n22302 & n22343 ;
  assign n22346 = ~n22344 & ~n22345 ;
  assign n22347 = ~n22291 & n22346 ;
  assign n22348 = n22291 & ~n22346 ;
  assign n22349 = ~n22347 & ~n22348 ;
  assign n22350 = x74 & n16076 ;
  assign n22351 = x72 & n16756 ;
  assign n22352 = x73 & n16071 ;
  assign n22353 = ~n22351 & ~n22352 ;
  assign n22354 = ~n22350 & n22353 ;
  assign n22355 = n994 & n16079 ;
  assign n22356 = n22354 & ~n22355 ;
  assign n22357 = x50 & ~n22356 ;
  assign n22358 = x50 & ~n22357 ;
  assign n22359 = ~n22356 & ~n22357 ;
  assign n22360 = ~n22358 & ~n22359 ;
  assign n22361 = n22349 & ~n22360 ;
  assign n22362 = n22349 & ~n22361 ;
  assign n22363 = ~n22360 & ~n22361 ;
  assign n22364 = ~n22362 & ~n22363 ;
  assign n22365 = ~n21682 & ~n21685 ;
  assign n22366 = n22364 & n22365 ;
  assign n22367 = ~n22364 & ~n22365 ;
  assign n22368 = ~n22366 & ~n22367 ;
  assign n22369 = x77 & n14233 ;
  assign n22370 = x75 & n14876 ;
  assign n22371 = x76 & n14228 ;
  assign n22372 = ~n22370 & ~n22371 ;
  assign n22373 = ~n22369 & n22372 ;
  assign n22374 = n1502 & n14236 ;
  assign n22375 = n22373 & ~n22374 ;
  assign n22376 = x47 & ~n22375 ;
  assign n22377 = x47 & ~n22376 ;
  assign n22378 = ~n22375 & ~n22376 ;
  assign n22379 = ~n22377 & ~n22378 ;
  assign n22380 = n22368 & ~n22379 ;
  assign n22381 = ~n22368 & n22379 ;
  assign n22382 = ~n22289 & ~n22381 ;
  assign n22383 = ~n22380 & n22382 ;
  assign n22384 = ~n22289 & ~n22383 ;
  assign n22385 = ~n22380 & ~n22383 ;
  assign n22386 = ~n22381 & n22385 ;
  assign n22387 = ~n22384 & ~n22386 ;
  assign n22388 = x80 & n12506 ;
  assign n22389 = x78 & n13131 ;
  assign n22390 = x79 & n12501 ;
  assign n22391 = ~n22389 & ~n22390 ;
  assign n22392 = ~n22388 & n22391 ;
  assign n22393 = n2028 & n12509 ;
  assign n22394 = n22392 & ~n22393 ;
  assign n22395 = x44 & ~n22394 ;
  assign n22396 = x44 & ~n22395 ;
  assign n22397 = ~n22394 & ~n22395 ;
  assign n22398 = ~n22396 & ~n22397 ;
  assign n22399 = ~n22387 & ~n22398 ;
  assign n22400 = ~n22387 & ~n22399 ;
  assign n22401 = ~n22398 & ~n22399 ;
  assign n22402 = ~n22400 & ~n22401 ;
  assign n22403 = ~n21694 & ~n21697 ;
  assign n22404 = n22402 & n22403 ;
  assign n22405 = ~n22402 & ~n22403 ;
  assign n22406 = ~n22404 & ~n22405 ;
  assign n22407 = x83 & n10905 ;
  assign n22408 = x81 & n11466 ;
  assign n22409 = x82 & n10900 ;
  assign n22410 = ~n22408 & ~n22409 ;
  assign n22411 = ~n22407 & n22410 ;
  assign n22412 = n2843 & n10908 ;
  assign n22413 = n22411 & ~n22412 ;
  assign n22414 = x41 & ~n22413 ;
  assign n22415 = x41 & ~n22414 ;
  assign n22416 = ~n22413 & ~n22414 ;
  assign n22417 = ~n22415 & ~n22416 ;
  assign n22418 = n22406 & ~n22417 ;
  assign n22419 = ~n22406 & n22417 ;
  assign n22420 = ~n22288 & ~n22419 ;
  assign n22421 = ~n22418 & n22420 ;
  assign n22422 = ~n22288 & ~n22421 ;
  assign n22423 = ~n22418 & ~n22421 ;
  assign n22424 = ~n22419 & n22423 ;
  assign n22425 = ~n22422 & ~n22424 ;
  assign n22426 = x86 & n9433 ;
  assign n22427 = x84 & n9915 ;
  assign n22428 = x85 & n9428 ;
  assign n22429 = ~n22427 & ~n22428 ;
  assign n22430 = ~n22426 & n22429 ;
  assign n22431 = n3686 & n9436 ;
  assign n22432 = n22430 & ~n22431 ;
  assign n22433 = x38 & ~n22432 ;
  assign n22434 = x38 & ~n22433 ;
  assign n22435 = ~n22432 & ~n22433 ;
  assign n22436 = ~n22434 & ~n22435 ;
  assign n22437 = ~n22425 & ~n22436 ;
  assign n22438 = ~n22425 & ~n22437 ;
  assign n22439 = ~n22436 & ~n22437 ;
  assign n22440 = ~n22438 & ~n22439 ;
  assign n22441 = ~n21708 & ~n21711 ;
  assign n22442 = n22440 & n22441 ;
  assign n22443 = ~n22440 & ~n22441 ;
  assign n22444 = ~n22442 & ~n22443 ;
  assign n22445 = x89 & n8006 ;
  assign n22446 = x87 & n8474 ;
  assign n22447 = x88 & n8001 ;
  assign n22448 = ~n22446 & ~n22447 ;
  assign n22449 = ~n22445 & n22448 ;
  assign n22450 = n4488 & n8009 ;
  assign n22451 = n22449 & ~n22450 ;
  assign n22452 = x35 & ~n22451 ;
  assign n22453 = x35 & ~n22452 ;
  assign n22454 = ~n22451 & ~n22452 ;
  assign n22455 = ~n22453 & ~n22454 ;
  assign n22456 = n22444 & ~n22455 ;
  assign n22457 = n22444 & ~n22456 ;
  assign n22458 = ~n22455 & ~n22456 ;
  assign n22459 = ~n22457 & ~n22458 ;
  assign n22460 = ~n21725 & ~n21731 ;
  assign n22461 = n22459 & n22460 ;
  assign n22462 = ~n22459 & ~n22460 ;
  assign n22463 = ~n22461 & ~n22462 ;
  assign n22464 = x92 & n6725 ;
  assign n22465 = x90 & n7129 ;
  assign n22466 = x91 & n6720 ;
  assign n22467 = ~n22465 & ~n22466 ;
  assign n22468 = ~n22464 & n22467 ;
  assign n22469 = n5710 & n6728 ;
  assign n22470 = n22468 & ~n22469 ;
  assign n22471 = x32 & ~n22470 ;
  assign n22472 = x32 & ~n22471 ;
  assign n22473 = ~n22470 & ~n22471 ;
  assign n22474 = ~n22472 & ~n22473 ;
  assign n22475 = n22463 & ~n22474 ;
  assign n22476 = n22463 & ~n22475 ;
  assign n22477 = ~n22474 & ~n22475 ;
  assign n22478 = ~n22476 & ~n22477 ;
  assign n22479 = ~n22287 & n22478 ;
  assign n22480 = n22287 & ~n22478 ;
  assign n22481 = ~n22479 & ~n22480 ;
  assign n22482 = x95 & n5560 ;
  assign n22483 = x93 & n5943 ;
  assign n22484 = x94 & n5555 ;
  assign n22485 = ~n22483 & ~n22484 ;
  assign n22486 = ~n22482 & n22485 ;
  assign n22487 = n5563 & n6894 ;
  assign n22488 = n22486 & ~n22487 ;
  assign n22489 = x29 & ~n22488 ;
  assign n22490 = x29 & ~n22489 ;
  assign n22491 = ~n22488 & ~n22489 ;
  assign n22492 = ~n22490 & ~n22491 ;
  assign n22493 = ~n22481 & ~n22492 ;
  assign n22494 = n22481 & n22492 ;
  assign n22495 = ~n22493 & ~n22494 ;
  assign n22496 = n22286 & ~n22495 ;
  assign n22497 = ~n22286 & n22495 ;
  assign n22498 = ~n22496 & ~n22497 ;
  assign n22499 = x98 & n4531 ;
  assign n22500 = x96 & n4847 ;
  assign n22501 = x97 & n4526 ;
  assign n22502 = ~n22500 & ~n22501 ;
  assign n22503 = ~n22499 & n22502 ;
  assign n22504 = n4534 & n8196 ;
  assign n22505 = n22503 & ~n22504 ;
  assign n22506 = x26 & ~n22505 ;
  assign n22507 = x26 & ~n22506 ;
  assign n22508 = ~n22505 & ~n22506 ;
  assign n22509 = ~n22507 & ~n22508 ;
  assign n22510 = n22498 & ~n22509 ;
  assign n22511 = n22498 & ~n22510 ;
  assign n22512 = ~n22509 & ~n22510 ;
  assign n22513 = ~n22511 & ~n22512 ;
  assign n22514 = ~n21569 & ~n21770 ;
  assign n22515 = ~n21767 & ~n22514 ;
  assign n22516 = n22513 & n22515 ;
  assign n22517 = ~n22513 & ~n22515 ;
  assign n22518 = ~n22516 & ~n22517 ;
  assign n22519 = x101 & n3589 ;
  assign n22520 = x99 & n3878 ;
  assign n22521 = x100 & n3584 ;
  assign n22522 = ~n22520 & ~n22521 ;
  assign n22523 = ~n22519 & n22522 ;
  assign n22524 = n3592 & n9601 ;
  assign n22525 = n22523 & ~n22524 ;
  assign n22526 = x23 & ~n22525 ;
  assign n22527 = x23 & ~n22526 ;
  assign n22528 = ~n22525 & ~n22526 ;
  assign n22529 = ~n22527 & ~n22528 ;
  assign n22530 = n22518 & ~n22529 ;
  assign n22531 = n22518 & ~n22530 ;
  assign n22532 = ~n22529 & ~n22530 ;
  assign n22533 = ~n22531 & ~n22532 ;
  assign n22534 = ~n21785 & ~n21789 ;
  assign n22535 = n22533 & n22534 ;
  assign n22536 = ~n22533 & ~n22534 ;
  assign n22537 = ~n22535 & ~n22536 ;
  assign n22538 = x104 & n2751 ;
  assign n22539 = x102 & n3020 ;
  assign n22540 = x103 & n2746 ;
  assign n22541 = ~n22539 & ~n22540 ;
  assign n22542 = ~n22538 & n22541 ;
  assign n22543 = n2754 & n11116 ;
  assign n22544 = n22542 & ~n22543 ;
  assign n22545 = x20 & ~n22544 ;
  assign n22546 = x20 & ~n22545 ;
  assign n22547 = ~n22544 & ~n22545 ;
  assign n22548 = ~n22546 & ~n22547 ;
  assign n22549 = n22537 & ~n22548 ;
  assign n22550 = n22537 & ~n22549 ;
  assign n22551 = ~n22548 & ~n22549 ;
  assign n22552 = ~n22550 & ~n22551 ;
  assign n22553 = ~n21802 & ~n21808 ;
  assign n22554 = n22552 & n22553 ;
  assign n22555 = ~n22552 & ~n22553 ;
  assign n22556 = ~n22554 & ~n22555 ;
  assign n22557 = x107 & n2093 ;
  assign n22558 = x105 & n2275 ;
  assign n22559 = x106 & n2088 ;
  assign n22560 = ~n22558 & ~n22559 ;
  assign n22561 = ~n22557 & n22560 ;
  assign n22562 = n2096 & n12749 ;
  assign n22563 = n22561 & ~n22562 ;
  assign n22564 = x17 & ~n22563 ;
  assign n22565 = x17 & ~n22564 ;
  assign n22566 = ~n22563 & ~n22564 ;
  assign n22567 = ~n22565 & ~n22566 ;
  assign n22568 = n22556 & ~n22567 ;
  assign n22569 = ~n22556 & n22567 ;
  assign n22570 = ~n22285 & ~n22569 ;
  assign n22571 = ~n22568 & n22570 ;
  assign n22572 = ~n22285 & ~n22571 ;
  assign n22573 = ~n22568 & ~n22571 ;
  assign n22574 = ~n22569 & n22573 ;
  assign n22575 = ~n22572 & ~n22574 ;
  assign n22576 = x110 & n1434 ;
  assign n22577 = x108 & n1646 ;
  assign n22578 = x109 & n1429 ;
  assign n22579 = ~n22577 & ~n22578 ;
  assign n22580 = ~n22576 & n22579 ;
  assign n22581 = n1437 & n14497 ;
  assign n22582 = n22580 & ~n22581 ;
  assign n22583 = x14 & ~n22582 ;
  assign n22584 = x14 & ~n22583 ;
  assign n22585 = ~n22582 & ~n22583 ;
  assign n22586 = ~n22584 & ~n22585 ;
  assign n22587 = n22575 & n22586 ;
  assign n22588 = ~n22575 & ~n22586 ;
  assign n22589 = ~n22587 & ~n22588 ;
  assign n22590 = ~n22284 & n22589 ;
  assign n22591 = n22284 & ~n22589 ;
  assign n22592 = ~n22590 & ~n22591 ;
  assign n22593 = n22283 & ~n22592 ;
  assign n22594 = ~n22283 & n22592 ;
  assign n22595 = ~n22593 & ~n22594 ;
  assign n22596 = ~n22272 & n22595 ;
  assign n22597 = n22272 & ~n22595 ;
  assign n22598 = ~n22596 & ~n22597 ;
  assign n22599 = n22271 & ~n22598 ;
  assign n22600 = ~n22271 & n22598 ;
  assign n22601 = ~n22599 & ~n22600 ;
  assign n22602 = ~n22260 & n22601 ;
  assign n22603 = n22260 & ~n22601 ;
  assign n22604 = ~n22602 & ~n22603 ;
  assign n22605 = n22259 & ~n22604 ;
  assign n22606 = ~n22259 & n22604 ;
  assign n22607 = ~n22605 & ~n22606 ;
  assign n22608 = ~n22248 & n22607 ;
  assign n22609 = n22248 & ~n22607 ;
  assign n22610 = ~n22608 & ~n22609 ;
  assign n22611 = x122 & n146 ;
  assign n22612 = x120 & n182 ;
  assign n22613 = x121 & n141 ;
  assign n22614 = ~n22612 & ~n22613 ;
  assign n22615 = ~n22611 & n22614 ;
  assign n22616 = ~n21866 & ~n21868 ;
  assign n22617 = ~x121 & ~x122 ;
  assign n22618 = x121 & x122 ;
  assign n22619 = ~n22617 & ~n22618 ;
  assign n22620 = ~n22616 & n22619 ;
  assign n22621 = n22616 & ~n22619 ;
  assign n22622 = ~n22620 & ~n22621 ;
  assign n22623 = n149 & n22622 ;
  assign n22624 = n22615 & ~n22623 ;
  assign n22625 = x2 & ~n22624 ;
  assign n22626 = x2 & ~n22625 ;
  assign n22627 = ~n22624 & ~n22625 ;
  assign n22628 = ~n22626 & ~n22627 ;
  assign n22629 = n22610 & ~n22628 ;
  assign n22630 = n22610 & ~n22629 ;
  assign n22631 = ~n22628 & ~n22629 ;
  assign n22632 = ~n22630 & ~n22631 ;
  assign n22633 = ~n21877 & ~n21882 ;
  assign n22634 = ~n22632 & ~n22633 ;
  assign n22635 = n22632 & n22633 ;
  assign n22636 = ~n22634 & ~n22635 ;
  assign n23014 = n22636 & x186 ;
  assign n22637 = ~n22213 & ~n22217 ;
  assign n22638 = ~x119 & n293 ;
  assign n22639 = ~x117 & n373 ;
  assign n22640 = ~x118 & n288 ;
  assign n22641 = ~n22639 & ~n22640 ;
  assign n22642 = ~n22638 & n22641 ;
  assign n22643 = n296 & n20778 ;
  assign n22644 = n22642 & ~n22643 ;
  assign n22645 = ~x5 & ~n22644 ;
  assign n22646 = ~x5 & ~n22645 ;
  assign n22647 = ~n22644 & ~n22645 ;
  assign n22648 = ~n22646 & ~n22647 ;
  assign n22649 = ~n22205 & ~n22209 ;
  assign n22650 = ~x116 & n574 ;
  assign n22651 = ~x114 & n673 ;
  assign n22652 = ~x115 & n569 ;
  assign n22653 = ~n22651 & ~n22652 ;
  assign n22654 = ~n22650 & n22653 ;
  assign n22655 = n577 & n18678 ;
  assign n22656 = n22654 & ~n22655 ;
  assign n22657 = ~x8 & ~n22656 ;
  assign n22658 = ~x8 & ~n22657 ;
  assign n22659 = ~n22656 & ~n22657 ;
  assign n22660 = ~n22658 & ~n22659 ;
  assign n22661 = ~n22197 & ~n22201 ;
  assign n22662 = ~x113 & n945 ;
  assign n22663 = ~x111 & n1099 ;
  assign n22664 = ~x112 & n940 ;
  assign n22665 = ~n22663 & ~n22664 ;
  assign n22666 = ~n22662 & n22665 ;
  assign n22667 = n948 & n16684 ;
  assign n22668 = n22666 & ~n22667 ;
  assign n22669 = ~x11 & ~n22668 ;
  assign n22670 = ~x11 & ~n22669 ;
  assign n22671 = ~n22668 & ~n22669 ;
  assign n22672 = ~n22670 & ~n22671 ;
  assign n22673 = ~n22189 & ~n22193 ;
  assign n22674 = ~n22184 & ~n22186 ;
  assign n22675 = ~n22112 & ~n22115 ;
  assign n22676 = ~n22107 & ~n22109 ;
  assign n22677 = ~n22062 & ~n22066 ;
  assign n22678 = ~n22051 & ~n22053 ;
  assign n22679 = ~n21245 & ~n22029 ;
  assign n22680 = ~n22026 & ~n22679 ;
  assign n22681 = ~x71 & n18025 ;
  assign n22682 = ~x69 & n18764 ;
  assign n22683 = ~x70 & n18020 ;
  assign n22684 = ~n22682 & ~n22683 ;
  assign n22685 = ~n22681 & n22684 ;
  assign n22686 = n622 & n18028 ;
  assign n22687 = n22685 & ~n22686 ;
  assign n22688 = ~x53 & ~n22687 ;
  assign n22689 = ~x53 & ~n22688 ;
  assign n22690 = ~n22687 & ~n22688 ;
  assign n22691 = ~n22689 & ~n22690 ;
  assign n22692 = n21227 & n21997 ;
  assign n22693 = ~n22012 & ~n22692 ;
  assign n22694 = ~x68 & n20143 ;
  assign n22695 = ~x66 & n20854 ;
  assign n22696 = ~x67 & n20138 ;
  assign n22697 = ~n22695 & ~n22696 ;
  assign n22698 = ~n22694 & n22697 ;
  assign n22699 = n352 & n20146 ;
  assign n22700 = n22698 & ~n22699 ;
  assign n22701 = ~x56 & ~n22700 ;
  assign n22702 = ~x56 & ~n22701 ;
  assign n22703 = ~n22700 & ~n22701 ;
  assign n22704 = ~n22702 & ~n22703 ;
  assign n22705 = ~x59 & ~n21997 ;
  assign n22706 = ~x64 & n22320 ;
  assign n22707 = ~x65 & n22325 ;
  assign n22708 = ~n22706 & ~n22707 ;
  assign n22709 = ~n22329 & n22708 ;
  assign n22710 = ~x59 & ~n22709 ;
  assign n22711 = ~x59 & ~n22710 ;
  assign n22712 = ~n22709 & ~n22710 ;
  assign n22713 = ~n22711 & ~n22712 ;
  assign n22714 = n22705 & ~n22713 ;
  assign n22715 = ~n22705 & n22713 ;
  assign n22716 = ~n22714 & ~n22715 ;
  assign n22717 = n22704 & ~n22716 ;
  assign n22718 = ~n22704 & n22716 ;
  assign n22719 = ~n22717 & ~n22718 ;
  assign n22720 = ~n22693 & n22719 ;
  assign n22721 = n22693 & ~n22719 ;
  assign n22722 = ~n22720 & ~n22721 ;
  assign n22723 = n22691 & ~n22722 ;
  assign n22724 = ~n22691 & n22722 ;
  assign n22725 = ~n22723 & ~n22724 ;
  assign n22726 = ~n22680 & n22725 ;
  assign n22727 = n22680 & ~n22725 ;
  assign n22728 = ~n22726 & ~n22727 ;
  assign n22729 = ~x74 & n16076 ;
  assign n22730 = ~x72 & n16756 ;
  assign n22731 = ~x73 & n16071 ;
  assign n22732 = ~n22730 & ~n22731 ;
  assign n22733 = ~n22729 & n22732 ;
  assign n22734 = n1066 & n16079 ;
  assign n22735 = n22733 & ~n22734 ;
  assign n22736 = ~x50 & ~n22735 ;
  assign n22737 = ~x50 & ~n22736 ;
  assign n22738 = ~n22735 & ~n22736 ;
  assign n22739 = ~n22737 & ~n22738 ;
  assign n22740 = n22728 & ~n22739 ;
  assign n22741 = n22728 & ~n22740 ;
  assign n22742 = ~n22739 & ~n22740 ;
  assign n22743 = ~n22741 & ~n22742 ;
  assign n22744 = ~n22044 & ~n22047 ;
  assign n22745 = n22743 & n22744 ;
  assign n22746 = ~n22743 & ~n22744 ;
  assign n22747 = ~n22745 & ~n22746 ;
  assign n22748 = ~x77 & n14233 ;
  assign n22749 = ~x75 & n14876 ;
  assign n22750 = ~x76 & n14228 ;
  assign n22751 = ~n22749 & ~n22750 ;
  assign n22752 = ~n22748 & n22751 ;
  assign n22753 = n1594 & n14236 ;
  assign n22754 = n22752 & ~n22753 ;
  assign n22755 = ~x47 & ~n22754 ;
  assign n22756 = ~x47 & ~n22755 ;
  assign n22757 = ~n22754 & ~n22755 ;
  assign n22758 = ~n22756 & ~n22757 ;
  assign n22759 = n22747 & ~n22758 ;
  assign n22760 = ~n22747 & n22758 ;
  assign n22761 = ~n22678 & ~n22760 ;
  assign n22762 = ~n22759 & n22761 ;
  assign n22763 = ~n22678 & ~n22762 ;
  assign n22764 = ~n22759 & ~n22762 ;
  assign n22765 = ~n22760 & n22764 ;
  assign n22766 = ~n22763 & ~n22765 ;
  assign n22767 = ~x80 & n12506 ;
  assign n22768 = ~x78 & n13131 ;
  assign n22769 = ~x79 & n12501 ;
  assign n22770 = ~n22768 & ~n22769 ;
  assign n22771 = ~n22767 & n22770 ;
  assign n22772 = n2145 & n12509 ;
  assign n22773 = n22771 & ~n22772 ;
  assign n22774 = ~x44 & ~n22773 ;
  assign n22775 = ~x44 & ~n22774 ;
  assign n22776 = ~n22773 & ~n22774 ;
  assign n22777 = ~n22775 & ~n22776 ;
  assign n22778 = ~n22766 & ~n22777 ;
  assign n22779 = ~n22766 & ~n22778 ;
  assign n22780 = ~n22777 & ~n22778 ;
  assign n22781 = ~n22779 & ~n22780 ;
  assign n22782 = ~n22056 & ~n22059 ;
  assign n22783 = n22781 & n22782 ;
  assign n22784 = ~n22781 & ~n22782 ;
  assign n22785 = ~n22783 & ~n22784 ;
  assign n22786 = ~x83 & n10905 ;
  assign n22787 = ~x81 & n11466 ;
  assign n22788 = ~x82 & n10900 ;
  assign n22789 = ~n22787 & ~n22788 ;
  assign n22790 = ~n22786 & n22789 ;
  assign n22791 = n2972 & n10908 ;
  assign n22792 = n22790 & ~n22791 ;
  assign n22793 = ~x41 & ~n22792 ;
  assign n22794 = ~x41 & ~n22793 ;
  assign n22795 = ~n22792 & ~n22793 ;
  assign n22796 = ~n22794 & ~n22795 ;
  assign n22797 = n22785 & ~n22796 ;
  assign n22798 = ~n22785 & n22796 ;
  assign n22799 = ~n22677 & ~n22798 ;
  assign n22800 = ~n22797 & n22799 ;
  assign n22801 = ~n22677 & ~n22800 ;
  assign n22802 = ~n22797 & ~n22800 ;
  assign n22803 = ~n22798 & n22802 ;
  assign n22804 = ~n22801 & ~n22803 ;
  assign n22805 = ~x86 & n9433 ;
  assign n22806 = ~x84 & n9915 ;
  assign n22807 = ~x85 & n9428 ;
  assign n22808 = ~n22806 & ~n22807 ;
  assign n22809 = ~n22805 & n22808 ;
  assign n22810 = n3832 & n9436 ;
  assign n22811 = n22809 & ~n22810 ;
  assign n22812 = ~x38 & ~n22811 ;
  assign n22813 = ~x38 & ~n22812 ;
  assign n22814 = ~n22811 & ~n22812 ;
  assign n22815 = ~n22813 & ~n22814 ;
  assign n22816 = ~n22804 & ~n22815 ;
  assign n22817 = ~n22804 & ~n22816 ;
  assign n22818 = ~n22815 & ~n22816 ;
  assign n22819 = ~n22817 & ~n22818 ;
  assign n22820 = ~n22070 & ~n22073 ;
  assign n22821 = n22819 & n22820 ;
  assign n22822 = ~n22819 & ~n22820 ;
  assign n22823 = ~n22821 & ~n22822 ;
  assign n22824 = ~x89 & n8006 ;
  assign n22825 = ~x87 & n8474 ;
  assign n22826 = ~x88 & n8001 ;
  assign n22827 = ~n22825 & ~n22826 ;
  assign n22828 = ~n22824 & n22827 ;
  assign n22829 = n4664 & n8009 ;
  assign n22830 = n22828 & ~n22829 ;
  assign n22831 = ~x35 & ~n22830 ;
  assign n22832 = ~x35 & ~n22831 ;
  assign n22833 = ~n22830 & ~n22831 ;
  assign n22834 = ~n22832 & ~n22833 ;
  assign n22835 = n22823 & ~n22834 ;
  assign n22836 = n22823 & ~n22835 ;
  assign n22837 = ~n22834 & ~n22835 ;
  assign n22838 = ~n22836 & ~n22837 ;
  assign n22839 = ~n22087 & ~n22093 ;
  assign n22840 = n22838 & n22839 ;
  assign n22841 = ~n22838 & ~n22839 ;
  assign n22842 = ~n22840 & ~n22841 ;
  assign n22843 = ~x92 & n6725 ;
  assign n22844 = ~x90 & n7129 ;
  assign n22845 = ~x91 & n6720 ;
  assign n22846 = ~n22844 & ~n22845 ;
  assign n22847 = ~n22843 & n22846 ;
  assign n22848 = n5896 & n6728 ;
  assign n22849 = n22847 & ~n22848 ;
  assign n22850 = ~x32 & ~n22849 ;
  assign n22851 = ~x32 & ~n22850 ;
  assign n22852 = ~n22849 & ~n22850 ;
  assign n22853 = ~n22851 & ~n22852 ;
  assign n22854 = n22842 & ~n22853 ;
  assign n22855 = n22842 & ~n22854 ;
  assign n22856 = ~n22853 & ~n22854 ;
  assign n22857 = ~n22855 & ~n22856 ;
  assign n22858 = ~n22676 & n22857 ;
  assign n22859 = n22676 & ~n22857 ;
  assign n22860 = ~n22858 & ~n22859 ;
  assign n22861 = ~x95 & n5560 ;
  assign n22862 = ~x93 & n5943 ;
  assign n22863 = ~x94 & n5555 ;
  assign n22864 = ~n22862 & ~n22863 ;
  assign n22865 = ~n22861 & n22864 ;
  assign n22866 = n5563 & n7100 ;
  assign n22867 = n22865 & ~n22866 ;
  assign n22868 = ~x29 & ~n22867 ;
  assign n22869 = ~x29 & ~n22868 ;
  assign n22870 = ~n22867 & ~n22868 ;
  assign n22871 = ~n22869 & ~n22870 ;
  assign n22872 = ~n22860 & ~n22871 ;
  assign n22873 = n22860 & n22871 ;
  assign n22874 = ~n22872 & ~n22873 ;
  assign n22875 = n22675 & ~n22874 ;
  assign n22876 = ~n22675 & n22874 ;
  assign n22877 = ~n22875 & ~n22876 ;
  assign n22878 = ~x98 & n4531 ;
  assign n22879 = ~x96 & n4847 ;
  assign n22880 = ~x97 & n4526 ;
  assign n22881 = ~n22879 & ~n22880 ;
  assign n22882 = ~n22878 & n22881 ;
  assign n22883 = n4534 & n8426 ;
  assign n22884 = n22882 & ~n22883 ;
  assign n22885 = ~x26 & ~n22884 ;
  assign n22886 = ~x26 & ~n22885 ;
  assign n22887 = ~n22884 & ~n22885 ;
  assign n22888 = ~n22886 & ~n22887 ;
  assign n22889 = n22877 & ~n22888 ;
  assign n22890 = n22877 & ~n22889 ;
  assign n22891 = ~n22888 & ~n22889 ;
  assign n22892 = ~n22890 & ~n22891 ;
  assign n22893 = ~n21934 & ~n22132 ;
  assign n22894 = ~n22129 & ~n22893 ;
  assign n22895 = n22892 & n22894 ;
  assign n22896 = ~n22892 & ~n22894 ;
  assign n22897 = ~n22895 & ~n22896 ;
  assign n22898 = ~x101 & n3589 ;
  assign n22899 = ~x99 & n3878 ;
  assign n22900 = ~x100 & n3584 ;
  assign n22901 = ~n22899 & ~n22900 ;
  assign n22902 = ~n22898 & n22901 ;
  assign n22903 = n3592 & n9844 ;
  assign n22904 = n22902 & ~n22903 ;
  assign n22905 = ~x23 & ~n22904 ;
  assign n22906 = ~x23 & ~n22905 ;
  assign n22907 = ~n22904 & ~n22905 ;
  assign n22908 = ~n22906 & ~n22907 ;
  assign n22909 = n22897 & ~n22908 ;
  assign n22910 = n22897 & ~n22909 ;
  assign n22911 = ~n22908 & ~n22909 ;
  assign n22912 = ~n22910 & ~n22911 ;
  assign n22913 = ~n22147 & ~n22151 ;
  assign n22914 = n22912 & n22913 ;
  assign n22915 = ~n22912 & ~n22913 ;
  assign n22916 = ~n22914 & ~n22915 ;
  assign n22917 = ~x104 & n2751 ;
  assign n22918 = ~x102 & n3020 ;
  assign n22919 = ~x103 & n2746 ;
  assign n22920 = ~n22918 & ~n22919 ;
  assign n22921 = ~n22917 & n22920 ;
  assign n22922 = n2754 & n11380 ;
  assign n22923 = n22921 & ~n22922 ;
  assign n22924 = ~x20 & ~n22923 ;
  assign n22925 = ~x20 & ~n22924 ;
  assign n22926 = ~n22923 & ~n22924 ;
  assign n22927 = ~n22925 & ~n22926 ;
  assign n22928 = n22916 & ~n22927 ;
  assign n22929 = n22916 & ~n22928 ;
  assign n22930 = ~n22927 & ~n22928 ;
  assign n22931 = ~n22929 & ~n22930 ;
  assign n22932 = ~n22164 & ~n22170 ;
  assign n22933 = n22931 & n22932 ;
  assign n22934 = ~n22931 & ~n22932 ;
  assign n22935 = ~n22933 & ~n22934 ;
  assign n22936 = ~x107 & n2093 ;
  assign n22937 = ~x105 & n2275 ;
  assign n22938 = ~x106 & n2088 ;
  assign n22939 = ~n22937 & ~n22938 ;
  assign n22940 = ~n22936 & n22939 ;
  assign n22941 = n2096 & n13034 ;
  assign n22942 = n22940 & ~n22941 ;
  assign n22943 = ~x17 & ~n22942 ;
  assign n22944 = ~x17 & ~n22943 ;
  assign n22945 = ~n22942 & ~n22943 ;
  assign n22946 = ~n22944 & ~n22945 ;
  assign n22947 = n22935 & ~n22946 ;
  assign n22948 = ~n22935 & n22946 ;
  assign n22949 = ~n22674 & ~n22948 ;
  assign n22950 = ~n22947 & n22949 ;
  assign n22951 = ~n22674 & ~n22950 ;
  assign n22952 = ~n22947 & ~n22950 ;
  assign n22953 = ~n22948 & n22952 ;
  assign n22954 = ~n22951 & ~n22953 ;
  assign n22955 = ~x110 & n1434 ;
  assign n22956 = ~x108 & n1646 ;
  assign n22957 = ~x109 & n1429 ;
  assign n22958 = ~n22956 & ~n22957 ;
  assign n22959 = ~n22955 & n22958 ;
  assign n22960 = n1437 & n14802 ;
  assign n22961 = n22959 & ~n22960 ;
  assign n22962 = ~x14 & ~n22961 ;
  assign n22963 = ~x14 & ~n22962 ;
  assign n22964 = ~n22961 & ~n22962 ;
  assign n22965 = ~n22963 & ~n22964 ;
  assign n22966 = n22954 & n22965 ;
  assign n22967 = ~n22954 & ~n22965 ;
  assign n22968 = ~n22966 & ~n22967 ;
  assign n22969 = ~n22673 & n22968 ;
  assign n22970 = n22673 & ~n22968 ;
  assign n22971 = ~n22969 & ~n22970 ;
  assign n22972 = n22672 & ~n22971 ;
  assign n22973 = ~n22672 & n22971 ;
  assign n22974 = ~n22972 & ~n22973 ;
  assign n22975 = ~n22661 & n22974 ;
  assign n22976 = n22661 & ~n22974 ;
  assign n22977 = ~n22975 & ~n22976 ;
  assign n22978 = n22660 & ~n22977 ;
  assign n22979 = ~n22660 & n22977 ;
  assign n22980 = ~n22978 & ~n22979 ;
  assign n22981 = ~n22649 & n22980 ;
  assign n22982 = n22649 & ~n22980 ;
  assign n22983 = ~n22981 & ~n22982 ;
  assign n22984 = n22648 & ~n22983 ;
  assign n22985 = ~n22648 & n22983 ;
  assign n22986 = ~n22984 & ~n22985 ;
  assign n22987 = ~n22637 & n22986 ;
  assign n22988 = n22637 & ~n22986 ;
  assign n22989 = ~n22987 & ~n22988 ;
  assign n22990 = ~x122 & n164 ;
  assign n22991 = ~x120 & n205 ;
  assign n22992 = ~x121 & n162 ;
  assign n22993 = ~n22991 & ~n22992 ;
  assign n22994 = ~n22990 & n22993 ;
  assign n22995 = ~n21865 & ~n22227 ;
  assign n22996 = n22619 & ~n22995 ;
  assign n22997 = ~n22619 & n22995 ;
  assign n22998 = ~n22996 & ~n22997 ;
  assign n22999 = n167 & n22998 ;
  assign n23000 = n22994 & ~n22999 ;
  assign n23001 = ~x2 & ~n23000 ;
  assign n23002 = ~x2 & ~n23001 ;
  assign n23003 = ~n23000 & ~n23001 ;
  assign n23004 = ~n23002 & ~n23003 ;
  assign n23005 = n22989 & ~n23004 ;
  assign n23006 = n22989 & ~n23005 ;
  assign n23007 = ~n23004 & ~n23005 ;
  assign n23008 = ~n23006 & ~n23007 ;
  assign n23009 = ~n22236 & ~n22241 ;
  assign n23010 = ~n23008 & ~n23009 ;
  assign n23011 = n23008 & n23009 ;
  assign n23012 = ~n23010 & ~n23011 ;
  assign n23015 = ~n23012 & ~x186 ;
  assign n23016 = ~n23014 & ~n23015 ;
  assign n23017 = ~n22629 & ~n22634 ;
  assign n23018 = ~n22606 & ~n22608 ;
  assign n23019 = ~n22600 & ~n22602 ;
  assign n23020 = x117 & n574 ;
  assign n23021 = x115 & n673 ;
  assign n23022 = x116 & n569 ;
  assign n23023 = ~n23021 & ~n23022 ;
  assign n23024 = ~n23020 & n23023 ;
  assign n23025 = n577 & n19026 ;
  assign n23026 = n23024 & ~n23025 ;
  assign n23027 = x8 & ~n23026 ;
  assign n23028 = x8 & ~n23027 ;
  assign n23029 = ~n23026 & ~n23027 ;
  assign n23030 = ~n23028 & ~n23029 ;
  assign n23031 = ~n22594 & ~n22596 ;
  assign n23032 = ~n22588 & ~n22590 ;
  assign n23033 = ~n22549 & ~n22555 ;
  assign n23034 = ~n22493 & ~n22497 ;
  assign n23035 = ~n22287 & ~n22478 ;
  assign n23036 = ~n22475 & ~n23035 ;
  assign n23037 = ~n22437 & ~n22443 ;
  assign n23038 = ~n22399 & ~n22405 ;
  assign n23039 = x81 & n12506 ;
  assign n23040 = x79 & n13131 ;
  assign n23041 = x80 & n12501 ;
  assign n23042 = ~n23040 & ~n23041 ;
  assign n23043 = ~n23039 & n23042 ;
  assign n23044 = n2348 & n12509 ;
  assign n23045 = n23043 & ~n23044 ;
  assign n23046 = x44 & ~n23045 ;
  assign n23047 = x44 & ~n23046 ;
  assign n23048 = ~n23045 & ~n23046 ;
  assign n23049 = ~n23047 & ~n23048 ;
  assign n23050 = ~n22361 & ~n22367 ;
  assign n23051 = x75 & n16076 ;
  assign n23052 = x73 & n16756 ;
  assign n23053 = x74 & n16071 ;
  assign n23054 = ~n23052 & ~n23053 ;
  assign n23055 = ~n23051 & n23054 ;
  assign n23056 = n1150 & n16079 ;
  assign n23057 = n23055 & ~n23056 ;
  assign n23058 = x50 & ~n23057 ;
  assign n23059 = x50 & ~n23058 ;
  assign n23060 = ~n23057 & ~n23058 ;
  assign n23061 = ~n23059 & ~n23060 ;
  assign n23062 = ~n22345 & ~n22347 ;
  assign n23063 = ~n22339 & ~n22341 ;
  assign n23064 = x66 & n22325 ;
  assign n23065 = n21634 & ~n22324 ;
  assign n23066 = n22319 & n23065 ;
  assign n23067 = x64 & n23066 ;
  assign n23068 = x65 & n22320 ;
  assign n23069 = ~n23067 & ~n23068 ;
  assign n23070 = ~n23064 & n23069 ;
  assign n23071 = n194 & n22328 ;
  assign n23072 = n23070 & ~n23071 ;
  assign n23073 = x59 & ~n23072 ;
  assign n23074 = x59 & ~n23073 ;
  assign n23075 = ~n23072 & ~n23073 ;
  assign n23076 = ~n23074 & ~n23075 ;
  assign n23077 = ~n22335 & n23076 ;
  assign n23078 = n22335 & ~n23076 ;
  assign n23079 = ~n23077 & ~n23078 ;
  assign n23080 = x69 & n20143 ;
  assign n23081 = x67 & n20854 ;
  assign n23082 = x68 & n20138 ;
  assign n23083 = ~n23081 & ~n23082 ;
  assign n23084 = ~n23080 & n23083 ;
  assign n23085 = n398 & n20146 ;
  assign n23086 = n23084 & ~n23085 ;
  assign n23087 = x56 & ~n23086 ;
  assign n23088 = x56 & ~n23087 ;
  assign n23089 = ~n23086 & ~n23087 ;
  assign n23090 = ~n23088 & ~n23089 ;
  assign n23091 = n23079 & ~n23090 ;
  assign n23092 = ~n23079 & n23090 ;
  assign n23093 = ~n23063 & ~n23092 ;
  assign n23094 = ~n23091 & n23093 ;
  assign n23095 = ~n23063 & ~n23094 ;
  assign n23096 = ~n23091 & ~n23094 ;
  assign n23097 = ~n23092 & n23096 ;
  assign n23098 = ~n23095 & ~n23097 ;
  assign n23099 = x72 & n18025 ;
  assign n23100 = x70 & n18764 ;
  assign n23101 = x71 & n18020 ;
  assign n23102 = ~n23100 & ~n23101 ;
  assign n23103 = ~n23099 & n23102 ;
  assign n23104 = n717 & n18028 ;
  assign n23105 = n23103 & ~n23104 ;
  assign n23106 = x53 & ~n23105 ;
  assign n23107 = x53 & ~n23106 ;
  assign n23108 = ~n23105 & ~n23106 ;
  assign n23109 = ~n23107 & ~n23108 ;
  assign n23110 = n23098 & n23109 ;
  assign n23111 = ~n23098 & ~n23109 ;
  assign n23112 = ~n23110 & ~n23111 ;
  assign n23113 = ~n23062 & n23112 ;
  assign n23114 = n23062 & ~n23112 ;
  assign n23115 = ~n23113 & ~n23114 ;
  assign n23116 = n23061 & ~n23115 ;
  assign n23117 = ~n23061 & n23115 ;
  assign n23118 = ~n23116 & ~n23117 ;
  assign n23119 = ~n23050 & n23118 ;
  assign n23120 = n23050 & ~n23118 ;
  assign n23121 = ~n23119 & ~n23120 ;
  assign n23122 = x78 & n14233 ;
  assign n23123 = x76 & n14876 ;
  assign n23124 = x77 & n14228 ;
  assign n23125 = ~n23123 & ~n23124 ;
  assign n23126 = ~n23122 & n23125 ;
  assign n23127 = n1624 & n14236 ;
  assign n23128 = n23126 & ~n23127 ;
  assign n23129 = x47 & ~n23128 ;
  assign n23130 = x47 & ~n23129 ;
  assign n23131 = ~n23128 & ~n23129 ;
  assign n23132 = ~n23130 & ~n23131 ;
  assign n23133 = n23121 & ~n23132 ;
  assign n23134 = n23121 & ~n23133 ;
  assign n23135 = ~n23132 & ~n23133 ;
  assign n23136 = ~n23134 & ~n23135 ;
  assign n23137 = ~n22385 & ~n23136 ;
  assign n23138 = n22385 & n23136 ;
  assign n23139 = ~n23137 & ~n23138 ;
  assign n23140 = ~n23049 & n23139 ;
  assign n23141 = ~n23049 & ~n23140 ;
  assign n23142 = n23139 & ~n23140 ;
  assign n23143 = ~n23141 & ~n23142 ;
  assign n23144 = ~n23038 & ~n23143 ;
  assign n23145 = ~n23038 & ~n23144 ;
  assign n23146 = ~n23143 & ~n23144 ;
  assign n23147 = ~n23145 & ~n23146 ;
  assign n23148 = x84 & n10905 ;
  assign n23149 = x82 & n11466 ;
  assign n23150 = x83 & n10900 ;
  assign n23151 = ~n23149 & ~n23150 ;
  assign n23152 = ~n23148 & n23151 ;
  assign n23153 = n3114 & n10908 ;
  assign n23154 = n23152 & ~n23153 ;
  assign n23155 = x41 & ~n23154 ;
  assign n23156 = x41 & ~n23155 ;
  assign n23157 = ~n23154 & ~n23155 ;
  assign n23158 = ~n23156 & ~n23157 ;
  assign n23159 = ~n23147 & ~n23158 ;
  assign n23160 = ~n23147 & ~n23159 ;
  assign n23161 = ~n23158 & ~n23159 ;
  assign n23162 = ~n23160 & ~n23161 ;
  assign n23163 = ~n22423 & n23162 ;
  assign n23164 = n22423 & ~n23162 ;
  assign n23165 = ~n23163 & ~n23164 ;
  assign n23166 = x87 & n9433 ;
  assign n23167 = x85 & n9915 ;
  assign n23168 = x86 & n9428 ;
  assign n23169 = ~n23167 & ~n23168 ;
  assign n23170 = ~n23166 & n23169 ;
  assign n23171 = n3991 & n9436 ;
  assign n23172 = n23170 & ~n23171 ;
  assign n23173 = x38 & ~n23172 ;
  assign n23174 = x38 & ~n23173 ;
  assign n23175 = ~n23172 & ~n23173 ;
  assign n23176 = ~n23174 & ~n23175 ;
  assign n23177 = ~n23165 & ~n23176 ;
  assign n23178 = n23165 & n23176 ;
  assign n23179 = ~n23177 & ~n23178 ;
  assign n23180 = n23037 & ~n23179 ;
  assign n23181 = ~n23037 & n23179 ;
  assign n23182 = ~n23180 & ~n23181 ;
  assign n23183 = x90 & n8006 ;
  assign n23184 = x88 & n8474 ;
  assign n23185 = x89 & n8001 ;
  assign n23186 = ~n23184 & ~n23185 ;
  assign n23187 = ~n23183 & n23186 ;
  assign n23188 = n4986 & n8009 ;
  assign n23189 = n23187 & ~n23188 ;
  assign n23190 = x35 & ~n23189 ;
  assign n23191 = x35 & ~n23190 ;
  assign n23192 = ~n23189 & ~n23190 ;
  assign n23193 = ~n23191 & ~n23192 ;
  assign n23194 = n23182 & ~n23193 ;
  assign n23195 = n23182 & ~n23194 ;
  assign n23196 = ~n23193 & ~n23194 ;
  assign n23197 = ~n23195 & ~n23196 ;
  assign n23198 = ~n22456 & ~n22462 ;
  assign n23199 = n23197 & n23198 ;
  assign n23200 = ~n23197 & ~n23198 ;
  assign n23201 = ~n23199 & ~n23200 ;
  assign n23202 = x93 & n6725 ;
  assign n23203 = x91 & n7129 ;
  assign n23204 = x92 & n6720 ;
  assign n23205 = ~n23203 & ~n23204 ;
  assign n23206 = ~n23202 & n23205 ;
  assign n23207 = n6094 & n6728 ;
  assign n23208 = n23206 & ~n23207 ;
  assign n23209 = x32 & ~n23208 ;
  assign n23210 = x32 & ~n23209 ;
  assign n23211 = ~n23208 & ~n23209 ;
  assign n23212 = ~n23210 & ~n23211 ;
  assign n23213 = n23201 & ~n23212 ;
  assign n23214 = ~n23201 & n23212 ;
  assign n23215 = ~n23036 & ~n23214 ;
  assign n23216 = ~n23213 & n23215 ;
  assign n23217 = ~n23036 & ~n23216 ;
  assign n23218 = ~n23213 & ~n23216 ;
  assign n23219 = ~n23214 & n23218 ;
  assign n23220 = ~n23217 & ~n23219 ;
  assign n23221 = x96 & n5560 ;
  assign n23222 = x94 & n5943 ;
  assign n23223 = x95 & n5555 ;
  assign n23224 = ~n23222 & ~n23223 ;
  assign n23225 = ~n23221 & n23224 ;
  assign n23226 = n5563 & n7321 ;
  assign n23227 = n23225 & ~n23226 ;
  assign n23228 = x29 & ~n23227 ;
  assign n23229 = x29 & ~n23228 ;
  assign n23230 = ~n23227 & ~n23228 ;
  assign n23231 = ~n23229 & ~n23230 ;
  assign n23232 = n23220 & n23231 ;
  assign n23233 = ~n23220 & ~n23231 ;
  assign n23234 = ~n23232 & ~n23233 ;
  assign n23235 = ~n23034 & n23234 ;
  assign n23236 = n23034 & ~n23234 ;
  assign n23237 = ~n23235 & ~n23236 ;
  assign n23238 = x99 & n4531 ;
  assign n23239 = x97 & n4847 ;
  assign n23240 = x98 & n4526 ;
  assign n23241 = ~n23239 & ~n23240 ;
  assign n23242 = ~n23238 & n23241 ;
  assign n23243 = n4534 & n8660 ;
  assign n23244 = n23242 & ~n23243 ;
  assign n23245 = x26 & ~n23244 ;
  assign n23246 = x26 & ~n23245 ;
  assign n23247 = ~n23244 & ~n23245 ;
  assign n23248 = ~n23246 & ~n23247 ;
  assign n23249 = n23237 & ~n23248 ;
  assign n23250 = n23237 & ~n23249 ;
  assign n23251 = ~n23248 & ~n23249 ;
  assign n23252 = ~n23250 & ~n23251 ;
  assign n23253 = ~n22510 & ~n22517 ;
  assign n23254 = n23252 & n23253 ;
  assign n23255 = ~n23252 & ~n23253 ;
  assign n23256 = ~n23254 & ~n23255 ;
  assign n23257 = x102 & n3589 ;
  assign n23258 = x100 & n3878 ;
  assign n23259 = x101 & n3584 ;
  assign n23260 = ~n23258 & ~n23259 ;
  assign n23261 = ~n23257 & n23260 ;
  assign n23262 = n3592 & n10092 ;
  assign n23263 = n23261 & ~n23262 ;
  assign n23264 = x23 & ~n23263 ;
  assign n23265 = x23 & ~n23264 ;
  assign n23266 = ~n23263 & ~n23264 ;
  assign n23267 = ~n23265 & ~n23266 ;
  assign n23268 = n23256 & ~n23267 ;
  assign n23269 = n23256 & ~n23268 ;
  assign n23270 = ~n23267 & ~n23268 ;
  assign n23271 = ~n23269 & ~n23270 ;
  assign n23272 = ~n22530 & ~n22536 ;
  assign n23273 = n23271 & n23272 ;
  assign n23274 = ~n23271 & ~n23272 ;
  assign n23275 = ~n23273 & ~n23274 ;
  assign n23276 = x105 & n2751 ;
  assign n23277 = x103 & n3020 ;
  assign n23278 = x104 & n2746 ;
  assign n23279 = ~n23277 & ~n23278 ;
  assign n23280 = ~n23276 & n23279 ;
  assign n23281 = n2754 & n11648 ;
  assign n23282 = n23280 & ~n23281 ;
  assign n23283 = x20 & ~n23282 ;
  assign n23284 = x20 & ~n23283 ;
  assign n23285 = ~n23282 & ~n23283 ;
  assign n23286 = ~n23284 & ~n23285 ;
  assign n23287 = n23275 & ~n23286 ;
  assign n23288 = ~n23275 & n23286 ;
  assign n23289 = ~n23033 & ~n23288 ;
  assign n23290 = ~n23287 & n23289 ;
  assign n23291 = ~n23033 & ~n23290 ;
  assign n23292 = ~n23287 & ~n23290 ;
  assign n23293 = ~n23288 & n23292 ;
  assign n23294 = ~n23291 & ~n23293 ;
  assign n23295 = x108 & n2093 ;
  assign n23296 = x106 & n2275 ;
  assign n23297 = x107 & n2088 ;
  assign n23298 = ~n23296 & ~n23297 ;
  assign n23299 = ~n23295 & n23298 ;
  assign n23300 = n2096 & n13323 ;
  assign n23301 = n23299 & ~n23300 ;
  assign n23302 = x17 & ~n23301 ;
  assign n23303 = x17 & ~n23302 ;
  assign n23304 = ~n23301 & ~n23302 ;
  assign n23305 = ~n23303 & ~n23304 ;
  assign n23306 = ~n23294 & ~n23305 ;
  assign n23307 = ~n23294 & ~n23306 ;
  assign n23308 = ~n23305 & ~n23306 ;
  assign n23309 = ~n23307 & ~n23308 ;
  assign n23310 = ~n22573 & n23309 ;
  assign n23311 = n22573 & ~n23309 ;
  assign n23312 = ~n23310 & ~n23311 ;
  assign n23313 = x111 & n1434 ;
  assign n23314 = x109 & n1646 ;
  assign n23315 = x110 & n1429 ;
  assign n23316 = ~n23314 & ~n23315 ;
  assign n23317 = ~n23313 & n23316 ;
  assign n23318 = n1437 & n15111 ;
  assign n23319 = n23317 & ~n23318 ;
  assign n23320 = x14 & ~n23319 ;
  assign n23321 = x14 & ~n23320 ;
  assign n23322 = ~n23319 & ~n23320 ;
  assign n23323 = ~n23321 & ~n23322 ;
  assign n23324 = ~n23312 & ~n23323 ;
  assign n23325 = n23312 & n23323 ;
  assign n23326 = ~n23324 & ~n23325 ;
  assign n23327 = ~n23032 & n23326 ;
  assign n23328 = n23032 & ~n23326 ;
  assign n23329 = ~n23327 & ~n23328 ;
  assign n23330 = x114 & n945 ;
  assign n23331 = x112 & n1099 ;
  assign n23332 = x113 & n940 ;
  assign n23333 = ~n23331 & ~n23332 ;
  assign n23334 = ~n23330 & n23333 ;
  assign n23335 = n948 & n17012 ;
  assign n23336 = n23334 & ~n23335 ;
  assign n23337 = x11 & ~n23336 ;
  assign n23338 = x11 & ~n23337 ;
  assign n23339 = ~n23336 & ~n23337 ;
  assign n23340 = ~n23338 & ~n23339 ;
  assign n23341 = n23329 & ~n23340 ;
  assign n23342 = n23329 & ~n23341 ;
  assign n23343 = ~n23340 & ~n23341 ;
  assign n23344 = ~n23342 & ~n23343 ;
  assign n23345 = ~n23031 & ~n23344 ;
  assign n23346 = n23031 & n23344 ;
  assign n23347 = ~n23345 & ~n23346 ;
  assign n23348 = ~n23030 & n23347 ;
  assign n23349 = ~n23030 & ~n23348 ;
  assign n23350 = n23347 & ~n23348 ;
  assign n23351 = ~n23349 & ~n23350 ;
  assign n23352 = ~n23019 & ~n23351 ;
  assign n23353 = ~n23019 & ~n23352 ;
  assign n23354 = ~n23351 & ~n23352 ;
  assign n23355 = ~n23353 & ~n23354 ;
  assign n23356 = x120 & n293 ;
  assign n23357 = x118 & n373 ;
  assign n23358 = x119 & n288 ;
  assign n23359 = ~n23357 & ~n23358 ;
  assign n23360 = ~n23356 & n23359 ;
  assign n23361 = n296 & n21143 ;
  assign n23362 = n23360 & ~n23361 ;
  assign n23363 = x5 & ~n23362 ;
  assign n23364 = x5 & ~n23363 ;
  assign n23365 = ~n23362 & ~n23363 ;
  assign n23366 = ~n23364 & ~n23365 ;
  assign n23367 = ~n23355 & ~n23366 ;
  assign n23368 = ~n23355 & ~n23367 ;
  assign n23369 = ~n23366 & ~n23367 ;
  assign n23370 = ~n23368 & ~n23369 ;
  assign n23371 = x123 & n146 ;
  assign n23372 = x121 & n182 ;
  assign n23373 = x122 & n141 ;
  assign n23374 = ~n23372 & ~n23373 ;
  assign n23375 = ~n23371 & n23374 ;
  assign n23376 = ~n22618 & ~n22620 ;
  assign n23377 = ~x122 & ~x123 ;
  assign n23378 = x122 & x123 ;
  assign n23379 = ~n23377 & ~n23378 ;
  assign n23380 = ~n23376 & n23379 ;
  assign n23381 = n23376 & ~n23379 ;
  assign n23382 = ~n23380 & ~n23381 ;
  assign n23383 = n149 & n23382 ;
  assign n23384 = n23375 & ~n23383 ;
  assign n23385 = x2 & ~n23384 ;
  assign n23386 = x2 & ~n23385 ;
  assign n23387 = ~n23384 & ~n23385 ;
  assign n23388 = ~n23386 & ~n23387 ;
  assign n23389 = ~n23370 & n23388 ;
  assign n23390 = n23370 & ~n23388 ;
  assign n23391 = ~n23389 & ~n23390 ;
  assign n23392 = ~n23018 & ~n23391 ;
  assign n23393 = ~n23018 & ~n23392 ;
  assign n23394 = ~n23391 & ~n23392 ;
  assign n23395 = ~n23393 & ~n23394 ;
  assign n23396 = ~n23017 & ~n23395 ;
  assign n23397 = n23017 & ~n23394 ;
  assign n23398 = ~n23393 & n23397 ;
  assign n23399 = ~n23396 & ~n23398 ;
  assign n23779 = n23399 & x187 ;
  assign n23400 = ~n23005 & ~n23010 ;
  assign n23401 = ~n22985 & ~n22987 ;
  assign n23402 = ~n22979 & ~n22981 ;
  assign n23403 = ~x117 & n574 ;
  assign n23404 = ~x115 & n673 ;
  assign n23405 = ~x116 & n569 ;
  assign n23406 = ~n23404 & ~n23405 ;
  assign n23407 = ~n23403 & n23406 ;
  assign n23408 = n577 & n19365 ;
  assign n23409 = n23407 & ~n23408 ;
  assign n23410 = ~x8 & ~n23409 ;
  assign n23411 = ~x8 & ~n23410 ;
  assign n23412 = ~n23409 & ~n23410 ;
  assign n23413 = ~n23411 & ~n23412 ;
  assign n23414 = ~n22973 & ~n22975 ;
  assign n23415 = ~n22967 & ~n22969 ;
  assign n23416 = ~n22928 & ~n22934 ;
  assign n23417 = ~n22872 & ~n22876 ;
  assign n23418 = ~n22676 & ~n22857 ;
  assign n23419 = ~n22854 & ~n23418 ;
  assign n23420 = ~n22816 & ~n22822 ;
  assign n23421 = ~n22778 & ~n22784 ;
  assign n23422 = ~x81 & n12506 ;
  assign n23423 = ~x79 & n13131 ;
  assign n23424 = ~x80 & n12501 ;
  assign n23425 = ~n23423 & ~n23424 ;
  assign n23426 = ~n23422 & n23425 ;
  assign n23427 = n2460 & n12509 ;
  assign n23428 = n23426 & ~n23427 ;
  assign n23429 = ~x44 & ~n23428 ;
  assign n23430 = ~x44 & ~n23429 ;
  assign n23431 = ~n23428 & ~n23429 ;
  assign n23432 = ~n23430 & ~n23431 ;
  assign n23433 = ~n22740 & ~n22746 ;
  assign n23434 = ~x75 & n16076 ;
  assign n23435 = ~x73 & n16756 ;
  assign n23436 = ~x74 & n16071 ;
  assign n23437 = ~n23435 & ~n23436 ;
  assign n23438 = ~n23434 & n23437 ;
  assign n23439 = n1225 & n16079 ;
  assign n23440 = n23438 & ~n23439 ;
  assign n23441 = ~x50 & ~n23440 ;
  assign n23442 = ~x50 & ~n23441 ;
  assign n23443 = ~n23440 & ~n23441 ;
  assign n23444 = ~n23442 & ~n23443 ;
  assign n23445 = ~n22724 & ~n22726 ;
  assign n23446 = ~n22718 & ~n22720 ;
  assign n23447 = ~x66 & n22325 ;
  assign n23448 = ~x64 & n23066 ;
  assign n23449 = ~x65 & n22320 ;
  assign n23450 = ~n23448 & ~n23449 ;
  assign n23451 = ~n23447 & n23450 ;
  assign n23452 = n214 & n22328 ;
  assign n23453 = n23451 & ~n23452 ;
  assign n23454 = ~x59 & ~n23453 ;
  assign n23455 = ~x59 & ~n23454 ;
  assign n23456 = ~n23453 & ~n23454 ;
  assign n23457 = ~n23455 & ~n23456 ;
  assign n23458 = ~n22714 & n23457 ;
  assign n23459 = n22714 & ~n23457 ;
  assign n23460 = ~n23458 & ~n23459 ;
  assign n23461 = ~x69 & n20143 ;
  assign n23462 = ~x67 & n20854 ;
  assign n23463 = ~x68 & n20138 ;
  assign n23464 = ~n23462 & ~n23463 ;
  assign n23465 = ~n23461 & n23464 ;
  assign n23466 = n435 & n20146 ;
  assign n23467 = n23465 & ~n23466 ;
  assign n23468 = ~x56 & ~n23467 ;
  assign n23469 = ~x56 & ~n23468 ;
  assign n23470 = ~n23467 & ~n23468 ;
  assign n23471 = ~n23469 & ~n23470 ;
  assign n23472 = n23460 & ~n23471 ;
  assign n23473 = ~n23460 & n23471 ;
  assign n23474 = ~n23446 & ~n23473 ;
  assign n23475 = ~n23472 & n23474 ;
  assign n23476 = ~n23446 & ~n23475 ;
  assign n23477 = ~n23472 & ~n23475 ;
  assign n23478 = ~n23473 & n23477 ;
  assign n23479 = ~n23476 & ~n23478 ;
  assign n23480 = ~x72 & n18025 ;
  assign n23481 = ~x70 & n18764 ;
  assign n23482 = ~x71 & n18020 ;
  assign n23483 = ~n23481 & ~n23482 ;
  assign n23484 = ~n23480 & n23483 ;
  assign n23485 = n773 & n18028 ;
  assign n23486 = n23484 & ~n23485 ;
  assign n23487 = ~x53 & ~n23486 ;
  assign n23488 = ~x53 & ~n23487 ;
  assign n23489 = ~n23486 & ~n23487 ;
  assign n23490 = ~n23488 & ~n23489 ;
  assign n23491 = n23479 & n23490 ;
  assign n23492 = ~n23479 & ~n23490 ;
  assign n23493 = ~n23491 & ~n23492 ;
  assign n23494 = ~n23445 & n23493 ;
  assign n23495 = n23445 & ~n23493 ;
  assign n23496 = ~n23494 & ~n23495 ;
  assign n23497 = n23444 & ~n23496 ;
  assign n23498 = ~n23444 & n23496 ;
  assign n23499 = ~n23497 & ~n23498 ;
  assign n23500 = ~n23433 & n23499 ;
  assign n23501 = n23433 & ~n23499 ;
  assign n23502 = ~n23500 & ~n23501 ;
  assign n23503 = ~x78 & n14233 ;
  assign n23504 = ~x76 & n14876 ;
  assign n23505 = ~x77 & n14228 ;
  assign n23506 = ~n23504 & ~n23505 ;
  assign n23507 = ~n23503 & n23506 ;
  assign n23508 = n1718 & n14236 ;
  assign n23509 = n23507 & ~n23508 ;
  assign n23510 = ~x47 & ~n23509 ;
  assign n23511 = ~x47 & ~n23510 ;
  assign n23512 = ~n23509 & ~n23510 ;
  assign n23513 = ~n23511 & ~n23512 ;
  assign n23514 = n23502 & ~n23513 ;
  assign n23515 = n23502 & ~n23514 ;
  assign n23516 = ~n23513 & ~n23514 ;
  assign n23517 = ~n23515 & ~n23516 ;
  assign n23518 = ~n22764 & ~n23517 ;
  assign n23519 = n22764 & n23517 ;
  assign n23520 = ~n23518 & ~n23519 ;
  assign n23521 = ~n23432 & n23520 ;
  assign n23522 = ~n23432 & ~n23521 ;
  assign n23523 = n23520 & ~n23521 ;
  assign n23524 = ~n23522 & ~n23523 ;
  assign n23525 = ~n23421 & ~n23524 ;
  assign n23526 = ~n23421 & ~n23525 ;
  assign n23527 = ~n23524 & ~n23525 ;
  assign n23528 = ~n23526 & ~n23527 ;
  assign n23529 = ~x84 & n10905 ;
  assign n23530 = ~x82 & n11466 ;
  assign n23531 = ~x83 & n10900 ;
  assign n23532 = ~n23530 & ~n23531 ;
  assign n23533 = ~n23529 & n23532 ;
  assign n23534 = n3247 & n10908 ;
  assign n23535 = n23533 & ~n23534 ;
  assign n23536 = ~x41 & ~n23535 ;
  assign n23537 = ~x41 & ~n23536 ;
  assign n23538 = ~n23535 & ~n23536 ;
  assign n23539 = ~n23537 & ~n23538 ;
  assign n23540 = ~n23528 & ~n23539 ;
  assign n23541 = ~n23528 & ~n23540 ;
  assign n23542 = ~n23539 & ~n23540 ;
  assign n23543 = ~n23541 & ~n23542 ;
  assign n23544 = ~n22802 & n23543 ;
  assign n23545 = n22802 & ~n23543 ;
  assign n23546 = ~n23544 & ~n23545 ;
  assign n23547 = ~x87 & n9433 ;
  assign n23548 = ~x85 & n9915 ;
  assign n23549 = ~x86 & n9428 ;
  assign n23550 = ~n23548 & ~n23549 ;
  assign n23551 = ~n23547 & n23550 ;
  assign n23552 = n4143 & n9436 ;
  assign n23553 = n23551 & ~n23552 ;
  assign n23554 = ~x38 & ~n23553 ;
  assign n23555 = ~x38 & ~n23554 ;
  assign n23556 = ~n23553 & ~n23554 ;
  assign n23557 = ~n23555 & ~n23556 ;
  assign n23558 = ~n23546 & ~n23557 ;
  assign n23559 = n23546 & n23557 ;
  assign n23560 = ~n23558 & ~n23559 ;
  assign n23561 = n23420 & ~n23560 ;
  assign n23562 = ~n23420 & n23560 ;
  assign n23563 = ~n23561 & ~n23562 ;
  assign n23564 = ~x90 & n8006 ;
  assign n23565 = ~x88 & n8474 ;
  assign n23566 = ~x89 & n8001 ;
  assign n23567 = ~n23565 & ~n23566 ;
  assign n23568 = ~n23564 & n23567 ;
  assign n23569 = n5155 & n8009 ;
  assign n23570 = n23568 & ~n23569 ;
  assign n23571 = ~x35 & ~n23570 ;
  assign n23572 = ~x35 & ~n23571 ;
  assign n23573 = ~n23570 & ~n23571 ;
  assign n23574 = ~n23572 & ~n23573 ;
  assign n23575 = n23563 & ~n23574 ;
  assign n23576 = n23563 & ~n23575 ;
  assign n23577 = ~n23574 & ~n23575 ;
  assign n23578 = ~n23576 & ~n23577 ;
  assign n23579 = ~n22835 & ~n22841 ;
  assign n23580 = n23578 & n23579 ;
  assign n23581 = ~n23578 & ~n23579 ;
  assign n23582 = ~n23580 & ~n23581 ;
  assign n23583 = ~x93 & n6725 ;
  assign n23584 = ~x91 & n7129 ;
  assign n23585 = ~x92 & n6720 ;
  assign n23586 = ~n23584 & ~n23585 ;
  assign n23587 = ~n23583 & n23586 ;
  assign n23588 = n6285 & n6728 ;
  assign n23589 = n23587 & ~n23588 ;
  assign n23590 = ~x32 & ~n23589 ;
  assign n23591 = ~x32 & ~n23590 ;
  assign n23592 = ~n23589 & ~n23590 ;
  assign n23593 = ~n23591 & ~n23592 ;
  assign n23594 = n23582 & ~n23593 ;
  assign n23595 = ~n23582 & n23593 ;
  assign n23596 = ~n23419 & ~n23595 ;
  assign n23597 = ~n23594 & n23596 ;
  assign n23598 = ~n23419 & ~n23597 ;
  assign n23599 = ~n23594 & ~n23597 ;
  assign n23600 = ~n23595 & n23599 ;
  assign n23601 = ~n23598 & ~n23600 ;
  assign n23602 = ~x96 & n5560 ;
  assign n23603 = ~x94 & n5943 ;
  assign n23604 = ~x95 & n5555 ;
  assign n23605 = ~n23603 & ~n23604 ;
  assign n23606 = ~n23602 & n23605 ;
  assign n23607 = n5563 & n7531 ;
  assign n23608 = n23606 & ~n23607 ;
  assign n23609 = ~x29 & ~n23608 ;
  assign n23610 = ~x29 & ~n23609 ;
  assign n23611 = ~n23608 & ~n23609 ;
  assign n23612 = ~n23610 & ~n23611 ;
  assign n23613 = n23601 & n23612 ;
  assign n23614 = ~n23601 & ~n23612 ;
  assign n23615 = ~n23613 & ~n23614 ;
  assign n23616 = ~n23417 & n23615 ;
  assign n23617 = n23417 & ~n23615 ;
  assign n23618 = ~n23616 & ~n23617 ;
  assign n23619 = ~x99 & n4531 ;
  assign n23620 = ~x97 & n4847 ;
  assign n23621 = ~x98 & n4526 ;
  assign n23622 = ~n23620 & ~n23621 ;
  assign n23623 = ~n23619 & n23622 ;
  assign n23624 = n4534 & n8885 ;
  assign n23625 = n23623 & ~n23624 ;
  assign n23626 = ~x26 & ~n23625 ;
  assign n23627 = ~x26 & ~n23626 ;
  assign n23628 = ~n23625 & ~n23626 ;
  assign n23629 = ~n23627 & ~n23628 ;
  assign n23630 = n23618 & ~n23629 ;
  assign n23631 = n23618 & ~n23630 ;
  assign n23632 = ~n23629 & ~n23630 ;
  assign n23633 = ~n23631 & ~n23632 ;
  assign n23634 = ~n22889 & ~n22896 ;
  assign n23635 = n23633 & n23634 ;
  assign n23636 = ~n23633 & ~n23634 ;
  assign n23637 = ~n23635 & ~n23636 ;
  assign n23638 = ~x102 & n3589 ;
  assign n23639 = ~x100 & n3878 ;
  assign n23640 = ~x101 & n3584 ;
  assign n23641 = ~n23639 & ~n23640 ;
  assign n23642 = ~n23638 & n23641 ;
  assign n23643 = n3592 & n10333 ;
  assign n23644 = n23642 & ~n23643 ;
  assign n23645 = ~x23 & ~n23644 ;
  assign n23646 = ~x23 & ~n23645 ;
  assign n23647 = ~n23644 & ~n23645 ;
  assign n23648 = ~n23646 & ~n23647 ;
  assign n23649 = n23637 & ~n23648 ;
  assign n23650 = n23637 & ~n23649 ;
  assign n23651 = ~n23648 & ~n23649 ;
  assign n23652 = ~n23650 & ~n23651 ;
  assign n23653 = ~n22909 & ~n22915 ;
  assign n23654 = n23652 & n23653 ;
  assign n23655 = ~n23652 & ~n23653 ;
  assign n23656 = ~n23654 & ~n23655 ;
  assign n23657 = ~x105 & n2751 ;
  assign n23658 = ~x103 & n3020 ;
  assign n23659 = ~x104 & n2746 ;
  assign n23660 = ~n23658 & ~n23659 ;
  assign n23661 = ~n23657 & n23660 ;
  assign n23662 = n2754 & n11907 ;
  assign n23663 = n23661 & ~n23662 ;
  assign n23664 = ~x20 & ~n23663 ;
  assign n23665 = ~x20 & ~n23664 ;
  assign n23666 = ~n23663 & ~n23664 ;
  assign n23667 = ~n23665 & ~n23666 ;
  assign n23668 = n23656 & ~n23667 ;
  assign n23669 = ~n23656 & n23667 ;
  assign n23670 = ~n23416 & ~n23669 ;
  assign n23671 = ~n23668 & n23670 ;
  assign n23672 = ~n23416 & ~n23671 ;
  assign n23673 = ~n23668 & ~n23671 ;
  assign n23674 = ~n23669 & n23673 ;
  assign n23675 = ~n23672 & ~n23674 ;
  assign n23676 = ~x108 & n2093 ;
  assign n23677 = ~x106 & n2275 ;
  assign n23678 = ~x107 & n2088 ;
  assign n23679 = ~n23677 & ~n23678 ;
  assign n23680 = ~n23676 & n23679 ;
  assign n23681 = n2096 & n13601 ;
  assign n23682 = n23680 & ~n23681 ;
  assign n23683 = ~x17 & ~n23682 ;
  assign n23684 = ~x17 & ~n23683 ;
  assign n23685 = ~n23682 & ~n23683 ;
  assign n23686 = ~n23684 & ~n23685 ;
  assign n23687 = ~n23675 & ~n23686 ;
  assign n23688 = ~n23675 & ~n23687 ;
  assign n23689 = ~n23686 & ~n23687 ;
  assign n23690 = ~n23688 & ~n23689 ;
  assign n23691 = ~n22952 & n23690 ;
  assign n23692 = n22952 & ~n23690 ;
  assign n23693 = ~n23691 & ~n23692 ;
  assign n23694 = ~x111 & n1434 ;
  assign n23695 = ~x109 & n1646 ;
  assign n23696 = ~x110 & n1429 ;
  assign n23697 = ~n23695 & ~n23696 ;
  assign n23698 = ~n23694 & n23697 ;
  assign n23699 = n1437 & n15411 ;
  assign n23700 = n23698 & ~n23699 ;
  assign n23701 = ~x14 & ~n23700 ;
  assign n23702 = ~x14 & ~n23701 ;
  assign n23703 = ~n23700 & ~n23701 ;
  assign n23704 = ~n23702 & ~n23703 ;
  assign n23705 = ~n23693 & ~n23704 ;
  assign n23706 = n23693 & n23704 ;
  assign n23707 = ~n23705 & ~n23706 ;
  assign n23708 = ~n23415 & n23707 ;
  assign n23709 = n23415 & ~n23707 ;
  assign n23710 = ~n23708 & ~n23709 ;
  assign n23711 = ~x114 & n945 ;
  assign n23712 = ~x112 & n1099 ;
  assign n23713 = ~x113 & n940 ;
  assign n23714 = ~n23712 & ~n23713 ;
  assign n23715 = ~n23711 & n23714 ;
  assign n23716 = n948 & n17333 ;
  assign n23717 = n23715 & ~n23716 ;
  assign n23718 = ~x11 & ~n23717 ;
  assign n23719 = ~x11 & ~n23718 ;
  assign n23720 = ~n23717 & ~n23718 ;
  assign n23721 = ~n23719 & ~n23720 ;
  assign n23722 = n23710 & ~n23721 ;
  assign n23723 = n23710 & ~n23722 ;
  assign n23724 = ~n23721 & ~n23722 ;
  assign n23725 = ~n23723 & ~n23724 ;
  assign n23726 = ~n23414 & ~n23725 ;
  assign n23727 = n23414 & n23725 ;
  assign n23728 = ~n23726 & ~n23727 ;
  assign n23729 = ~n23413 & n23728 ;
  assign n23730 = ~n23413 & ~n23729 ;
  assign n23731 = n23728 & ~n23729 ;
  assign n23732 = ~n23730 & ~n23731 ;
  assign n23733 = ~n23402 & ~n23732 ;
  assign n23734 = ~n23402 & ~n23733 ;
  assign n23735 = ~n23732 & ~n23733 ;
  assign n23736 = ~n23734 & ~n23735 ;
  assign n23737 = ~x120 & n293 ;
  assign n23738 = ~x118 & n373 ;
  assign n23739 = ~x119 & n288 ;
  assign n23740 = ~n23738 & ~n23739 ;
  assign n23741 = ~n23737 & n23740 ;
  assign n23742 = n296 & n21501 ;
  assign n23743 = n23741 & ~n23742 ;
  assign n23744 = ~x5 & ~n23743 ;
  assign n23745 = ~x5 & ~n23744 ;
  assign n23746 = ~n23743 & ~n23744 ;
  assign n23747 = ~n23745 & ~n23746 ;
  assign n23748 = ~n23736 & ~n23747 ;
  assign n23749 = ~n23736 & ~n23748 ;
  assign n23750 = ~n23747 & ~n23748 ;
  assign n23751 = ~n23749 & ~n23750 ;
  assign n23752 = ~x123 & n164 ;
  assign n23753 = ~x121 & n205 ;
  assign n23754 = ~x122 & n162 ;
  assign n23755 = ~n23753 & ~n23754 ;
  assign n23756 = ~n23752 & n23755 ;
  assign n23757 = ~n22617 & ~n22996 ;
  assign n23758 = n23379 & ~n23757 ;
  assign n23759 = ~n23379 & n23757 ;
  assign n23760 = ~n23758 & ~n23759 ;
  assign n23761 = n167 & n23760 ;
  assign n23762 = n23756 & ~n23761 ;
  assign n23763 = ~x2 & ~n23762 ;
  assign n23764 = ~x2 & ~n23763 ;
  assign n23765 = ~n23762 & ~n23763 ;
  assign n23766 = ~n23764 & ~n23765 ;
  assign n23767 = ~n23751 & n23766 ;
  assign n23768 = n23751 & ~n23766 ;
  assign n23769 = ~n23767 & ~n23768 ;
  assign n23770 = ~n23401 & ~n23769 ;
  assign n23771 = ~n23401 & ~n23770 ;
  assign n23772 = ~n23769 & ~n23770 ;
  assign n23773 = ~n23771 & ~n23772 ;
  assign n23774 = ~n23400 & ~n23773 ;
  assign n23775 = n23400 & ~n23772 ;
  assign n23776 = ~n23771 & n23775 ;
  assign n23777 = ~n23774 & ~n23776 ;
  assign n23780 = ~n23777 & ~x187 ;
  assign n23781 = ~n23779 & ~n23780 ;
  assign n23782 = ~n23392 & ~n23396 ;
  assign n23783 = ~n23370 & ~n23388 ;
  assign n23784 = ~n23367 & ~n23783 ;
  assign n23785 = x124 & n146 ;
  assign n23786 = x122 & n182 ;
  assign n23787 = x123 & n141 ;
  assign n23788 = ~n23786 & ~n23787 ;
  assign n23789 = ~n23785 & n23788 ;
  assign n23790 = ~n23378 & ~n23380 ;
  assign n23791 = ~x123 & ~x124 ;
  assign n23792 = x123 & x124 ;
  assign n23793 = ~n23791 & ~n23792 ;
  assign n23794 = ~n23790 & n23793 ;
  assign n23795 = n23790 & ~n23793 ;
  assign n23796 = ~n23794 & ~n23795 ;
  assign n23797 = n149 & n23796 ;
  assign n23798 = n23789 & ~n23797 ;
  assign n23799 = x2 & ~n23798 ;
  assign n23800 = x2 & ~n23799 ;
  assign n23801 = ~n23798 & ~n23799 ;
  assign n23802 = ~n23800 & ~n23801 ;
  assign n23803 = x121 & n293 ;
  assign n23804 = x119 & n373 ;
  assign n23805 = x120 & n288 ;
  assign n23806 = ~n23804 & ~n23805 ;
  assign n23807 = ~n23803 & n23806 ;
  assign n23808 = n296 & n21870 ;
  assign n23809 = n23807 & ~n23808 ;
  assign n23810 = x5 & ~n23809 ;
  assign n23811 = x5 & ~n23810 ;
  assign n23812 = ~n23809 & ~n23810 ;
  assign n23813 = ~n23811 & ~n23812 ;
  assign n23814 = ~n23348 & ~n23352 ;
  assign n23815 = x118 & n574 ;
  assign n23816 = x116 & n673 ;
  assign n23817 = x117 & n569 ;
  assign n23818 = ~n23816 & ~n23817 ;
  assign n23819 = ~n23815 & n23818 ;
  assign n23820 = n577 & n19395 ;
  assign n23821 = n23819 & ~n23820 ;
  assign n23822 = x8 & ~n23821 ;
  assign n23823 = x8 & ~n23822 ;
  assign n23824 = ~n23821 & ~n23822 ;
  assign n23825 = ~n23823 & ~n23824 ;
  assign n23826 = ~n23341 & ~n23345 ;
  assign n23827 = x115 & n945 ;
  assign n23828 = x113 & n1099 ;
  assign n23829 = x114 & n940 ;
  assign n23830 = ~n23828 & ~n23829 ;
  assign n23831 = ~n23827 & n23830 ;
  assign n23832 = n948 & n17364 ;
  assign n23833 = n23831 & ~n23832 ;
  assign n23834 = x11 & ~n23833 ;
  assign n23835 = x11 & ~n23834 ;
  assign n23836 = ~n23833 & ~n23834 ;
  assign n23837 = ~n23835 & ~n23836 ;
  assign n23838 = ~n23324 & ~n23327 ;
  assign n23839 = x112 & n1434 ;
  assign n23840 = x110 & n1646 ;
  assign n23841 = x111 & n1429 ;
  assign n23842 = ~n23840 & ~n23841 ;
  assign n23843 = ~n23839 & n23842 ;
  assign n23844 = n1437 & n15442 ;
  assign n23845 = n23843 & ~n23844 ;
  assign n23846 = x14 & ~n23845 ;
  assign n23847 = x14 & ~n23846 ;
  assign n23848 = ~n23845 & ~n23846 ;
  assign n23849 = ~n23847 & ~n23848 ;
  assign n23850 = ~n22573 & ~n23309 ;
  assign n23851 = ~n23306 & ~n23850 ;
  assign n23852 = x109 & n2093 ;
  assign n23853 = x107 & n2275 ;
  assign n23854 = x108 & n2088 ;
  assign n23855 = ~n23853 & ~n23854 ;
  assign n23856 = ~n23852 & n23855 ;
  assign n23857 = n2096 & n13894 ;
  assign n23858 = n23856 & ~n23857 ;
  assign n23859 = x17 & ~n23858 ;
  assign n23860 = x17 & ~n23859 ;
  assign n23861 = ~n23858 & ~n23859 ;
  assign n23862 = ~n23860 & ~n23861 ;
  assign n23863 = ~n23249 & ~n23255 ;
  assign n23864 = ~n23233 & ~n23235 ;
  assign n23865 = ~n22423 & ~n23162 ;
  assign n23866 = ~n23159 & ~n23865 ;
  assign n23867 = x85 & n10905 ;
  assign n23868 = x83 & n11466 ;
  assign n23869 = x84 & n10900 ;
  assign n23870 = ~n23868 & ~n23869 ;
  assign n23871 = ~n23867 & n23870 ;
  assign n23872 = n3389 & n10908 ;
  assign n23873 = n23871 & ~n23872 ;
  assign n23874 = x41 & ~n23873 ;
  assign n23875 = x41 & ~n23874 ;
  assign n23876 = ~n23873 & ~n23874 ;
  assign n23877 = ~n23875 & ~n23876 ;
  assign n23878 = ~n23140 & ~n23144 ;
  assign n23879 = x82 & n12506 ;
  assign n23880 = x80 & n13131 ;
  assign n23881 = x81 & n12501 ;
  assign n23882 = ~n23880 & ~n23881 ;
  assign n23883 = ~n23879 & n23882 ;
  assign n23884 = n2584 & n12509 ;
  assign n23885 = n23883 & ~n23884 ;
  assign n23886 = x44 & ~n23885 ;
  assign n23887 = x44 & ~n23886 ;
  assign n23888 = ~n23885 & ~n23886 ;
  assign n23889 = ~n23887 & ~n23888 ;
  assign n23890 = ~n23133 & ~n23137 ;
  assign n23891 = x79 & n14233 ;
  assign n23892 = x77 & n14876 ;
  assign n23893 = x78 & n14228 ;
  assign n23894 = ~n23892 & ~n23893 ;
  assign n23895 = ~n23891 & n23894 ;
  assign n23896 = n1817 & n14236 ;
  assign n23897 = n23895 & ~n23896 ;
  assign n23898 = x47 & ~n23897 ;
  assign n23899 = x47 & ~n23898 ;
  assign n23900 = ~n23897 & ~n23898 ;
  assign n23901 = ~n23899 & ~n23900 ;
  assign n23902 = ~n23117 & ~n23119 ;
  assign n23903 = x76 & n16076 ;
  assign n23904 = x74 & n16756 ;
  assign n23905 = x75 & n16071 ;
  assign n23906 = ~n23904 & ~n23905 ;
  assign n23907 = ~n23903 & n23906 ;
  assign n23908 = n1311 & n16079 ;
  assign n23909 = n23907 & ~n23908 ;
  assign n23910 = x50 & ~n23909 ;
  assign n23911 = x50 & ~n23910 ;
  assign n23912 = ~n23909 & ~n23910 ;
  assign n23913 = ~n23911 & ~n23912 ;
  assign n23914 = ~n23111 & ~n23113 ;
  assign n23915 = x59 & ~x60 ;
  assign n23916 = ~x59 & x60 ;
  assign n23917 = ~n23915 & ~n23916 ;
  assign n23918 = x64 & ~n23917 ;
  assign n23919 = ~n23078 & n23918 ;
  assign n23920 = n23078 & ~n23918 ;
  assign n23921 = ~n23919 & ~n23920 ;
  assign n23922 = x67 & n22325 ;
  assign n23923 = x65 & n23066 ;
  assign n23924 = x66 & n22320 ;
  assign n23925 = ~n23923 & ~n23924 ;
  assign n23926 = ~n23922 & n23925 ;
  assign n23927 = n240 & n22328 ;
  assign n23928 = n23926 & ~n23927 ;
  assign n23929 = x59 & ~n23928 ;
  assign n23930 = x59 & ~n23929 ;
  assign n23931 = ~n23928 & ~n23929 ;
  assign n23932 = ~n23930 & ~n23931 ;
  assign n23933 = ~n23921 & ~n23932 ;
  assign n23934 = n23921 & n23932 ;
  assign n23935 = ~n23933 & ~n23934 ;
  assign n23936 = x70 & n20143 ;
  assign n23937 = x68 & n20854 ;
  assign n23938 = x69 & n20138 ;
  assign n23939 = ~n23937 & ~n23938 ;
  assign n23940 = ~n23936 & n23939 ;
  assign n23941 = n488 & n20146 ;
  assign n23942 = n23940 & ~n23941 ;
  assign n23943 = x56 & ~n23942 ;
  assign n23944 = x56 & ~n23943 ;
  assign n23945 = ~n23942 & ~n23943 ;
  assign n23946 = ~n23944 & ~n23945 ;
  assign n23947 = n23935 & ~n23946 ;
  assign n23948 = n23935 & ~n23947 ;
  assign n23949 = ~n23946 & ~n23947 ;
  assign n23950 = ~n23948 & ~n23949 ;
  assign n23951 = ~n23096 & n23950 ;
  assign n23952 = n23096 & ~n23950 ;
  assign n23953 = ~n23951 & ~n23952 ;
  assign n23954 = x73 & n18025 ;
  assign n23955 = x71 & n18764 ;
  assign n23956 = x72 & n18020 ;
  assign n23957 = ~n23955 & ~n23956 ;
  assign n23958 = ~n23954 & n23957 ;
  assign n23959 = n843 & n18028 ;
  assign n23960 = n23958 & ~n23959 ;
  assign n23961 = x53 & ~n23960 ;
  assign n23962 = x53 & ~n23961 ;
  assign n23963 = ~n23960 & ~n23961 ;
  assign n23964 = ~n23962 & ~n23963 ;
  assign n23965 = ~n23953 & ~n23964 ;
  assign n23966 = n23953 & n23964 ;
  assign n23967 = ~n23965 & ~n23966 ;
  assign n23968 = ~n23914 & n23967 ;
  assign n23969 = n23914 & ~n23967 ;
  assign n23970 = ~n23968 & ~n23969 ;
  assign n23971 = n23913 & ~n23970 ;
  assign n23972 = ~n23913 & n23970 ;
  assign n23973 = ~n23971 & ~n23972 ;
  assign n23974 = ~n23902 & n23973 ;
  assign n23975 = n23902 & ~n23973 ;
  assign n23976 = ~n23974 & ~n23975 ;
  assign n23977 = ~n23901 & n23976 ;
  assign n23978 = n23901 & ~n23976 ;
  assign n23979 = ~n23977 & ~n23978 ;
  assign n23980 = ~n23890 & n23979 ;
  assign n23981 = n23890 & ~n23979 ;
  assign n23982 = ~n23980 & ~n23981 ;
  assign n23983 = ~n23889 & n23982 ;
  assign n23984 = ~n23889 & ~n23983 ;
  assign n23985 = n23982 & ~n23983 ;
  assign n23986 = ~n23984 & ~n23985 ;
  assign n23987 = ~n23878 & ~n23986 ;
  assign n23988 = n23878 & ~n23985 ;
  assign n23989 = ~n23984 & n23988 ;
  assign n23990 = ~n23987 & ~n23989 ;
  assign n23991 = ~n23877 & n23990 ;
  assign n23992 = n23877 & ~n23990 ;
  assign n23993 = ~n23991 & ~n23992 ;
  assign n23994 = ~n23866 & n23993 ;
  assign n23995 = n23866 & ~n23993 ;
  assign n23996 = ~n23994 & ~n23995 ;
  assign n23997 = x88 & n9433 ;
  assign n23998 = x86 & n9915 ;
  assign n23999 = x87 & n9428 ;
  assign n24000 = ~n23998 & ~n23999 ;
  assign n24001 = ~n23997 & n24000 ;
  assign n24002 = n4305 & n9436 ;
  assign n24003 = n24001 & ~n24002 ;
  assign n24004 = x38 & ~n24003 ;
  assign n24005 = x38 & ~n24004 ;
  assign n24006 = ~n24003 & ~n24004 ;
  assign n24007 = ~n24005 & ~n24006 ;
  assign n24008 = n23996 & ~n24007 ;
  assign n24009 = n23996 & ~n24008 ;
  assign n24010 = ~n24007 & ~n24008 ;
  assign n24011 = ~n24009 & ~n24010 ;
  assign n24012 = ~n23177 & ~n23181 ;
  assign n24013 = n24011 & n24012 ;
  assign n24014 = ~n24011 & ~n24012 ;
  assign n24015 = ~n24013 & ~n24014 ;
  assign n24016 = x91 & n8006 ;
  assign n24017 = x89 & n8474 ;
  assign n24018 = x90 & n8001 ;
  assign n24019 = ~n24017 & ~n24018 ;
  assign n24020 = ~n24016 & n24019 ;
  assign n24021 = n5336 & n8009 ;
  assign n24022 = n24020 & ~n24021 ;
  assign n24023 = x35 & ~n24022 ;
  assign n24024 = x35 & ~n24023 ;
  assign n24025 = ~n24022 & ~n24023 ;
  assign n24026 = ~n24024 & ~n24025 ;
  assign n24027 = n24015 & ~n24026 ;
  assign n24028 = n24015 & ~n24027 ;
  assign n24029 = ~n24026 & ~n24027 ;
  assign n24030 = ~n24028 & ~n24029 ;
  assign n24031 = ~n23194 & ~n23200 ;
  assign n24032 = n24030 & n24031 ;
  assign n24033 = ~n24030 & ~n24031 ;
  assign n24034 = ~n24032 & ~n24033 ;
  assign n24035 = x94 & n6725 ;
  assign n24036 = x92 & n7129 ;
  assign n24037 = x93 & n6720 ;
  assign n24038 = ~n24036 & ~n24037 ;
  assign n24039 = ~n24035 & n24038 ;
  assign n24040 = n6483 & n6728 ;
  assign n24041 = n24039 & ~n24040 ;
  assign n24042 = x32 & ~n24041 ;
  assign n24043 = x32 & ~n24042 ;
  assign n24044 = ~n24041 & ~n24042 ;
  assign n24045 = ~n24043 & ~n24044 ;
  assign n24046 = ~n24034 & n24045 ;
  assign n24047 = n24034 & ~n24045 ;
  assign n24048 = ~n24046 & ~n24047 ;
  assign n24049 = ~n23218 & n24048 ;
  assign n24050 = n23218 & ~n24048 ;
  assign n24051 = ~n24049 & ~n24050 ;
  assign n24052 = x97 & n5560 ;
  assign n24053 = x95 & n5943 ;
  assign n24054 = x96 & n5555 ;
  assign n24055 = ~n24053 & ~n24054 ;
  assign n24056 = ~n24052 & n24055 ;
  assign n24057 = n5563 & n7745 ;
  assign n24058 = n24056 & ~n24057 ;
  assign n24059 = x29 & ~n24058 ;
  assign n24060 = x29 & ~n24059 ;
  assign n24061 = ~n24058 & ~n24059 ;
  assign n24062 = ~n24060 & ~n24061 ;
  assign n24063 = n24051 & ~n24062 ;
  assign n24064 = n24051 & ~n24063 ;
  assign n24065 = ~n24062 & ~n24063 ;
  assign n24066 = ~n24064 & ~n24065 ;
  assign n24067 = ~n23864 & n24066 ;
  assign n24068 = n23864 & ~n24066 ;
  assign n24069 = ~n24067 & ~n24068 ;
  assign n24070 = x100 & n4531 ;
  assign n24071 = x98 & n4847 ;
  assign n24072 = x99 & n4526 ;
  assign n24073 = ~n24071 & ~n24072 ;
  assign n24074 = ~n24070 & n24073 ;
  assign n24075 = n4534 & n9115 ;
  assign n24076 = n24074 & ~n24075 ;
  assign n24077 = x26 & ~n24076 ;
  assign n24078 = x26 & ~n24077 ;
  assign n24079 = ~n24076 & ~n24077 ;
  assign n24080 = ~n24078 & ~n24079 ;
  assign n24081 = ~n24069 & ~n24080 ;
  assign n24082 = n24069 & n24080 ;
  assign n24083 = ~n24081 & ~n24082 ;
  assign n24084 = n23863 & ~n24083 ;
  assign n24085 = ~n23863 & n24083 ;
  assign n24086 = ~n24084 & ~n24085 ;
  assign n24087 = x103 & n3589 ;
  assign n24088 = x101 & n3878 ;
  assign n24089 = x102 & n3584 ;
  assign n24090 = ~n24088 & ~n24089 ;
  assign n24091 = ~n24087 & n24090 ;
  assign n24092 = n3592 & n10588 ;
  assign n24093 = n24091 & ~n24092 ;
  assign n24094 = x23 & ~n24093 ;
  assign n24095 = x23 & ~n24094 ;
  assign n24096 = ~n24093 & ~n24094 ;
  assign n24097 = ~n24095 & ~n24096 ;
  assign n24098 = n24086 & ~n24097 ;
  assign n24099 = n24086 & ~n24098 ;
  assign n24100 = ~n24097 & ~n24098 ;
  assign n24101 = ~n24099 & ~n24100 ;
  assign n24102 = ~n23268 & ~n23274 ;
  assign n24103 = n24101 & n24102 ;
  assign n24104 = ~n24101 & ~n24102 ;
  assign n24105 = ~n24103 & ~n24104 ;
  assign n24106 = x106 & n2751 ;
  assign n24107 = x104 & n3020 ;
  assign n24108 = x105 & n2746 ;
  assign n24109 = ~n24107 & ~n24108 ;
  assign n24110 = ~n24106 & n24109 ;
  assign n24111 = n2754 & n12181 ;
  assign n24112 = n24110 & ~n24111 ;
  assign n24113 = x20 & ~n24112 ;
  assign n24114 = x20 & ~n24113 ;
  assign n24115 = ~n24112 & ~n24113 ;
  assign n24116 = ~n24114 & ~n24115 ;
  assign n24117 = ~n24105 & n24116 ;
  assign n24118 = n24105 & ~n24116 ;
  assign n24119 = ~n24117 & ~n24118 ;
  assign n24120 = ~n23292 & n24119 ;
  assign n24121 = n23292 & ~n24119 ;
  assign n24122 = ~n24120 & ~n24121 ;
  assign n24123 = ~n23862 & n24122 ;
  assign n24124 = ~n23862 & ~n24123 ;
  assign n24125 = n24122 & ~n24123 ;
  assign n24126 = ~n24124 & ~n24125 ;
  assign n24127 = ~n23851 & ~n24126 ;
  assign n24128 = n23851 & ~n24125 ;
  assign n24129 = ~n24124 & n24128 ;
  assign n24130 = ~n24127 & ~n24129 ;
  assign n24131 = ~n23849 & n24130 ;
  assign n24132 = ~n23849 & ~n24131 ;
  assign n24133 = n24130 & ~n24131 ;
  assign n24134 = ~n24132 & ~n24133 ;
  assign n24135 = ~n23838 & ~n24134 ;
  assign n24136 = n23838 & ~n24133 ;
  assign n24137 = ~n24132 & n24136 ;
  assign n24138 = ~n24135 & ~n24137 ;
  assign n24139 = ~n23837 & n24138 ;
  assign n24140 = ~n23837 & ~n24139 ;
  assign n24141 = n24138 & ~n24139 ;
  assign n24142 = ~n24140 & ~n24141 ;
  assign n24143 = ~n23826 & ~n24142 ;
  assign n24144 = n23826 & ~n24141 ;
  assign n24145 = ~n24140 & n24144 ;
  assign n24146 = ~n24143 & ~n24145 ;
  assign n24147 = ~n23825 & n24146 ;
  assign n24148 = n23825 & ~n24146 ;
  assign n24149 = ~n24147 & ~n24148 ;
  assign n24150 = ~n23814 & n24149 ;
  assign n24151 = n23814 & ~n24149 ;
  assign n24152 = ~n24150 & ~n24151 ;
  assign n24153 = ~n23813 & n24152 ;
  assign n24154 = n23813 & ~n24152 ;
  assign n24155 = ~n24153 & ~n24154 ;
  assign n24156 = ~n23802 & n24155 ;
  assign n24157 = n23802 & ~n24155 ;
  assign n24158 = ~n24156 & ~n24157 ;
  assign n24159 = ~n23784 & n24158 ;
  assign n24160 = n23784 & ~n24158 ;
  assign n24161 = ~n24159 & ~n24160 ;
  assign n24162 = ~n23782 & n24161 ;
  assign n24163 = n23782 & ~n24161 ;
  assign n24164 = ~n24162 & ~n24163 ;
  assign n24543 = n24164 & x188 ;
  assign n24165 = ~n23770 & ~n23774 ;
  assign n24166 = ~n23751 & ~n23766 ;
  assign n24167 = ~n23748 & ~n24166 ;
  assign n24168 = ~x124 & n164 ;
  assign n24169 = ~x122 & n205 ;
  assign n24170 = ~x123 & n162 ;
  assign n24171 = ~n24169 & ~n24170 ;
  assign n24172 = ~n24168 & n24171 ;
  assign n24173 = ~n23377 & ~n23758 ;
  assign n24174 = n23793 & ~n24173 ;
  assign n24175 = ~n23793 & n24173 ;
  assign n24176 = ~n24174 & ~n24175 ;
  assign n24177 = n167 & n24176 ;
  assign n24178 = n24172 & ~n24177 ;
  assign n24179 = ~x2 & ~n24178 ;
  assign n24180 = ~x2 & ~n24179 ;
  assign n24181 = ~n24178 & ~n24179 ;
  assign n24182 = ~n24180 & ~n24181 ;
  assign n24183 = ~x121 & n293 ;
  assign n24184 = ~x119 & n373 ;
  assign n24185 = ~x120 & n288 ;
  assign n24186 = ~n24184 & ~n24185 ;
  assign n24187 = ~n24183 & n24186 ;
  assign n24188 = n296 & n22229 ;
  assign n24189 = n24187 & ~n24188 ;
  assign n24190 = ~x5 & ~n24189 ;
  assign n24191 = ~x5 & ~n24190 ;
  assign n24192 = ~n24189 & ~n24190 ;
  assign n24193 = ~n24191 & ~n24192 ;
  assign n24194 = ~n23729 & ~n23733 ;
  assign n24195 = ~x118 & n574 ;
  assign n24196 = ~x116 & n673 ;
  assign n24197 = ~x117 & n569 ;
  assign n24198 = ~n24196 & ~n24197 ;
  assign n24199 = ~n24195 & n24198 ;
  assign n24200 = n577 & n19736 ;
  assign n24201 = n24199 & ~n24200 ;
  assign n24202 = ~x8 & ~n24201 ;
  assign n24203 = ~x8 & ~n24202 ;
  assign n24204 = ~n24201 & ~n24202 ;
  assign n24205 = ~n24203 & ~n24204 ;
  assign n24206 = ~n23722 & ~n23726 ;
  assign n24207 = ~x115 & n945 ;
  assign n24208 = ~x113 & n1099 ;
  assign n24209 = ~x114 & n940 ;
  assign n24210 = ~n24208 & ~n24209 ;
  assign n24211 = ~n24207 & n24210 ;
  assign n24212 = n948 & n17683 ;
  assign n24213 = n24211 & ~n24212 ;
  assign n24214 = ~x11 & ~n24213 ;
  assign n24215 = ~x11 & ~n24214 ;
  assign n24216 = ~n24213 & ~n24214 ;
  assign n24217 = ~n24215 & ~n24216 ;
  assign n24218 = ~n23705 & ~n23708 ;
  assign n24219 = ~x112 & n1434 ;
  assign n24220 = ~x110 & n1646 ;
  assign n24221 = ~x111 & n1429 ;
  assign n24222 = ~n24220 & ~n24221 ;
  assign n24223 = ~n24219 & n24222 ;
  assign n24224 = n1437 & n15744 ;
  assign n24225 = n24223 & ~n24224 ;
  assign n24226 = ~x14 & ~n24225 ;
  assign n24227 = ~x14 & ~n24226 ;
  assign n24228 = ~n24225 & ~n24226 ;
  assign n24229 = ~n24227 & ~n24228 ;
  assign n24230 = ~n22952 & ~n23690 ;
  assign n24231 = ~n23687 & ~n24230 ;
  assign n24232 = ~x109 & n2093 ;
  assign n24233 = ~x107 & n2275 ;
  assign n24234 = ~x108 & n2088 ;
  assign n24235 = ~n24233 & ~n24234 ;
  assign n24236 = ~n24232 & n24235 ;
  assign n24237 = n2096 & n14177 ;
  assign n24238 = n24236 & ~n24237 ;
  assign n24239 = ~x17 & ~n24238 ;
  assign n24240 = ~x17 & ~n24239 ;
  assign n24241 = ~n24238 & ~n24239 ;
  assign n24242 = ~n24240 & ~n24241 ;
  assign n24243 = ~n23630 & ~n23636 ;
  assign n24244 = ~n23614 & ~n23616 ;
  assign n24245 = ~n22802 & ~n23543 ;
  assign n24246 = ~n23540 & ~n24245 ;
  assign n24247 = ~x85 & n10905 ;
  assign n24248 = ~x83 & n11466 ;
  assign n24249 = ~x84 & n10900 ;
  assign n24250 = ~n24248 & ~n24249 ;
  assign n24251 = ~n24247 & n24250 ;
  assign n24252 = n3521 & n10908 ;
  assign n24253 = n24251 & ~n24252 ;
  assign n24254 = ~x41 & ~n24253 ;
  assign n24255 = ~x41 & ~n24254 ;
  assign n24256 = ~n24253 & ~n24254 ;
  assign n24257 = ~n24255 & ~n24256 ;
  assign n24258 = ~n23521 & ~n23525 ;
  assign n24259 = ~x82 & n12506 ;
  assign n24260 = ~x80 & n13131 ;
  assign n24261 = ~x81 & n12501 ;
  assign n24262 = ~n24260 & ~n24261 ;
  assign n24263 = ~n24259 & n24262 ;
  assign n24264 = n2697 & n12509 ;
  assign n24265 = n24263 & ~n24264 ;
  assign n24266 = ~x44 & ~n24265 ;
  assign n24267 = ~x44 & ~n24266 ;
  assign n24268 = ~n24265 & ~n24266 ;
  assign n24269 = ~n24267 & ~n24268 ;
  assign n24270 = ~n23514 & ~n23518 ;
  assign n24271 = ~x79 & n14233 ;
  assign n24272 = ~x77 & n14876 ;
  assign n24273 = ~x78 & n14228 ;
  assign n24274 = ~n24272 & ~n24273 ;
  assign n24275 = ~n24271 & n24274 ;
  assign n24276 = n1921 & n14236 ;
  assign n24277 = n24275 & ~n24276 ;
  assign n24278 = ~x47 & ~n24277 ;
  assign n24279 = ~x47 & ~n24278 ;
  assign n24280 = ~n24277 & ~n24278 ;
  assign n24281 = ~n24279 & ~n24280 ;
  assign n24282 = ~n23498 & ~n23500 ;
  assign n24283 = ~x76 & n16076 ;
  assign n24284 = ~x74 & n16756 ;
  assign n24285 = ~x75 & n16071 ;
  assign n24286 = ~n24284 & ~n24285 ;
  assign n24287 = ~n24283 & n24286 ;
  assign n24288 = n1390 & n16079 ;
  assign n24289 = n24287 & ~n24288 ;
  assign n24290 = ~x50 & ~n24289 ;
  assign n24291 = ~x50 & ~n24290 ;
  assign n24292 = ~n24289 & ~n24290 ;
  assign n24293 = ~n24291 & ~n24292 ;
  assign n24294 = ~n23492 & ~n23494 ;
  assign n24295 = ~x64 & ~n23917 ;
  assign n24296 = ~n23459 & n24295 ;
  assign n24297 = n23459 & ~n24295 ;
  assign n24298 = ~n24296 & ~n24297 ;
  assign n24299 = ~x67 & n22325 ;
  assign n24300 = ~x65 & n23066 ;
  assign n24301 = ~x66 & n22320 ;
  assign n24302 = ~n24300 & ~n24301 ;
  assign n24303 = ~n24299 & n24302 ;
  assign n24304 = n266 & n22328 ;
  assign n24305 = n24303 & ~n24304 ;
  assign n24306 = ~x59 & ~n24305 ;
  assign n24307 = ~x59 & ~n24306 ;
  assign n24308 = ~n24305 & ~n24306 ;
  assign n24309 = ~n24307 & ~n24308 ;
  assign n24310 = ~n24298 & ~n24309 ;
  assign n24311 = n24298 & n24309 ;
  assign n24312 = ~n24310 & ~n24311 ;
  assign n24313 = ~x70 & n20143 ;
  assign n24314 = ~x68 & n20854 ;
  assign n24315 = ~x69 & n20138 ;
  assign n24316 = ~n24314 & ~n24315 ;
  assign n24317 = ~n24313 & n24316 ;
  assign n24318 = n529 & n20146 ;
  assign n24319 = n24317 & ~n24318 ;
  assign n24320 = ~x56 & ~n24319 ;
  assign n24321 = ~x56 & ~n24320 ;
  assign n24322 = ~n24319 & ~n24320 ;
  assign n24323 = ~n24321 & ~n24322 ;
  assign n24324 = n24312 & ~n24323 ;
  assign n24325 = n24312 & ~n24324 ;
  assign n24326 = ~n24323 & ~n24324 ;
  assign n24327 = ~n24325 & ~n24326 ;
  assign n24328 = ~n23477 & n24327 ;
  assign n24329 = n23477 & ~n24327 ;
  assign n24330 = ~n24328 & ~n24329 ;
  assign n24331 = ~x73 & n18025 ;
  assign n24332 = ~x71 & n18764 ;
  assign n24333 = ~x72 & n18020 ;
  assign n24334 = ~n24332 & ~n24333 ;
  assign n24335 = ~n24331 & n24334 ;
  assign n24336 = n903 & n18028 ;
  assign n24337 = n24335 & ~n24336 ;
  assign n24338 = ~x53 & ~n24337 ;
  assign n24339 = ~x53 & ~n24338 ;
  assign n24340 = ~n24337 & ~n24338 ;
  assign n24341 = ~n24339 & ~n24340 ;
  assign n24342 = ~n24330 & ~n24341 ;
  assign n24343 = n24330 & n24341 ;
  assign n24344 = ~n24342 & ~n24343 ;
  assign n24345 = ~n24294 & n24344 ;
  assign n24346 = n24294 & ~n24344 ;
  assign n24347 = ~n24345 & ~n24346 ;
  assign n24348 = n24293 & ~n24347 ;
  assign n24349 = ~n24293 & n24347 ;
  assign n24350 = ~n24348 & ~n24349 ;
  assign n24351 = ~n24282 & n24350 ;
  assign n24352 = n24282 & ~n24350 ;
  assign n24353 = ~n24351 & ~n24352 ;
  assign n24354 = ~n24281 & n24353 ;
  assign n24355 = n24281 & ~n24353 ;
  assign n24356 = ~n24354 & ~n24355 ;
  assign n24357 = ~n24270 & n24356 ;
  assign n24358 = n24270 & ~n24356 ;
  assign n24359 = ~n24357 & ~n24358 ;
  assign n24360 = ~n24269 & n24359 ;
  assign n24361 = ~n24269 & ~n24360 ;
  assign n24362 = n24359 & ~n24360 ;
  assign n24363 = ~n24361 & ~n24362 ;
  assign n24364 = ~n24258 & ~n24363 ;
  assign n24365 = n24258 & ~n24362 ;
  assign n24366 = ~n24361 & n24365 ;
  assign n24367 = ~n24364 & ~n24366 ;
  assign n24368 = ~n24257 & n24367 ;
  assign n24369 = n24257 & ~n24367 ;
  assign n24370 = ~n24368 & ~n24369 ;
  assign n24371 = ~n24246 & n24370 ;
  assign n24372 = n24246 & ~n24370 ;
  assign n24373 = ~n24371 & ~n24372 ;
  assign n24374 = ~x88 & n9433 ;
  assign n24375 = ~x86 & n9915 ;
  assign n24376 = ~x87 & n9428 ;
  assign n24377 = ~n24375 & ~n24376 ;
  assign n24378 = ~n24374 & n24377 ;
  assign n24379 = n4457 & n9436 ;
  assign n24380 = n24378 & ~n24379 ;
  assign n24381 = ~x38 & ~n24380 ;
  assign n24382 = ~x38 & ~n24381 ;
  assign n24383 = ~n24380 & ~n24381 ;
  assign n24384 = ~n24382 & ~n24383 ;
  assign n24385 = n24373 & ~n24384 ;
  assign n24386 = n24373 & ~n24385 ;
  assign n24387 = ~n24384 & ~n24385 ;
  assign n24388 = ~n24386 & ~n24387 ;
  assign n24389 = ~n23558 & ~n23562 ;
  assign n24390 = n24388 & n24389 ;
  assign n24391 = ~n24388 & ~n24389 ;
  assign n24392 = ~n24390 & ~n24391 ;
  assign n24393 = ~x91 & n8006 ;
  assign n24394 = ~x89 & n8474 ;
  assign n24395 = ~x90 & n8001 ;
  assign n24396 = ~n24394 & ~n24395 ;
  assign n24397 = ~n24393 & n24396 ;
  assign n24398 = n5507 & n8009 ;
  assign n24399 = n24397 & ~n24398 ;
  assign n24400 = ~x35 & ~n24399 ;
  assign n24401 = ~x35 & ~n24400 ;
  assign n24402 = ~n24399 & ~n24400 ;
  assign n24403 = ~n24401 & ~n24402 ;
  assign n24404 = n24392 & ~n24403 ;
  assign n24405 = n24392 & ~n24404 ;
  assign n24406 = ~n24403 & ~n24404 ;
  assign n24407 = ~n24405 & ~n24406 ;
  assign n24408 = ~n23575 & ~n23581 ;
  assign n24409 = n24407 & n24408 ;
  assign n24410 = ~n24407 & ~n24408 ;
  assign n24411 = ~n24409 & ~n24410 ;
  assign n24412 = ~x94 & n6725 ;
  assign n24413 = ~x92 & n7129 ;
  assign n24414 = ~x93 & n6720 ;
  assign n24415 = ~n24413 & ~n24414 ;
  assign n24416 = ~n24412 & n24415 ;
  assign n24417 = n6671 & n6728 ;
  assign n24418 = n24416 & ~n24417 ;
  assign n24419 = ~x32 & ~n24418 ;
  assign n24420 = ~x32 & ~n24419 ;
  assign n24421 = ~n24418 & ~n24419 ;
  assign n24422 = ~n24420 & ~n24421 ;
  assign n24423 = ~n24411 & n24422 ;
  assign n24424 = n24411 & ~n24422 ;
  assign n24425 = ~n24423 & ~n24424 ;
  assign n24426 = ~n23599 & n24425 ;
  assign n24427 = n23599 & ~n24425 ;
  assign n24428 = ~n24426 & ~n24427 ;
  assign n24429 = ~x97 & n5560 ;
  assign n24430 = ~x95 & n5943 ;
  assign n24431 = ~x96 & n5555 ;
  assign n24432 = ~n24430 & ~n24431 ;
  assign n24433 = ~n24429 & n24432 ;
  assign n24434 = n5563 & n7949 ;
  assign n24435 = n24433 & ~n24434 ;
  assign n24436 = ~x29 & ~n24435 ;
  assign n24437 = ~x29 & ~n24436 ;
  assign n24438 = ~n24435 & ~n24436 ;
  assign n24439 = ~n24437 & ~n24438 ;
  assign n24440 = n24428 & ~n24439 ;
  assign n24441 = n24428 & ~n24440 ;
  assign n24442 = ~n24439 & ~n24440 ;
  assign n24443 = ~n24441 & ~n24442 ;
  assign n24444 = ~n24244 & n24443 ;
  assign n24445 = n24244 & ~n24443 ;
  assign n24446 = ~n24444 & ~n24445 ;
  assign n24447 = ~x100 & n4531 ;
  assign n24448 = ~x98 & n4847 ;
  assign n24449 = ~x99 & n4526 ;
  assign n24450 = ~n24448 & ~n24449 ;
  assign n24451 = ~n24447 & n24450 ;
  assign n24452 = n4534 & n9338 ;
  assign n24453 = n24451 & ~n24452 ;
  assign n24454 = ~x26 & ~n24453 ;
  assign n24455 = ~x26 & ~n24454 ;
  assign n24456 = ~n24453 & ~n24454 ;
  assign n24457 = ~n24455 & ~n24456 ;
  assign n24458 = ~n24446 & ~n24457 ;
  assign n24459 = n24446 & n24457 ;
  assign n24460 = ~n24458 & ~n24459 ;
  assign n24461 = n24243 & ~n24460 ;
  assign n24462 = ~n24243 & n24460 ;
  assign n24463 = ~n24461 & ~n24462 ;
  assign n24464 = ~x103 & n3589 ;
  assign n24465 = ~x101 & n3878 ;
  assign n24466 = ~x102 & n3584 ;
  assign n24467 = ~n24465 & ~n24466 ;
  assign n24468 = ~n24464 & n24467 ;
  assign n24469 = n3592 & n10833 ;
  assign n24470 = n24468 & ~n24469 ;
  assign n24471 = ~x23 & ~n24470 ;
  assign n24472 = ~x23 & ~n24471 ;
  assign n24473 = ~n24470 & ~n24471 ;
  assign n24474 = ~n24472 & ~n24473 ;
  assign n24475 = n24463 & ~n24474 ;
  assign n24476 = n24463 & ~n24475 ;
  assign n24477 = ~n24474 & ~n24475 ;
  assign n24478 = ~n24476 & ~n24477 ;
  assign n24479 = ~n23649 & ~n23655 ;
  assign n24480 = n24478 & n24479 ;
  assign n24481 = ~n24478 & ~n24479 ;
  assign n24482 = ~n24480 & ~n24481 ;
  assign n24483 = ~x106 & n2751 ;
  assign n24484 = ~x104 & n3020 ;
  assign n24485 = ~x105 & n2746 ;
  assign n24486 = ~n24484 & ~n24485 ;
  assign n24487 = ~n24483 & n24486 ;
  assign n24488 = n2754 & n12447 ;
  assign n24489 = n24487 & ~n24488 ;
  assign n24490 = ~x20 & ~n24489 ;
  assign n24491 = ~x20 & ~n24490 ;
  assign n24492 = ~n24489 & ~n24490 ;
  assign n24493 = ~n24491 & ~n24492 ;
  assign n24494 = ~n24482 & n24493 ;
  assign n24495 = n24482 & ~n24493 ;
  assign n24496 = ~n24494 & ~n24495 ;
  assign n24497 = ~n23673 & n24496 ;
  assign n24498 = n23673 & ~n24496 ;
  assign n24499 = ~n24497 & ~n24498 ;
  assign n24500 = ~n24242 & n24499 ;
  assign n24501 = ~n24242 & ~n24500 ;
  assign n24502 = n24499 & ~n24500 ;
  assign n24503 = ~n24501 & ~n24502 ;
  assign n24504 = ~n24231 & ~n24503 ;
  assign n24505 = n24231 & ~n24502 ;
  assign n24506 = ~n24501 & n24505 ;
  assign n24507 = ~n24504 & ~n24506 ;
  assign n24508 = ~n24229 & n24507 ;
  assign n24509 = ~n24229 & ~n24508 ;
  assign n24510 = n24507 & ~n24508 ;
  assign n24511 = ~n24509 & ~n24510 ;
  assign n24512 = ~n24218 & ~n24511 ;
  assign n24513 = n24218 & ~n24510 ;
  assign n24514 = ~n24509 & n24513 ;
  assign n24515 = ~n24512 & ~n24514 ;
  assign n24516 = ~n24217 & n24515 ;
  assign n24517 = ~n24217 & ~n24516 ;
  assign n24518 = n24515 & ~n24516 ;
  assign n24519 = ~n24517 & ~n24518 ;
  assign n24520 = ~n24206 & ~n24519 ;
  assign n24521 = n24206 & ~n24518 ;
  assign n24522 = ~n24517 & n24521 ;
  assign n24523 = ~n24520 & ~n24522 ;
  assign n24524 = ~n24205 & n24523 ;
  assign n24525 = n24205 & ~n24523 ;
  assign n24526 = ~n24524 & ~n24525 ;
  assign n24527 = ~n24194 & n24526 ;
  assign n24528 = n24194 & ~n24526 ;
  assign n24529 = ~n24527 & ~n24528 ;
  assign n24530 = ~n24193 & n24529 ;
  assign n24531 = n24193 & ~n24529 ;
  assign n24532 = ~n24530 & ~n24531 ;
  assign n24533 = ~n24182 & n24532 ;
  assign n24534 = n24182 & ~n24532 ;
  assign n24535 = ~n24533 & ~n24534 ;
  assign n24536 = ~n24167 & n24535 ;
  assign n24537 = n24167 & ~n24535 ;
  assign n24538 = ~n24536 & ~n24537 ;
  assign n24539 = ~n24165 & n24538 ;
  assign n24540 = n24165 & ~n24538 ;
  assign n24541 = ~n24539 & ~n24540 ;
  assign n24544 = ~n24541 & ~x188 ;
  assign n24545 = ~n24543 & ~n24544 ;
  assign n24546 = ~n24139 & ~n24143 ;
  assign n24547 = x116 & n945 ;
  assign n24548 = x114 & n1099 ;
  assign n24549 = x115 & n940 ;
  assign n24550 = ~n24548 & ~n24549 ;
  assign n24551 = ~n24547 & n24550 ;
  assign n24552 = n948 & n18336 ;
  assign n24553 = n24551 & ~n24552 ;
  assign n24554 = x11 & ~n24553 ;
  assign n24555 = x11 & ~n24554 ;
  assign n24556 = ~n24553 & ~n24554 ;
  assign n24557 = ~n24555 & ~n24556 ;
  assign n24558 = ~n24131 & ~n24135 ;
  assign n24559 = x113 & n1434 ;
  assign n24560 = x111 & n1646 ;
  assign n24561 = x112 & n1429 ;
  assign n24562 = ~n24560 & ~n24561 ;
  assign n24563 = ~n24559 & n24562 ;
  assign n24564 = n1437 & n16361 ;
  assign n24565 = n24563 & ~n24564 ;
  assign n24566 = x14 & ~n24565 ;
  assign n24567 = x14 & ~n24566 ;
  assign n24568 = ~n24565 & ~n24566 ;
  assign n24569 = ~n24567 & ~n24568 ;
  assign n24570 = ~n24123 & ~n24127 ;
  assign n24571 = ~n24118 & ~n24120 ;
  assign n24572 = ~n23864 & ~n24066 ;
  assign n24573 = ~n24063 & ~n24572 ;
  assign n24574 = ~n24047 & ~n24049 ;
  assign n24575 = ~n23983 & ~n23987 ;
  assign n24576 = ~n23972 & ~n23974 ;
  assign n24577 = ~n23096 & ~n23950 ;
  assign n24578 = ~n23947 & ~n24577 ;
  assign n24579 = x71 & n20143 ;
  assign n24580 = x69 & n20854 ;
  assign n24581 = x70 & n20138 ;
  assign n24582 = ~n24580 & ~n24581 ;
  assign n24583 = ~n24579 & n24582 ;
  assign n24584 = n558 & n20146 ;
  assign n24585 = n24583 & ~n24584 ;
  assign n24586 = x56 & ~n24585 ;
  assign n24587 = x56 & ~n24586 ;
  assign n24588 = ~n24585 & ~n24586 ;
  assign n24589 = ~n24587 & ~n24588 ;
  assign n24590 = n23078 & n23918 ;
  assign n24591 = ~n23933 & ~n24590 ;
  assign n24592 = x68 & n22325 ;
  assign n24593 = x66 & n23066 ;
  assign n24594 = x67 & n22320 ;
  assign n24595 = ~n24593 & ~n24594 ;
  assign n24596 = ~n24592 & n24595 ;
  assign n24597 = n317 & n22328 ;
  assign n24598 = n24596 & ~n24597 ;
  assign n24599 = x59 & ~n24598 ;
  assign n24600 = x59 & ~n24599 ;
  assign n24601 = ~n24598 & ~n24599 ;
  assign n24602 = ~n24600 & ~n24601 ;
  assign n24603 = x62 & ~n23918 ;
  assign n24604 = ~x60 & x61 ;
  assign n24605 = x60 & ~x61 ;
  assign n24606 = ~n24604 & ~n24605 ;
  assign n24607 = n23917 & ~n24606 ;
  assign n24608 = x64 & n24607 ;
  assign n24609 = ~x61 & x62 ;
  assign n24610 = x61 & ~x62 ;
  assign n24611 = ~n24609 & ~n24610 ;
  assign n24612 = ~n23917 & n24611 ;
  assign n24613 = x65 & n24612 ;
  assign n24614 = ~n24608 & ~n24613 ;
  assign n24615 = ~n23917 & ~n24611 ;
  assign n24616 = ~n152 & n24615 ;
  assign n24617 = n24614 & ~n24616 ;
  assign n24618 = x62 & ~n24617 ;
  assign n24619 = x62 & ~n24618 ;
  assign n24620 = ~n24617 & ~n24618 ;
  assign n24621 = ~n24619 & ~n24620 ;
  assign n24622 = n24603 & ~n24621 ;
  assign n24623 = ~n24603 & n24621 ;
  assign n24624 = ~n24622 & ~n24623 ;
  assign n24625 = n24602 & ~n24624 ;
  assign n24626 = ~n24602 & n24624 ;
  assign n24627 = ~n24625 & ~n24626 ;
  assign n24628 = ~n24591 & n24627 ;
  assign n24629 = n24591 & ~n24627 ;
  assign n24630 = ~n24628 & ~n24629 ;
  assign n24631 = n24589 & ~n24630 ;
  assign n24632 = ~n24589 & n24630 ;
  assign n24633 = ~n24631 & ~n24632 ;
  assign n24634 = ~n24578 & n24633 ;
  assign n24635 = n24578 & ~n24633 ;
  assign n24636 = ~n24634 & ~n24635 ;
  assign n24637 = x74 & n18025 ;
  assign n24638 = x72 & n18764 ;
  assign n24639 = x73 & n18020 ;
  assign n24640 = ~n24638 & ~n24639 ;
  assign n24641 = ~n24637 & n24640 ;
  assign n24642 = n994 & n18028 ;
  assign n24643 = n24641 & ~n24642 ;
  assign n24644 = x53 & ~n24643 ;
  assign n24645 = x53 & ~n24644 ;
  assign n24646 = ~n24643 & ~n24644 ;
  assign n24647 = ~n24645 & ~n24646 ;
  assign n24648 = n24636 & ~n24647 ;
  assign n24649 = n24636 & ~n24648 ;
  assign n24650 = ~n24647 & ~n24648 ;
  assign n24651 = ~n24649 & ~n24650 ;
  assign n24652 = ~n23965 & ~n23968 ;
  assign n24653 = n24651 & n24652 ;
  assign n24654 = ~n24651 & ~n24652 ;
  assign n24655 = ~n24653 & ~n24654 ;
  assign n24656 = x77 & n16076 ;
  assign n24657 = x75 & n16756 ;
  assign n24658 = x76 & n16071 ;
  assign n24659 = ~n24657 & ~n24658 ;
  assign n24660 = ~n24656 & n24659 ;
  assign n24661 = n1502 & n16079 ;
  assign n24662 = n24660 & ~n24661 ;
  assign n24663 = x50 & ~n24662 ;
  assign n24664 = x50 & ~n24663 ;
  assign n24665 = ~n24662 & ~n24663 ;
  assign n24666 = ~n24664 & ~n24665 ;
  assign n24667 = n24655 & ~n24666 ;
  assign n24668 = ~n24655 & n24666 ;
  assign n24669 = ~n24576 & ~n24668 ;
  assign n24670 = ~n24667 & n24669 ;
  assign n24671 = ~n24576 & ~n24670 ;
  assign n24672 = ~n24667 & ~n24670 ;
  assign n24673 = ~n24668 & n24672 ;
  assign n24674 = ~n24671 & ~n24673 ;
  assign n24675 = x80 & n14233 ;
  assign n24676 = x78 & n14876 ;
  assign n24677 = x79 & n14228 ;
  assign n24678 = ~n24676 & ~n24677 ;
  assign n24679 = ~n24675 & n24678 ;
  assign n24680 = n2028 & n14236 ;
  assign n24681 = n24679 & ~n24680 ;
  assign n24682 = x47 & ~n24681 ;
  assign n24683 = x47 & ~n24682 ;
  assign n24684 = ~n24681 & ~n24682 ;
  assign n24685 = ~n24683 & ~n24684 ;
  assign n24686 = ~n24674 & ~n24685 ;
  assign n24687 = ~n24674 & ~n24686 ;
  assign n24688 = ~n24685 & ~n24686 ;
  assign n24689 = ~n24687 & ~n24688 ;
  assign n24690 = ~n23977 & ~n23980 ;
  assign n24691 = n24689 & n24690 ;
  assign n24692 = ~n24689 & ~n24690 ;
  assign n24693 = ~n24691 & ~n24692 ;
  assign n24694 = x83 & n12506 ;
  assign n24695 = x81 & n13131 ;
  assign n24696 = x82 & n12501 ;
  assign n24697 = ~n24695 & ~n24696 ;
  assign n24698 = ~n24694 & n24697 ;
  assign n24699 = n2843 & n12509 ;
  assign n24700 = n24698 & ~n24699 ;
  assign n24701 = x44 & ~n24700 ;
  assign n24702 = x44 & ~n24701 ;
  assign n24703 = ~n24700 & ~n24701 ;
  assign n24704 = ~n24702 & ~n24703 ;
  assign n24705 = n24693 & ~n24704 ;
  assign n24706 = ~n24693 & n24704 ;
  assign n24707 = ~n24575 & ~n24706 ;
  assign n24708 = ~n24705 & n24707 ;
  assign n24709 = ~n24575 & ~n24708 ;
  assign n24710 = ~n24705 & ~n24708 ;
  assign n24711 = ~n24706 & n24710 ;
  assign n24712 = ~n24709 & ~n24711 ;
  assign n24713 = x86 & n10905 ;
  assign n24714 = x84 & n11466 ;
  assign n24715 = x85 & n10900 ;
  assign n24716 = ~n24714 & ~n24715 ;
  assign n24717 = ~n24713 & n24716 ;
  assign n24718 = n3686 & n10908 ;
  assign n24719 = n24717 & ~n24718 ;
  assign n24720 = x41 & ~n24719 ;
  assign n24721 = x41 & ~n24720 ;
  assign n24722 = ~n24719 & ~n24720 ;
  assign n24723 = ~n24721 & ~n24722 ;
  assign n24724 = ~n24712 & ~n24723 ;
  assign n24725 = ~n24712 & ~n24724 ;
  assign n24726 = ~n24723 & ~n24724 ;
  assign n24727 = ~n24725 & ~n24726 ;
  assign n24728 = ~n23991 & ~n23994 ;
  assign n24729 = n24727 & n24728 ;
  assign n24730 = ~n24727 & ~n24728 ;
  assign n24731 = ~n24729 & ~n24730 ;
  assign n24732 = x89 & n9433 ;
  assign n24733 = x87 & n9915 ;
  assign n24734 = x88 & n9428 ;
  assign n24735 = ~n24733 & ~n24734 ;
  assign n24736 = ~n24732 & n24735 ;
  assign n24737 = n4488 & n9436 ;
  assign n24738 = n24736 & ~n24737 ;
  assign n24739 = x38 & ~n24738 ;
  assign n24740 = x38 & ~n24739 ;
  assign n24741 = ~n24738 & ~n24739 ;
  assign n24742 = ~n24740 & ~n24741 ;
  assign n24743 = n24731 & ~n24742 ;
  assign n24744 = n24731 & ~n24743 ;
  assign n24745 = ~n24742 & ~n24743 ;
  assign n24746 = ~n24744 & ~n24745 ;
  assign n24747 = ~n24008 & ~n24014 ;
  assign n24748 = n24746 & n24747 ;
  assign n24749 = ~n24746 & ~n24747 ;
  assign n24750 = ~n24748 & ~n24749 ;
  assign n24751 = x92 & n8006 ;
  assign n24752 = x90 & n8474 ;
  assign n24753 = x91 & n8001 ;
  assign n24754 = ~n24752 & ~n24753 ;
  assign n24755 = ~n24751 & n24754 ;
  assign n24756 = n5710 & n8009 ;
  assign n24757 = n24755 & ~n24756 ;
  assign n24758 = x35 & ~n24757 ;
  assign n24759 = x35 & ~n24758 ;
  assign n24760 = ~n24757 & ~n24758 ;
  assign n24761 = ~n24759 & ~n24760 ;
  assign n24762 = n24750 & ~n24761 ;
  assign n24763 = n24750 & ~n24762 ;
  assign n24764 = ~n24761 & ~n24762 ;
  assign n24765 = ~n24763 & ~n24764 ;
  assign n24766 = ~n24027 & ~n24033 ;
  assign n24767 = n24765 & n24766 ;
  assign n24768 = ~n24765 & ~n24766 ;
  assign n24769 = ~n24767 & ~n24768 ;
  assign n24770 = x95 & n6725 ;
  assign n24771 = x93 & n7129 ;
  assign n24772 = x94 & n6720 ;
  assign n24773 = ~n24771 & ~n24772 ;
  assign n24774 = ~n24770 & n24773 ;
  assign n24775 = n6728 & n6894 ;
  assign n24776 = n24774 & ~n24775 ;
  assign n24777 = x32 & ~n24776 ;
  assign n24778 = x32 & ~n24777 ;
  assign n24779 = ~n24776 & ~n24777 ;
  assign n24780 = ~n24778 & ~n24779 ;
  assign n24781 = n24769 & ~n24780 ;
  assign n24782 = n24769 & ~n24781 ;
  assign n24783 = ~n24780 & ~n24781 ;
  assign n24784 = ~n24782 & ~n24783 ;
  assign n24785 = ~n24574 & n24784 ;
  assign n24786 = n24574 & ~n24784 ;
  assign n24787 = ~n24785 & ~n24786 ;
  assign n24788 = x98 & n5560 ;
  assign n24789 = x96 & n5943 ;
  assign n24790 = x97 & n5555 ;
  assign n24791 = ~n24789 & ~n24790 ;
  assign n24792 = ~n24788 & n24791 ;
  assign n24793 = n5563 & n8196 ;
  assign n24794 = n24792 & ~n24793 ;
  assign n24795 = x29 & ~n24794 ;
  assign n24796 = x29 & ~n24795 ;
  assign n24797 = ~n24794 & ~n24795 ;
  assign n24798 = ~n24796 & ~n24797 ;
  assign n24799 = ~n24787 & ~n24798 ;
  assign n24800 = n24787 & n24798 ;
  assign n24801 = ~n24799 & ~n24800 ;
  assign n24802 = n24573 & ~n24801 ;
  assign n24803 = ~n24573 & n24801 ;
  assign n24804 = ~n24802 & ~n24803 ;
  assign n24805 = x101 & n4531 ;
  assign n24806 = x99 & n4847 ;
  assign n24807 = x100 & n4526 ;
  assign n24808 = ~n24806 & ~n24807 ;
  assign n24809 = ~n24805 & n24808 ;
  assign n24810 = n4534 & n9601 ;
  assign n24811 = n24809 & ~n24810 ;
  assign n24812 = x26 & ~n24811 ;
  assign n24813 = x26 & ~n24812 ;
  assign n24814 = ~n24811 & ~n24812 ;
  assign n24815 = ~n24813 & ~n24814 ;
  assign n24816 = n24804 & ~n24815 ;
  assign n24817 = n24804 & ~n24816 ;
  assign n24818 = ~n24815 & ~n24816 ;
  assign n24819 = ~n24817 & ~n24818 ;
  assign n24820 = ~n24081 & ~n24085 ;
  assign n24821 = n24819 & n24820 ;
  assign n24822 = ~n24819 & ~n24820 ;
  assign n24823 = ~n24821 & ~n24822 ;
  assign n24824 = x104 & n3589 ;
  assign n24825 = x102 & n3878 ;
  assign n24826 = x103 & n3584 ;
  assign n24827 = ~n24825 & ~n24826 ;
  assign n24828 = ~n24824 & n24827 ;
  assign n24829 = n3592 & n11116 ;
  assign n24830 = n24828 & ~n24829 ;
  assign n24831 = x23 & ~n24830 ;
  assign n24832 = x23 & ~n24831 ;
  assign n24833 = ~n24830 & ~n24831 ;
  assign n24834 = ~n24832 & ~n24833 ;
  assign n24835 = n24823 & ~n24834 ;
  assign n24836 = n24823 & ~n24835 ;
  assign n24837 = ~n24834 & ~n24835 ;
  assign n24838 = ~n24836 & ~n24837 ;
  assign n24839 = ~n24098 & ~n24104 ;
  assign n24840 = n24838 & n24839 ;
  assign n24841 = ~n24838 & ~n24839 ;
  assign n24842 = ~n24840 & ~n24841 ;
  assign n24843 = x107 & n2751 ;
  assign n24844 = x105 & n3020 ;
  assign n24845 = x106 & n2746 ;
  assign n24846 = ~n24844 & ~n24845 ;
  assign n24847 = ~n24843 & n24846 ;
  assign n24848 = n2754 & n12749 ;
  assign n24849 = n24847 & ~n24848 ;
  assign n24850 = x20 & ~n24849 ;
  assign n24851 = x20 & ~n24850 ;
  assign n24852 = ~n24849 & ~n24850 ;
  assign n24853 = ~n24851 & ~n24852 ;
  assign n24854 = n24842 & ~n24853 ;
  assign n24855 = ~n24842 & n24853 ;
  assign n24856 = ~n24571 & ~n24855 ;
  assign n24857 = ~n24854 & n24856 ;
  assign n24858 = ~n24571 & ~n24857 ;
  assign n24859 = ~n24854 & ~n24857 ;
  assign n24860 = ~n24855 & n24859 ;
  assign n24861 = ~n24858 & ~n24860 ;
  assign n24862 = x110 & n2093 ;
  assign n24863 = x108 & n2275 ;
  assign n24864 = x109 & n2088 ;
  assign n24865 = ~n24863 & ~n24864 ;
  assign n24866 = ~n24862 & n24865 ;
  assign n24867 = n2096 & n14497 ;
  assign n24868 = n24866 & ~n24867 ;
  assign n24869 = x17 & ~n24868 ;
  assign n24870 = x17 & ~n24869 ;
  assign n24871 = ~n24868 & ~n24869 ;
  assign n24872 = ~n24870 & ~n24871 ;
  assign n24873 = n24861 & n24872 ;
  assign n24874 = ~n24861 & ~n24872 ;
  assign n24875 = ~n24873 & ~n24874 ;
  assign n24876 = ~n24570 & n24875 ;
  assign n24877 = n24570 & ~n24875 ;
  assign n24878 = ~n24876 & ~n24877 ;
  assign n24879 = n24569 & ~n24878 ;
  assign n24880 = ~n24569 & n24878 ;
  assign n24881 = ~n24879 & ~n24880 ;
  assign n24882 = ~n24558 & n24881 ;
  assign n24883 = n24558 & ~n24881 ;
  assign n24884 = ~n24882 & ~n24883 ;
  assign n24885 = n24557 & ~n24884 ;
  assign n24886 = ~n24557 & n24884 ;
  assign n24887 = ~n24885 & ~n24886 ;
  assign n24888 = ~n24546 & n24887 ;
  assign n24889 = n24546 & ~n24887 ;
  assign n24890 = ~n24888 & ~n24889 ;
  assign n24891 = x119 & n574 ;
  assign n24892 = x117 & n673 ;
  assign n24893 = x118 & n569 ;
  assign n24894 = ~n24892 & ~n24893 ;
  assign n24895 = ~n24891 & n24894 ;
  assign n24896 = n577 & n20423 ;
  assign n24897 = n24895 & ~n24896 ;
  assign n24898 = x8 & ~n24897 ;
  assign n24899 = x8 & ~n24898 ;
  assign n24900 = ~n24897 & ~n24898 ;
  assign n24901 = ~n24899 & ~n24900 ;
  assign n24902 = n24890 & ~n24901 ;
  assign n24903 = n24890 & ~n24902 ;
  assign n24904 = ~n24901 & ~n24902 ;
  assign n24905 = ~n24903 & ~n24904 ;
  assign n24906 = ~n24147 & ~n24150 ;
  assign n24907 = n24905 & n24906 ;
  assign n24908 = ~n24905 & ~n24906 ;
  assign n24909 = ~n24907 & ~n24908 ;
  assign n24910 = x122 & n293 ;
  assign n24911 = x120 & n373 ;
  assign n24912 = x121 & n288 ;
  assign n24913 = ~n24911 & ~n24912 ;
  assign n24914 = ~n24910 & n24913 ;
  assign n24915 = n296 & n22622 ;
  assign n24916 = n24914 & ~n24915 ;
  assign n24917 = x5 & ~n24916 ;
  assign n24918 = x5 & ~n24917 ;
  assign n24919 = ~n24916 & ~n24917 ;
  assign n24920 = ~n24918 & ~n24919 ;
  assign n24921 = ~n24909 & n24920 ;
  assign n24922 = n24909 & ~n24920 ;
  assign n24923 = ~n24921 & ~n24922 ;
  assign n24924 = x125 & n146 ;
  assign n24925 = x123 & n182 ;
  assign n24926 = x124 & n141 ;
  assign n24927 = ~n24925 & ~n24926 ;
  assign n24928 = ~n24924 & n24927 ;
  assign n24929 = ~n23792 & ~n23794 ;
  assign n24930 = ~x124 & ~x125 ;
  assign n24931 = x124 & x125 ;
  assign n24932 = ~n24930 & ~n24931 ;
  assign n24933 = ~n24929 & n24932 ;
  assign n24934 = n24929 & ~n24932 ;
  assign n24935 = ~n24933 & ~n24934 ;
  assign n24936 = n149 & n24935 ;
  assign n24937 = n24928 & ~n24936 ;
  assign n24938 = x2 & ~n24937 ;
  assign n24939 = x2 & ~n24938 ;
  assign n24940 = ~n24937 & ~n24938 ;
  assign n24941 = ~n24939 & ~n24940 ;
  assign n24942 = n24923 & ~n24941 ;
  assign n24943 = n24923 & ~n24942 ;
  assign n24944 = ~n24941 & ~n24942 ;
  assign n24945 = ~n24943 & ~n24944 ;
  assign n24946 = ~n24153 & ~n24156 ;
  assign n24947 = n24945 & n24946 ;
  assign n24948 = ~n24945 & ~n24946 ;
  assign n24949 = ~n24947 & ~n24948 ;
  assign n24950 = ~n24159 & ~n24162 ;
  assign n24951 = n24949 & ~n24950 ;
  assign n24952 = ~n24949 & n24950 ;
  assign n24953 = ~n24951 & ~n24952 ;
  assign n25350 = n24953 & x189 ;
  assign n24954 = ~n24516 & ~n24520 ;
  assign n24955 = ~x116 & n945 ;
  assign n24956 = ~x114 & n1099 ;
  assign n24957 = ~x115 & n940 ;
  assign n24958 = ~n24956 & ~n24957 ;
  assign n24959 = ~n24955 & n24958 ;
  assign n24960 = n948 & n18678 ;
  assign n24961 = n24959 & ~n24960 ;
  assign n24962 = ~x11 & ~n24961 ;
  assign n24963 = ~x11 & ~n24962 ;
  assign n24964 = ~n24961 & ~n24962 ;
  assign n24965 = ~n24963 & ~n24964 ;
  assign n24966 = ~n24508 & ~n24512 ;
  assign n24967 = ~x113 & n1434 ;
  assign n24968 = ~x111 & n1646 ;
  assign n24969 = ~x112 & n1429 ;
  assign n24970 = ~n24968 & ~n24969 ;
  assign n24971 = ~n24967 & n24970 ;
  assign n24972 = n1437 & n16684 ;
  assign n24973 = n24971 & ~n24972 ;
  assign n24974 = ~x14 & ~n24973 ;
  assign n24975 = ~x14 & ~n24974 ;
  assign n24976 = ~n24973 & ~n24974 ;
  assign n24977 = ~n24975 & ~n24976 ;
  assign n24978 = ~n24500 & ~n24504 ;
  assign n24979 = ~n24495 & ~n24497 ;
  assign n24980 = ~n24244 & ~n24443 ;
  assign n24981 = ~n24440 & ~n24980 ;
  assign n24982 = ~n24424 & ~n24426 ;
  assign n24983 = ~n24360 & ~n24364 ;
  assign n24984 = ~n24349 & ~n24351 ;
  assign n24985 = ~n23477 & ~n24327 ;
  assign n24986 = ~n24324 & ~n24985 ;
  assign n24987 = ~x71 & n20143 ;
  assign n24988 = ~x69 & n20854 ;
  assign n24989 = ~x70 & n20138 ;
  assign n24990 = ~n24988 & ~n24989 ;
  assign n24991 = ~n24987 & n24990 ;
  assign n24992 = n622 & n20146 ;
  assign n24993 = n24991 & ~n24992 ;
  assign n24994 = ~x56 & ~n24993 ;
  assign n24995 = ~x56 & ~n24994 ;
  assign n24996 = ~n24993 & ~n24994 ;
  assign n24997 = ~n24995 & ~n24996 ;
  assign n24998 = n23459 & n24295 ;
  assign n24999 = ~n24310 & ~n24998 ;
  assign n25000 = ~x68 & n22325 ;
  assign n25001 = ~x66 & n23066 ;
  assign n25002 = ~x67 & n22320 ;
  assign n25003 = ~n25001 & ~n25002 ;
  assign n25004 = ~n25000 & n25003 ;
  assign n25005 = n352 & n22328 ;
  assign n25006 = n25004 & ~n25005 ;
  assign n25007 = ~x59 & ~n25006 ;
  assign n25008 = ~x59 & ~n25007 ;
  assign n25009 = ~n25006 & ~n25007 ;
  assign n25010 = ~n25008 & ~n25009 ;
  assign n25011 = ~x62 & ~n24295 ;
  assign n25012 = ~x64 & n24607 ;
  assign n25013 = ~x65 & n24612 ;
  assign n25014 = ~n25012 & ~n25013 ;
  assign n25015 = ~n24616 & n25014 ;
  assign n25016 = ~x62 & ~n25015 ;
  assign n25017 = ~x62 & ~n25016 ;
  assign n25018 = ~n25015 & ~n25016 ;
  assign n25019 = ~n25017 & ~n25018 ;
  assign n25020 = n25011 & ~n25019 ;
  assign n25021 = ~n25011 & n25019 ;
  assign n25022 = ~n25020 & ~n25021 ;
  assign n25023 = n25010 & ~n25022 ;
  assign n25024 = ~n25010 & n25022 ;
  assign n25025 = ~n25023 & ~n25024 ;
  assign n25026 = ~n24999 & n25025 ;
  assign n25027 = n24999 & ~n25025 ;
  assign n25028 = ~n25026 & ~n25027 ;
  assign n25029 = n24997 & ~n25028 ;
  assign n25030 = ~n24997 & n25028 ;
  assign n25031 = ~n25029 & ~n25030 ;
  assign n25032 = ~n24986 & n25031 ;
  assign n25033 = n24986 & ~n25031 ;
  assign n25034 = ~n25032 & ~n25033 ;
  assign n25035 = ~x74 & n18025 ;
  assign n25036 = ~x72 & n18764 ;
  assign n25037 = ~x73 & n18020 ;
  assign n25038 = ~n25036 & ~n25037 ;
  assign n25039 = ~n25035 & n25038 ;
  assign n25040 = n1066 & n18028 ;
  assign n25041 = n25039 & ~n25040 ;
  assign n25042 = ~x53 & ~n25041 ;
  assign n25043 = ~x53 & ~n25042 ;
  assign n25044 = ~n25041 & ~n25042 ;
  assign n25045 = ~n25043 & ~n25044 ;
  assign n25046 = n25034 & ~n25045 ;
  assign n25047 = n25034 & ~n25046 ;
  assign n25048 = ~n25045 & ~n25046 ;
  assign n25049 = ~n25047 & ~n25048 ;
  assign n25050 = ~n24342 & ~n24345 ;
  assign n25051 = n25049 & n25050 ;
  assign n25052 = ~n25049 & ~n25050 ;
  assign n25053 = ~n25051 & ~n25052 ;
  assign n25054 = ~x77 & n16076 ;
  assign n25055 = ~x75 & n16756 ;
  assign n25056 = ~x76 & n16071 ;
  assign n25057 = ~n25055 & ~n25056 ;
  assign n25058 = ~n25054 & n25057 ;
  assign n25059 = n1594 & n16079 ;
  assign n25060 = n25058 & ~n25059 ;
  assign n25061 = ~x50 & ~n25060 ;
  assign n25062 = ~x50 & ~n25061 ;
  assign n25063 = ~n25060 & ~n25061 ;
  assign n25064 = ~n25062 & ~n25063 ;
  assign n25065 = n25053 & ~n25064 ;
  assign n25066 = ~n25053 & n25064 ;
  assign n25067 = ~n24984 & ~n25066 ;
  assign n25068 = ~n25065 & n25067 ;
  assign n25069 = ~n24984 & ~n25068 ;
  assign n25070 = ~n25065 & ~n25068 ;
  assign n25071 = ~n25066 & n25070 ;
  assign n25072 = ~n25069 & ~n25071 ;
  assign n25073 = ~x80 & n14233 ;
  assign n25074 = ~x78 & n14876 ;
  assign n25075 = ~x79 & n14228 ;
  assign n25076 = ~n25074 & ~n25075 ;
  assign n25077 = ~n25073 & n25076 ;
  assign n25078 = n2145 & n14236 ;
  assign n25079 = n25077 & ~n25078 ;
  assign n25080 = ~x47 & ~n25079 ;
  assign n25081 = ~x47 & ~n25080 ;
  assign n25082 = ~n25079 & ~n25080 ;
  assign n25083 = ~n25081 & ~n25082 ;
  assign n25084 = ~n25072 & ~n25083 ;
  assign n25085 = ~n25072 & ~n25084 ;
  assign n25086 = ~n25083 & ~n25084 ;
  assign n25087 = ~n25085 & ~n25086 ;
  assign n25088 = ~n24354 & ~n24357 ;
  assign n25089 = n25087 & n25088 ;
  assign n25090 = ~n25087 & ~n25088 ;
  assign n25091 = ~n25089 & ~n25090 ;
  assign n25092 = ~x83 & n12506 ;
  assign n25093 = ~x81 & n13131 ;
  assign n25094 = ~x82 & n12501 ;
  assign n25095 = ~n25093 & ~n25094 ;
  assign n25096 = ~n25092 & n25095 ;
  assign n25097 = n2972 & n12509 ;
  assign n25098 = n25096 & ~n25097 ;
  assign n25099 = ~x44 & ~n25098 ;
  assign n25100 = ~x44 & ~n25099 ;
  assign n25101 = ~n25098 & ~n25099 ;
  assign n25102 = ~n25100 & ~n25101 ;
  assign n25103 = n25091 & ~n25102 ;
  assign n25104 = ~n25091 & n25102 ;
  assign n25105 = ~n24983 & ~n25104 ;
  assign n25106 = ~n25103 & n25105 ;
  assign n25107 = ~n24983 & ~n25106 ;
  assign n25108 = ~n25103 & ~n25106 ;
  assign n25109 = ~n25104 & n25108 ;
  assign n25110 = ~n25107 & ~n25109 ;
  assign n25111 = ~x86 & n10905 ;
  assign n25112 = ~x84 & n11466 ;
  assign n25113 = ~x85 & n10900 ;
  assign n25114 = ~n25112 & ~n25113 ;
  assign n25115 = ~n25111 & n25114 ;
  assign n25116 = n3832 & n10908 ;
  assign n25117 = n25115 & ~n25116 ;
  assign n25118 = ~x41 & ~n25117 ;
  assign n25119 = ~x41 & ~n25118 ;
  assign n25120 = ~n25117 & ~n25118 ;
  assign n25121 = ~n25119 & ~n25120 ;
  assign n25122 = ~n25110 & ~n25121 ;
  assign n25123 = ~n25110 & ~n25122 ;
  assign n25124 = ~n25121 & ~n25122 ;
  assign n25125 = ~n25123 & ~n25124 ;
  assign n25126 = ~n24368 & ~n24371 ;
  assign n25127 = n25125 & n25126 ;
  assign n25128 = ~n25125 & ~n25126 ;
  assign n25129 = ~n25127 & ~n25128 ;
  assign n25130 = ~x89 & n9433 ;
  assign n25131 = ~x87 & n9915 ;
  assign n25132 = ~x88 & n9428 ;
  assign n25133 = ~n25131 & ~n25132 ;
  assign n25134 = ~n25130 & n25133 ;
  assign n25135 = n4664 & n9436 ;
  assign n25136 = n25134 & ~n25135 ;
  assign n25137 = ~x38 & ~n25136 ;
  assign n25138 = ~x38 & ~n25137 ;
  assign n25139 = ~n25136 & ~n25137 ;
  assign n25140 = ~n25138 & ~n25139 ;
  assign n25141 = n25129 & ~n25140 ;
  assign n25142 = n25129 & ~n25141 ;
  assign n25143 = ~n25140 & ~n25141 ;
  assign n25144 = ~n25142 & ~n25143 ;
  assign n25145 = ~n24385 & ~n24391 ;
  assign n25146 = n25144 & n25145 ;
  assign n25147 = ~n25144 & ~n25145 ;
  assign n25148 = ~n25146 & ~n25147 ;
  assign n25149 = ~x92 & n8006 ;
  assign n25150 = ~x90 & n8474 ;
  assign n25151 = ~x91 & n8001 ;
  assign n25152 = ~n25150 & ~n25151 ;
  assign n25153 = ~n25149 & n25152 ;
  assign n25154 = n5896 & n8009 ;
  assign n25155 = n25153 & ~n25154 ;
  assign n25156 = ~x35 & ~n25155 ;
  assign n25157 = ~x35 & ~n25156 ;
  assign n25158 = ~n25155 & ~n25156 ;
  assign n25159 = ~n25157 & ~n25158 ;
  assign n25160 = n25148 & ~n25159 ;
  assign n25161 = n25148 & ~n25160 ;
  assign n25162 = ~n25159 & ~n25160 ;
  assign n25163 = ~n25161 & ~n25162 ;
  assign n25164 = ~n24404 & ~n24410 ;
  assign n25165 = n25163 & n25164 ;
  assign n25166 = ~n25163 & ~n25164 ;
  assign n25167 = ~n25165 & ~n25166 ;
  assign n25168 = ~x95 & n6725 ;
  assign n25169 = ~x93 & n7129 ;
  assign n25170 = ~x94 & n6720 ;
  assign n25171 = ~n25169 & ~n25170 ;
  assign n25172 = ~n25168 & n25171 ;
  assign n25173 = n6728 & n7100 ;
  assign n25174 = n25172 & ~n25173 ;
  assign n25175 = ~x32 & ~n25174 ;
  assign n25176 = ~x32 & ~n25175 ;
  assign n25177 = ~n25174 & ~n25175 ;
  assign n25178 = ~n25176 & ~n25177 ;
  assign n25179 = n25167 & ~n25178 ;
  assign n25180 = n25167 & ~n25179 ;
  assign n25181 = ~n25178 & ~n25179 ;
  assign n25182 = ~n25180 & ~n25181 ;
  assign n25183 = ~n24982 & n25182 ;
  assign n25184 = n24982 & ~n25182 ;
  assign n25185 = ~n25183 & ~n25184 ;
  assign n25186 = ~x98 & n5560 ;
  assign n25187 = ~x96 & n5943 ;
  assign n25188 = ~x97 & n5555 ;
  assign n25189 = ~n25187 & ~n25188 ;
  assign n25190 = ~n25186 & n25189 ;
  assign n25191 = n5563 & n8426 ;
  assign n25192 = n25190 & ~n25191 ;
  assign n25193 = ~x29 & ~n25192 ;
  assign n25194 = ~x29 & ~n25193 ;
  assign n25195 = ~n25192 & ~n25193 ;
  assign n25196 = ~n25194 & ~n25195 ;
  assign n25197 = ~n25185 & ~n25196 ;
  assign n25198 = n25185 & n25196 ;
  assign n25199 = ~n25197 & ~n25198 ;
  assign n25200 = n24981 & ~n25199 ;
  assign n25201 = ~n24981 & n25199 ;
  assign n25202 = ~n25200 & ~n25201 ;
  assign n25203 = ~x101 & n4531 ;
  assign n25204 = ~x99 & n4847 ;
  assign n25205 = ~x100 & n4526 ;
  assign n25206 = ~n25204 & ~n25205 ;
  assign n25207 = ~n25203 & n25206 ;
  assign n25208 = n4534 & n9844 ;
  assign n25209 = n25207 & ~n25208 ;
  assign n25210 = ~x26 & ~n25209 ;
  assign n25211 = ~x26 & ~n25210 ;
  assign n25212 = ~n25209 & ~n25210 ;
  assign n25213 = ~n25211 & ~n25212 ;
  assign n25214 = n25202 & ~n25213 ;
  assign n25215 = n25202 & ~n25214 ;
  assign n25216 = ~n25213 & ~n25214 ;
  assign n25217 = ~n25215 & ~n25216 ;
  assign n25218 = ~n24458 & ~n24462 ;
  assign n25219 = n25217 & n25218 ;
  assign n25220 = ~n25217 & ~n25218 ;
  assign n25221 = ~n25219 & ~n25220 ;
  assign n25222 = ~x104 & n3589 ;
  assign n25223 = ~x102 & n3878 ;
  assign n25224 = ~x103 & n3584 ;
  assign n25225 = ~n25223 & ~n25224 ;
  assign n25226 = ~n25222 & n25225 ;
  assign n25227 = n3592 & n11380 ;
  assign n25228 = n25226 & ~n25227 ;
  assign n25229 = ~x23 & ~n25228 ;
  assign n25230 = ~x23 & ~n25229 ;
  assign n25231 = ~n25228 & ~n25229 ;
  assign n25232 = ~n25230 & ~n25231 ;
  assign n25233 = n25221 & ~n25232 ;
  assign n25234 = n25221 & ~n25233 ;
  assign n25235 = ~n25232 & ~n25233 ;
  assign n25236 = ~n25234 & ~n25235 ;
  assign n25237 = ~n24475 & ~n24481 ;
  assign n25238 = n25236 & n25237 ;
  assign n25239 = ~n25236 & ~n25237 ;
  assign n25240 = ~n25238 & ~n25239 ;
  assign n25241 = ~x107 & n2751 ;
  assign n25242 = ~x105 & n3020 ;
  assign n25243 = ~x106 & n2746 ;
  assign n25244 = ~n25242 & ~n25243 ;
  assign n25245 = ~n25241 & n25244 ;
  assign n25246 = n2754 & n13034 ;
  assign n25247 = n25245 & ~n25246 ;
  assign n25248 = ~x20 & ~n25247 ;
  assign n25249 = ~x20 & ~n25248 ;
  assign n25250 = ~n25247 & ~n25248 ;
  assign n25251 = ~n25249 & ~n25250 ;
  assign n25252 = n25240 & ~n25251 ;
  assign n25253 = ~n25240 & n25251 ;
  assign n25254 = ~n24979 & ~n25253 ;
  assign n25255 = ~n25252 & n25254 ;
  assign n25256 = ~n24979 & ~n25255 ;
  assign n25257 = ~n25252 & ~n25255 ;
  assign n25258 = ~n25253 & n25257 ;
  assign n25259 = ~n25256 & ~n25258 ;
  assign n25260 = ~x110 & n2093 ;
  assign n25261 = ~x108 & n2275 ;
  assign n25262 = ~x109 & n2088 ;
  assign n25263 = ~n25261 & ~n25262 ;
  assign n25264 = ~n25260 & n25263 ;
  assign n25265 = n2096 & n14802 ;
  assign n25266 = n25264 & ~n25265 ;
  assign n25267 = ~x17 & ~n25266 ;
  assign n25268 = ~x17 & ~n25267 ;
  assign n25269 = ~n25266 & ~n25267 ;
  assign n25270 = ~n25268 & ~n25269 ;
  assign n25271 = n25259 & n25270 ;
  assign n25272 = ~n25259 & ~n25270 ;
  assign n25273 = ~n25271 & ~n25272 ;
  assign n25274 = ~n24978 & n25273 ;
  assign n25275 = n24978 & ~n25273 ;
  assign n25276 = ~n25274 & ~n25275 ;
  assign n25277 = n24977 & ~n25276 ;
  assign n25278 = ~n24977 & n25276 ;
  assign n25279 = ~n25277 & ~n25278 ;
  assign n25280 = ~n24966 & n25279 ;
  assign n25281 = n24966 & ~n25279 ;
  assign n25282 = ~n25280 & ~n25281 ;
  assign n25283 = n24965 & ~n25282 ;
  assign n25284 = ~n24965 & n25282 ;
  assign n25285 = ~n25283 & ~n25284 ;
  assign n25286 = ~n24954 & n25285 ;
  assign n25287 = n24954 & ~n25285 ;
  assign n25288 = ~n25286 & ~n25287 ;
  assign n25289 = ~x119 & n574 ;
  assign n25290 = ~x117 & n673 ;
  assign n25291 = ~x118 & n569 ;
  assign n25292 = ~n25290 & ~n25291 ;
  assign n25293 = ~n25289 & n25292 ;
  assign n25294 = n577 & n20778 ;
  assign n25295 = n25293 & ~n25294 ;
  assign n25296 = ~x8 & ~n25295 ;
  assign n25297 = ~x8 & ~n25296 ;
  assign n25298 = ~n25295 & ~n25296 ;
  assign n25299 = ~n25297 & ~n25298 ;
  assign n25300 = n25288 & ~n25299 ;
  assign n25301 = n25288 & ~n25300 ;
  assign n25302 = ~n25299 & ~n25300 ;
  assign n25303 = ~n25301 & ~n25302 ;
  assign n25304 = ~n24524 & ~n24527 ;
  assign n25305 = n25303 & n25304 ;
  assign n25306 = ~n25303 & ~n25304 ;
  assign n25307 = ~n25305 & ~n25306 ;
  assign n25308 = ~x122 & n293 ;
  assign n25309 = ~x120 & n373 ;
  assign n25310 = ~x121 & n288 ;
  assign n25311 = ~n25309 & ~n25310 ;
  assign n25312 = ~n25308 & n25311 ;
  assign n25313 = n296 & n22998 ;
  assign n25314 = n25312 & ~n25313 ;
  assign n25315 = ~x5 & ~n25314 ;
  assign n25316 = ~x5 & ~n25315 ;
  assign n25317 = ~n25314 & ~n25315 ;
  assign n25318 = ~n25316 & ~n25317 ;
  assign n25319 = ~n25307 & n25318 ;
  assign n25320 = n25307 & ~n25318 ;
  assign n25321 = ~n25319 & ~n25320 ;
  assign n25322 = ~x125 & n164 ;
  assign n25323 = ~x123 & n205 ;
  assign n25324 = ~x124 & n162 ;
  assign n25325 = ~n25323 & ~n25324 ;
  assign n25326 = ~n25322 & n25325 ;
  assign n25327 = ~n23791 & ~n24174 ;
  assign n25328 = n24932 & ~n25327 ;
  assign n25329 = ~n24932 & n25327 ;
  assign n25330 = ~n25328 & ~n25329 ;
  assign n25331 = n167 & n25330 ;
  assign n25332 = n25326 & ~n25331 ;
  assign n25333 = ~x2 & ~n25332 ;
  assign n25334 = ~x2 & ~n25333 ;
  assign n25335 = ~n25332 & ~n25333 ;
  assign n25336 = ~n25334 & ~n25335 ;
  assign n25337 = n25321 & ~n25336 ;
  assign n25338 = n25321 & ~n25337 ;
  assign n25339 = ~n25336 & ~n25337 ;
  assign n25340 = ~n25338 & ~n25339 ;
  assign n25341 = ~n24530 & ~n24533 ;
  assign n25342 = n25340 & n25341 ;
  assign n25343 = ~n25340 & ~n25341 ;
  assign n25344 = ~n25342 & ~n25343 ;
  assign n25345 = ~n24536 & ~n24539 ;
  assign n25346 = n25344 & ~n25345 ;
  assign n25347 = ~n25344 & n25345 ;
  assign n25348 = ~n25346 & ~n25347 ;
  assign n25351 = ~n25348 & ~x189 ;
  assign n25352 = ~n25350 & ~n25351 ;
  assign n25353 = ~n24948 & ~n24951 ;
  assign n25354 = ~n24922 & ~n24942 ;
  assign n25355 = ~n24886 & ~n24888 ;
  assign n25356 = ~n24880 & ~n24882 ;
  assign n25357 = ~n24874 & ~n24876 ;
  assign n25358 = ~n24835 & ~n24841 ;
  assign n25359 = ~n24574 & ~n24784 ;
  assign n25360 = ~n24781 & ~n25359 ;
  assign n25361 = ~n24724 & ~n24730 ;
  assign n25362 = ~n24686 & ~n24692 ;
  assign n25363 = x81 & n14233 ;
  assign n25364 = x79 & n14876 ;
  assign n25365 = x80 & n14228 ;
  assign n25366 = ~n25364 & ~n25365 ;
  assign n25367 = ~n25363 & n25366 ;
  assign n25368 = n2348 & n14236 ;
  assign n25369 = n25367 & ~n25368 ;
  assign n25370 = x47 & ~n25369 ;
  assign n25371 = x47 & ~n25370 ;
  assign n25372 = ~n25369 & ~n25370 ;
  assign n25373 = ~n25371 & ~n25372 ;
  assign n25374 = ~n24648 & ~n24654 ;
  assign n25375 = x75 & n18025 ;
  assign n25376 = x73 & n18764 ;
  assign n25377 = x74 & n18020 ;
  assign n25378 = ~n25376 & ~n25377 ;
  assign n25379 = ~n25375 & n25378 ;
  assign n25380 = n1150 & n18028 ;
  assign n25381 = n25379 & ~n25380 ;
  assign n25382 = x53 & ~n25381 ;
  assign n25383 = x53 & ~n25382 ;
  assign n25384 = ~n25381 & ~n25382 ;
  assign n25385 = ~n25383 & ~n25384 ;
  assign n25386 = ~n24632 & ~n24634 ;
  assign n25387 = ~n24626 & ~n24628 ;
  assign n25388 = x66 & n24612 ;
  assign n25389 = n23917 & ~n24611 ;
  assign n25390 = n24606 & n25389 ;
  assign n25391 = x64 & n25390 ;
  assign n25392 = x65 & n24607 ;
  assign n25393 = ~n25391 & ~n25392 ;
  assign n25394 = ~n25388 & n25393 ;
  assign n25395 = n194 & n24615 ;
  assign n25396 = n25394 & ~n25395 ;
  assign n25397 = x62 & ~n25396 ;
  assign n25398 = x62 & ~n25397 ;
  assign n25399 = ~n25396 & ~n25397 ;
  assign n25400 = ~n25398 & ~n25399 ;
  assign n25401 = ~n24622 & n25400 ;
  assign n25402 = n24622 & ~n25400 ;
  assign n25403 = ~n25401 & ~n25402 ;
  assign n25404 = x69 & n22325 ;
  assign n25405 = x67 & n23066 ;
  assign n25406 = x68 & n22320 ;
  assign n25407 = ~n25405 & ~n25406 ;
  assign n25408 = ~n25404 & n25407 ;
  assign n25409 = n398 & n22328 ;
  assign n25410 = n25408 & ~n25409 ;
  assign n25411 = x59 & ~n25410 ;
  assign n25412 = x59 & ~n25411 ;
  assign n25413 = ~n25410 & ~n25411 ;
  assign n25414 = ~n25412 & ~n25413 ;
  assign n25415 = n25403 & ~n25414 ;
  assign n25416 = ~n25403 & n25414 ;
  assign n25417 = ~n25387 & ~n25416 ;
  assign n25418 = ~n25415 & n25417 ;
  assign n25419 = ~n25387 & ~n25418 ;
  assign n25420 = ~n25415 & ~n25418 ;
  assign n25421 = ~n25416 & n25420 ;
  assign n25422 = ~n25419 & ~n25421 ;
  assign n25423 = x72 & n20143 ;
  assign n25424 = x70 & n20854 ;
  assign n25425 = x71 & n20138 ;
  assign n25426 = ~n25424 & ~n25425 ;
  assign n25427 = ~n25423 & n25426 ;
  assign n25428 = n717 & n20146 ;
  assign n25429 = n25427 & ~n25428 ;
  assign n25430 = x56 & ~n25429 ;
  assign n25431 = x56 & ~n25430 ;
  assign n25432 = ~n25429 & ~n25430 ;
  assign n25433 = ~n25431 & ~n25432 ;
  assign n25434 = n25422 & n25433 ;
  assign n25435 = ~n25422 & ~n25433 ;
  assign n25436 = ~n25434 & ~n25435 ;
  assign n25437 = ~n25386 & n25436 ;
  assign n25438 = n25386 & ~n25436 ;
  assign n25439 = ~n25437 & ~n25438 ;
  assign n25440 = n25385 & ~n25439 ;
  assign n25441 = ~n25385 & n25439 ;
  assign n25442 = ~n25440 & ~n25441 ;
  assign n25443 = ~n25374 & n25442 ;
  assign n25444 = n25374 & ~n25442 ;
  assign n25445 = ~n25443 & ~n25444 ;
  assign n25446 = x78 & n16076 ;
  assign n25447 = x76 & n16756 ;
  assign n25448 = x77 & n16071 ;
  assign n25449 = ~n25447 & ~n25448 ;
  assign n25450 = ~n25446 & n25449 ;
  assign n25451 = n1624 & n16079 ;
  assign n25452 = n25450 & ~n25451 ;
  assign n25453 = x50 & ~n25452 ;
  assign n25454 = x50 & ~n25453 ;
  assign n25455 = ~n25452 & ~n25453 ;
  assign n25456 = ~n25454 & ~n25455 ;
  assign n25457 = n25445 & ~n25456 ;
  assign n25458 = n25445 & ~n25457 ;
  assign n25459 = ~n25456 & ~n25457 ;
  assign n25460 = ~n25458 & ~n25459 ;
  assign n25461 = ~n24672 & ~n25460 ;
  assign n25462 = n24672 & n25460 ;
  assign n25463 = ~n25461 & ~n25462 ;
  assign n25464 = ~n25373 & n25463 ;
  assign n25465 = ~n25373 & ~n25464 ;
  assign n25466 = n25463 & ~n25464 ;
  assign n25467 = ~n25465 & ~n25466 ;
  assign n25468 = ~n25362 & ~n25467 ;
  assign n25469 = ~n25362 & ~n25468 ;
  assign n25470 = ~n25467 & ~n25468 ;
  assign n25471 = ~n25469 & ~n25470 ;
  assign n25472 = x84 & n12506 ;
  assign n25473 = x82 & n13131 ;
  assign n25474 = x83 & n12501 ;
  assign n25475 = ~n25473 & ~n25474 ;
  assign n25476 = ~n25472 & n25475 ;
  assign n25477 = n3114 & n12509 ;
  assign n25478 = n25476 & ~n25477 ;
  assign n25479 = x44 & ~n25478 ;
  assign n25480 = x44 & ~n25479 ;
  assign n25481 = ~n25478 & ~n25479 ;
  assign n25482 = ~n25480 & ~n25481 ;
  assign n25483 = ~n25471 & ~n25482 ;
  assign n25484 = ~n25471 & ~n25483 ;
  assign n25485 = ~n25482 & ~n25483 ;
  assign n25486 = ~n25484 & ~n25485 ;
  assign n25487 = ~n24710 & n25486 ;
  assign n25488 = n24710 & ~n25486 ;
  assign n25489 = ~n25487 & ~n25488 ;
  assign n25490 = x87 & n10905 ;
  assign n25491 = x85 & n11466 ;
  assign n25492 = x86 & n10900 ;
  assign n25493 = ~n25491 & ~n25492 ;
  assign n25494 = ~n25490 & n25493 ;
  assign n25495 = n3991 & n10908 ;
  assign n25496 = n25494 & ~n25495 ;
  assign n25497 = x41 & ~n25496 ;
  assign n25498 = x41 & ~n25497 ;
  assign n25499 = ~n25496 & ~n25497 ;
  assign n25500 = ~n25498 & ~n25499 ;
  assign n25501 = ~n25489 & ~n25500 ;
  assign n25502 = n25489 & n25500 ;
  assign n25503 = ~n25501 & ~n25502 ;
  assign n25504 = n25361 & ~n25503 ;
  assign n25505 = ~n25361 & n25503 ;
  assign n25506 = ~n25504 & ~n25505 ;
  assign n25507 = x90 & n9433 ;
  assign n25508 = x88 & n9915 ;
  assign n25509 = x89 & n9428 ;
  assign n25510 = ~n25508 & ~n25509 ;
  assign n25511 = ~n25507 & n25510 ;
  assign n25512 = n4986 & n9436 ;
  assign n25513 = n25511 & ~n25512 ;
  assign n25514 = x38 & ~n25513 ;
  assign n25515 = x38 & ~n25514 ;
  assign n25516 = ~n25513 & ~n25514 ;
  assign n25517 = ~n25515 & ~n25516 ;
  assign n25518 = n25506 & ~n25517 ;
  assign n25519 = n25506 & ~n25518 ;
  assign n25520 = ~n25517 & ~n25518 ;
  assign n25521 = ~n25519 & ~n25520 ;
  assign n25522 = ~n24743 & ~n24749 ;
  assign n25523 = n25521 & n25522 ;
  assign n25524 = ~n25521 & ~n25522 ;
  assign n25525 = ~n25523 & ~n25524 ;
  assign n25526 = x93 & n8006 ;
  assign n25527 = x91 & n8474 ;
  assign n25528 = x92 & n8001 ;
  assign n25529 = ~n25527 & ~n25528 ;
  assign n25530 = ~n25526 & n25529 ;
  assign n25531 = n6094 & n8009 ;
  assign n25532 = n25530 & ~n25531 ;
  assign n25533 = x35 & ~n25532 ;
  assign n25534 = x35 & ~n25533 ;
  assign n25535 = ~n25532 & ~n25533 ;
  assign n25536 = ~n25534 & ~n25535 ;
  assign n25537 = n25525 & ~n25536 ;
  assign n25538 = n25525 & ~n25537 ;
  assign n25539 = ~n25536 & ~n25537 ;
  assign n25540 = ~n25538 & ~n25539 ;
  assign n25541 = ~n24762 & ~n24768 ;
  assign n25542 = n25540 & n25541 ;
  assign n25543 = ~n25540 & ~n25541 ;
  assign n25544 = ~n25542 & ~n25543 ;
  assign n25545 = x96 & n6725 ;
  assign n25546 = x94 & n7129 ;
  assign n25547 = x95 & n6720 ;
  assign n25548 = ~n25546 & ~n25547 ;
  assign n25549 = ~n25545 & n25548 ;
  assign n25550 = n6728 & n7321 ;
  assign n25551 = n25549 & ~n25550 ;
  assign n25552 = x32 & ~n25551 ;
  assign n25553 = x32 & ~n25552 ;
  assign n25554 = ~n25551 & ~n25552 ;
  assign n25555 = ~n25553 & ~n25554 ;
  assign n25556 = n25544 & ~n25555 ;
  assign n25557 = ~n25544 & n25555 ;
  assign n25558 = ~n25360 & ~n25557 ;
  assign n25559 = ~n25556 & n25558 ;
  assign n25560 = ~n25360 & ~n25559 ;
  assign n25561 = ~n25556 & ~n25559 ;
  assign n25562 = ~n25557 & n25561 ;
  assign n25563 = ~n25560 & ~n25562 ;
  assign n25564 = x99 & n5560 ;
  assign n25565 = x97 & n5943 ;
  assign n25566 = x98 & n5555 ;
  assign n25567 = ~n25565 & ~n25566 ;
  assign n25568 = ~n25564 & n25567 ;
  assign n25569 = n5563 & n8660 ;
  assign n25570 = n25568 & ~n25569 ;
  assign n25571 = x29 & ~n25570 ;
  assign n25572 = x29 & ~n25571 ;
  assign n25573 = ~n25570 & ~n25571 ;
  assign n25574 = ~n25572 & ~n25573 ;
  assign n25575 = ~n25563 & ~n25574 ;
  assign n25576 = ~n25563 & ~n25575 ;
  assign n25577 = ~n25574 & ~n25575 ;
  assign n25578 = ~n25576 & ~n25577 ;
  assign n25579 = ~n24799 & ~n24803 ;
  assign n25580 = n25578 & n25579 ;
  assign n25581 = ~n25578 & ~n25579 ;
  assign n25582 = ~n25580 & ~n25581 ;
  assign n25583 = x102 & n4531 ;
  assign n25584 = x100 & n4847 ;
  assign n25585 = x101 & n4526 ;
  assign n25586 = ~n25584 & ~n25585 ;
  assign n25587 = ~n25583 & n25586 ;
  assign n25588 = n4534 & n10092 ;
  assign n25589 = n25587 & ~n25588 ;
  assign n25590 = x26 & ~n25589 ;
  assign n25591 = x26 & ~n25590 ;
  assign n25592 = ~n25589 & ~n25590 ;
  assign n25593 = ~n25591 & ~n25592 ;
  assign n25594 = n25582 & ~n25593 ;
  assign n25595 = n25582 & ~n25594 ;
  assign n25596 = ~n25593 & ~n25594 ;
  assign n25597 = ~n25595 & ~n25596 ;
  assign n25598 = ~n24816 & ~n24822 ;
  assign n25599 = n25597 & n25598 ;
  assign n25600 = ~n25597 & ~n25598 ;
  assign n25601 = ~n25599 & ~n25600 ;
  assign n25602 = x105 & n3589 ;
  assign n25603 = x103 & n3878 ;
  assign n25604 = x104 & n3584 ;
  assign n25605 = ~n25603 & ~n25604 ;
  assign n25606 = ~n25602 & n25605 ;
  assign n25607 = n3592 & n11648 ;
  assign n25608 = n25606 & ~n25607 ;
  assign n25609 = x23 & ~n25608 ;
  assign n25610 = x23 & ~n25609 ;
  assign n25611 = ~n25608 & ~n25609 ;
  assign n25612 = ~n25610 & ~n25611 ;
  assign n25613 = n25601 & ~n25612 ;
  assign n25614 = ~n25601 & n25612 ;
  assign n25615 = ~n25358 & ~n25614 ;
  assign n25616 = ~n25613 & n25615 ;
  assign n25617 = ~n25358 & ~n25616 ;
  assign n25618 = ~n25613 & ~n25616 ;
  assign n25619 = ~n25614 & n25618 ;
  assign n25620 = ~n25617 & ~n25619 ;
  assign n25621 = x108 & n2751 ;
  assign n25622 = x106 & n3020 ;
  assign n25623 = x107 & n2746 ;
  assign n25624 = ~n25622 & ~n25623 ;
  assign n25625 = ~n25621 & n25624 ;
  assign n25626 = n2754 & n13323 ;
  assign n25627 = n25625 & ~n25626 ;
  assign n25628 = x20 & ~n25627 ;
  assign n25629 = x20 & ~n25628 ;
  assign n25630 = ~n25627 & ~n25628 ;
  assign n25631 = ~n25629 & ~n25630 ;
  assign n25632 = ~n25620 & ~n25631 ;
  assign n25633 = ~n25620 & ~n25632 ;
  assign n25634 = ~n25631 & ~n25632 ;
  assign n25635 = ~n25633 & ~n25634 ;
  assign n25636 = ~n24859 & n25635 ;
  assign n25637 = n24859 & ~n25635 ;
  assign n25638 = ~n25636 & ~n25637 ;
  assign n25639 = x111 & n2093 ;
  assign n25640 = x109 & n2275 ;
  assign n25641 = x110 & n2088 ;
  assign n25642 = ~n25640 & ~n25641 ;
  assign n25643 = ~n25639 & n25642 ;
  assign n25644 = n2096 & n15111 ;
  assign n25645 = n25643 & ~n25644 ;
  assign n25646 = x17 & ~n25645 ;
  assign n25647 = x17 & ~n25646 ;
  assign n25648 = ~n25645 & ~n25646 ;
  assign n25649 = ~n25647 & ~n25648 ;
  assign n25650 = ~n25638 & ~n25649 ;
  assign n25651 = n25638 & n25649 ;
  assign n25652 = ~n25650 & ~n25651 ;
  assign n25653 = ~n25357 & n25652 ;
  assign n25654 = n25357 & ~n25652 ;
  assign n25655 = ~n25653 & ~n25654 ;
  assign n25656 = x114 & n1434 ;
  assign n25657 = x112 & n1646 ;
  assign n25658 = x113 & n1429 ;
  assign n25659 = ~n25657 & ~n25658 ;
  assign n25660 = ~n25656 & n25659 ;
  assign n25661 = n1437 & n17012 ;
  assign n25662 = n25660 & ~n25661 ;
  assign n25663 = x14 & ~n25662 ;
  assign n25664 = x14 & ~n25663 ;
  assign n25665 = ~n25662 & ~n25663 ;
  assign n25666 = ~n25664 & ~n25665 ;
  assign n25667 = n25655 & ~n25666 ;
  assign n25668 = n25655 & ~n25667 ;
  assign n25669 = ~n25666 & ~n25667 ;
  assign n25670 = ~n25668 & ~n25669 ;
  assign n25671 = ~n25356 & n25670 ;
  assign n25672 = n25356 & ~n25670 ;
  assign n25673 = ~n25671 & ~n25672 ;
  assign n25674 = x117 & n945 ;
  assign n25675 = x115 & n1099 ;
  assign n25676 = x116 & n940 ;
  assign n25677 = ~n25675 & ~n25676 ;
  assign n25678 = ~n25674 & n25677 ;
  assign n25679 = n948 & n19026 ;
  assign n25680 = n25678 & ~n25679 ;
  assign n25681 = x11 & ~n25680 ;
  assign n25682 = x11 & ~n25681 ;
  assign n25683 = ~n25680 & ~n25681 ;
  assign n25684 = ~n25682 & ~n25683 ;
  assign n25685 = ~n25673 & ~n25684 ;
  assign n25686 = n25673 & n25684 ;
  assign n25687 = ~n25685 & ~n25686 ;
  assign n25688 = ~n25355 & n25687 ;
  assign n25689 = n25355 & ~n25687 ;
  assign n25690 = ~n25688 & ~n25689 ;
  assign n25691 = x120 & n574 ;
  assign n25692 = x118 & n673 ;
  assign n25693 = x119 & n569 ;
  assign n25694 = ~n25692 & ~n25693 ;
  assign n25695 = ~n25691 & n25694 ;
  assign n25696 = n577 & n21143 ;
  assign n25697 = n25695 & ~n25696 ;
  assign n25698 = x8 & ~n25697 ;
  assign n25699 = x8 & ~n25698 ;
  assign n25700 = ~n25697 & ~n25698 ;
  assign n25701 = ~n25699 & ~n25700 ;
  assign n25702 = ~n25690 & n25701 ;
  assign n25703 = n25690 & ~n25701 ;
  assign n25704 = ~n25702 & ~n25703 ;
  assign n25705 = x123 & n293 ;
  assign n25706 = x121 & n373 ;
  assign n25707 = x122 & n288 ;
  assign n25708 = ~n25706 & ~n25707 ;
  assign n25709 = ~n25705 & n25708 ;
  assign n25710 = n296 & n23382 ;
  assign n25711 = n25709 & ~n25710 ;
  assign n25712 = x5 & ~n25711 ;
  assign n25713 = x5 & ~n25712 ;
  assign n25714 = ~n25711 & ~n25712 ;
  assign n25715 = ~n25713 & ~n25714 ;
  assign n25716 = n25704 & ~n25715 ;
  assign n25717 = n25704 & ~n25716 ;
  assign n25718 = ~n25715 & ~n25716 ;
  assign n25719 = ~n25717 & ~n25718 ;
  assign n25720 = ~n24902 & ~n24908 ;
  assign n25721 = n25719 & n25720 ;
  assign n25722 = ~n25719 & ~n25720 ;
  assign n25723 = ~n25721 & ~n25722 ;
  assign n25724 = x126 & n146 ;
  assign n25725 = x124 & n182 ;
  assign n25726 = x125 & n141 ;
  assign n25727 = ~n25725 & ~n25726 ;
  assign n25728 = ~n25724 & n25727 ;
  assign n25729 = ~n24931 & ~n24933 ;
  assign n25730 = ~x125 & ~x126 ;
  assign n25731 = x125 & x126 ;
  assign n25732 = ~n25730 & ~n25731 ;
  assign n25733 = ~n25729 & n25732 ;
  assign n25734 = n25729 & ~n25732 ;
  assign n25735 = ~n25733 & ~n25734 ;
  assign n25736 = n149 & n25735 ;
  assign n25737 = n25728 & ~n25736 ;
  assign n25738 = x2 & ~n25737 ;
  assign n25739 = x2 & ~n25738 ;
  assign n25740 = ~n25737 & ~n25738 ;
  assign n25741 = ~n25739 & ~n25740 ;
  assign n25742 = ~n25723 & n25741 ;
  assign n25743 = n25723 & ~n25741 ;
  assign n25744 = ~n25742 & ~n25743 ;
  assign n25745 = ~n25354 & n25744 ;
  assign n25746 = n25354 & ~n25744 ;
  assign n25747 = ~n25745 & ~n25746 ;
  assign n25748 = ~n25353 & n25747 ;
  assign n25749 = n25353 & ~n25747 ;
  assign n25750 = ~n25748 & ~n25749 ;
  assign n26145 = n25750 & x190 ;
  assign n25751 = ~n25343 & ~n25346 ;
  assign n25752 = ~n25320 & ~n25337 ;
  assign n25753 = ~n25284 & ~n25286 ;
  assign n25754 = ~n25278 & ~n25280 ;
  assign n25755 = ~n25272 & ~n25274 ;
  assign n25756 = ~n25233 & ~n25239 ;
  assign n25757 = ~n24982 & ~n25182 ;
  assign n25758 = ~n25179 & ~n25757 ;
  assign n25759 = ~n25122 & ~n25128 ;
  assign n25760 = ~n25084 & ~n25090 ;
  assign n25761 = ~x81 & n14233 ;
  assign n25762 = ~x79 & n14876 ;
  assign n25763 = ~x80 & n14228 ;
  assign n25764 = ~n25762 & ~n25763 ;
  assign n25765 = ~n25761 & n25764 ;
  assign n25766 = n2460 & n14236 ;
  assign n25767 = n25765 & ~n25766 ;
  assign n25768 = ~x47 & ~n25767 ;
  assign n25769 = ~x47 & ~n25768 ;
  assign n25770 = ~n25767 & ~n25768 ;
  assign n25771 = ~n25769 & ~n25770 ;
  assign n25772 = ~n25046 & ~n25052 ;
  assign n25773 = ~x75 & n18025 ;
  assign n25774 = ~x73 & n18764 ;
  assign n25775 = ~x74 & n18020 ;
  assign n25776 = ~n25774 & ~n25775 ;
  assign n25777 = ~n25773 & n25776 ;
  assign n25778 = n1225 & n18028 ;
  assign n25779 = n25777 & ~n25778 ;
  assign n25780 = ~x53 & ~n25779 ;
  assign n25781 = ~x53 & ~n25780 ;
  assign n25782 = ~n25779 & ~n25780 ;
  assign n25783 = ~n25781 & ~n25782 ;
  assign n25784 = ~n25030 & ~n25032 ;
  assign n25785 = ~n25024 & ~n25026 ;
  assign n25786 = ~x66 & n24612 ;
  assign n25787 = ~x64 & n25390 ;
  assign n25788 = ~x65 & n24607 ;
  assign n25789 = ~n25787 & ~n25788 ;
  assign n25790 = ~n25786 & n25789 ;
  assign n25791 = n214 & n24615 ;
  assign n25792 = n25790 & ~n25791 ;
  assign n25793 = ~x62 & ~n25792 ;
  assign n25794 = ~x62 & ~n25793 ;
  assign n25795 = ~n25792 & ~n25793 ;
  assign n25796 = ~n25794 & ~n25795 ;
  assign n25797 = ~n25020 & n25796 ;
  assign n25798 = n25020 & ~n25796 ;
  assign n25799 = ~n25797 & ~n25798 ;
  assign n25800 = ~x69 & n22325 ;
  assign n25801 = ~x67 & n23066 ;
  assign n25802 = ~x68 & n22320 ;
  assign n25803 = ~n25801 & ~n25802 ;
  assign n25804 = ~n25800 & n25803 ;
  assign n25805 = n435 & n22328 ;
  assign n25806 = n25804 & ~n25805 ;
  assign n25807 = ~x59 & ~n25806 ;
  assign n25808 = ~x59 & ~n25807 ;
  assign n25809 = ~n25806 & ~n25807 ;
  assign n25810 = ~n25808 & ~n25809 ;
  assign n25811 = n25799 & ~n25810 ;
  assign n25812 = ~n25799 & n25810 ;
  assign n25813 = ~n25785 & ~n25812 ;
  assign n25814 = ~n25811 & n25813 ;
  assign n25815 = ~n25785 & ~n25814 ;
  assign n25816 = ~n25811 & ~n25814 ;
  assign n25817 = ~n25812 & n25816 ;
  assign n25818 = ~n25815 & ~n25817 ;
  assign n25819 = ~x72 & n20143 ;
  assign n25820 = ~x70 & n20854 ;
  assign n25821 = ~x71 & n20138 ;
  assign n25822 = ~n25820 & ~n25821 ;
  assign n25823 = ~n25819 & n25822 ;
  assign n25824 = n773 & n20146 ;
  assign n25825 = n25823 & ~n25824 ;
  assign n25826 = ~x56 & ~n25825 ;
  assign n25827 = ~x56 & ~n25826 ;
  assign n25828 = ~n25825 & ~n25826 ;
  assign n25829 = ~n25827 & ~n25828 ;
  assign n25830 = n25818 & n25829 ;
  assign n25831 = ~n25818 & ~n25829 ;
  assign n25832 = ~n25830 & ~n25831 ;
  assign n25833 = ~n25784 & n25832 ;
  assign n25834 = n25784 & ~n25832 ;
  assign n25835 = ~n25833 & ~n25834 ;
  assign n25836 = n25783 & ~n25835 ;
  assign n25837 = ~n25783 & n25835 ;
  assign n25838 = ~n25836 & ~n25837 ;
  assign n25839 = ~n25772 & n25838 ;
  assign n25840 = n25772 & ~n25838 ;
  assign n25841 = ~n25839 & ~n25840 ;
  assign n25842 = ~x78 & n16076 ;
  assign n25843 = ~x76 & n16756 ;
  assign n25844 = ~x77 & n16071 ;
  assign n25845 = ~n25843 & ~n25844 ;
  assign n25846 = ~n25842 & n25845 ;
  assign n25847 = n1718 & n16079 ;
  assign n25848 = n25846 & ~n25847 ;
  assign n25849 = ~x50 & ~n25848 ;
  assign n25850 = ~x50 & ~n25849 ;
  assign n25851 = ~n25848 & ~n25849 ;
  assign n25852 = ~n25850 & ~n25851 ;
  assign n25853 = n25841 & ~n25852 ;
  assign n25854 = n25841 & ~n25853 ;
  assign n25855 = ~n25852 & ~n25853 ;
  assign n25856 = ~n25854 & ~n25855 ;
  assign n25857 = ~n25070 & ~n25856 ;
  assign n25858 = n25070 & n25856 ;
  assign n25859 = ~n25857 & ~n25858 ;
  assign n25860 = ~n25771 & n25859 ;
  assign n25861 = ~n25771 & ~n25860 ;
  assign n25862 = n25859 & ~n25860 ;
  assign n25863 = ~n25861 & ~n25862 ;
  assign n25864 = ~n25760 & ~n25863 ;
  assign n25865 = ~n25760 & ~n25864 ;
  assign n25866 = ~n25863 & ~n25864 ;
  assign n25867 = ~n25865 & ~n25866 ;
  assign n25868 = ~x84 & n12506 ;
  assign n25869 = ~x82 & n13131 ;
  assign n25870 = ~x83 & n12501 ;
  assign n25871 = ~n25869 & ~n25870 ;
  assign n25872 = ~n25868 & n25871 ;
  assign n25873 = n3247 & n12509 ;
  assign n25874 = n25872 & ~n25873 ;
  assign n25875 = ~x44 & ~n25874 ;
  assign n25876 = ~x44 & ~n25875 ;
  assign n25877 = ~n25874 & ~n25875 ;
  assign n25878 = ~n25876 & ~n25877 ;
  assign n25879 = ~n25867 & ~n25878 ;
  assign n25880 = ~n25867 & ~n25879 ;
  assign n25881 = ~n25878 & ~n25879 ;
  assign n25882 = ~n25880 & ~n25881 ;
  assign n25883 = ~n25108 & n25882 ;
  assign n25884 = n25108 & ~n25882 ;
  assign n25885 = ~n25883 & ~n25884 ;
  assign n25886 = ~x87 & n10905 ;
  assign n25887 = ~x85 & n11466 ;
  assign n25888 = ~x86 & n10900 ;
  assign n25889 = ~n25887 & ~n25888 ;
  assign n25890 = ~n25886 & n25889 ;
  assign n25891 = n4143 & n10908 ;
  assign n25892 = n25890 & ~n25891 ;
  assign n25893 = ~x41 & ~n25892 ;
  assign n25894 = ~x41 & ~n25893 ;
  assign n25895 = ~n25892 & ~n25893 ;
  assign n25896 = ~n25894 & ~n25895 ;
  assign n25897 = ~n25885 & ~n25896 ;
  assign n25898 = n25885 & n25896 ;
  assign n25899 = ~n25897 & ~n25898 ;
  assign n25900 = n25759 & ~n25899 ;
  assign n25901 = ~n25759 & n25899 ;
  assign n25902 = ~n25900 & ~n25901 ;
  assign n25903 = ~x90 & n9433 ;
  assign n25904 = ~x88 & n9915 ;
  assign n25905 = ~x89 & n9428 ;
  assign n25906 = ~n25904 & ~n25905 ;
  assign n25907 = ~n25903 & n25906 ;
  assign n25908 = n5155 & n9436 ;
  assign n25909 = n25907 & ~n25908 ;
  assign n25910 = ~x38 & ~n25909 ;
  assign n25911 = ~x38 & ~n25910 ;
  assign n25912 = ~n25909 & ~n25910 ;
  assign n25913 = ~n25911 & ~n25912 ;
  assign n25914 = n25902 & ~n25913 ;
  assign n25915 = n25902 & ~n25914 ;
  assign n25916 = ~n25913 & ~n25914 ;
  assign n25917 = ~n25915 & ~n25916 ;
  assign n25918 = ~n25141 & ~n25147 ;
  assign n25919 = n25917 & n25918 ;
  assign n25920 = ~n25917 & ~n25918 ;
  assign n25921 = ~n25919 & ~n25920 ;
  assign n25922 = ~x93 & n8006 ;
  assign n25923 = ~x91 & n8474 ;
  assign n25924 = ~x92 & n8001 ;
  assign n25925 = ~n25923 & ~n25924 ;
  assign n25926 = ~n25922 & n25925 ;
  assign n25927 = n6285 & n8009 ;
  assign n25928 = n25926 & ~n25927 ;
  assign n25929 = ~x35 & ~n25928 ;
  assign n25930 = ~x35 & ~n25929 ;
  assign n25931 = ~n25928 & ~n25929 ;
  assign n25932 = ~n25930 & ~n25931 ;
  assign n25933 = n25921 & ~n25932 ;
  assign n25934 = n25921 & ~n25933 ;
  assign n25935 = ~n25932 & ~n25933 ;
  assign n25936 = ~n25934 & ~n25935 ;
  assign n25937 = ~n25160 & ~n25166 ;
  assign n25938 = n25936 & n25937 ;
  assign n25939 = ~n25936 & ~n25937 ;
  assign n25940 = ~n25938 & ~n25939 ;
  assign n25941 = ~x96 & n6725 ;
  assign n25942 = ~x94 & n7129 ;
  assign n25943 = ~x95 & n6720 ;
  assign n25944 = ~n25942 & ~n25943 ;
  assign n25945 = ~n25941 & n25944 ;
  assign n25946 = n6728 & n7531 ;
  assign n25947 = n25945 & ~n25946 ;
  assign n25948 = ~x32 & ~n25947 ;
  assign n25949 = ~x32 & ~n25948 ;
  assign n25950 = ~n25947 & ~n25948 ;
  assign n25951 = ~n25949 & ~n25950 ;
  assign n25952 = n25940 & ~n25951 ;
  assign n25953 = ~n25940 & n25951 ;
  assign n25954 = ~n25758 & ~n25953 ;
  assign n25955 = ~n25952 & n25954 ;
  assign n25956 = ~n25758 & ~n25955 ;
  assign n25957 = ~n25952 & ~n25955 ;
  assign n25958 = ~n25953 & n25957 ;
  assign n25959 = ~n25956 & ~n25958 ;
  assign n25960 = ~x99 & n5560 ;
  assign n25961 = ~x97 & n5943 ;
  assign n25962 = ~x98 & n5555 ;
  assign n25963 = ~n25961 & ~n25962 ;
  assign n25964 = ~n25960 & n25963 ;
  assign n25965 = n5563 & n8885 ;
  assign n25966 = n25964 & ~n25965 ;
  assign n25967 = ~x29 & ~n25966 ;
  assign n25968 = ~x29 & ~n25967 ;
  assign n25969 = ~n25966 & ~n25967 ;
  assign n25970 = ~n25968 & ~n25969 ;
  assign n25971 = ~n25959 & ~n25970 ;
  assign n25972 = ~n25959 & ~n25971 ;
  assign n25973 = ~n25970 & ~n25971 ;
  assign n25974 = ~n25972 & ~n25973 ;
  assign n25975 = ~n25197 & ~n25201 ;
  assign n25976 = n25974 & n25975 ;
  assign n25977 = ~n25974 & ~n25975 ;
  assign n25978 = ~n25976 & ~n25977 ;
  assign n25979 = ~x102 & n4531 ;
  assign n25980 = ~x100 & n4847 ;
  assign n25981 = ~x101 & n4526 ;
  assign n25982 = ~n25980 & ~n25981 ;
  assign n25983 = ~n25979 & n25982 ;
  assign n25984 = n4534 & n10333 ;
  assign n25985 = n25983 & ~n25984 ;
  assign n25986 = ~x26 & ~n25985 ;
  assign n25987 = ~x26 & ~n25986 ;
  assign n25988 = ~n25985 & ~n25986 ;
  assign n25989 = ~n25987 & ~n25988 ;
  assign n25990 = n25978 & ~n25989 ;
  assign n25991 = n25978 & ~n25990 ;
  assign n25992 = ~n25989 & ~n25990 ;
  assign n25993 = ~n25991 & ~n25992 ;
  assign n25994 = ~n25214 & ~n25220 ;
  assign n25995 = n25993 & n25994 ;
  assign n25996 = ~n25993 & ~n25994 ;
  assign n25997 = ~n25995 & ~n25996 ;
  assign n25998 = ~x105 & n3589 ;
  assign n25999 = ~x103 & n3878 ;
  assign n26000 = ~x104 & n3584 ;
  assign n26001 = ~n25999 & ~n26000 ;
  assign n26002 = ~n25998 & n26001 ;
  assign n26003 = n3592 & n11907 ;
  assign n26004 = n26002 & ~n26003 ;
  assign n26005 = ~x23 & ~n26004 ;
  assign n26006 = ~x23 & ~n26005 ;
  assign n26007 = ~n26004 & ~n26005 ;
  assign n26008 = ~n26006 & ~n26007 ;
  assign n26009 = n25997 & ~n26008 ;
  assign n26010 = ~n25997 & n26008 ;
  assign n26011 = ~n25756 & ~n26010 ;
  assign n26012 = ~n26009 & n26011 ;
  assign n26013 = ~n25756 & ~n26012 ;
  assign n26014 = ~n26009 & ~n26012 ;
  assign n26015 = ~n26010 & n26014 ;
  assign n26016 = ~n26013 & ~n26015 ;
  assign n26017 = ~x108 & n2751 ;
  assign n26018 = ~x106 & n3020 ;
  assign n26019 = ~x107 & n2746 ;
  assign n26020 = ~n26018 & ~n26019 ;
  assign n26021 = ~n26017 & n26020 ;
  assign n26022 = n2754 & n13601 ;
  assign n26023 = n26021 & ~n26022 ;
  assign n26024 = ~x20 & ~n26023 ;
  assign n26025 = ~x20 & ~n26024 ;
  assign n26026 = ~n26023 & ~n26024 ;
  assign n26027 = ~n26025 & ~n26026 ;
  assign n26028 = ~n26016 & ~n26027 ;
  assign n26029 = ~n26016 & ~n26028 ;
  assign n26030 = ~n26027 & ~n26028 ;
  assign n26031 = ~n26029 & ~n26030 ;
  assign n26032 = ~n25257 & n26031 ;
  assign n26033 = n25257 & ~n26031 ;
  assign n26034 = ~n26032 & ~n26033 ;
  assign n26035 = ~x111 & n2093 ;
  assign n26036 = ~x109 & n2275 ;
  assign n26037 = ~x110 & n2088 ;
  assign n26038 = ~n26036 & ~n26037 ;
  assign n26039 = ~n26035 & n26038 ;
  assign n26040 = n2096 & n15411 ;
  assign n26041 = n26039 & ~n26040 ;
  assign n26042 = ~x17 & ~n26041 ;
  assign n26043 = ~x17 & ~n26042 ;
  assign n26044 = ~n26041 & ~n26042 ;
  assign n26045 = ~n26043 & ~n26044 ;
  assign n26046 = ~n26034 & ~n26045 ;
  assign n26047 = n26034 & n26045 ;
  assign n26048 = ~n26046 & ~n26047 ;
  assign n26049 = ~n25755 & n26048 ;
  assign n26050 = n25755 & ~n26048 ;
  assign n26051 = ~n26049 & ~n26050 ;
  assign n26052 = ~x114 & n1434 ;
  assign n26053 = ~x112 & n1646 ;
  assign n26054 = ~x113 & n1429 ;
  assign n26055 = ~n26053 & ~n26054 ;
  assign n26056 = ~n26052 & n26055 ;
  assign n26057 = n1437 & n17333 ;
  assign n26058 = n26056 & ~n26057 ;
  assign n26059 = ~x14 & ~n26058 ;
  assign n26060 = ~x14 & ~n26059 ;
  assign n26061 = ~n26058 & ~n26059 ;
  assign n26062 = ~n26060 & ~n26061 ;
  assign n26063 = n26051 & ~n26062 ;
  assign n26064 = n26051 & ~n26063 ;
  assign n26065 = ~n26062 & ~n26063 ;
  assign n26066 = ~n26064 & ~n26065 ;
  assign n26067 = ~n25754 & n26066 ;
  assign n26068 = n25754 & ~n26066 ;
  assign n26069 = ~n26067 & ~n26068 ;
  assign n26070 = ~x117 & n945 ;
  assign n26071 = ~x115 & n1099 ;
  assign n26072 = ~x116 & n940 ;
  assign n26073 = ~n26071 & ~n26072 ;
  assign n26074 = ~n26070 & n26073 ;
  assign n26075 = n948 & n19365 ;
  assign n26076 = n26074 & ~n26075 ;
  assign n26077 = ~x11 & ~n26076 ;
  assign n26078 = ~x11 & ~n26077 ;
  assign n26079 = ~n26076 & ~n26077 ;
  assign n26080 = ~n26078 & ~n26079 ;
  assign n26081 = ~n26069 & ~n26080 ;
  assign n26082 = n26069 & n26080 ;
  assign n26083 = ~n26081 & ~n26082 ;
  assign n26084 = ~n25753 & n26083 ;
  assign n26085 = n25753 & ~n26083 ;
  assign n26086 = ~n26084 & ~n26085 ;
  assign n26087 = ~x120 & n574 ;
  assign n26088 = ~x118 & n673 ;
  assign n26089 = ~x119 & n569 ;
  assign n26090 = ~n26088 & ~n26089 ;
  assign n26091 = ~n26087 & n26090 ;
  assign n26092 = n577 & n21501 ;
  assign n26093 = n26091 & ~n26092 ;
  assign n26094 = ~x8 & ~n26093 ;
  assign n26095 = ~x8 & ~n26094 ;
  assign n26096 = ~n26093 & ~n26094 ;
  assign n26097 = ~n26095 & ~n26096 ;
  assign n26098 = ~n26086 & n26097 ;
  assign n26099 = n26086 & ~n26097 ;
  assign n26100 = ~n26098 & ~n26099 ;
  assign n26101 = ~x123 & n293 ;
  assign n26102 = ~x121 & n373 ;
  assign n26103 = ~x122 & n288 ;
  assign n26104 = ~n26102 & ~n26103 ;
  assign n26105 = ~n26101 & n26104 ;
  assign n26106 = n296 & n23760 ;
  assign n26107 = n26105 & ~n26106 ;
  assign n26108 = ~x5 & ~n26107 ;
  assign n26109 = ~x5 & ~n26108 ;
  assign n26110 = ~n26107 & ~n26108 ;
  assign n26111 = ~n26109 & ~n26110 ;
  assign n26112 = n26100 & ~n26111 ;
  assign n26113 = n26100 & ~n26112 ;
  assign n26114 = ~n26111 & ~n26112 ;
  assign n26115 = ~n26113 & ~n26114 ;
  assign n26116 = ~n25300 & ~n25306 ;
  assign n26117 = n26115 & n26116 ;
  assign n26118 = ~n26115 & ~n26116 ;
  assign n26119 = ~n26117 & ~n26118 ;
  assign n26120 = ~x126 & n164 ;
  assign n26121 = ~x124 & n205 ;
  assign n26122 = ~x125 & n162 ;
  assign n26123 = ~n26121 & ~n26122 ;
  assign n26124 = ~n26120 & n26123 ;
  assign n26125 = ~n24930 & ~n25328 ;
  assign n26126 = n25732 & ~n26125 ;
  assign n26127 = ~n25732 & n26125 ;
  assign n26128 = ~n26126 & ~n26127 ;
  assign n26129 = n167 & n26128 ;
  assign n26130 = n26124 & ~n26129 ;
  assign n26131 = ~x2 & ~n26130 ;
  assign n26132 = ~x2 & ~n26131 ;
  assign n26133 = ~n26130 & ~n26131 ;
  assign n26134 = ~n26132 & ~n26133 ;
  assign n26135 = ~n26119 & n26134 ;
  assign n26136 = n26119 & ~n26134 ;
  assign n26137 = ~n26135 & ~n26136 ;
  assign n26138 = ~n25752 & n26137 ;
  assign n26139 = n25752 & ~n26137 ;
  assign n26140 = ~n26138 & ~n26139 ;
  assign n26141 = ~n25751 & n26140 ;
  assign n26142 = n25751 & ~n26140 ;
  assign n26143 = ~n26141 & ~n26142 ;
  assign n26146 = ~n26143 & ~x190 ;
  assign n26147 = ~n26145 & ~n26146 ;
  assign n26148 = ~n25356 & ~n25670 ;
  assign n26149 = ~n25667 & ~n26148 ;
  assign n26150 = x115 & n1434 ;
  assign n26151 = x113 & n1646 ;
  assign n26152 = x114 & n1429 ;
  assign n26153 = ~n26151 & ~n26152 ;
  assign n26154 = ~n26150 & n26153 ;
  assign n26155 = n1437 & n17364 ;
  assign n26156 = n26154 & ~n26155 ;
  assign n26157 = x14 & ~n26156 ;
  assign n26158 = x14 & ~n26157 ;
  assign n26159 = ~n26156 & ~n26157 ;
  assign n26160 = ~n26158 & ~n26159 ;
  assign n26161 = ~n25650 & ~n25653 ;
  assign n26162 = x112 & n2093 ;
  assign n26163 = x110 & n2275 ;
  assign n26164 = x111 & n2088 ;
  assign n26165 = ~n26163 & ~n26164 ;
  assign n26166 = ~n26162 & n26165 ;
  assign n26167 = n2096 & n15442 ;
  assign n26168 = n26166 & ~n26167 ;
  assign n26169 = x17 & ~n26168 ;
  assign n26170 = x17 & ~n26169 ;
  assign n26171 = ~n26168 & ~n26169 ;
  assign n26172 = ~n26170 & ~n26171 ;
  assign n26173 = ~n24859 & ~n25635 ;
  assign n26174 = ~n25632 & ~n26173 ;
  assign n26175 = x109 & n2751 ;
  assign n26176 = x107 & n3020 ;
  assign n26177 = x108 & n2746 ;
  assign n26178 = ~n26176 & ~n26177 ;
  assign n26179 = ~n26175 & n26178 ;
  assign n26180 = n2754 & n13894 ;
  assign n26181 = n26179 & ~n26180 ;
  assign n26182 = x20 & ~n26181 ;
  assign n26183 = x20 & ~n26182 ;
  assign n26184 = ~n26181 & ~n26182 ;
  assign n26185 = ~n26183 & ~n26184 ;
  assign n26186 = x106 & n3589 ;
  assign n26187 = x104 & n3878 ;
  assign n26188 = x105 & n3584 ;
  assign n26189 = ~n26187 & ~n26188 ;
  assign n26190 = ~n26186 & n26189 ;
  assign n26191 = n3592 & n12181 ;
  assign n26192 = n26190 & ~n26191 ;
  assign n26193 = x23 & ~n26192 ;
  assign n26194 = x23 & ~n26193 ;
  assign n26195 = ~n26192 & ~n26193 ;
  assign n26196 = ~n26194 & ~n26195 ;
  assign n26197 = ~n25594 & ~n25600 ;
  assign n26198 = ~n25575 & ~n25581 ;
  assign n26199 = ~n24710 & ~n25486 ;
  assign n26200 = ~n25483 & ~n26199 ;
  assign n26201 = x85 & n12506 ;
  assign n26202 = x83 & n13131 ;
  assign n26203 = x84 & n12501 ;
  assign n26204 = ~n26202 & ~n26203 ;
  assign n26205 = ~n26201 & n26204 ;
  assign n26206 = n3389 & n12509 ;
  assign n26207 = n26205 & ~n26206 ;
  assign n26208 = x44 & ~n26207 ;
  assign n26209 = x44 & ~n26208 ;
  assign n26210 = ~n26207 & ~n26208 ;
  assign n26211 = ~n26209 & ~n26210 ;
  assign n26212 = ~n25464 & ~n25468 ;
  assign n26213 = ~n25441 & ~n25443 ;
  assign n26214 = ~n25435 & ~n25437 ;
  assign n26215 = x62 & ~x63 ;
  assign n26216 = ~x62 & x63 ;
  assign n26217 = ~n26215 & ~n26216 ;
  assign n26218 = x64 & ~n26217 ;
  assign n26219 = n25402 & n26218 ;
  assign n26220 = n25402 & ~n26219 ;
  assign n26221 = n26218 & ~n26219 ;
  assign n26222 = ~n26220 & ~n26221 ;
  assign n26223 = x67 & n24612 ;
  assign n26224 = x65 & n25390 ;
  assign n26225 = x66 & n24607 ;
  assign n26226 = ~n26224 & ~n26225 ;
  assign n26227 = ~n26223 & n26226 ;
  assign n26228 = n240 & n24615 ;
  assign n26229 = n26227 & ~n26228 ;
  assign n26230 = x62 & ~n26229 ;
  assign n26231 = x62 & ~n26230 ;
  assign n26232 = ~n26229 & ~n26230 ;
  assign n26233 = ~n26231 & ~n26232 ;
  assign n26234 = ~n26222 & ~n26233 ;
  assign n26235 = ~n26222 & ~n26234 ;
  assign n26236 = ~n26233 & ~n26234 ;
  assign n26237 = ~n26235 & ~n26236 ;
  assign n26238 = x70 & n22325 ;
  assign n26239 = x68 & n23066 ;
  assign n26240 = x69 & n22320 ;
  assign n26241 = ~n26239 & ~n26240 ;
  assign n26242 = ~n26238 & n26241 ;
  assign n26243 = n488 & n22328 ;
  assign n26244 = n26242 & ~n26243 ;
  assign n26245 = x59 & ~n26244 ;
  assign n26246 = x59 & ~n26245 ;
  assign n26247 = ~n26244 & ~n26245 ;
  assign n26248 = ~n26246 & ~n26247 ;
  assign n26249 = n26237 & n26248 ;
  assign n26250 = ~n26237 & ~n26248 ;
  assign n26251 = ~n26249 & ~n26250 ;
  assign n26252 = ~n25420 & n26251 ;
  assign n26253 = n25420 & ~n26251 ;
  assign n26254 = ~n26252 & ~n26253 ;
  assign n26255 = x73 & n20143 ;
  assign n26256 = x71 & n20854 ;
  assign n26257 = x72 & n20138 ;
  assign n26258 = ~n26256 & ~n26257 ;
  assign n26259 = ~n26255 & n26258 ;
  assign n26260 = n843 & n20146 ;
  assign n26261 = n26259 & ~n26260 ;
  assign n26262 = x56 & ~n26261 ;
  assign n26263 = x56 & ~n26262 ;
  assign n26264 = ~n26261 & ~n26262 ;
  assign n26265 = ~n26263 & ~n26264 ;
  assign n26266 = n26254 & ~n26265 ;
  assign n26267 = n26254 & ~n26266 ;
  assign n26268 = ~n26265 & ~n26266 ;
  assign n26269 = ~n26267 & ~n26268 ;
  assign n26270 = ~n26214 & n26269 ;
  assign n26271 = n26214 & ~n26269 ;
  assign n26272 = ~n26270 & ~n26271 ;
  assign n26273 = x76 & n18025 ;
  assign n26274 = x74 & n18764 ;
  assign n26275 = x75 & n18020 ;
  assign n26276 = ~n26274 & ~n26275 ;
  assign n26277 = ~n26273 & n26276 ;
  assign n26278 = n1311 & n18028 ;
  assign n26279 = n26277 & ~n26278 ;
  assign n26280 = x53 & ~n26279 ;
  assign n26281 = x53 & ~n26280 ;
  assign n26282 = ~n26279 & ~n26280 ;
  assign n26283 = ~n26281 & ~n26282 ;
  assign n26284 = n26272 & n26283 ;
  assign n26285 = ~n26272 & ~n26283 ;
  assign n26286 = ~n26284 & ~n26285 ;
  assign n26287 = ~n26213 & n26286 ;
  assign n26288 = n26213 & ~n26286 ;
  assign n26289 = ~n26287 & ~n26288 ;
  assign n26290 = x79 & n16076 ;
  assign n26291 = x77 & n16756 ;
  assign n26292 = x78 & n16071 ;
  assign n26293 = ~n26291 & ~n26292 ;
  assign n26294 = ~n26290 & n26293 ;
  assign n26295 = n1817 & n16079 ;
  assign n26296 = n26294 & ~n26295 ;
  assign n26297 = x50 & ~n26296 ;
  assign n26298 = x50 & ~n26297 ;
  assign n26299 = ~n26296 & ~n26297 ;
  assign n26300 = ~n26298 & ~n26299 ;
  assign n26301 = n26289 & ~n26300 ;
  assign n26302 = n26289 & ~n26301 ;
  assign n26303 = ~n26300 & ~n26301 ;
  assign n26304 = ~n26302 & ~n26303 ;
  assign n26305 = ~n25457 & ~n25461 ;
  assign n26306 = n26304 & n26305 ;
  assign n26307 = ~n26304 & ~n26305 ;
  assign n26308 = ~n26306 & ~n26307 ;
  assign n26309 = x82 & n14233 ;
  assign n26310 = x80 & n14876 ;
  assign n26311 = x81 & n14228 ;
  assign n26312 = ~n26310 & ~n26311 ;
  assign n26313 = ~n26309 & n26312 ;
  assign n26314 = n2584 & n14236 ;
  assign n26315 = n26313 & ~n26314 ;
  assign n26316 = x47 & ~n26315 ;
  assign n26317 = x47 & ~n26316 ;
  assign n26318 = ~n26315 & ~n26316 ;
  assign n26319 = ~n26317 & ~n26318 ;
  assign n26320 = ~n26308 & n26319 ;
  assign n26321 = n26308 & ~n26319 ;
  assign n26322 = ~n26320 & ~n26321 ;
  assign n26323 = ~n26212 & n26322 ;
  assign n26324 = n26212 & ~n26322 ;
  assign n26325 = ~n26323 & ~n26324 ;
  assign n26326 = ~n26211 & n26325 ;
  assign n26327 = n26211 & ~n26325 ;
  assign n26328 = ~n26326 & ~n26327 ;
  assign n26329 = ~n26200 & n26328 ;
  assign n26330 = n26200 & ~n26328 ;
  assign n26331 = ~n26329 & ~n26330 ;
  assign n26332 = x88 & n10905 ;
  assign n26333 = x86 & n11466 ;
  assign n26334 = x87 & n10900 ;
  assign n26335 = ~n26333 & ~n26334 ;
  assign n26336 = ~n26332 & n26335 ;
  assign n26337 = n4305 & n10908 ;
  assign n26338 = n26336 & ~n26337 ;
  assign n26339 = x41 & ~n26338 ;
  assign n26340 = x41 & ~n26339 ;
  assign n26341 = ~n26338 & ~n26339 ;
  assign n26342 = ~n26340 & ~n26341 ;
  assign n26343 = n26331 & ~n26342 ;
  assign n26344 = n26331 & ~n26343 ;
  assign n26345 = ~n26342 & ~n26343 ;
  assign n26346 = ~n26344 & ~n26345 ;
  assign n26347 = ~n25501 & ~n25505 ;
  assign n26348 = n26346 & n26347 ;
  assign n26349 = ~n26346 & ~n26347 ;
  assign n26350 = ~n26348 & ~n26349 ;
  assign n26351 = x91 & n9433 ;
  assign n26352 = x89 & n9915 ;
  assign n26353 = x90 & n9428 ;
  assign n26354 = ~n26352 & ~n26353 ;
  assign n26355 = ~n26351 & n26354 ;
  assign n26356 = n5336 & n9436 ;
  assign n26357 = n26355 & ~n26356 ;
  assign n26358 = x38 & ~n26357 ;
  assign n26359 = x38 & ~n26358 ;
  assign n26360 = ~n26357 & ~n26358 ;
  assign n26361 = ~n26359 & ~n26360 ;
  assign n26362 = n26350 & ~n26361 ;
  assign n26363 = n26350 & ~n26362 ;
  assign n26364 = ~n26361 & ~n26362 ;
  assign n26365 = ~n26363 & ~n26364 ;
  assign n26366 = ~n25518 & ~n25524 ;
  assign n26367 = n26365 & n26366 ;
  assign n26368 = ~n26365 & ~n26366 ;
  assign n26369 = ~n26367 & ~n26368 ;
  assign n26370 = x94 & n8006 ;
  assign n26371 = x92 & n8474 ;
  assign n26372 = x93 & n8001 ;
  assign n26373 = ~n26371 & ~n26372 ;
  assign n26374 = ~n26370 & n26373 ;
  assign n26375 = n6483 & n8009 ;
  assign n26376 = n26374 & ~n26375 ;
  assign n26377 = x35 & ~n26376 ;
  assign n26378 = x35 & ~n26377 ;
  assign n26379 = ~n26376 & ~n26377 ;
  assign n26380 = ~n26378 & ~n26379 ;
  assign n26381 = ~n26369 & n26380 ;
  assign n26382 = n26369 & ~n26380 ;
  assign n26383 = ~n26381 & ~n26382 ;
  assign n26384 = ~n25537 & ~n25543 ;
  assign n26385 = n26383 & ~n26384 ;
  assign n26386 = ~n26383 & n26384 ;
  assign n26387 = ~n26385 & ~n26386 ;
  assign n26388 = x97 & n6725 ;
  assign n26389 = x95 & n7129 ;
  assign n26390 = x96 & n6720 ;
  assign n26391 = ~n26389 & ~n26390 ;
  assign n26392 = ~n26388 & n26391 ;
  assign n26393 = n6728 & n7745 ;
  assign n26394 = n26392 & ~n26393 ;
  assign n26395 = x32 & ~n26394 ;
  assign n26396 = x32 & ~n26395 ;
  assign n26397 = ~n26394 & ~n26395 ;
  assign n26398 = ~n26396 & ~n26397 ;
  assign n26399 = n26387 & ~n26398 ;
  assign n26400 = n26387 & ~n26399 ;
  assign n26401 = ~n26398 & ~n26399 ;
  assign n26402 = ~n26400 & ~n26401 ;
  assign n26403 = ~n25561 & n26402 ;
  assign n26404 = n25561 & ~n26402 ;
  assign n26405 = ~n26403 & ~n26404 ;
  assign n26406 = x100 & n5560 ;
  assign n26407 = x98 & n5943 ;
  assign n26408 = x99 & n5555 ;
  assign n26409 = ~n26407 & ~n26408 ;
  assign n26410 = ~n26406 & n26409 ;
  assign n26411 = n5563 & n9115 ;
  assign n26412 = n26410 & ~n26411 ;
  assign n26413 = x29 & ~n26412 ;
  assign n26414 = x29 & ~n26413 ;
  assign n26415 = ~n26412 & ~n26413 ;
  assign n26416 = ~n26414 & ~n26415 ;
  assign n26417 = ~n26405 & ~n26416 ;
  assign n26418 = n26405 & n26416 ;
  assign n26419 = ~n26417 & ~n26418 ;
  assign n26420 = n26198 & ~n26419 ;
  assign n26421 = ~n26198 & n26419 ;
  assign n26422 = ~n26420 & ~n26421 ;
  assign n26423 = x103 & n4531 ;
  assign n26424 = x101 & n4847 ;
  assign n26425 = x102 & n4526 ;
  assign n26426 = ~n26424 & ~n26425 ;
  assign n26427 = ~n26423 & n26426 ;
  assign n26428 = n4534 & n10588 ;
  assign n26429 = n26427 & ~n26428 ;
  assign n26430 = x26 & ~n26429 ;
  assign n26431 = x26 & ~n26430 ;
  assign n26432 = ~n26429 & ~n26430 ;
  assign n26433 = ~n26431 & ~n26432 ;
  assign n26434 = ~n26422 & n26433 ;
  assign n26435 = n26422 & ~n26433 ;
  assign n26436 = ~n26434 & ~n26435 ;
  assign n26437 = ~n26197 & n26436 ;
  assign n26438 = n26197 & ~n26436 ;
  assign n26439 = ~n26437 & ~n26438 ;
  assign n26440 = ~n26196 & n26439 ;
  assign n26441 = ~n26196 & ~n26440 ;
  assign n26442 = n26439 & ~n26440 ;
  assign n26443 = ~n26441 & ~n26442 ;
  assign n26444 = ~n25618 & ~n26443 ;
  assign n26445 = n25618 & ~n26442 ;
  assign n26446 = ~n26441 & n26445 ;
  assign n26447 = ~n26444 & ~n26446 ;
  assign n26448 = ~n26185 & n26447 ;
  assign n26449 = ~n26185 & ~n26448 ;
  assign n26450 = n26447 & ~n26448 ;
  assign n26451 = ~n26449 & ~n26450 ;
  assign n26452 = ~n26174 & ~n26451 ;
  assign n26453 = n26174 & ~n26450 ;
  assign n26454 = ~n26449 & n26453 ;
  assign n26455 = ~n26452 & ~n26454 ;
  assign n26456 = ~n26172 & n26455 ;
  assign n26457 = ~n26172 & ~n26456 ;
  assign n26458 = n26455 & ~n26456 ;
  assign n26459 = ~n26457 & ~n26458 ;
  assign n26460 = ~n26161 & ~n26459 ;
  assign n26461 = n26161 & ~n26458 ;
  assign n26462 = ~n26457 & n26461 ;
  assign n26463 = ~n26460 & ~n26462 ;
  assign n26464 = ~n26160 & n26463 ;
  assign n26465 = n26160 & ~n26463 ;
  assign n26466 = ~n26464 & ~n26465 ;
  assign n26467 = ~n26149 & n26466 ;
  assign n26468 = n26149 & ~n26466 ;
  assign n26469 = ~n26467 & ~n26468 ;
  assign n26470 = x118 & n945 ;
  assign n26471 = x116 & n1099 ;
  assign n26472 = x117 & n940 ;
  assign n26473 = ~n26471 & ~n26472 ;
  assign n26474 = ~n26470 & n26473 ;
  assign n26475 = n948 & n19395 ;
  assign n26476 = n26474 & ~n26475 ;
  assign n26477 = x11 & ~n26476 ;
  assign n26478 = x11 & ~n26477 ;
  assign n26479 = ~n26476 & ~n26477 ;
  assign n26480 = ~n26478 & ~n26479 ;
  assign n26481 = n26469 & ~n26480 ;
  assign n26482 = n26469 & ~n26481 ;
  assign n26483 = ~n26480 & ~n26481 ;
  assign n26484 = ~n26482 & ~n26483 ;
  assign n26485 = ~n25685 & ~n25688 ;
  assign n26486 = n26484 & n26485 ;
  assign n26487 = ~n26484 & ~n26485 ;
  assign n26488 = ~n26486 & ~n26487 ;
  assign n26489 = x121 & n574 ;
  assign n26490 = x119 & n673 ;
  assign n26491 = x120 & n569 ;
  assign n26492 = ~n26490 & ~n26491 ;
  assign n26493 = ~n26489 & n26492 ;
  assign n26494 = n577 & n21870 ;
  assign n26495 = n26493 & ~n26494 ;
  assign n26496 = x8 & ~n26495 ;
  assign n26497 = x8 & ~n26496 ;
  assign n26498 = ~n26495 & ~n26496 ;
  assign n26499 = ~n26497 & ~n26498 ;
  assign n26500 = n26488 & ~n26499 ;
  assign n26501 = n26488 & ~n26500 ;
  assign n26502 = ~n26499 & ~n26500 ;
  assign n26503 = ~n26501 & ~n26502 ;
  assign n26504 = x124 & n293 ;
  assign n26505 = x122 & n373 ;
  assign n26506 = x123 & n288 ;
  assign n26507 = ~n26505 & ~n26506 ;
  assign n26508 = ~n26504 & n26507 ;
  assign n26509 = n296 & n23796 ;
  assign n26510 = n26508 & ~n26509 ;
  assign n26511 = x5 & ~n26510 ;
  assign n26512 = x5 & ~n26511 ;
  assign n26513 = ~n26510 & ~n26511 ;
  assign n26514 = ~n26512 & ~n26513 ;
  assign n26515 = ~n26503 & n26514 ;
  assign n26516 = n26503 & ~n26514 ;
  assign n26517 = ~n26515 & ~n26516 ;
  assign n26518 = ~n25703 & ~n25716 ;
  assign n26519 = n26517 & n26518 ;
  assign n26520 = ~n26517 & ~n26518 ;
  assign n26521 = ~n26519 & ~n26520 ;
  assign n26522 = x127 & n146 ;
  assign n26523 = x125 & n182 ;
  assign n26524 = x126 & n141 ;
  assign n26525 = ~n26523 & ~n26524 ;
  assign n26526 = ~n26522 & n26525 ;
  assign n26527 = ~n25731 & ~n25733 ;
  assign n26528 = x126 & ~x127 ;
  assign n26529 = ~x126 & x127 ;
  assign n26530 = ~n26528 & ~n26529 ;
  assign n26531 = ~n26527 & ~n26530 ;
  assign n26532 = n26527 & n26530 ;
  assign n26533 = ~n26531 & ~n26532 ;
  assign n26534 = n149 & n26533 ;
  assign n26535 = n26526 & ~n26534 ;
  assign n26536 = x2 & ~n26535 ;
  assign n26537 = x2 & ~n26536 ;
  assign n26538 = ~n26535 & ~n26536 ;
  assign n26539 = ~n26537 & ~n26538 ;
  assign n26540 = n26521 & ~n26539 ;
  assign n26541 = n26521 & ~n26540 ;
  assign n26542 = ~n26539 & ~n26540 ;
  assign n26543 = ~n26541 & ~n26542 ;
  assign n26544 = ~n25722 & ~n25743 ;
  assign n26545 = ~n26543 & ~n26544 ;
  assign n26546 = ~n26543 & ~n26545 ;
  assign n26547 = ~n26544 & ~n26545 ;
  assign n26548 = ~n26546 & ~n26547 ;
  assign n26549 = ~n25745 & ~n25748 ;
  assign n26550 = ~n26548 & ~n26549 ;
  assign n26551 = n26548 & n26549 ;
  assign n26552 = ~n26550 & ~n26551 ;
  assign n26953 = n26552 & x191 ;
  assign n26553 = ~n25754 & ~n26066 ;
  assign n26554 = ~n26063 & ~n26553 ;
  assign n26555 = ~x115 & n1434 ;
  assign n26556 = ~x113 & n1646 ;
  assign n26557 = ~x114 & n1429 ;
  assign n26558 = ~n26556 & ~n26557 ;
  assign n26559 = ~n26555 & n26558 ;
  assign n26560 = n1437 & n17683 ;
  assign n26561 = n26559 & ~n26560 ;
  assign n26562 = ~x14 & ~n26561 ;
  assign n26563 = ~x14 & ~n26562 ;
  assign n26564 = ~n26561 & ~n26562 ;
  assign n26565 = ~n26563 & ~n26564 ;
  assign n26566 = ~n26046 & ~n26049 ;
  assign n26567 = ~x112 & n2093 ;
  assign n26568 = ~x110 & n2275 ;
  assign n26569 = ~x111 & n2088 ;
  assign n26570 = ~n26568 & ~n26569 ;
  assign n26571 = ~n26567 & n26570 ;
  assign n26572 = n2096 & n15744 ;
  assign n26573 = n26571 & ~n26572 ;
  assign n26574 = ~x17 & ~n26573 ;
  assign n26575 = ~x17 & ~n26574 ;
  assign n26576 = ~n26573 & ~n26574 ;
  assign n26577 = ~n26575 & ~n26576 ;
  assign n26578 = ~n25257 & ~n26031 ;
  assign n26579 = ~n26028 & ~n26578 ;
  assign n26580 = ~x109 & n2751 ;
  assign n26581 = ~x107 & n3020 ;
  assign n26582 = ~x108 & n2746 ;
  assign n26583 = ~n26581 & ~n26582 ;
  assign n26584 = ~n26580 & n26583 ;
  assign n26585 = n2754 & n14177 ;
  assign n26586 = n26584 & ~n26585 ;
  assign n26587 = ~x20 & ~n26586 ;
  assign n26588 = ~x20 & ~n26587 ;
  assign n26589 = ~n26586 & ~n26587 ;
  assign n26590 = ~n26588 & ~n26589 ;
  assign n26591 = ~x106 & n3589 ;
  assign n26592 = ~x104 & n3878 ;
  assign n26593 = ~x105 & n3584 ;
  assign n26594 = ~n26592 & ~n26593 ;
  assign n26595 = ~n26591 & n26594 ;
  assign n26596 = n3592 & n12447 ;
  assign n26597 = n26595 & ~n26596 ;
  assign n26598 = ~x23 & ~n26597 ;
  assign n26599 = ~x23 & ~n26598 ;
  assign n26600 = ~n26597 & ~n26598 ;
  assign n26601 = ~n26599 & ~n26600 ;
  assign n26602 = ~n25990 & ~n25996 ;
  assign n26603 = ~n25971 & ~n25977 ;
  assign n26604 = ~n25108 & ~n25882 ;
  assign n26605 = ~n25879 & ~n26604 ;
  assign n26606 = ~x85 & n12506 ;
  assign n26607 = ~x83 & n13131 ;
  assign n26608 = ~x84 & n12501 ;
  assign n26609 = ~n26607 & ~n26608 ;
  assign n26610 = ~n26606 & n26609 ;
  assign n26611 = n3521 & n12509 ;
  assign n26612 = n26610 & ~n26611 ;
  assign n26613 = ~x44 & ~n26612 ;
  assign n26614 = ~x44 & ~n26613 ;
  assign n26615 = ~n26612 & ~n26613 ;
  assign n26616 = ~n26614 & ~n26615 ;
  assign n26617 = ~n25860 & ~n25864 ;
  assign n26618 = ~n25837 & ~n25839 ;
  assign n26619 = ~n25831 & ~n25833 ;
  assign n26620 = ~x64 & ~n26217 ;
  assign n26621 = n25798 & n26620 ;
  assign n26622 = n25798 & ~n26621 ;
  assign n26623 = n26620 & ~n26621 ;
  assign n26624 = ~n26622 & ~n26623 ;
  assign n26625 = ~x67 & n24612 ;
  assign n26626 = ~x65 & n25390 ;
  assign n26627 = ~x66 & n24607 ;
  assign n26628 = ~n26626 & ~n26627 ;
  assign n26629 = ~n26625 & n26628 ;
  assign n26630 = n266 & n24615 ;
  assign n26631 = n26629 & ~n26630 ;
  assign n26632 = ~x62 & ~n26631 ;
  assign n26633 = ~x62 & ~n26632 ;
  assign n26634 = ~n26631 & ~n26632 ;
  assign n26635 = ~n26633 & ~n26634 ;
  assign n26636 = ~n26624 & ~n26635 ;
  assign n26637 = ~n26624 & ~n26636 ;
  assign n26638 = ~n26635 & ~n26636 ;
  assign n26639 = ~n26637 & ~n26638 ;
  assign n26640 = ~x70 & n22325 ;
  assign n26641 = ~x68 & n23066 ;
  assign n26642 = ~x69 & n22320 ;
  assign n26643 = ~n26641 & ~n26642 ;
  assign n26644 = ~n26640 & n26643 ;
  assign n26645 = n529 & n22328 ;
  assign n26646 = n26644 & ~n26645 ;
  assign n26647 = ~x59 & ~n26646 ;
  assign n26648 = ~x59 & ~n26647 ;
  assign n26649 = ~n26646 & ~n26647 ;
  assign n26650 = ~n26648 & ~n26649 ;
  assign n26651 = n26639 & n26650 ;
  assign n26652 = ~n26639 & ~n26650 ;
  assign n26653 = ~n26651 & ~n26652 ;
  assign n26654 = ~n25816 & n26653 ;
  assign n26655 = n25816 & ~n26653 ;
  assign n26656 = ~n26654 & ~n26655 ;
  assign n26657 = ~x73 & n20143 ;
  assign n26658 = ~x71 & n20854 ;
  assign n26659 = ~x72 & n20138 ;
  assign n26660 = ~n26658 & ~n26659 ;
  assign n26661 = ~n26657 & n26660 ;
  assign n26662 = n903 & n20146 ;
  assign n26663 = n26661 & ~n26662 ;
  assign n26664 = ~x56 & ~n26663 ;
  assign n26665 = ~x56 & ~n26664 ;
  assign n26666 = ~n26663 & ~n26664 ;
  assign n26667 = ~n26665 & ~n26666 ;
  assign n26668 = n26656 & ~n26667 ;
  assign n26669 = n26656 & ~n26668 ;
  assign n26670 = ~n26667 & ~n26668 ;
  assign n26671 = ~n26669 & ~n26670 ;
  assign n26672 = ~n26619 & n26671 ;
  assign n26673 = n26619 & ~n26671 ;
  assign n26674 = ~n26672 & ~n26673 ;
  assign n26675 = ~x76 & n18025 ;
  assign n26676 = ~x74 & n18764 ;
  assign n26677 = ~x75 & n18020 ;
  assign n26678 = ~n26676 & ~n26677 ;
  assign n26679 = ~n26675 & n26678 ;
  assign n26680 = n1390 & n18028 ;
  assign n26681 = n26679 & ~n26680 ;
  assign n26682 = ~x53 & ~n26681 ;
  assign n26683 = ~x53 & ~n26682 ;
  assign n26684 = ~n26681 & ~n26682 ;
  assign n26685 = ~n26683 & ~n26684 ;
  assign n26686 = n26674 & n26685 ;
  assign n26687 = ~n26674 & ~n26685 ;
  assign n26688 = ~n26686 & ~n26687 ;
  assign n26689 = ~n26618 & n26688 ;
  assign n26690 = n26618 & ~n26688 ;
  assign n26691 = ~n26689 & ~n26690 ;
  assign n26692 = ~x79 & n16076 ;
  assign n26693 = ~x77 & n16756 ;
  assign n26694 = ~x78 & n16071 ;
  assign n26695 = ~n26693 & ~n26694 ;
  assign n26696 = ~n26692 & n26695 ;
  assign n26697 = n1921 & n16079 ;
  assign n26698 = n26696 & ~n26697 ;
  assign n26699 = ~x50 & ~n26698 ;
  assign n26700 = ~x50 & ~n26699 ;
  assign n26701 = ~n26698 & ~n26699 ;
  assign n26702 = ~n26700 & ~n26701 ;
  assign n26703 = n26691 & ~n26702 ;
  assign n26704 = n26691 & ~n26703 ;
  assign n26705 = ~n26702 & ~n26703 ;
  assign n26706 = ~n26704 & ~n26705 ;
  assign n26707 = ~n25853 & ~n25857 ;
  assign n26708 = n26706 & n26707 ;
  assign n26709 = ~n26706 & ~n26707 ;
  assign n26710 = ~n26708 & ~n26709 ;
  assign n26711 = ~x82 & n14233 ;
  assign n26712 = ~x80 & n14876 ;
  assign n26713 = ~x81 & n14228 ;
  assign n26714 = ~n26712 & ~n26713 ;
  assign n26715 = ~n26711 & n26714 ;
  assign n26716 = n2697 & n14236 ;
  assign n26717 = n26715 & ~n26716 ;
  assign n26718 = ~x47 & ~n26717 ;
  assign n26719 = ~x47 & ~n26718 ;
  assign n26720 = ~n26717 & ~n26718 ;
  assign n26721 = ~n26719 & ~n26720 ;
  assign n26722 = ~n26710 & n26721 ;
  assign n26723 = n26710 & ~n26721 ;
  assign n26724 = ~n26722 & ~n26723 ;
  assign n26725 = ~n26617 & n26724 ;
  assign n26726 = n26617 & ~n26724 ;
  assign n26727 = ~n26725 & ~n26726 ;
  assign n26728 = ~n26616 & n26727 ;
  assign n26729 = n26616 & ~n26727 ;
  assign n26730 = ~n26728 & ~n26729 ;
  assign n26731 = ~n26605 & n26730 ;
  assign n26732 = n26605 & ~n26730 ;
  assign n26733 = ~n26731 & ~n26732 ;
  assign n26734 = ~x88 & n10905 ;
  assign n26735 = ~x86 & n11466 ;
  assign n26736 = ~x87 & n10900 ;
  assign n26737 = ~n26735 & ~n26736 ;
  assign n26738 = ~n26734 & n26737 ;
  assign n26739 = n4457 & n10908 ;
  assign n26740 = n26738 & ~n26739 ;
  assign n26741 = ~x41 & ~n26740 ;
  assign n26742 = ~x41 & ~n26741 ;
  assign n26743 = ~n26740 & ~n26741 ;
  assign n26744 = ~n26742 & ~n26743 ;
  assign n26745 = n26733 & ~n26744 ;
  assign n26746 = n26733 & ~n26745 ;
  assign n26747 = ~n26744 & ~n26745 ;
  assign n26748 = ~n26746 & ~n26747 ;
  assign n26749 = ~n25897 & ~n25901 ;
  assign n26750 = n26748 & n26749 ;
  assign n26751 = ~n26748 & ~n26749 ;
  assign n26752 = ~n26750 & ~n26751 ;
  assign n26753 = ~x91 & n9433 ;
  assign n26754 = ~x89 & n9915 ;
  assign n26755 = ~x90 & n9428 ;
  assign n26756 = ~n26754 & ~n26755 ;
  assign n26757 = ~n26753 & n26756 ;
  assign n26758 = n5507 & n9436 ;
  assign n26759 = n26757 & ~n26758 ;
  assign n26760 = ~x38 & ~n26759 ;
  assign n26761 = ~x38 & ~n26760 ;
  assign n26762 = ~n26759 & ~n26760 ;
  assign n26763 = ~n26761 & ~n26762 ;
  assign n26764 = n26752 & ~n26763 ;
  assign n26765 = n26752 & ~n26764 ;
  assign n26766 = ~n26763 & ~n26764 ;
  assign n26767 = ~n26765 & ~n26766 ;
  assign n26768 = ~n25914 & ~n25920 ;
  assign n26769 = n26767 & n26768 ;
  assign n26770 = ~n26767 & ~n26768 ;
  assign n26771 = ~n26769 & ~n26770 ;
  assign n26772 = ~x94 & n8006 ;
  assign n26773 = ~x92 & n8474 ;
  assign n26774 = ~x93 & n8001 ;
  assign n26775 = ~n26773 & ~n26774 ;
  assign n26776 = ~n26772 & n26775 ;
  assign n26777 = n6671 & n8009 ;
  assign n26778 = n26776 & ~n26777 ;
  assign n26779 = ~x35 & ~n26778 ;
  assign n26780 = ~x35 & ~n26779 ;
  assign n26781 = ~n26778 & ~n26779 ;
  assign n26782 = ~n26780 & ~n26781 ;
  assign n26783 = ~n26771 & n26782 ;
  assign n26784 = n26771 & ~n26782 ;
  assign n26785 = ~n26783 & ~n26784 ;
  assign n26786 = ~n25933 & ~n25939 ;
  assign n26787 = n26785 & ~n26786 ;
  assign n26788 = ~n26785 & n26786 ;
  assign n26789 = ~n26787 & ~n26788 ;
  assign n26790 = ~x97 & n6725 ;
  assign n26791 = ~x95 & n7129 ;
  assign n26792 = ~x96 & n6720 ;
  assign n26793 = ~n26791 & ~n26792 ;
  assign n26794 = ~n26790 & n26793 ;
  assign n26795 = n6728 & n7949 ;
  assign n26796 = n26794 & ~n26795 ;
  assign n26797 = ~x32 & ~n26796 ;
  assign n26798 = ~x32 & ~n26797 ;
  assign n26799 = ~n26796 & ~n26797 ;
  assign n26800 = ~n26798 & ~n26799 ;
  assign n26801 = n26789 & ~n26800 ;
  assign n26802 = n26789 & ~n26801 ;
  assign n26803 = ~n26800 & ~n26801 ;
  assign n26804 = ~n26802 & ~n26803 ;
  assign n26805 = ~n25957 & n26804 ;
  assign n26806 = n25957 & ~n26804 ;
  assign n26807 = ~n26805 & ~n26806 ;
  assign n26808 = ~x100 & n5560 ;
  assign n26809 = ~x98 & n5943 ;
  assign n26810 = ~x99 & n5555 ;
  assign n26811 = ~n26809 & ~n26810 ;
  assign n26812 = ~n26808 & n26811 ;
  assign n26813 = n5563 & n9338 ;
  assign n26814 = n26812 & ~n26813 ;
  assign n26815 = ~x29 & ~n26814 ;
  assign n26816 = ~x29 & ~n26815 ;
  assign n26817 = ~n26814 & ~n26815 ;
  assign n26818 = ~n26816 & ~n26817 ;
  assign n26819 = ~n26807 & ~n26818 ;
  assign n26820 = n26807 & n26818 ;
  assign n26821 = ~n26819 & ~n26820 ;
  assign n26822 = n26603 & ~n26821 ;
  assign n26823 = ~n26603 & n26821 ;
  assign n26824 = ~n26822 & ~n26823 ;
  assign n26825 = ~x103 & n4531 ;
  assign n26826 = ~x101 & n4847 ;
  assign n26827 = ~x102 & n4526 ;
  assign n26828 = ~n26826 & ~n26827 ;
  assign n26829 = ~n26825 & n26828 ;
  assign n26830 = n4534 & n10833 ;
  assign n26831 = n26829 & ~n26830 ;
  assign n26832 = ~x26 & ~n26831 ;
  assign n26833 = ~x26 & ~n26832 ;
  assign n26834 = ~n26831 & ~n26832 ;
  assign n26835 = ~n26833 & ~n26834 ;
  assign n26836 = ~n26824 & n26835 ;
  assign n26837 = n26824 & ~n26835 ;
  assign n26838 = ~n26836 & ~n26837 ;
  assign n26839 = ~n26602 & n26838 ;
  assign n26840 = n26602 & ~n26838 ;
  assign n26841 = ~n26839 & ~n26840 ;
  assign n26842 = ~n26601 & n26841 ;
  assign n26843 = ~n26601 & ~n26842 ;
  assign n26844 = n26841 & ~n26842 ;
  assign n26845 = ~n26843 & ~n26844 ;
  assign n26846 = ~n26014 & ~n26845 ;
  assign n26847 = n26014 & ~n26844 ;
  assign n26848 = ~n26843 & n26847 ;
  assign n26849 = ~n26846 & ~n26848 ;
  assign n26850 = ~n26590 & n26849 ;
  assign n26851 = ~n26590 & ~n26850 ;
  assign n26852 = n26849 & ~n26850 ;
  assign n26853 = ~n26851 & ~n26852 ;
  assign n26854 = ~n26579 & ~n26853 ;
  assign n26855 = n26579 & ~n26852 ;
  assign n26856 = ~n26851 & n26855 ;
  assign n26857 = ~n26854 & ~n26856 ;
  assign n26858 = ~n26577 & n26857 ;
  assign n26859 = ~n26577 & ~n26858 ;
  assign n26860 = n26857 & ~n26858 ;
  assign n26861 = ~n26859 & ~n26860 ;
  assign n26862 = ~n26566 & ~n26861 ;
  assign n26863 = n26566 & ~n26860 ;
  assign n26864 = ~n26859 & n26863 ;
  assign n26865 = ~n26862 & ~n26864 ;
  assign n26866 = ~n26565 & n26865 ;
  assign n26867 = n26565 & ~n26865 ;
  assign n26868 = ~n26866 & ~n26867 ;
  assign n26869 = ~n26554 & n26868 ;
  assign n26870 = n26554 & ~n26868 ;
  assign n26871 = ~n26869 & ~n26870 ;
  assign n26872 = ~x118 & n945 ;
  assign n26873 = ~x116 & n1099 ;
  assign n26874 = ~x117 & n940 ;
  assign n26875 = ~n26873 & ~n26874 ;
  assign n26876 = ~n26872 & n26875 ;
  assign n26877 = n948 & n19736 ;
  assign n26878 = n26876 & ~n26877 ;
  assign n26879 = ~x11 & ~n26878 ;
  assign n26880 = ~x11 & ~n26879 ;
  assign n26881 = ~n26878 & ~n26879 ;
  assign n26882 = ~n26880 & ~n26881 ;
  assign n26883 = n26871 & ~n26882 ;
  assign n26884 = n26871 & ~n26883 ;
  assign n26885 = ~n26882 & ~n26883 ;
  assign n26886 = ~n26884 & ~n26885 ;
  assign n26887 = ~n26081 & ~n26084 ;
  assign n26888 = n26886 & n26887 ;
  assign n26889 = ~n26886 & ~n26887 ;
  assign n26890 = ~n26888 & ~n26889 ;
  assign n26891 = ~x121 & n574 ;
  assign n26892 = ~x119 & n673 ;
  assign n26893 = ~x120 & n569 ;
  assign n26894 = ~n26892 & ~n26893 ;
  assign n26895 = ~n26891 & n26894 ;
  assign n26896 = n577 & n22229 ;
  assign n26897 = n26895 & ~n26896 ;
  assign n26898 = ~x8 & ~n26897 ;
  assign n26899 = ~x8 & ~n26898 ;
  assign n26900 = ~n26897 & ~n26898 ;
  assign n26901 = ~n26899 & ~n26900 ;
  assign n26902 = n26890 & ~n26901 ;
  assign n26903 = n26890 & ~n26902 ;
  assign n26904 = ~n26901 & ~n26902 ;
  assign n26905 = ~n26903 & ~n26904 ;
  assign n26906 = ~x124 & n293 ;
  assign n26907 = ~x122 & n373 ;
  assign n26908 = ~x123 & n288 ;
  assign n26909 = ~n26907 & ~n26908 ;
  assign n26910 = ~n26906 & n26909 ;
  assign n26911 = n296 & n24176 ;
  assign n26912 = n26910 & ~n26911 ;
  assign n26913 = ~x5 & ~n26912 ;
  assign n26914 = ~x5 & ~n26913 ;
  assign n26915 = ~n26912 & ~n26913 ;
  assign n26916 = ~n26914 & ~n26915 ;
  assign n26917 = ~n26905 & n26916 ;
  assign n26918 = n26905 & ~n26916 ;
  assign n26919 = ~n26917 & ~n26918 ;
  assign n26920 = ~n26099 & ~n26112 ;
  assign n26921 = n26919 & n26920 ;
  assign n26922 = ~n26919 & ~n26920 ;
  assign n26923 = ~n26921 & ~n26922 ;
  assign n26924 = ~x127 & n164 ;
  assign n26925 = ~x125 & n205 ;
  assign n26926 = ~x126 & n162 ;
  assign n26927 = ~n26925 & ~n26926 ;
  assign n26928 = ~n26924 & n26927 ;
  assign n26929 = ~n25730 & ~n26126 ;
  assign n26930 = ~n26530 & ~n26929 ;
  assign n26931 = n26530 & n26929 ;
  assign n26932 = ~n26930 & ~n26931 ;
  assign n26933 = n167 & n26932 ;
  assign n26934 = n26928 & ~n26933 ;
  assign n26935 = ~x2 & ~n26934 ;
  assign n26936 = ~x2 & ~n26935 ;
  assign n26937 = ~n26934 & ~n26935 ;
  assign n26938 = ~n26936 & ~n26937 ;
  assign n26939 = n26923 & ~n26938 ;
  assign n26940 = n26923 & ~n26939 ;
  assign n26941 = ~n26938 & ~n26939 ;
  assign n26942 = ~n26940 & ~n26941 ;
  assign n26943 = ~n26118 & ~n26136 ;
  assign n26944 = ~n26942 & ~n26943 ;
  assign n26945 = ~n26942 & ~n26944 ;
  assign n26946 = ~n26943 & ~n26944 ;
  assign n26947 = ~n26945 & ~n26946 ;
  assign n26948 = ~n26138 & ~n26141 ;
  assign n26949 = ~n26947 & ~n26948 ;
  assign n26950 = n26947 & n26948 ;
  assign n26951 = ~n26949 & ~n26950 ;
  assign n26954 = ~n26951 & ~x191 ;
  assign n26955 = ~n26953 & ~n26954 ;
  assign n26956 = ~n26545 & ~n26550 ;
  assign n26957 = ~n26520 & ~n26540 ;
  assign n26958 = x126 & n182 ;
  assign n26959 = x127 & n141 ;
  assign n26960 = ~n26958 & ~n26959 ;
  assign n26961 = ~x126 & ~n26531 ;
  assign n26962 = x127 & ~n26961 ;
  assign n26963 = x127 & ~n26962 ;
  assign n26964 = ~n26527 & n26528 ;
  assign n26965 = ~n26963 & ~n26964 ;
  assign n26966 = n149 & ~n26965 ;
  assign n26967 = n26960 & ~n26966 ;
  assign n26968 = x2 & ~n26967 ;
  assign n26969 = x2 & ~n26968 ;
  assign n26970 = ~n26967 & ~n26968 ;
  assign n26971 = ~n26969 & ~n26970 ;
  assign n26972 = ~n26503 & ~n26514 ;
  assign n26973 = ~n26500 & ~n26972 ;
  assign n26974 = ~n26481 & ~n26487 ;
  assign n26975 = x119 & n945 ;
  assign n26976 = x117 & n1099 ;
  assign n26977 = x118 & n940 ;
  assign n26978 = ~n26976 & ~n26977 ;
  assign n26979 = ~n26975 & n26978 ;
  assign n26980 = n948 & n20423 ;
  assign n26981 = n26979 & ~n26980 ;
  assign n26982 = x11 & ~n26981 ;
  assign n26983 = x11 & ~n26982 ;
  assign n26984 = ~n26981 & ~n26982 ;
  assign n26985 = ~n26983 & ~n26984 ;
  assign n26986 = ~n26464 & ~n26467 ;
  assign n26987 = x116 & n1434 ;
  assign n26988 = x114 & n1646 ;
  assign n26989 = x115 & n1429 ;
  assign n26990 = ~n26988 & ~n26989 ;
  assign n26991 = ~n26987 & n26990 ;
  assign n26992 = n1437 & n18336 ;
  assign n26993 = n26991 & ~n26992 ;
  assign n26994 = x14 & ~n26993 ;
  assign n26995 = x14 & ~n26994 ;
  assign n26996 = ~n26993 & ~n26994 ;
  assign n26997 = ~n26995 & ~n26996 ;
  assign n26998 = ~n26456 & ~n26460 ;
  assign n26999 = x113 & n2093 ;
  assign n27000 = x111 & n2275 ;
  assign n27001 = x112 & n2088 ;
  assign n27002 = ~n27000 & ~n27001 ;
  assign n27003 = ~n26999 & n27002 ;
  assign n27004 = n2096 & n16361 ;
  assign n27005 = n27003 & ~n27004 ;
  assign n27006 = x17 & ~n27005 ;
  assign n27007 = x17 & ~n27006 ;
  assign n27008 = ~n27005 & ~n27006 ;
  assign n27009 = ~n27007 & ~n27008 ;
  assign n27010 = ~n26448 & ~n26452 ;
  assign n27011 = x110 & n2751 ;
  assign n27012 = x108 & n3020 ;
  assign n27013 = x109 & n2746 ;
  assign n27014 = ~n27012 & ~n27013 ;
  assign n27015 = ~n27011 & n27014 ;
  assign n27016 = n2754 & n14497 ;
  assign n27017 = n27015 & ~n27016 ;
  assign n27018 = x20 & ~n27017 ;
  assign n27019 = x20 & ~n27018 ;
  assign n27020 = ~n27017 & ~n27018 ;
  assign n27021 = ~n27019 & ~n27020 ;
  assign n27022 = ~n26440 & ~n26444 ;
  assign n27023 = ~n26250 & ~n26252 ;
  assign n27024 = x63 & n26217 ;
  assign n27025 = x64 & n27024 ;
  assign n27026 = x65 & ~n26217 ;
  assign n27027 = ~n27025 & ~n27026 ;
  assign n27028 = x68 & n24612 ;
  assign n27029 = x66 & n25390 ;
  assign n27030 = x67 & n24607 ;
  assign n27031 = ~n27029 & ~n27030 ;
  assign n27032 = ~n27028 & n27031 ;
  assign n27033 = n317 & n24615 ;
  assign n27034 = n27032 & ~n27033 ;
  assign n27035 = x62 & ~n27034 ;
  assign n27036 = x62 & ~n27035 ;
  assign n27037 = ~n27034 & ~n27035 ;
  assign n27038 = ~n27036 & ~n27037 ;
  assign n27039 = ~n27027 & ~n27038 ;
  assign n27040 = ~n27027 & ~n27039 ;
  assign n27041 = ~n27038 & ~n27039 ;
  assign n27042 = ~n27040 & ~n27041 ;
  assign n27043 = ~n26219 & ~n26234 ;
  assign n27044 = n27042 & n27043 ;
  assign n27045 = ~n27042 & ~n27043 ;
  assign n27046 = ~n27044 & ~n27045 ;
  assign n27047 = x71 & n22325 ;
  assign n27048 = x69 & n23066 ;
  assign n27049 = x70 & n22320 ;
  assign n27050 = ~n27048 & ~n27049 ;
  assign n27051 = ~n27047 & n27050 ;
  assign n27052 = n558 & n22328 ;
  assign n27053 = n27051 & ~n27052 ;
  assign n27054 = x59 & ~n27053 ;
  assign n27055 = x59 & ~n27054 ;
  assign n27056 = ~n27053 & ~n27054 ;
  assign n27057 = ~n27055 & ~n27056 ;
  assign n27058 = ~n27046 & n27057 ;
  assign n27059 = n27046 & ~n27057 ;
  assign n27060 = ~n27058 & ~n27059 ;
  assign n27061 = ~n27023 & n27060 ;
  assign n27062 = n27023 & ~n27060 ;
  assign n27063 = ~n27061 & ~n27062 ;
  assign n27064 = x74 & n20143 ;
  assign n27065 = x72 & n20854 ;
  assign n27066 = x73 & n20138 ;
  assign n27067 = ~n27065 & ~n27066 ;
  assign n27068 = ~n27064 & n27067 ;
  assign n27069 = n994 & n20146 ;
  assign n27070 = n27068 & ~n27069 ;
  assign n27071 = x56 & ~n27070 ;
  assign n27072 = x56 & ~n27071 ;
  assign n27073 = ~n27070 & ~n27071 ;
  assign n27074 = ~n27072 & ~n27073 ;
  assign n27075 = n27063 & ~n27074 ;
  assign n27076 = n27063 & ~n27075 ;
  assign n27077 = ~n27074 & ~n27075 ;
  assign n27078 = ~n27076 & ~n27077 ;
  assign n27079 = ~n26214 & ~n26269 ;
  assign n27080 = ~n26266 & ~n27079 ;
  assign n27081 = n27078 & n27080 ;
  assign n27082 = ~n27078 & ~n27080 ;
  assign n27083 = ~n27081 & ~n27082 ;
  assign n27084 = x77 & n18025 ;
  assign n27085 = x75 & n18764 ;
  assign n27086 = x76 & n18020 ;
  assign n27087 = ~n27085 & ~n27086 ;
  assign n27088 = ~n27084 & n27087 ;
  assign n27089 = n1502 & n18028 ;
  assign n27090 = n27088 & ~n27089 ;
  assign n27091 = x53 & ~n27090 ;
  assign n27092 = x53 & ~n27091 ;
  assign n27093 = ~n27090 & ~n27091 ;
  assign n27094 = ~n27092 & ~n27093 ;
  assign n27095 = ~n27083 & n27094 ;
  assign n27096 = n27083 & ~n27094 ;
  assign n27097 = ~n27095 & ~n27096 ;
  assign n27098 = ~n26285 & ~n26287 ;
  assign n27099 = n27097 & ~n27098 ;
  assign n27100 = ~n27097 & n27098 ;
  assign n27101 = ~n27099 & ~n27100 ;
  assign n27102 = x80 & n16076 ;
  assign n27103 = x78 & n16756 ;
  assign n27104 = x79 & n16071 ;
  assign n27105 = ~n27103 & ~n27104 ;
  assign n27106 = ~n27102 & n27105 ;
  assign n27107 = n2028 & n16079 ;
  assign n27108 = n27106 & ~n27107 ;
  assign n27109 = x50 & ~n27108 ;
  assign n27110 = x50 & ~n27109 ;
  assign n27111 = ~n27108 & ~n27109 ;
  assign n27112 = ~n27110 & ~n27111 ;
  assign n27113 = n27101 & ~n27112 ;
  assign n27114 = n27101 & ~n27113 ;
  assign n27115 = ~n27112 & ~n27113 ;
  assign n27116 = ~n27114 & ~n27115 ;
  assign n27117 = ~n26301 & ~n26307 ;
  assign n27118 = n27116 & n27117 ;
  assign n27119 = ~n27116 & ~n27117 ;
  assign n27120 = ~n27118 & ~n27119 ;
  assign n27121 = x83 & n14233 ;
  assign n27122 = x81 & n14876 ;
  assign n27123 = x82 & n14228 ;
  assign n27124 = ~n27122 & ~n27123 ;
  assign n27125 = ~n27121 & n27124 ;
  assign n27126 = n2843 & n14236 ;
  assign n27127 = n27125 & ~n27126 ;
  assign n27128 = x47 & ~n27127 ;
  assign n27129 = x47 & ~n27128 ;
  assign n27130 = ~n27127 & ~n27128 ;
  assign n27131 = ~n27129 & ~n27130 ;
  assign n27132 = ~n27120 & n27131 ;
  assign n27133 = n27120 & ~n27131 ;
  assign n27134 = ~n27132 & ~n27133 ;
  assign n27135 = ~n26321 & ~n26323 ;
  assign n27136 = n27134 & ~n27135 ;
  assign n27137 = ~n27134 & n27135 ;
  assign n27138 = ~n27136 & ~n27137 ;
  assign n27139 = x86 & n12506 ;
  assign n27140 = x84 & n13131 ;
  assign n27141 = x85 & n12501 ;
  assign n27142 = ~n27140 & ~n27141 ;
  assign n27143 = ~n27139 & n27142 ;
  assign n27144 = n3686 & n12509 ;
  assign n27145 = n27143 & ~n27144 ;
  assign n27146 = x44 & ~n27145 ;
  assign n27147 = x44 & ~n27146 ;
  assign n27148 = ~n27145 & ~n27146 ;
  assign n27149 = ~n27147 & ~n27148 ;
  assign n27150 = n27138 & ~n27149 ;
  assign n27151 = n27138 & ~n27150 ;
  assign n27152 = ~n27149 & ~n27150 ;
  assign n27153 = ~n27151 & ~n27152 ;
  assign n27154 = ~n26326 & ~n26329 ;
  assign n27155 = n27153 & n27154 ;
  assign n27156 = ~n27153 & ~n27154 ;
  assign n27157 = ~n27155 & ~n27156 ;
  assign n27158 = x89 & n10905 ;
  assign n27159 = x87 & n11466 ;
  assign n27160 = x88 & n10900 ;
  assign n27161 = ~n27159 & ~n27160 ;
  assign n27162 = ~n27158 & n27161 ;
  assign n27163 = n4488 & n10908 ;
  assign n27164 = n27162 & ~n27163 ;
  assign n27165 = x41 & ~n27164 ;
  assign n27166 = x41 & ~n27165 ;
  assign n27167 = ~n27164 & ~n27165 ;
  assign n27168 = ~n27166 & ~n27167 ;
  assign n27169 = n27157 & ~n27168 ;
  assign n27170 = n27157 & ~n27169 ;
  assign n27171 = ~n27168 & ~n27169 ;
  assign n27172 = ~n27170 & ~n27171 ;
  assign n27173 = ~n26343 & ~n26349 ;
  assign n27174 = n27172 & n27173 ;
  assign n27175 = ~n27172 & ~n27173 ;
  assign n27176 = ~n27174 & ~n27175 ;
  assign n27177 = x92 & n9433 ;
  assign n27178 = x90 & n9915 ;
  assign n27179 = x91 & n9428 ;
  assign n27180 = ~n27178 & ~n27179 ;
  assign n27181 = ~n27177 & n27180 ;
  assign n27182 = n5710 & n9436 ;
  assign n27183 = n27181 & ~n27182 ;
  assign n27184 = x38 & ~n27183 ;
  assign n27185 = x38 & ~n27184 ;
  assign n27186 = ~n27183 & ~n27184 ;
  assign n27187 = ~n27185 & ~n27186 ;
  assign n27188 = n27176 & ~n27187 ;
  assign n27189 = n27176 & ~n27188 ;
  assign n27190 = ~n27187 & ~n27188 ;
  assign n27191 = ~n27189 & ~n27190 ;
  assign n27192 = ~n26362 & ~n26368 ;
  assign n27193 = n27191 & n27192 ;
  assign n27194 = ~n27191 & ~n27192 ;
  assign n27195 = ~n27193 & ~n27194 ;
  assign n27196 = x95 & n8006 ;
  assign n27197 = x93 & n8474 ;
  assign n27198 = x94 & n8001 ;
  assign n27199 = ~n27197 & ~n27198 ;
  assign n27200 = ~n27196 & n27199 ;
  assign n27201 = n6894 & n8009 ;
  assign n27202 = n27200 & ~n27201 ;
  assign n27203 = x35 & ~n27202 ;
  assign n27204 = x35 & ~n27203 ;
  assign n27205 = ~n27202 & ~n27203 ;
  assign n27206 = ~n27204 & ~n27205 ;
  assign n27207 = ~n27195 & n27206 ;
  assign n27208 = n27195 & ~n27206 ;
  assign n27209 = ~n27207 & ~n27208 ;
  assign n27210 = ~n26382 & ~n26385 ;
  assign n27211 = n27209 & ~n27210 ;
  assign n27212 = ~n27209 & n27210 ;
  assign n27213 = ~n27211 & ~n27212 ;
  assign n27214 = x98 & n6725 ;
  assign n27215 = x96 & n7129 ;
  assign n27216 = x97 & n6720 ;
  assign n27217 = ~n27215 & ~n27216 ;
  assign n27218 = ~n27214 & n27217 ;
  assign n27219 = n6728 & n8196 ;
  assign n27220 = n27218 & ~n27219 ;
  assign n27221 = x32 & ~n27220 ;
  assign n27222 = x32 & ~n27221 ;
  assign n27223 = ~n27220 & ~n27221 ;
  assign n27224 = ~n27222 & ~n27223 ;
  assign n27225 = n27213 & ~n27224 ;
  assign n27226 = n27213 & ~n27225 ;
  assign n27227 = ~n27224 & ~n27225 ;
  assign n27228 = ~n27226 & ~n27227 ;
  assign n27229 = ~n25561 & ~n26402 ;
  assign n27230 = ~n26399 & ~n27229 ;
  assign n27231 = n27228 & n27230 ;
  assign n27232 = ~n27228 & ~n27230 ;
  assign n27233 = ~n27231 & ~n27232 ;
  assign n27234 = x101 & n5560 ;
  assign n27235 = x99 & n5943 ;
  assign n27236 = x100 & n5555 ;
  assign n27237 = ~n27235 & ~n27236 ;
  assign n27238 = ~n27234 & n27237 ;
  assign n27239 = n5563 & n9601 ;
  assign n27240 = n27238 & ~n27239 ;
  assign n27241 = x29 & ~n27240 ;
  assign n27242 = x29 & ~n27241 ;
  assign n27243 = ~n27240 & ~n27241 ;
  assign n27244 = ~n27242 & ~n27243 ;
  assign n27245 = n27233 & ~n27244 ;
  assign n27246 = n27233 & ~n27245 ;
  assign n27247 = ~n27244 & ~n27245 ;
  assign n27248 = ~n27246 & ~n27247 ;
  assign n27249 = ~n26417 & ~n26421 ;
  assign n27250 = n27248 & n27249 ;
  assign n27251 = ~n27248 & ~n27249 ;
  assign n27252 = ~n27250 & ~n27251 ;
  assign n27253 = x104 & n4531 ;
  assign n27254 = x102 & n4847 ;
  assign n27255 = x103 & n4526 ;
  assign n27256 = ~n27254 & ~n27255 ;
  assign n27257 = ~n27253 & n27256 ;
  assign n27258 = n4534 & n11116 ;
  assign n27259 = n27257 & ~n27258 ;
  assign n27260 = x26 & ~n27259 ;
  assign n27261 = x26 & ~n27260 ;
  assign n27262 = ~n27259 & ~n27260 ;
  assign n27263 = ~n27261 & ~n27262 ;
  assign n27264 = n27252 & ~n27263 ;
  assign n27265 = n27252 & ~n27264 ;
  assign n27266 = ~n27263 & ~n27264 ;
  assign n27267 = ~n27265 & ~n27266 ;
  assign n27268 = ~n26435 & ~n26437 ;
  assign n27269 = ~n27267 & ~n27268 ;
  assign n27270 = ~n27267 & ~n27269 ;
  assign n27271 = ~n27268 & ~n27269 ;
  assign n27272 = ~n27270 & ~n27271 ;
  assign n27273 = x107 & n3589 ;
  assign n27274 = x105 & n3878 ;
  assign n27275 = x106 & n3584 ;
  assign n27276 = ~n27274 & ~n27275 ;
  assign n27277 = ~n27273 & n27276 ;
  assign n27278 = n3592 & n12749 ;
  assign n27279 = n27277 & ~n27278 ;
  assign n27280 = x23 & ~n27279 ;
  assign n27281 = x23 & ~n27280 ;
  assign n27282 = ~n27279 & ~n27280 ;
  assign n27283 = ~n27281 & ~n27282 ;
  assign n27284 = ~n27272 & n27283 ;
  assign n27285 = n27272 & ~n27283 ;
  assign n27286 = ~n27284 & ~n27285 ;
  assign n27287 = ~n27022 & ~n27286 ;
  assign n27288 = n27022 & n27286 ;
  assign n27289 = ~n27287 & ~n27288 ;
  assign n27290 = ~n27021 & n27289 ;
  assign n27291 = ~n27021 & ~n27290 ;
  assign n27292 = n27289 & ~n27290 ;
  assign n27293 = ~n27291 & ~n27292 ;
  assign n27294 = ~n27010 & ~n27293 ;
  assign n27295 = n27010 & ~n27292 ;
  assign n27296 = ~n27291 & n27295 ;
  assign n27297 = ~n27294 & ~n27296 ;
  assign n27298 = ~n27009 & n27297 ;
  assign n27299 = ~n27009 & ~n27298 ;
  assign n27300 = n27297 & ~n27298 ;
  assign n27301 = ~n27299 & ~n27300 ;
  assign n27302 = ~n26998 & ~n27301 ;
  assign n27303 = n26998 & ~n27300 ;
  assign n27304 = ~n27299 & n27303 ;
  assign n27305 = ~n27302 & ~n27304 ;
  assign n27306 = ~n26997 & n27305 ;
  assign n27307 = n26997 & ~n27305 ;
  assign n27308 = ~n27306 & ~n27307 ;
  assign n27309 = ~n26986 & n27308 ;
  assign n27310 = n26986 & ~n27308 ;
  assign n27311 = ~n27309 & ~n27310 ;
  assign n27312 = ~n26985 & n27311 ;
  assign n27313 = n26985 & ~n27311 ;
  assign n27314 = ~n27312 & ~n27313 ;
  assign n27315 = ~n26974 & n27314 ;
  assign n27316 = n26974 & ~n27314 ;
  assign n27317 = ~n27315 & ~n27316 ;
  assign n27318 = x122 & n574 ;
  assign n27319 = x120 & n673 ;
  assign n27320 = x121 & n569 ;
  assign n27321 = ~n27319 & ~n27320 ;
  assign n27322 = ~n27318 & n27321 ;
  assign n27323 = n577 & n22622 ;
  assign n27324 = n27322 & ~n27323 ;
  assign n27325 = x8 & ~n27324 ;
  assign n27326 = x8 & ~n27325 ;
  assign n27327 = ~n27324 & ~n27325 ;
  assign n27328 = ~n27326 & ~n27327 ;
  assign n27329 = n27317 & ~n27328 ;
  assign n27330 = n27317 & ~n27329 ;
  assign n27331 = ~n27328 & ~n27329 ;
  assign n27332 = ~n27330 & ~n27331 ;
  assign n27333 = x125 & n293 ;
  assign n27334 = x123 & n373 ;
  assign n27335 = x124 & n288 ;
  assign n27336 = ~n27334 & ~n27335 ;
  assign n27337 = ~n27333 & n27336 ;
  assign n27338 = n296 & n24935 ;
  assign n27339 = n27337 & ~n27338 ;
  assign n27340 = x5 & ~n27339 ;
  assign n27341 = x5 & ~n27340 ;
  assign n27342 = ~n27339 & ~n27340 ;
  assign n27343 = ~n27341 & ~n27342 ;
  assign n27344 = ~n27332 & n27343 ;
  assign n27345 = n27332 & ~n27343 ;
  assign n27346 = ~n27344 & ~n27345 ;
  assign n27347 = ~n26973 & ~n27346 ;
  assign n27348 = n26973 & n27346 ;
  assign n27349 = ~n27347 & ~n27348 ;
  assign n27350 = ~n26971 & n27349 ;
  assign n27351 = n26971 & ~n27349 ;
  assign n27352 = ~n27350 & ~n27351 ;
  assign n27353 = ~n26957 & n27352 ;
  assign n27354 = n26957 & ~n27352 ;
  assign n27355 = ~n27353 & ~n27354 ;
  assign n27356 = ~n26956 & n27355 ;
  assign n27357 = n26956 & ~n27355 ;
  assign n27358 = ~n27356 & ~n27357 ;
  assign n27763 = n27358 & x192 ;
  assign n27359 = ~n26944 & ~n26949 ;
  assign n27360 = ~n26922 & ~n26939 ;
  assign n27361 = ~x126 & n205 ;
  assign n27362 = ~x127 & n162 ;
  assign n27363 = ~n27361 & ~n27362 ;
  assign n27364 = x126 & ~n26930 ;
  assign n27365 = ~x127 & ~n27364 ;
  assign n27366 = ~x127 & ~n27365 ;
  assign n27367 = n26529 & ~n26929 ;
  assign n27368 = ~n27366 & ~n27367 ;
  assign n27369 = n167 & ~n27368 ;
  assign n27370 = n27363 & ~n27369 ;
  assign n27371 = ~x2 & ~n27370 ;
  assign n27372 = ~x2 & ~n27371 ;
  assign n27373 = ~n27370 & ~n27371 ;
  assign n27374 = ~n27372 & ~n27373 ;
  assign n27375 = ~n26905 & ~n26916 ;
  assign n27376 = ~n26902 & ~n27375 ;
  assign n27377 = ~n26883 & ~n26889 ;
  assign n27378 = ~x119 & n945 ;
  assign n27379 = ~x117 & n1099 ;
  assign n27380 = ~x118 & n940 ;
  assign n27381 = ~n27379 & ~n27380 ;
  assign n27382 = ~n27378 & n27381 ;
  assign n27383 = n948 & n20778 ;
  assign n27384 = n27382 & ~n27383 ;
  assign n27385 = ~x11 & ~n27384 ;
  assign n27386 = ~x11 & ~n27385 ;
  assign n27387 = ~n27384 & ~n27385 ;
  assign n27388 = ~n27386 & ~n27387 ;
  assign n27389 = ~n26866 & ~n26869 ;
  assign n27390 = ~x116 & n1434 ;
  assign n27391 = ~x114 & n1646 ;
  assign n27392 = ~x115 & n1429 ;
  assign n27393 = ~n27391 & ~n27392 ;
  assign n27394 = ~n27390 & n27393 ;
  assign n27395 = n1437 & n18678 ;
  assign n27396 = n27394 & ~n27395 ;
  assign n27397 = ~x14 & ~n27396 ;
  assign n27398 = ~x14 & ~n27397 ;
  assign n27399 = ~n27396 & ~n27397 ;
  assign n27400 = ~n27398 & ~n27399 ;
  assign n27401 = ~n26858 & ~n26862 ;
  assign n27402 = ~x113 & n2093 ;
  assign n27403 = ~x111 & n2275 ;
  assign n27404 = ~x112 & n2088 ;
  assign n27405 = ~n27403 & ~n27404 ;
  assign n27406 = ~n27402 & n27405 ;
  assign n27407 = n2096 & n16684 ;
  assign n27408 = n27406 & ~n27407 ;
  assign n27409 = ~x17 & ~n27408 ;
  assign n27410 = ~x17 & ~n27409 ;
  assign n27411 = ~n27408 & ~n27409 ;
  assign n27412 = ~n27410 & ~n27411 ;
  assign n27413 = ~n26850 & ~n26854 ;
  assign n27414 = ~x110 & n2751 ;
  assign n27415 = ~x108 & n3020 ;
  assign n27416 = ~x109 & n2746 ;
  assign n27417 = ~n27415 & ~n27416 ;
  assign n27418 = ~n27414 & n27417 ;
  assign n27419 = n2754 & n14802 ;
  assign n27420 = n27418 & ~n27419 ;
  assign n27421 = ~x20 & ~n27420 ;
  assign n27422 = ~x20 & ~n27421 ;
  assign n27423 = ~n27420 & ~n27421 ;
  assign n27424 = ~n27422 & ~n27423 ;
  assign n27425 = ~n26842 & ~n26846 ;
  assign n27426 = ~n26652 & ~n26654 ;
  assign n27427 = ~x63 & n26217 ;
  assign n27428 = ~x64 & n27427 ;
  assign n27429 = ~x65 & ~n26217 ;
  assign n27430 = ~n27428 & ~n27429 ;
  assign n27431 = ~x68 & n24612 ;
  assign n27432 = ~x66 & n25390 ;
  assign n27433 = ~x67 & n24607 ;
  assign n27434 = ~n27432 & ~n27433 ;
  assign n27435 = ~n27431 & n27434 ;
  assign n27436 = n352 & n24615 ;
  assign n27437 = n27435 & ~n27436 ;
  assign n27438 = ~x62 & ~n27437 ;
  assign n27439 = ~x62 & ~n27438 ;
  assign n27440 = ~n27437 & ~n27438 ;
  assign n27441 = ~n27439 & ~n27440 ;
  assign n27442 = ~n27430 & ~n27441 ;
  assign n27443 = ~n27430 & ~n27442 ;
  assign n27444 = ~n27441 & ~n27442 ;
  assign n27445 = ~n27443 & ~n27444 ;
  assign n27446 = ~n26621 & ~n26636 ;
  assign n27447 = n27445 & n27446 ;
  assign n27448 = ~n27445 & ~n27446 ;
  assign n27449 = ~n27447 & ~n27448 ;
  assign n27450 = ~x71 & n22325 ;
  assign n27451 = ~x69 & n23066 ;
  assign n27452 = ~x70 & n22320 ;
  assign n27453 = ~n27451 & ~n27452 ;
  assign n27454 = ~n27450 & n27453 ;
  assign n27455 = n622 & n22328 ;
  assign n27456 = n27454 & ~n27455 ;
  assign n27457 = ~x59 & ~n27456 ;
  assign n27458 = ~x59 & ~n27457 ;
  assign n27459 = ~n27456 & ~n27457 ;
  assign n27460 = ~n27458 & ~n27459 ;
  assign n27461 = ~n27449 & n27460 ;
  assign n27462 = n27449 & ~n27460 ;
  assign n27463 = ~n27461 & ~n27462 ;
  assign n27464 = ~n27426 & n27463 ;
  assign n27465 = n27426 & ~n27463 ;
  assign n27466 = ~n27464 & ~n27465 ;
  assign n27467 = ~x74 & n20143 ;
  assign n27468 = ~x72 & n20854 ;
  assign n27469 = ~x73 & n20138 ;
  assign n27470 = ~n27468 & ~n27469 ;
  assign n27471 = ~n27467 & n27470 ;
  assign n27472 = n1066 & n20146 ;
  assign n27473 = n27471 & ~n27472 ;
  assign n27474 = ~x56 & ~n27473 ;
  assign n27475 = ~x56 & ~n27474 ;
  assign n27476 = ~n27473 & ~n27474 ;
  assign n27477 = ~n27475 & ~n27476 ;
  assign n27478 = n27466 & ~n27477 ;
  assign n27479 = n27466 & ~n27478 ;
  assign n27480 = ~n27477 & ~n27478 ;
  assign n27481 = ~n27479 & ~n27480 ;
  assign n27482 = ~n26619 & ~n26671 ;
  assign n27483 = ~n26668 & ~n27482 ;
  assign n27484 = n27481 & n27483 ;
  assign n27485 = ~n27481 & ~n27483 ;
  assign n27486 = ~n27484 & ~n27485 ;
  assign n27487 = ~x77 & n18025 ;
  assign n27488 = ~x75 & n18764 ;
  assign n27489 = ~x76 & n18020 ;
  assign n27490 = ~n27488 & ~n27489 ;
  assign n27491 = ~n27487 & n27490 ;
  assign n27492 = n1594 & n18028 ;
  assign n27493 = n27491 & ~n27492 ;
  assign n27494 = ~x53 & ~n27493 ;
  assign n27495 = ~x53 & ~n27494 ;
  assign n27496 = ~n27493 & ~n27494 ;
  assign n27497 = ~n27495 & ~n27496 ;
  assign n27498 = ~n27486 & n27497 ;
  assign n27499 = n27486 & ~n27497 ;
  assign n27500 = ~n27498 & ~n27499 ;
  assign n27501 = ~n26687 & ~n26689 ;
  assign n27502 = n27500 & ~n27501 ;
  assign n27503 = ~n27500 & n27501 ;
  assign n27504 = ~n27502 & ~n27503 ;
  assign n27505 = ~x80 & n16076 ;
  assign n27506 = ~x78 & n16756 ;
  assign n27507 = ~x79 & n16071 ;
  assign n27508 = ~n27506 & ~n27507 ;
  assign n27509 = ~n27505 & n27508 ;
  assign n27510 = n2145 & n16079 ;
  assign n27511 = n27509 & ~n27510 ;
  assign n27512 = ~x50 & ~n27511 ;
  assign n27513 = ~x50 & ~n27512 ;
  assign n27514 = ~n27511 & ~n27512 ;
  assign n27515 = ~n27513 & ~n27514 ;
  assign n27516 = n27504 & ~n27515 ;
  assign n27517 = n27504 & ~n27516 ;
  assign n27518 = ~n27515 & ~n27516 ;
  assign n27519 = ~n27517 & ~n27518 ;
  assign n27520 = ~n26703 & ~n26709 ;
  assign n27521 = n27519 & n27520 ;
  assign n27522 = ~n27519 & ~n27520 ;
  assign n27523 = ~n27521 & ~n27522 ;
  assign n27524 = ~x83 & n14233 ;
  assign n27525 = ~x81 & n14876 ;
  assign n27526 = ~x82 & n14228 ;
  assign n27527 = ~n27525 & ~n27526 ;
  assign n27528 = ~n27524 & n27527 ;
  assign n27529 = n2972 & n14236 ;
  assign n27530 = n27528 & ~n27529 ;
  assign n27531 = ~x47 & ~n27530 ;
  assign n27532 = ~x47 & ~n27531 ;
  assign n27533 = ~n27530 & ~n27531 ;
  assign n27534 = ~n27532 & ~n27533 ;
  assign n27535 = ~n27523 & n27534 ;
  assign n27536 = n27523 & ~n27534 ;
  assign n27537 = ~n27535 & ~n27536 ;
  assign n27538 = ~n26723 & ~n26725 ;
  assign n27539 = n27537 & ~n27538 ;
  assign n27540 = ~n27537 & n27538 ;
  assign n27541 = ~n27539 & ~n27540 ;
  assign n27542 = ~x86 & n12506 ;
  assign n27543 = ~x84 & n13131 ;
  assign n27544 = ~x85 & n12501 ;
  assign n27545 = ~n27543 & ~n27544 ;
  assign n27546 = ~n27542 & n27545 ;
  assign n27547 = n3832 & n12509 ;
  assign n27548 = n27546 & ~n27547 ;
  assign n27549 = ~x44 & ~n27548 ;
  assign n27550 = ~x44 & ~n27549 ;
  assign n27551 = ~n27548 & ~n27549 ;
  assign n27552 = ~n27550 & ~n27551 ;
  assign n27553 = n27541 & ~n27552 ;
  assign n27554 = n27541 & ~n27553 ;
  assign n27555 = ~n27552 & ~n27553 ;
  assign n27556 = ~n27554 & ~n27555 ;
  assign n27557 = ~n26728 & ~n26731 ;
  assign n27558 = n27556 & n27557 ;
  assign n27559 = ~n27556 & ~n27557 ;
  assign n27560 = ~n27558 & ~n27559 ;
  assign n27561 = ~x89 & n10905 ;
  assign n27562 = ~x87 & n11466 ;
  assign n27563 = ~x88 & n10900 ;
  assign n27564 = ~n27562 & ~n27563 ;
  assign n27565 = ~n27561 & n27564 ;
  assign n27566 = n4664 & n10908 ;
  assign n27567 = n27565 & ~n27566 ;
  assign n27568 = ~x41 & ~n27567 ;
  assign n27569 = ~x41 & ~n27568 ;
  assign n27570 = ~n27567 & ~n27568 ;
  assign n27571 = ~n27569 & ~n27570 ;
  assign n27572 = n27560 & ~n27571 ;
  assign n27573 = n27560 & ~n27572 ;
  assign n27574 = ~n27571 & ~n27572 ;
  assign n27575 = ~n27573 & ~n27574 ;
  assign n27576 = ~n26745 & ~n26751 ;
  assign n27577 = n27575 & n27576 ;
  assign n27578 = ~n27575 & ~n27576 ;
  assign n27579 = ~n27577 & ~n27578 ;
  assign n27580 = ~x92 & n9433 ;
  assign n27581 = ~x90 & n9915 ;
  assign n27582 = ~x91 & n9428 ;
  assign n27583 = ~n27581 & ~n27582 ;
  assign n27584 = ~n27580 & n27583 ;
  assign n27585 = n5896 & n9436 ;
  assign n27586 = n27584 & ~n27585 ;
  assign n27587 = ~x38 & ~n27586 ;
  assign n27588 = ~x38 & ~n27587 ;
  assign n27589 = ~n27586 & ~n27587 ;
  assign n27590 = ~n27588 & ~n27589 ;
  assign n27591 = n27579 & ~n27590 ;
  assign n27592 = n27579 & ~n27591 ;
  assign n27593 = ~n27590 & ~n27591 ;
  assign n27594 = ~n27592 & ~n27593 ;
  assign n27595 = ~n26764 & ~n26770 ;
  assign n27596 = n27594 & n27595 ;
  assign n27597 = ~n27594 & ~n27595 ;
  assign n27598 = ~n27596 & ~n27597 ;
  assign n27599 = ~x95 & n8006 ;
  assign n27600 = ~x93 & n8474 ;
  assign n27601 = ~x94 & n8001 ;
  assign n27602 = ~n27600 & ~n27601 ;
  assign n27603 = ~n27599 & n27602 ;
  assign n27604 = n7100 & n8009 ;
  assign n27605 = n27603 & ~n27604 ;
  assign n27606 = ~x35 & ~n27605 ;
  assign n27607 = ~x35 & ~n27606 ;
  assign n27608 = ~n27605 & ~n27606 ;
  assign n27609 = ~n27607 & ~n27608 ;
  assign n27610 = ~n27598 & n27609 ;
  assign n27611 = n27598 & ~n27609 ;
  assign n27612 = ~n27610 & ~n27611 ;
  assign n27613 = ~n26784 & ~n26787 ;
  assign n27614 = n27612 & ~n27613 ;
  assign n27615 = ~n27612 & n27613 ;
  assign n27616 = ~n27614 & ~n27615 ;
  assign n27617 = ~x98 & n6725 ;
  assign n27618 = ~x96 & n7129 ;
  assign n27619 = ~x97 & n6720 ;
  assign n27620 = ~n27618 & ~n27619 ;
  assign n27621 = ~n27617 & n27620 ;
  assign n27622 = n6728 & n8426 ;
  assign n27623 = n27621 & ~n27622 ;
  assign n27624 = ~x32 & ~n27623 ;
  assign n27625 = ~x32 & ~n27624 ;
  assign n27626 = ~n27623 & ~n27624 ;
  assign n27627 = ~n27625 & ~n27626 ;
  assign n27628 = n27616 & ~n27627 ;
  assign n27629 = n27616 & ~n27628 ;
  assign n27630 = ~n27627 & ~n27628 ;
  assign n27631 = ~n27629 & ~n27630 ;
  assign n27632 = ~n25957 & ~n26804 ;
  assign n27633 = ~n26801 & ~n27632 ;
  assign n27634 = n27631 & n27633 ;
  assign n27635 = ~n27631 & ~n27633 ;
  assign n27636 = ~n27634 & ~n27635 ;
  assign n27637 = ~x101 & n5560 ;
  assign n27638 = ~x99 & n5943 ;
  assign n27639 = ~x100 & n5555 ;
  assign n27640 = ~n27638 & ~n27639 ;
  assign n27641 = ~n27637 & n27640 ;
  assign n27642 = n5563 & n9844 ;
  assign n27643 = n27641 & ~n27642 ;
  assign n27644 = ~x29 & ~n27643 ;
  assign n27645 = ~x29 & ~n27644 ;
  assign n27646 = ~n27643 & ~n27644 ;
  assign n27647 = ~n27645 & ~n27646 ;
  assign n27648 = n27636 & ~n27647 ;
  assign n27649 = n27636 & ~n27648 ;
  assign n27650 = ~n27647 & ~n27648 ;
  assign n27651 = ~n27649 & ~n27650 ;
  assign n27652 = ~n26819 & ~n26823 ;
  assign n27653 = n27651 & n27652 ;
  assign n27654 = ~n27651 & ~n27652 ;
  assign n27655 = ~n27653 & ~n27654 ;
  assign n27656 = ~x104 & n4531 ;
  assign n27657 = ~x102 & n4847 ;
  assign n27658 = ~x103 & n4526 ;
  assign n27659 = ~n27657 & ~n27658 ;
  assign n27660 = ~n27656 & n27659 ;
  assign n27661 = n4534 & n11380 ;
  assign n27662 = n27660 & ~n27661 ;
  assign n27663 = ~x26 & ~n27662 ;
  assign n27664 = ~x26 & ~n27663 ;
  assign n27665 = ~n27662 & ~n27663 ;
  assign n27666 = ~n27664 & ~n27665 ;
  assign n27667 = n27655 & ~n27666 ;
  assign n27668 = n27655 & ~n27667 ;
  assign n27669 = ~n27666 & ~n27667 ;
  assign n27670 = ~n27668 & ~n27669 ;
  assign n27671 = ~n26837 & ~n26839 ;
  assign n27672 = ~n27670 & ~n27671 ;
  assign n27673 = ~n27670 & ~n27672 ;
  assign n27674 = ~n27671 & ~n27672 ;
  assign n27675 = ~n27673 & ~n27674 ;
  assign n27676 = ~x107 & n3589 ;
  assign n27677 = ~x105 & n3878 ;
  assign n27678 = ~x106 & n3584 ;
  assign n27679 = ~n27677 & ~n27678 ;
  assign n27680 = ~n27676 & n27679 ;
  assign n27681 = n3592 & n13034 ;
  assign n27682 = n27680 & ~n27681 ;
  assign n27683 = ~x23 & ~n27682 ;
  assign n27684 = ~x23 & ~n27683 ;
  assign n27685 = ~n27682 & ~n27683 ;
  assign n27686 = ~n27684 & ~n27685 ;
  assign n27687 = ~n27675 & n27686 ;
  assign n27688 = n27675 & ~n27686 ;
  assign n27689 = ~n27687 & ~n27688 ;
  assign n27690 = ~n27425 & ~n27689 ;
  assign n27691 = n27425 & n27689 ;
  assign n27692 = ~n27690 & ~n27691 ;
  assign n27693 = ~n27424 & n27692 ;
  assign n27694 = ~n27424 & ~n27693 ;
  assign n27695 = n27692 & ~n27693 ;
  assign n27696 = ~n27694 & ~n27695 ;
  assign n27697 = ~n27413 & ~n27696 ;
  assign n27698 = n27413 & ~n27695 ;
  assign n27699 = ~n27694 & n27698 ;
  assign n27700 = ~n27697 & ~n27699 ;
  assign n27701 = ~n27412 & n27700 ;
  assign n27702 = ~n27412 & ~n27701 ;
  assign n27703 = n27700 & ~n27701 ;
  assign n27704 = ~n27702 & ~n27703 ;
  assign n27705 = ~n27401 & ~n27704 ;
  assign n27706 = n27401 & ~n27703 ;
  assign n27707 = ~n27702 & n27706 ;
  assign n27708 = ~n27705 & ~n27707 ;
  assign n27709 = ~n27400 & n27708 ;
  assign n27710 = n27400 & ~n27708 ;
  assign n27711 = ~n27709 & ~n27710 ;
  assign n27712 = ~n27389 & n27711 ;
  assign n27713 = n27389 & ~n27711 ;
  assign n27714 = ~n27712 & ~n27713 ;
  assign n27715 = ~n27388 & n27714 ;
  assign n27716 = n27388 & ~n27714 ;
  assign n27717 = ~n27715 & ~n27716 ;
  assign n27718 = ~n27377 & n27717 ;
  assign n27719 = n27377 & ~n27717 ;
  assign n27720 = ~n27718 & ~n27719 ;
  assign n27721 = ~x122 & n574 ;
  assign n27722 = ~x120 & n673 ;
  assign n27723 = ~x121 & n569 ;
  assign n27724 = ~n27722 & ~n27723 ;
  assign n27725 = ~n27721 & n27724 ;
  assign n27726 = n577 & n22998 ;
  assign n27727 = n27725 & ~n27726 ;
  assign n27728 = ~x8 & ~n27727 ;
  assign n27729 = ~x8 & ~n27728 ;
  assign n27730 = ~n27727 & ~n27728 ;
  assign n27731 = ~n27729 & ~n27730 ;
  assign n27732 = n27720 & ~n27731 ;
  assign n27733 = n27720 & ~n27732 ;
  assign n27734 = ~n27731 & ~n27732 ;
  assign n27735 = ~n27733 & ~n27734 ;
  assign n27736 = ~x125 & n293 ;
  assign n27737 = ~x123 & n373 ;
  assign n27738 = ~x124 & n288 ;
  assign n27739 = ~n27737 & ~n27738 ;
  assign n27740 = ~n27736 & n27739 ;
  assign n27741 = n296 & n25330 ;
  assign n27742 = n27740 & ~n27741 ;
  assign n27743 = ~x5 & ~n27742 ;
  assign n27744 = ~x5 & ~n27743 ;
  assign n27745 = ~n27742 & ~n27743 ;
  assign n27746 = ~n27744 & ~n27745 ;
  assign n27747 = ~n27735 & n27746 ;
  assign n27748 = n27735 & ~n27746 ;
  assign n27749 = ~n27747 & ~n27748 ;
  assign n27750 = ~n27376 & ~n27749 ;
  assign n27751 = n27376 & n27749 ;
  assign n27752 = ~n27750 & ~n27751 ;
  assign n27753 = ~n27374 & n27752 ;
  assign n27754 = n27374 & ~n27752 ;
  assign n27755 = ~n27753 & ~n27754 ;
  assign n27756 = ~n27360 & n27755 ;
  assign n27757 = n27360 & ~n27755 ;
  assign n27758 = ~n27756 & ~n27757 ;
  assign n27759 = ~n27359 & n27758 ;
  assign n27760 = n27359 & ~n27758 ;
  assign n27761 = ~n27759 & ~n27760 ;
  assign n27764 = ~n27761 & ~x192 ;
  assign n27765 = ~n27763 & ~n27764 ;
  assign n27766 = ~n27298 & ~n27302 ;
  assign n27767 = ~n27290 & ~n27294 ;
  assign n27768 = x111 & n2751 ;
  assign n27769 = x109 & n3020 ;
  assign n27770 = x110 & n2746 ;
  assign n27771 = ~n27769 & ~n27770 ;
  assign n27772 = ~n27768 & n27771 ;
  assign n27773 = n2754 & n15111 ;
  assign n27774 = n27772 & ~n27773 ;
  assign n27775 = x20 & ~n27774 ;
  assign n27776 = x20 & ~n27775 ;
  assign n27777 = ~n27774 & ~n27775 ;
  assign n27778 = ~n27776 & ~n27777 ;
  assign n27779 = ~n27264 & ~n27269 ;
  assign n27780 = ~n27208 & ~n27211 ;
  assign n27781 = ~n27150 & ~n27156 ;
  assign n27782 = ~n27133 & ~n27136 ;
  assign n27783 = ~n27113 & ~n27119 ;
  assign n27784 = ~n27096 & ~n27099 ;
  assign n27785 = ~n27075 & ~n27082 ;
  assign n27786 = ~n27059 & ~n27061 ;
  assign n27787 = x65 & n27024 ;
  assign n27788 = x66 & ~n26217 ;
  assign n27789 = ~n27787 & ~n27788 ;
  assign n27790 = x69 & n24612 ;
  assign n27791 = x67 & n25390 ;
  assign n27792 = x68 & n24607 ;
  assign n27793 = ~n27791 & ~n27792 ;
  assign n27794 = ~n27790 & n27793 ;
  assign n27795 = n398 & n24615 ;
  assign n27796 = n27794 & ~n27795 ;
  assign n27797 = x62 & ~n27796 ;
  assign n27798 = x62 & ~n27797 ;
  assign n27799 = ~n27796 & ~n27797 ;
  assign n27800 = ~n27798 & ~n27799 ;
  assign n27801 = ~n27789 & ~n27800 ;
  assign n27802 = ~n27789 & ~n27801 ;
  assign n27803 = ~n27800 & ~n27801 ;
  assign n27804 = ~n27802 & ~n27803 ;
  assign n27805 = ~n27039 & ~n27045 ;
  assign n27806 = n27804 & n27805 ;
  assign n27807 = ~n27804 & ~n27805 ;
  assign n27808 = ~n27806 & ~n27807 ;
  assign n27809 = x72 & n22325 ;
  assign n27810 = x70 & n23066 ;
  assign n27811 = x71 & n22320 ;
  assign n27812 = ~n27810 & ~n27811 ;
  assign n27813 = ~n27809 & n27812 ;
  assign n27814 = n717 & n22328 ;
  assign n27815 = n27813 & ~n27814 ;
  assign n27816 = x59 & ~n27815 ;
  assign n27817 = x59 & ~n27816 ;
  assign n27818 = ~n27815 & ~n27816 ;
  assign n27819 = ~n27817 & ~n27818 ;
  assign n27820 = n27808 & ~n27819 ;
  assign n27821 = ~n27808 & n27819 ;
  assign n27822 = ~n27786 & ~n27821 ;
  assign n27823 = ~n27820 & n27822 ;
  assign n27824 = ~n27786 & ~n27823 ;
  assign n27825 = ~n27820 & ~n27823 ;
  assign n27826 = ~n27821 & n27825 ;
  assign n27827 = ~n27824 & ~n27826 ;
  assign n27828 = x75 & n20143 ;
  assign n27829 = x73 & n20854 ;
  assign n27830 = x74 & n20138 ;
  assign n27831 = ~n27829 & ~n27830 ;
  assign n27832 = ~n27828 & n27831 ;
  assign n27833 = n1150 & n20146 ;
  assign n27834 = n27832 & ~n27833 ;
  assign n27835 = x56 & ~n27834 ;
  assign n27836 = x56 & ~n27835 ;
  assign n27837 = ~n27834 & ~n27835 ;
  assign n27838 = ~n27836 & ~n27837 ;
  assign n27839 = n27827 & n27838 ;
  assign n27840 = ~n27827 & ~n27838 ;
  assign n27841 = ~n27839 & ~n27840 ;
  assign n27842 = ~n27785 & n27841 ;
  assign n27843 = n27785 & ~n27841 ;
  assign n27844 = ~n27842 & ~n27843 ;
  assign n27845 = x78 & n18025 ;
  assign n27846 = x76 & n18764 ;
  assign n27847 = x77 & n18020 ;
  assign n27848 = ~n27846 & ~n27847 ;
  assign n27849 = ~n27845 & n27848 ;
  assign n27850 = n1624 & n18028 ;
  assign n27851 = n27849 & ~n27850 ;
  assign n27852 = x53 & ~n27851 ;
  assign n27853 = x53 & ~n27852 ;
  assign n27854 = ~n27851 & ~n27852 ;
  assign n27855 = ~n27853 & ~n27854 ;
  assign n27856 = n27844 & ~n27855 ;
  assign n27857 = n27844 & ~n27856 ;
  assign n27858 = ~n27855 & ~n27856 ;
  assign n27859 = ~n27857 & ~n27858 ;
  assign n27860 = ~n27784 & n27859 ;
  assign n27861 = n27784 & ~n27859 ;
  assign n27862 = ~n27860 & ~n27861 ;
  assign n27863 = x81 & n16076 ;
  assign n27864 = x79 & n16756 ;
  assign n27865 = x80 & n16071 ;
  assign n27866 = ~n27864 & ~n27865 ;
  assign n27867 = ~n27863 & n27866 ;
  assign n27868 = n2348 & n16079 ;
  assign n27869 = n27867 & ~n27868 ;
  assign n27870 = x50 & ~n27869 ;
  assign n27871 = x50 & ~n27870 ;
  assign n27872 = ~n27869 & ~n27870 ;
  assign n27873 = ~n27871 & ~n27872 ;
  assign n27874 = ~n27862 & ~n27873 ;
  assign n27875 = n27862 & n27873 ;
  assign n27876 = ~n27874 & ~n27875 ;
  assign n27877 = n27783 & ~n27876 ;
  assign n27878 = ~n27783 & n27876 ;
  assign n27879 = ~n27877 & ~n27878 ;
  assign n27880 = x84 & n14233 ;
  assign n27881 = x82 & n14876 ;
  assign n27882 = x83 & n14228 ;
  assign n27883 = ~n27881 & ~n27882 ;
  assign n27884 = ~n27880 & n27883 ;
  assign n27885 = n3114 & n14236 ;
  assign n27886 = n27884 & ~n27885 ;
  assign n27887 = x47 & ~n27886 ;
  assign n27888 = x47 & ~n27887 ;
  assign n27889 = ~n27886 & ~n27887 ;
  assign n27890 = ~n27888 & ~n27889 ;
  assign n27891 = n27879 & ~n27890 ;
  assign n27892 = n27879 & ~n27891 ;
  assign n27893 = ~n27890 & ~n27891 ;
  assign n27894 = ~n27892 & ~n27893 ;
  assign n27895 = ~n27782 & n27894 ;
  assign n27896 = n27782 & ~n27894 ;
  assign n27897 = ~n27895 & ~n27896 ;
  assign n27898 = x87 & n12506 ;
  assign n27899 = x85 & n13131 ;
  assign n27900 = x86 & n12501 ;
  assign n27901 = ~n27899 & ~n27900 ;
  assign n27902 = ~n27898 & n27901 ;
  assign n27903 = n3991 & n12509 ;
  assign n27904 = n27902 & ~n27903 ;
  assign n27905 = x44 & ~n27904 ;
  assign n27906 = x44 & ~n27905 ;
  assign n27907 = ~n27904 & ~n27905 ;
  assign n27908 = ~n27906 & ~n27907 ;
  assign n27909 = ~n27897 & ~n27908 ;
  assign n27910 = n27897 & n27908 ;
  assign n27911 = ~n27909 & ~n27910 ;
  assign n27912 = n27781 & ~n27911 ;
  assign n27913 = ~n27781 & n27911 ;
  assign n27914 = ~n27912 & ~n27913 ;
  assign n27915 = x90 & n10905 ;
  assign n27916 = x88 & n11466 ;
  assign n27917 = x89 & n10900 ;
  assign n27918 = ~n27916 & ~n27917 ;
  assign n27919 = ~n27915 & n27918 ;
  assign n27920 = n4986 & n10908 ;
  assign n27921 = n27919 & ~n27920 ;
  assign n27922 = x41 & ~n27921 ;
  assign n27923 = x41 & ~n27922 ;
  assign n27924 = ~n27921 & ~n27922 ;
  assign n27925 = ~n27923 & ~n27924 ;
  assign n27926 = n27914 & ~n27925 ;
  assign n27927 = n27914 & ~n27926 ;
  assign n27928 = ~n27925 & ~n27926 ;
  assign n27929 = ~n27927 & ~n27928 ;
  assign n27930 = ~n27169 & ~n27175 ;
  assign n27931 = n27929 & n27930 ;
  assign n27932 = ~n27929 & ~n27930 ;
  assign n27933 = ~n27931 & ~n27932 ;
  assign n27934 = x93 & n9433 ;
  assign n27935 = x91 & n9915 ;
  assign n27936 = x92 & n9428 ;
  assign n27937 = ~n27935 & ~n27936 ;
  assign n27938 = ~n27934 & n27937 ;
  assign n27939 = n6094 & n9436 ;
  assign n27940 = n27938 & ~n27939 ;
  assign n27941 = x38 & ~n27940 ;
  assign n27942 = x38 & ~n27941 ;
  assign n27943 = ~n27940 & ~n27941 ;
  assign n27944 = ~n27942 & ~n27943 ;
  assign n27945 = n27933 & ~n27944 ;
  assign n27946 = n27933 & ~n27945 ;
  assign n27947 = ~n27944 & ~n27945 ;
  assign n27948 = ~n27946 & ~n27947 ;
  assign n27949 = ~n27188 & ~n27194 ;
  assign n27950 = n27948 & n27949 ;
  assign n27951 = ~n27948 & ~n27949 ;
  assign n27952 = ~n27950 & ~n27951 ;
  assign n27953 = x96 & n8006 ;
  assign n27954 = x94 & n8474 ;
  assign n27955 = x95 & n8001 ;
  assign n27956 = ~n27954 & ~n27955 ;
  assign n27957 = ~n27953 & n27956 ;
  assign n27958 = n7321 & n8009 ;
  assign n27959 = n27957 & ~n27958 ;
  assign n27960 = x35 & ~n27959 ;
  assign n27961 = x35 & ~n27960 ;
  assign n27962 = ~n27959 & ~n27960 ;
  assign n27963 = ~n27961 & ~n27962 ;
  assign n27964 = n27952 & ~n27963 ;
  assign n27965 = ~n27952 & n27963 ;
  assign n27966 = ~n27780 & ~n27965 ;
  assign n27967 = ~n27964 & n27966 ;
  assign n27968 = ~n27780 & ~n27967 ;
  assign n27969 = ~n27964 & ~n27967 ;
  assign n27970 = ~n27965 & n27969 ;
  assign n27971 = ~n27968 & ~n27970 ;
  assign n27972 = x99 & n6725 ;
  assign n27973 = x97 & n7129 ;
  assign n27974 = x98 & n6720 ;
  assign n27975 = ~n27973 & ~n27974 ;
  assign n27976 = ~n27972 & n27975 ;
  assign n27977 = n6728 & n8660 ;
  assign n27978 = n27976 & ~n27977 ;
  assign n27979 = x32 & ~n27978 ;
  assign n27980 = x32 & ~n27979 ;
  assign n27981 = ~n27978 & ~n27979 ;
  assign n27982 = ~n27980 & ~n27981 ;
  assign n27983 = ~n27971 & ~n27982 ;
  assign n27984 = ~n27971 & ~n27983 ;
  assign n27985 = ~n27982 & ~n27983 ;
  assign n27986 = ~n27984 & ~n27985 ;
  assign n27987 = ~n27225 & ~n27232 ;
  assign n27988 = n27986 & n27987 ;
  assign n27989 = ~n27986 & ~n27987 ;
  assign n27990 = ~n27988 & ~n27989 ;
  assign n27991 = x102 & n5560 ;
  assign n27992 = x100 & n5943 ;
  assign n27993 = x101 & n5555 ;
  assign n27994 = ~n27992 & ~n27993 ;
  assign n27995 = ~n27991 & n27994 ;
  assign n27996 = n5563 & n10092 ;
  assign n27997 = n27995 & ~n27996 ;
  assign n27998 = x29 & ~n27997 ;
  assign n27999 = x29 & ~n27998 ;
  assign n28000 = ~n27997 & ~n27998 ;
  assign n28001 = ~n27999 & ~n28000 ;
  assign n28002 = n27990 & ~n28001 ;
  assign n28003 = n27990 & ~n28002 ;
  assign n28004 = ~n28001 & ~n28002 ;
  assign n28005 = ~n28003 & ~n28004 ;
  assign n28006 = ~n27245 & ~n27251 ;
  assign n28007 = n28005 & n28006 ;
  assign n28008 = ~n28005 & ~n28006 ;
  assign n28009 = ~n28007 & ~n28008 ;
  assign n28010 = x105 & n4531 ;
  assign n28011 = x103 & n4847 ;
  assign n28012 = x104 & n4526 ;
  assign n28013 = ~n28011 & ~n28012 ;
  assign n28014 = ~n28010 & n28013 ;
  assign n28015 = n4534 & n11648 ;
  assign n28016 = n28014 & ~n28015 ;
  assign n28017 = x26 & ~n28016 ;
  assign n28018 = x26 & ~n28017 ;
  assign n28019 = ~n28016 & ~n28017 ;
  assign n28020 = ~n28018 & ~n28019 ;
  assign n28021 = n28009 & ~n28020 ;
  assign n28022 = ~n28009 & n28020 ;
  assign n28023 = ~n27779 & ~n28022 ;
  assign n28024 = ~n28021 & n28023 ;
  assign n28025 = ~n27779 & ~n28024 ;
  assign n28026 = ~n28021 & ~n28024 ;
  assign n28027 = ~n28022 & n28026 ;
  assign n28028 = ~n28025 & ~n28027 ;
  assign n28029 = x108 & n3589 ;
  assign n28030 = x106 & n3878 ;
  assign n28031 = x107 & n3584 ;
  assign n28032 = ~n28030 & ~n28031 ;
  assign n28033 = ~n28029 & n28032 ;
  assign n28034 = n3592 & n13323 ;
  assign n28035 = n28033 & ~n28034 ;
  assign n28036 = x23 & ~n28035 ;
  assign n28037 = x23 & ~n28036 ;
  assign n28038 = ~n28035 & ~n28036 ;
  assign n28039 = ~n28037 & ~n28038 ;
  assign n28040 = ~n28028 & ~n28039 ;
  assign n28041 = ~n28028 & ~n28040 ;
  assign n28042 = ~n28039 & ~n28040 ;
  assign n28043 = ~n28041 & ~n28042 ;
  assign n28044 = ~n27272 & ~n27283 ;
  assign n28045 = ~n27287 & ~n28044 ;
  assign n28046 = ~n28043 & ~n28045 ;
  assign n28047 = n28043 & n28045 ;
  assign n28048 = ~n28046 & ~n28047 ;
  assign n28049 = ~n27778 & n28048 ;
  assign n28050 = ~n27778 & ~n28049 ;
  assign n28051 = n28048 & ~n28049 ;
  assign n28052 = ~n28050 & ~n28051 ;
  assign n28053 = ~n27767 & ~n28052 ;
  assign n28054 = ~n27767 & ~n28053 ;
  assign n28055 = ~n28052 & ~n28053 ;
  assign n28056 = ~n28054 & ~n28055 ;
  assign n28057 = x114 & n2093 ;
  assign n28058 = x112 & n2275 ;
  assign n28059 = x113 & n2088 ;
  assign n28060 = ~n28058 & ~n28059 ;
  assign n28061 = ~n28057 & n28060 ;
  assign n28062 = n2096 & n17012 ;
  assign n28063 = n28061 & ~n28062 ;
  assign n28064 = x17 & ~n28063 ;
  assign n28065 = x17 & ~n28064 ;
  assign n28066 = ~n28063 & ~n28064 ;
  assign n28067 = ~n28065 & ~n28066 ;
  assign n28068 = n28056 & n28067 ;
  assign n28069 = ~n28056 & ~n28067 ;
  assign n28070 = ~n28068 & ~n28069 ;
  assign n28071 = ~n27766 & n28070 ;
  assign n28072 = n27766 & ~n28070 ;
  assign n28073 = ~n28071 & ~n28072 ;
  assign n28074 = x117 & n1434 ;
  assign n28075 = x115 & n1646 ;
  assign n28076 = x116 & n1429 ;
  assign n28077 = ~n28075 & ~n28076 ;
  assign n28078 = ~n28074 & n28077 ;
  assign n28079 = n1437 & n19026 ;
  assign n28080 = n28078 & ~n28079 ;
  assign n28081 = x14 & ~n28080 ;
  assign n28082 = x14 & ~n28081 ;
  assign n28083 = ~n28080 & ~n28081 ;
  assign n28084 = ~n28082 & ~n28083 ;
  assign n28085 = n28073 & ~n28084 ;
  assign n28086 = n28073 & ~n28085 ;
  assign n28087 = ~n28084 & ~n28085 ;
  assign n28088 = ~n28086 & ~n28087 ;
  assign n28089 = ~n27306 & ~n27309 ;
  assign n28090 = n28088 & n28089 ;
  assign n28091 = ~n28088 & ~n28089 ;
  assign n28092 = ~n28090 & ~n28091 ;
  assign n28093 = x120 & n945 ;
  assign n28094 = x118 & n1099 ;
  assign n28095 = x119 & n940 ;
  assign n28096 = ~n28094 & ~n28095 ;
  assign n28097 = ~n28093 & n28096 ;
  assign n28098 = n948 & n21143 ;
  assign n28099 = n28097 & ~n28098 ;
  assign n28100 = x11 & ~n28099 ;
  assign n28101 = x11 & ~n28100 ;
  assign n28102 = ~n28099 & ~n28100 ;
  assign n28103 = ~n28101 & ~n28102 ;
  assign n28104 = ~n28092 & n28103 ;
  assign n28105 = n28092 & ~n28103 ;
  assign n28106 = ~n28104 & ~n28105 ;
  assign n28107 = x123 & n574 ;
  assign n28108 = x121 & n673 ;
  assign n28109 = x122 & n569 ;
  assign n28110 = ~n28108 & ~n28109 ;
  assign n28111 = ~n28107 & n28110 ;
  assign n28112 = n577 & n23382 ;
  assign n28113 = n28111 & ~n28112 ;
  assign n28114 = x8 & ~n28113 ;
  assign n28115 = x8 & ~n28114 ;
  assign n28116 = ~n28113 & ~n28114 ;
  assign n28117 = ~n28115 & ~n28116 ;
  assign n28118 = n28106 & ~n28117 ;
  assign n28119 = n28106 & ~n28118 ;
  assign n28120 = ~n28117 & ~n28118 ;
  assign n28121 = ~n28119 & ~n28120 ;
  assign n28122 = ~n27312 & ~n27315 ;
  assign n28123 = n28121 & n28122 ;
  assign n28124 = ~n28121 & ~n28122 ;
  assign n28125 = ~n28123 & ~n28124 ;
  assign n28126 = x126 & n293 ;
  assign n28127 = x124 & n373 ;
  assign n28128 = x125 & n288 ;
  assign n28129 = ~n28127 & ~n28128 ;
  assign n28130 = ~n28126 & n28129 ;
  assign n28131 = n296 & n25735 ;
  assign n28132 = n28130 & ~n28131 ;
  assign n28133 = x5 & ~n28132 ;
  assign n28134 = x5 & ~n28133 ;
  assign n28135 = ~n28132 & ~n28133 ;
  assign n28136 = ~n28134 & ~n28135 ;
  assign n28137 = n28125 & ~n28136 ;
  assign n28138 = n28125 & ~n28137 ;
  assign n28139 = ~n28136 & ~n28137 ;
  assign n28140 = ~n28138 & ~n28139 ;
  assign n28141 = ~n27332 & ~n27343 ;
  assign n28142 = ~n27329 & ~n28141 ;
  assign n28143 = n149 & n26962 ;
  assign n28144 = ~x2 & ~n28143 ;
  assign n28145 = x127 & n182 ;
  assign n28146 = ~n28143 & ~n28145 ;
  assign n28147 = x2 & ~n28146 ;
  assign n28148 = ~n28144 & ~n28147 ;
  assign n28149 = ~n28142 & n28148 ;
  assign n28150 = n28142 & ~n28148 ;
  assign n28151 = ~n28149 & ~n28150 ;
  assign n28152 = ~n28140 & n28151 ;
  assign n28153 = ~n28140 & ~n28152 ;
  assign n28154 = n28151 & ~n28152 ;
  assign n28155 = ~n28153 & ~n28154 ;
  assign n28156 = ~n27347 & ~n27350 ;
  assign n28157 = n28155 & n28156 ;
  assign n28158 = ~n28155 & ~n28156 ;
  assign n28159 = ~n28157 & ~n28158 ;
  assign n28160 = ~n27353 & ~n27356 ;
  assign n28161 = n28159 & ~n28160 ;
  assign n28162 = ~n28159 & n28160 ;
  assign n28163 = ~n28161 & ~n28162 ;
  assign n28563 = n28163 & x193 ;
  assign n28164 = ~n27701 & ~n27705 ;
  assign n28165 = ~n27693 & ~n27697 ;
  assign n28166 = ~x111 & n2751 ;
  assign n28167 = ~x109 & n3020 ;
  assign n28168 = ~x110 & n2746 ;
  assign n28169 = ~n28167 & ~n28168 ;
  assign n28170 = ~n28166 & n28169 ;
  assign n28171 = n2754 & n15411 ;
  assign n28172 = n28170 & ~n28171 ;
  assign n28173 = ~x20 & ~n28172 ;
  assign n28174 = ~x20 & ~n28173 ;
  assign n28175 = ~n28172 & ~n28173 ;
  assign n28176 = ~n28174 & ~n28175 ;
  assign n28177 = ~n27667 & ~n27672 ;
  assign n28178 = ~n27611 & ~n27614 ;
  assign n28179 = ~n27553 & ~n27559 ;
  assign n28180 = ~n27536 & ~n27539 ;
  assign n28181 = ~n27516 & ~n27522 ;
  assign n28182 = ~n27499 & ~n27502 ;
  assign n28183 = ~n27478 & ~n27485 ;
  assign n28184 = ~n27462 & ~n27464 ;
  assign n28185 = ~x65 & n27427 ;
  assign n28186 = ~x66 & ~n26217 ;
  assign n28187 = ~n28185 & ~n28186 ;
  assign n28188 = ~x69 & n24612 ;
  assign n28189 = ~x67 & n25390 ;
  assign n28190 = ~x68 & n24607 ;
  assign n28191 = ~n28189 & ~n28190 ;
  assign n28192 = ~n28188 & n28191 ;
  assign n28193 = n435 & n24615 ;
  assign n28194 = n28192 & ~n28193 ;
  assign n28195 = ~x62 & ~n28194 ;
  assign n28196 = ~x62 & ~n28195 ;
  assign n28197 = ~n28194 & ~n28195 ;
  assign n28198 = ~n28196 & ~n28197 ;
  assign n28199 = ~n28187 & ~n28198 ;
  assign n28200 = ~n28187 & ~n28199 ;
  assign n28201 = ~n28198 & ~n28199 ;
  assign n28202 = ~n28200 & ~n28201 ;
  assign n28203 = ~n27442 & ~n27448 ;
  assign n28204 = n28202 & n28203 ;
  assign n28205 = ~n28202 & ~n28203 ;
  assign n28206 = ~n28204 & ~n28205 ;
  assign n28207 = ~x72 & n22325 ;
  assign n28208 = ~x70 & n23066 ;
  assign n28209 = ~x71 & n22320 ;
  assign n28210 = ~n28208 & ~n28209 ;
  assign n28211 = ~n28207 & n28210 ;
  assign n28212 = n773 & n22328 ;
  assign n28213 = n28211 & ~n28212 ;
  assign n28214 = ~x59 & ~n28213 ;
  assign n28215 = ~x59 & ~n28214 ;
  assign n28216 = ~n28213 & ~n28214 ;
  assign n28217 = ~n28215 & ~n28216 ;
  assign n28218 = n28206 & ~n28217 ;
  assign n28219 = ~n28206 & n28217 ;
  assign n28220 = ~n28184 & ~n28219 ;
  assign n28221 = ~n28218 & n28220 ;
  assign n28222 = ~n28184 & ~n28221 ;
  assign n28223 = ~n28218 & ~n28221 ;
  assign n28224 = ~n28219 & n28223 ;
  assign n28225 = ~n28222 & ~n28224 ;
  assign n28226 = ~x75 & n20143 ;
  assign n28227 = ~x73 & n20854 ;
  assign n28228 = ~x74 & n20138 ;
  assign n28229 = ~n28227 & ~n28228 ;
  assign n28230 = ~n28226 & n28229 ;
  assign n28231 = n1225 & n20146 ;
  assign n28232 = n28230 & ~n28231 ;
  assign n28233 = ~x56 & ~n28232 ;
  assign n28234 = ~x56 & ~n28233 ;
  assign n28235 = ~n28232 & ~n28233 ;
  assign n28236 = ~n28234 & ~n28235 ;
  assign n28237 = n28225 & n28236 ;
  assign n28238 = ~n28225 & ~n28236 ;
  assign n28239 = ~n28237 & ~n28238 ;
  assign n28240 = ~n28183 & n28239 ;
  assign n28241 = n28183 & ~n28239 ;
  assign n28242 = ~n28240 & ~n28241 ;
  assign n28243 = ~x78 & n18025 ;
  assign n28244 = ~x76 & n18764 ;
  assign n28245 = ~x77 & n18020 ;
  assign n28246 = ~n28244 & ~n28245 ;
  assign n28247 = ~n28243 & n28246 ;
  assign n28248 = n1718 & n18028 ;
  assign n28249 = n28247 & ~n28248 ;
  assign n28250 = ~x53 & ~n28249 ;
  assign n28251 = ~x53 & ~n28250 ;
  assign n28252 = ~n28249 & ~n28250 ;
  assign n28253 = ~n28251 & ~n28252 ;
  assign n28254 = n28242 & ~n28253 ;
  assign n28255 = n28242 & ~n28254 ;
  assign n28256 = ~n28253 & ~n28254 ;
  assign n28257 = ~n28255 & ~n28256 ;
  assign n28258 = ~n28182 & n28257 ;
  assign n28259 = n28182 & ~n28257 ;
  assign n28260 = ~n28258 & ~n28259 ;
  assign n28261 = ~x81 & n16076 ;
  assign n28262 = ~x79 & n16756 ;
  assign n28263 = ~x80 & n16071 ;
  assign n28264 = ~n28262 & ~n28263 ;
  assign n28265 = ~n28261 & n28264 ;
  assign n28266 = n2460 & n16079 ;
  assign n28267 = n28265 & ~n28266 ;
  assign n28268 = ~x50 & ~n28267 ;
  assign n28269 = ~x50 & ~n28268 ;
  assign n28270 = ~n28267 & ~n28268 ;
  assign n28271 = ~n28269 & ~n28270 ;
  assign n28272 = ~n28260 & ~n28271 ;
  assign n28273 = n28260 & n28271 ;
  assign n28274 = ~n28272 & ~n28273 ;
  assign n28275 = n28181 & ~n28274 ;
  assign n28276 = ~n28181 & n28274 ;
  assign n28277 = ~n28275 & ~n28276 ;
  assign n28278 = ~x84 & n14233 ;
  assign n28279 = ~x82 & n14876 ;
  assign n28280 = ~x83 & n14228 ;
  assign n28281 = ~n28279 & ~n28280 ;
  assign n28282 = ~n28278 & n28281 ;
  assign n28283 = n3247 & n14236 ;
  assign n28284 = n28282 & ~n28283 ;
  assign n28285 = ~x47 & ~n28284 ;
  assign n28286 = ~x47 & ~n28285 ;
  assign n28287 = ~n28284 & ~n28285 ;
  assign n28288 = ~n28286 & ~n28287 ;
  assign n28289 = n28277 & ~n28288 ;
  assign n28290 = n28277 & ~n28289 ;
  assign n28291 = ~n28288 & ~n28289 ;
  assign n28292 = ~n28290 & ~n28291 ;
  assign n28293 = ~n28180 & n28292 ;
  assign n28294 = n28180 & ~n28292 ;
  assign n28295 = ~n28293 & ~n28294 ;
  assign n28296 = ~x87 & n12506 ;
  assign n28297 = ~x85 & n13131 ;
  assign n28298 = ~x86 & n12501 ;
  assign n28299 = ~n28297 & ~n28298 ;
  assign n28300 = ~n28296 & n28299 ;
  assign n28301 = n4143 & n12509 ;
  assign n28302 = n28300 & ~n28301 ;
  assign n28303 = ~x44 & ~n28302 ;
  assign n28304 = ~x44 & ~n28303 ;
  assign n28305 = ~n28302 & ~n28303 ;
  assign n28306 = ~n28304 & ~n28305 ;
  assign n28307 = ~n28295 & ~n28306 ;
  assign n28308 = n28295 & n28306 ;
  assign n28309 = ~n28307 & ~n28308 ;
  assign n28310 = n28179 & ~n28309 ;
  assign n28311 = ~n28179 & n28309 ;
  assign n28312 = ~n28310 & ~n28311 ;
  assign n28313 = ~x90 & n10905 ;
  assign n28314 = ~x88 & n11466 ;
  assign n28315 = ~x89 & n10900 ;
  assign n28316 = ~n28314 & ~n28315 ;
  assign n28317 = ~n28313 & n28316 ;
  assign n28318 = n5155 & n10908 ;
  assign n28319 = n28317 & ~n28318 ;
  assign n28320 = ~x41 & ~n28319 ;
  assign n28321 = ~x41 & ~n28320 ;
  assign n28322 = ~n28319 & ~n28320 ;
  assign n28323 = ~n28321 & ~n28322 ;
  assign n28324 = n28312 & ~n28323 ;
  assign n28325 = n28312 & ~n28324 ;
  assign n28326 = ~n28323 & ~n28324 ;
  assign n28327 = ~n28325 & ~n28326 ;
  assign n28328 = ~n27572 & ~n27578 ;
  assign n28329 = n28327 & n28328 ;
  assign n28330 = ~n28327 & ~n28328 ;
  assign n28331 = ~n28329 & ~n28330 ;
  assign n28332 = ~x93 & n9433 ;
  assign n28333 = ~x91 & n9915 ;
  assign n28334 = ~x92 & n9428 ;
  assign n28335 = ~n28333 & ~n28334 ;
  assign n28336 = ~n28332 & n28335 ;
  assign n28337 = n6285 & n9436 ;
  assign n28338 = n28336 & ~n28337 ;
  assign n28339 = ~x38 & ~n28338 ;
  assign n28340 = ~x38 & ~n28339 ;
  assign n28341 = ~n28338 & ~n28339 ;
  assign n28342 = ~n28340 & ~n28341 ;
  assign n28343 = n28331 & ~n28342 ;
  assign n28344 = n28331 & ~n28343 ;
  assign n28345 = ~n28342 & ~n28343 ;
  assign n28346 = ~n28344 & ~n28345 ;
  assign n28347 = ~n27591 & ~n27597 ;
  assign n28348 = n28346 & n28347 ;
  assign n28349 = ~n28346 & ~n28347 ;
  assign n28350 = ~n28348 & ~n28349 ;
  assign n28351 = ~x96 & n8006 ;
  assign n28352 = ~x94 & n8474 ;
  assign n28353 = ~x95 & n8001 ;
  assign n28354 = ~n28352 & ~n28353 ;
  assign n28355 = ~n28351 & n28354 ;
  assign n28356 = n7531 & n8009 ;
  assign n28357 = n28355 & ~n28356 ;
  assign n28358 = ~x35 & ~n28357 ;
  assign n28359 = ~x35 & ~n28358 ;
  assign n28360 = ~n28357 & ~n28358 ;
  assign n28361 = ~n28359 & ~n28360 ;
  assign n28362 = n28350 & ~n28361 ;
  assign n28363 = ~n28350 & n28361 ;
  assign n28364 = ~n28178 & ~n28363 ;
  assign n28365 = ~n28362 & n28364 ;
  assign n28366 = ~n28178 & ~n28365 ;
  assign n28367 = ~n28362 & ~n28365 ;
  assign n28368 = ~n28363 & n28367 ;
  assign n28369 = ~n28366 & ~n28368 ;
  assign n28370 = ~x99 & n6725 ;
  assign n28371 = ~x97 & n7129 ;
  assign n28372 = ~x98 & n6720 ;
  assign n28373 = ~n28371 & ~n28372 ;
  assign n28374 = ~n28370 & n28373 ;
  assign n28375 = n6728 & n8885 ;
  assign n28376 = n28374 & ~n28375 ;
  assign n28377 = ~x32 & ~n28376 ;
  assign n28378 = ~x32 & ~n28377 ;
  assign n28379 = ~n28376 & ~n28377 ;
  assign n28380 = ~n28378 & ~n28379 ;
  assign n28381 = ~n28369 & ~n28380 ;
  assign n28382 = ~n28369 & ~n28381 ;
  assign n28383 = ~n28380 & ~n28381 ;
  assign n28384 = ~n28382 & ~n28383 ;
  assign n28385 = ~n27628 & ~n27635 ;
  assign n28386 = n28384 & n28385 ;
  assign n28387 = ~n28384 & ~n28385 ;
  assign n28388 = ~n28386 & ~n28387 ;
  assign n28389 = ~x102 & n5560 ;
  assign n28390 = ~x100 & n5943 ;
  assign n28391 = ~x101 & n5555 ;
  assign n28392 = ~n28390 & ~n28391 ;
  assign n28393 = ~n28389 & n28392 ;
  assign n28394 = n5563 & n10333 ;
  assign n28395 = n28393 & ~n28394 ;
  assign n28396 = ~x29 & ~n28395 ;
  assign n28397 = ~x29 & ~n28396 ;
  assign n28398 = ~n28395 & ~n28396 ;
  assign n28399 = ~n28397 & ~n28398 ;
  assign n28400 = n28388 & ~n28399 ;
  assign n28401 = n28388 & ~n28400 ;
  assign n28402 = ~n28399 & ~n28400 ;
  assign n28403 = ~n28401 & ~n28402 ;
  assign n28404 = ~n27648 & ~n27654 ;
  assign n28405 = n28403 & n28404 ;
  assign n28406 = ~n28403 & ~n28404 ;
  assign n28407 = ~n28405 & ~n28406 ;
  assign n28408 = ~x105 & n4531 ;
  assign n28409 = ~x103 & n4847 ;
  assign n28410 = ~x104 & n4526 ;
  assign n28411 = ~n28409 & ~n28410 ;
  assign n28412 = ~n28408 & n28411 ;
  assign n28413 = n4534 & n11907 ;
  assign n28414 = n28412 & ~n28413 ;
  assign n28415 = ~x26 & ~n28414 ;
  assign n28416 = ~x26 & ~n28415 ;
  assign n28417 = ~n28414 & ~n28415 ;
  assign n28418 = ~n28416 & ~n28417 ;
  assign n28419 = n28407 & ~n28418 ;
  assign n28420 = ~n28407 & n28418 ;
  assign n28421 = ~n28177 & ~n28420 ;
  assign n28422 = ~n28419 & n28421 ;
  assign n28423 = ~n28177 & ~n28422 ;
  assign n28424 = ~n28419 & ~n28422 ;
  assign n28425 = ~n28420 & n28424 ;
  assign n28426 = ~n28423 & ~n28425 ;
  assign n28427 = ~x108 & n3589 ;
  assign n28428 = ~x106 & n3878 ;
  assign n28429 = ~x107 & n3584 ;
  assign n28430 = ~n28428 & ~n28429 ;
  assign n28431 = ~n28427 & n28430 ;
  assign n28432 = n3592 & n13601 ;
  assign n28433 = n28431 & ~n28432 ;
  assign n28434 = ~x23 & ~n28433 ;
  assign n28435 = ~x23 & ~n28434 ;
  assign n28436 = ~n28433 & ~n28434 ;
  assign n28437 = ~n28435 & ~n28436 ;
  assign n28438 = ~n28426 & ~n28437 ;
  assign n28439 = ~n28426 & ~n28438 ;
  assign n28440 = ~n28437 & ~n28438 ;
  assign n28441 = ~n28439 & ~n28440 ;
  assign n28442 = ~n27675 & ~n27686 ;
  assign n28443 = ~n27690 & ~n28442 ;
  assign n28444 = ~n28441 & ~n28443 ;
  assign n28445 = n28441 & n28443 ;
  assign n28446 = ~n28444 & ~n28445 ;
  assign n28447 = ~n28176 & n28446 ;
  assign n28448 = ~n28176 & ~n28447 ;
  assign n28449 = n28446 & ~n28447 ;
  assign n28450 = ~n28448 & ~n28449 ;
  assign n28451 = ~n28165 & ~n28450 ;
  assign n28452 = ~n28165 & ~n28451 ;
  assign n28453 = ~n28450 & ~n28451 ;
  assign n28454 = ~n28452 & ~n28453 ;
  assign n28455 = ~x114 & n2093 ;
  assign n28456 = ~x112 & n2275 ;
  assign n28457 = ~x113 & n2088 ;
  assign n28458 = ~n28456 & ~n28457 ;
  assign n28459 = ~n28455 & n28458 ;
  assign n28460 = n2096 & n17333 ;
  assign n28461 = n28459 & ~n28460 ;
  assign n28462 = ~x17 & ~n28461 ;
  assign n28463 = ~x17 & ~n28462 ;
  assign n28464 = ~n28461 & ~n28462 ;
  assign n28465 = ~n28463 & ~n28464 ;
  assign n28466 = n28454 & n28465 ;
  assign n28467 = ~n28454 & ~n28465 ;
  assign n28468 = ~n28466 & ~n28467 ;
  assign n28469 = ~n28164 & n28468 ;
  assign n28470 = n28164 & ~n28468 ;
  assign n28471 = ~n28469 & ~n28470 ;
  assign n28472 = ~x117 & n1434 ;
  assign n28473 = ~x115 & n1646 ;
  assign n28474 = ~x116 & n1429 ;
  assign n28475 = ~n28473 & ~n28474 ;
  assign n28476 = ~n28472 & n28475 ;
  assign n28477 = n1437 & n19365 ;
  assign n28478 = n28476 & ~n28477 ;
  assign n28479 = ~x14 & ~n28478 ;
  assign n28480 = ~x14 & ~n28479 ;
  assign n28481 = ~n28478 & ~n28479 ;
  assign n28482 = ~n28480 & ~n28481 ;
  assign n28483 = n28471 & ~n28482 ;
  assign n28484 = n28471 & ~n28483 ;
  assign n28485 = ~n28482 & ~n28483 ;
  assign n28486 = ~n28484 & ~n28485 ;
  assign n28487 = ~n27709 & ~n27712 ;
  assign n28488 = n28486 & n28487 ;
  assign n28489 = ~n28486 & ~n28487 ;
  assign n28490 = ~n28488 & ~n28489 ;
  assign n28491 = ~x120 & n945 ;
  assign n28492 = ~x118 & n1099 ;
  assign n28493 = ~x119 & n940 ;
  assign n28494 = ~n28492 & ~n28493 ;
  assign n28495 = ~n28491 & n28494 ;
  assign n28496 = n948 & n21501 ;
  assign n28497 = n28495 & ~n28496 ;
  assign n28498 = ~x11 & ~n28497 ;
  assign n28499 = ~x11 & ~n28498 ;
  assign n28500 = ~n28497 & ~n28498 ;
  assign n28501 = ~n28499 & ~n28500 ;
  assign n28502 = ~n28490 & n28501 ;
  assign n28503 = n28490 & ~n28501 ;
  assign n28504 = ~n28502 & ~n28503 ;
  assign n28505 = ~x123 & n574 ;
  assign n28506 = ~x121 & n673 ;
  assign n28507 = ~x122 & n569 ;
  assign n28508 = ~n28506 & ~n28507 ;
  assign n28509 = ~n28505 & n28508 ;
  assign n28510 = n577 & n23760 ;
  assign n28511 = n28509 & ~n28510 ;
  assign n28512 = ~x8 & ~n28511 ;
  assign n28513 = ~x8 & ~n28512 ;
  assign n28514 = ~n28511 & ~n28512 ;
  assign n28515 = ~n28513 & ~n28514 ;
  assign n28516 = n28504 & ~n28515 ;
  assign n28517 = n28504 & ~n28516 ;
  assign n28518 = ~n28515 & ~n28516 ;
  assign n28519 = ~n28517 & ~n28518 ;
  assign n28520 = ~n27715 & ~n27718 ;
  assign n28521 = n28519 & n28520 ;
  assign n28522 = ~n28519 & ~n28520 ;
  assign n28523 = ~n28521 & ~n28522 ;
  assign n28524 = ~x126 & n293 ;
  assign n28525 = ~x124 & n373 ;
  assign n28526 = ~x125 & n288 ;
  assign n28527 = ~n28525 & ~n28526 ;
  assign n28528 = ~n28524 & n28527 ;
  assign n28529 = n296 & n26128 ;
  assign n28530 = n28528 & ~n28529 ;
  assign n28531 = ~x5 & ~n28530 ;
  assign n28532 = ~x5 & ~n28531 ;
  assign n28533 = ~n28530 & ~n28531 ;
  assign n28534 = ~n28532 & ~n28533 ;
  assign n28535 = n28523 & ~n28534 ;
  assign n28536 = n28523 & ~n28535 ;
  assign n28537 = ~n28534 & ~n28535 ;
  assign n28538 = ~n28536 & ~n28537 ;
  assign n28539 = ~n27735 & ~n27746 ;
  assign n28540 = ~n27732 & ~n28539 ;
  assign n28541 = n167 & n27365 ;
  assign n28542 = x2 & ~n28541 ;
  assign n28543 = ~x127 & n205 ;
  assign n28544 = ~n28541 & ~n28543 ;
  assign n28545 = ~x2 & ~n28544 ;
  assign n28546 = ~n28542 & ~n28545 ;
  assign n28547 = ~n28540 & n28546 ;
  assign n28548 = n28540 & ~n28546 ;
  assign n28549 = ~n28547 & ~n28548 ;
  assign n28550 = ~n28538 & n28549 ;
  assign n28551 = ~n28538 & ~n28550 ;
  assign n28552 = n28549 & ~n28550 ;
  assign n28553 = ~n28551 & ~n28552 ;
  assign n28554 = ~n27750 & ~n27753 ;
  assign n28555 = n28553 & n28554 ;
  assign n28556 = ~n28553 & ~n28554 ;
  assign n28557 = ~n28555 & ~n28556 ;
  assign n28558 = ~n27756 & ~n27759 ;
  assign n28559 = n28557 & ~n28558 ;
  assign n28560 = ~n28557 & n28558 ;
  assign n28561 = ~n28559 & ~n28560 ;
  assign n28564 = ~n28561 & ~x193 ;
  assign n28565 = ~n28563 & ~n28564 ;
  assign n28566 = ~n28124 & ~n28137 ;
  assign n28567 = x127 & n293 ;
  assign n28568 = x125 & n373 ;
  assign n28569 = x126 & n288 ;
  assign n28570 = ~n28568 & ~n28569 ;
  assign n28571 = ~n28567 & n28570 ;
  assign n28572 = n296 & n26533 ;
  assign n28573 = n28571 & ~n28572 ;
  assign n28574 = x5 & ~n28573 ;
  assign n28575 = x5 & ~n28574 ;
  assign n28576 = ~n28573 & ~n28574 ;
  assign n28577 = ~n28575 & ~n28576 ;
  assign n28578 = ~n28566 & ~n28577 ;
  assign n28579 = ~n28566 & ~n28578 ;
  assign n28580 = ~n28577 & ~n28578 ;
  assign n28581 = ~n28579 & ~n28580 ;
  assign n28582 = x121 & n945 ;
  assign n28583 = x119 & n1099 ;
  assign n28584 = x120 & n940 ;
  assign n28585 = ~n28583 & ~n28584 ;
  assign n28586 = ~n28582 & n28585 ;
  assign n28587 = n948 & n21870 ;
  assign n28588 = n28586 & ~n28587 ;
  assign n28589 = x11 & ~n28588 ;
  assign n28590 = x11 & ~n28589 ;
  assign n28591 = ~n28588 & ~n28589 ;
  assign n28592 = ~n28590 & ~n28591 ;
  assign n28593 = ~n28085 & ~n28091 ;
  assign n28594 = n28592 & n28593 ;
  assign n28595 = ~n28592 & ~n28593 ;
  assign n28596 = ~n28594 & ~n28595 ;
  assign n28597 = x115 & n2093 ;
  assign n28598 = x113 & n2275 ;
  assign n28599 = x114 & n2088 ;
  assign n28600 = ~n28598 & ~n28599 ;
  assign n28601 = ~n28597 & n28600 ;
  assign n28602 = n2096 & n17364 ;
  assign n28603 = n28601 & ~n28602 ;
  assign n28604 = x17 & ~n28603 ;
  assign n28605 = x17 & ~n28604 ;
  assign n28606 = ~n28603 & ~n28604 ;
  assign n28607 = ~n28605 & ~n28606 ;
  assign n28608 = ~n28049 & ~n28053 ;
  assign n28609 = n28607 & n28608 ;
  assign n28610 = ~n28607 & ~n28608 ;
  assign n28611 = ~n28609 & ~n28610 ;
  assign n28612 = x112 & n2751 ;
  assign n28613 = x110 & n3020 ;
  assign n28614 = x111 & n2746 ;
  assign n28615 = ~n28613 & ~n28614 ;
  assign n28616 = ~n28612 & n28615 ;
  assign n28617 = n2754 & n15442 ;
  assign n28618 = n28616 & ~n28617 ;
  assign n28619 = x20 & ~n28618 ;
  assign n28620 = x20 & ~n28619 ;
  assign n28621 = ~n28618 & ~n28619 ;
  assign n28622 = ~n28620 & ~n28621 ;
  assign n28623 = ~n28040 & ~n28046 ;
  assign n28624 = n28622 & n28623 ;
  assign n28625 = ~n28622 & ~n28623 ;
  assign n28626 = ~n28624 & ~n28625 ;
  assign n28627 = x109 & n3589 ;
  assign n28628 = x107 & n3878 ;
  assign n28629 = x108 & n3584 ;
  assign n28630 = ~n28628 & ~n28629 ;
  assign n28631 = ~n28627 & n28630 ;
  assign n28632 = n3592 & n13894 ;
  assign n28633 = n28631 & ~n28632 ;
  assign n28634 = x23 & ~n28633 ;
  assign n28635 = x23 & ~n28634 ;
  assign n28636 = ~n28633 & ~n28634 ;
  assign n28637 = ~n28635 & ~n28636 ;
  assign n28638 = ~n28026 & n28637 ;
  assign n28639 = n28026 & ~n28637 ;
  assign n28640 = ~n28638 & ~n28639 ;
  assign n28641 = x106 & n4531 ;
  assign n28642 = x104 & n4847 ;
  assign n28643 = x105 & n4526 ;
  assign n28644 = ~n28642 & ~n28643 ;
  assign n28645 = ~n28641 & n28644 ;
  assign n28646 = n4534 & n12181 ;
  assign n28647 = n28645 & ~n28646 ;
  assign n28648 = x26 & ~n28647 ;
  assign n28649 = x26 & ~n28648 ;
  assign n28650 = ~n28647 & ~n28648 ;
  assign n28651 = ~n28649 & ~n28650 ;
  assign n28652 = ~n28002 & ~n28008 ;
  assign n28653 = n28651 & n28652 ;
  assign n28654 = ~n28651 & ~n28652 ;
  assign n28655 = ~n28653 & ~n28654 ;
  assign n28656 = ~n27983 & ~n27989 ;
  assign n28657 = x103 & n5560 ;
  assign n28658 = x101 & n5943 ;
  assign n28659 = x102 & n5555 ;
  assign n28660 = ~n28658 & ~n28659 ;
  assign n28661 = ~n28657 & n28660 ;
  assign n28662 = ~n5563 & n28661 ;
  assign n28663 = ~n10588 & n28661 ;
  assign n28664 = ~n28662 & ~n28663 ;
  assign n28665 = x29 & ~n28664 ;
  assign n28666 = ~x29 & n28664 ;
  assign n28667 = ~n28665 & ~n28666 ;
  assign n28668 = ~n28656 & ~n28667 ;
  assign n28669 = n28656 & n28667 ;
  assign n28670 = ~n28668 & ~n28669 ;
  assign n28671 = ~n27840 & ~n27842 ;
  assign n28672 = ~n27801 & ~n27807 ;
  assign n28673 = x66 & n27024 ;
  assign n28674 = x67 & ~n26217 ;
  assign n28675 = ~n28673 & ~n28674 ;
  assign n28676 = x2 & ~n28675 ;
  assign n28677 = ~x2 & n28675 ;
  assign n28678 = ~n28676 & ~n28677 ;
  assign n28679 = x70 & n24612 ;
  assign n28680 = x68 & n25390 ;
  assign n28681 = x69 & n24607 ;
  assign n28682 = ~n28680 & ~n28681 ;
  assign n28683 = ~n28679 & n28682 ;
  assign n28684 = ~n24615 & n28683 ;
  assign n28685 = ~n488 & n28683 ;
  assign n28686 = ~n28684 & ~n28685 ;
  assign n28687 = x62 & ~n28686 ;
  assign n28688 = ~x62 & n28686 ;
  assign n28689 = ~n28687 & ~n28688 ;
  assign n28690 = n28678 & ~n28689 ;
  assign n28691 = ~n28678 & n28689 ;
  assign n28692 = ~n28690 & ~n28691 ;
  assign n28693 = ~n28672 & n28692 ;
  assign n28694 = n28672 & ~n28692 ;
  assign n28695 = ~n28693 & ~n28694 ;
  assign n28696 = x73 & n22325 ;
  assign n28697 = x71 & n23066 ;
  assign n28698 = x72 & n22320 ;
  assign n28699 = ~n28697 & ~n28698 ;
  assign n28700 = ~n28696 & n28699 ;
  assign n28701 = n843 & n22328 ;
  assign n28702 = n28700 & ~n28701 ;
  assign n28703 = x59 & ~n28702 ;
  assign n28704 = x59 & ~n28703 ;
  assign n28705 = ~n28702 & ~n28703 ;
  assign n28706 = ~n28704 & ~n28705 ;
  assign n28707 = n28695 & ~n28706 ;
  assign n28708 = n28695 & ~n28707 ;
  assign n28709 = ~n28706 & ~n28707 ;
  assign n28710 = ~n28708 & ~n28709 ;
  assign n28711 = ~n27825 & n28710 ;
  assign n28712 = n27825 & ~n28710 ;
  assign n28713 = ~n28711 & ~n28712 ;
  assign n28714 = x76 & n20143 ;
  assign n28715 = x74 & n20854 ;
  assign n28716 = x75 & n20138 ;
  assign n28717 = ~n28715 & ~n28716 ;
  assign n28718 = ~n28714 & n28717 ;
  assign n28719 = n1311 & n20146 ;
  assign n28720 = n28718 & ~n28719 ;
  assign n28721 = x56 & ~n28720 ;
  assign n28722 = x56 & ~n28721 ;
  assign n28723 = ~n28720 & ~n28721 ;
  assign n28724 = ~n28722 & ~n28723 ;
  assign n28725 = n28713 & n28724 ;
  assign n28726 = ~n28713 & ~n28724 ;
  assign n28727 = ~n28725 & ~n28726 ;
  assign n28728 = ~n28671 & n28727 ;
  assign n28729 = n28671 & ~n28727 ;
  assign n28730 = ~n28728 & ~n28729 ;
  assign n28731 = x79 & n18025 ;
  assign n28732 = x77 & n18764 ;
  assign n28733 = x78 & n18020 ;
  assign n28734 = ~n28732 & ~n28733 ;
  assign n28735 = ~n28731 & n28734 ;
  assign n28736 = n1817 & n18028 ;
  assign n28737 = n28735 & ~n28736 ;
  assign n28738 = x53 & ~n28737 ;
  assign n28739 = x53 & ~n28738 ;
  assign n28740 = ~n28737 & ~n28738 ;
  assign n28741 = ~n28739 & ~n28740 ;
  assign n28742 = n28730 & ~n28741 ;
  assign n28743 = n28730 & ~n28742 ;
  assign n28744 = ~n28741 & ~n28742 ;
  assign n28745 = ~n28743 & ~n28744 ;
  assign n28746 = ~n27784 & ~n27859 ;
  assign n28747 = ~n27856 & ~n28746 ;
  assign n28748 = n28745 & n28747 ;
  assign n28749 = ~n28745 & ~n28747 ;
  assign n28750 = ~n28748 & ~n28749 ;
  assign n28751 = x82 & n16076 ;
  assign n28752 = x80 & n16756 ;
  assign n28753 = x81 & n16071 ;
  assign n28754 = ~n28752 & ~n28753 ;
  assign n28755 = ~n28751 & n28754 ;
  assign n28756 = n2584 & n16079 ;
  assign n28757 = n28755 & ~n28756 ;
  assign n28758 = x50 & ~n28757 ;
  assign n28759 = x50 & ~n28758 ;
  assign n28760 = ~n28757 & ~n28758 ;
  assign n28761 = ~n28759 & ~n28760 ;
  assign n28762 = n28750 & ~n28761 ;
  assign n28763 = n28750 & ~n28762 ;
  assign n28764 = ~n28761 & ~n28762 ;
  assign n28765 = ~n28763 & ~n28764 ;
  assign n28766 = ~n27874 & ~n27878 ;
  assign n28767 = n28765 & n28766 ;
  assign n28768 = ~n28765 & ~n28766 ;
  assign n28769 = ~n28767 & ~n28768 ;
  assign n28770 = x85 & n14233 ;
  assign n28771 = x83 & n14876 ;
  assign n28772 = x84 & n14228 ;
  assign n28773 = ~n28771 & ~n28772 ;
  assign n28774 = ~n28770 & n28773 ;
  assign n28775 = n3389 & n14236 ;
  assign n28776 = n28774 & ~n28775 ;
  assign n28777 = x47 & ~n28776 ;
  assign n28778 = x47 & ~n28777 ;
  assign n28779 = ~n28776 & ~n28777 ;
  assign n28780 = ~n28778 & ~n28779 ;
  assign n28781 = ~n28769 & n28780 ;
  assign n28782 = n28769 & ~n28780 ;
  assign n28783 = ~n28781 & ~n28782 ;
  assign n28784 = ~n27782 & ~n27894 ;
  assign n28785 = ~n27891 & ~n28784 ;
  assign n28786 = n28783 & ~n28785 ;
  assign n28787 = ~n28783 & n28785 ;
  assign n28788 = ~n28786 & ~n28787 ;
  assign n28789 = x88 & n12506 ;
  assign n28790 = x86 & n13131 ;
  assign n28791 = x87 & n12501 ;
  assign n28792 = ~n28790 & ~n28791 ;
  assign n28793 = ~n28789 & n28792 ;
  assign n28794 = n4305 & n12509 ;
  assign n28795 = n28793 & ~n28794 ;
  assign n28796 = x44 & ~n28795 ;
  assign n28797 = x44 & ~n28796 ;
  assign n28798 = ~n28795 & ~n28796 ;
  assign n28799 = ~n28797 & ~n28798 ;
  assign n28800 = n28788 & ~n28799 ;
  assign n28801 = n28788 & ~n28800 ;
  assign n28802 = ~n28799 & ~n28800 ;
  assign n28803 = ~n28801 & ~n28802 ;
  assign n28804 = ~n27909 & ~n27913 ;
  assign n28805 = n28803 & n28804 ;
  assign n28806 = ~n28803 & ~n28804 ;
  assign n28807 = ~n28805 & ~n28806 ;
  assign n28808 = x91 & n10905 ;
  assign n28809 = x89 & n11466 ;
  assign n28810 = x90 & n10900 ;
  assign n28811 = ~n28809 & ~n28810 ;
  assign n28812 = ~n28808 & n28811 ;
  assign n28813 = n5336 & n10908 ;
  assign n28814 = n28812 & ~n28813 ;
  assign n28815 = x41 & ~n28814 ;
  assign n28816 = x41 & ~n28815 ;
  assign n28817 = ~n28814 & ~n28815 ;
  assign n28818 = ~n28816 & ~n28817 ;
  assign n28819 = n28807 & ~n28818 ;
  assign n28820 = n28807 & ~n28819 ;
  assign n28821 = ~n28818 & ~n28819 ;
  assign n28822 = ~n28820 & ~n28821 ;
  assign n28823 = ~n27926 & ~n27932 ;
  assign n28824 = n28822 & n28823 ;
  assign n28825 = ~n28822 & ~n28823 ;
  assign n28826 = ~n28824 & ~n28825 ;
  assign n28827 = x94 & n9433 ;
  assign n28828 = x92 & n9915 ;
  assign n28829 = x93 & n9428 ;
  assign n28830 = ~n28828 & ~n28829 ;
  assign n28831 = ~n28827 & n28830 ;
  assign n28832 = n6483 & n9436 ;
  assign n28833 = n28831 & ~n28832 ;
  assign n28834 = x38 & ~n28833 ;
  assign n28835 = x38 & ~n28834 ;
  assign n28836 = ~n28833 & ~n28834 ;
  assign n28837 = ~n28835 & ~n28836 ;
  assign n28838 = ~n28826 & n28837 ;
  assign n28839 = n28826 & ~n28837 ;
  assign n28840 = ~n28838 & ~n28839 ;
  assign n28841 = ~n27945 & ~n27951 ;
  assign n28842 = n28840 & ~n28841 ;
  assign n28843 = ~n28840 & n28841 ;
  assign n28844 = ~n28842 & ~n28843 ;
  assign n28845 = x97 & n8006 ;
  assign n28846 = x95 & n8474 ;
  assign n28847 = x96 & n8001 ;
  assign n28848 = ~n28846 & ~n28847 ;
  assign n28849 = ~n28845 & n28848 ;
  assign n28850 = n7745 & n8009 ;
  assign n28851 = n28849 & ~n28850 ;
  assign n28852 = x35 & ~n28851 ;
  assign n28853 = x35 & ~n28852 ;
  assign n28854 = ~n28851 & ~n28852 ;
  assign n28855 = ~n28853 & ~n28854 ;
  assign n28856 = n28844 & ~n28855 ;
  assign n28857 = n28844 & ~n28856 ;
  assign n28858 = ~n28855 & ~n28856 ;
  assign n28859 = ~n28857 & ~n28858 ;
  assign n28860 = x100 & n6725 ;
  assign n28861 = x98 & n7129 ;
  assign n28862 = x99 & n6720 ;
  assign n28863 = ~n28861 & ~n28862 ;
  assign n28864 = ~n28860 & n28863 ;
  assign n28865 = ~n6728 & n28864 ;
  assign n28866 = ~n9115 & n28864 ;
  assign n28867 = ~n28865 & ~n28866 ;
  assign n28868 = x32 & ~n28867 ;
  assign n28869 = ~x32 & n28867 ;
  assign n28870 = ~n28868 & ~n28869 ;
  assign n28871 = ~n27969 & ~n28870 ;
  assign n28872 = ~n27969 & ~n28871 ;
  assign n28873 = ~n28870 & ~n28871 ;
  assign n28874 = ~n28872 & ~n28873 ;
  assign n28875 = ~n28859 & ~n28874 ;
  assign n28876 = ~n28859 & ~n28875 ;
  assign n28877 = ~n28874 & ~n28875 ;
  assign n28878 = ~n28876 & ~n28877 ;
  assign n28879 = n28670 & ~n28878 ;
  assign n28880 = n28670 & ~n28879 ;
  assign n28881 = ~n28878 & ~n28879 ;
  assign n28882 = ~n28880 & ~n28881 ;
  assign n28883 = n28655 & ~n28882 ;
  assign n28884 = ~n28655 & n28882 ;
  assign n28885 = ~n28640 & ~n28884 ;
  assign n28886 = ~n28883 & n28885 ;
  assign n28887 = ~n28640 & ~n28886 ;
  assign n28888 = ~n28884 & ~n28886 ;
  assign n28889 = ~n28883 & n28888 ;
  assign n28890 = ~n28887 & ~n28889 ;
  assign n28891 = n28626 & ~n28890 ;
  assign n28892 = ~n28626 & n28890 ;
  assign n28893 = n28611 & ~n28892 ;
  assign n28894 = ~n28891 & n28893 ;
  assign n28895 = n28611 & ~n28894 ;
  assign n28896 = ~n28892 & ~n28894 ;
  assign n28897 = ~n28891 & n28896 ;
  assign n28898 = ~n28895 & ~n28897 ;
  assign n28899 = ~n28069 & ~n28071 ;
  assign n28900 = x118 & n1434 ;
  assign n28901 = x116 & n1646 ;
  assign n28902 = x117 & n1429 ;
  assign n28903 = ~n28901 & ~n28902 ;
  assign n28904 = ~n28900 & n28903 ;
  assign n28905 = ~n1437 & n28904 ;
  assign n28906 = ~n19395 & n28904 ;
  assign n28907 = ~n28905 & ~n28906 ;
  assign n28908 = x14 & ~n28907 ;
  assign n28909 = ~x14 & n28907 ;
  assign n28910 = ~n28908 & ~n28909 ;
  assign n28911 = ~n28899 & ~n28910 ;
  assign n28912 = ~n28899 & ~n28911 ;
  assign n28913 = ~n28910 & ~n28911 ;
  assign n28914 = ~n28912 & ~n28913 ;
  assign n28915 = ~n28898 & ~n28914 ;
  assign n28916 = ~n28898 & ~n28915 ;
  assign n28917 = ~n28914 & ~n28915 ;
  assign n28918 = ~n28916 & ~n28917 ;
  assign n28919 = n28596 & ~n28918 ;
  assign n28920 = n28596 & ~n28919 ;
  assign n28921 = ~n28918 & ~n28919 ;
  assign n28922 = ~n28920 & ~n28921 ;
  assign n28923 = x124 & n574 ;
  assign n28924 = x122 & n673 ;
  assign n28925 = x123 & n569 ;
  assign n28926 = ~n28924 & ~n28925 ;
  assign n28927 = ~n28923 & n28926 ;
  assign n28928 = n577 & n23796 ;
  assign n28929 = n28927 & ~n28928 ;
  assign n28930 = x8 & ~n28929 ;
  assign n28931 = x8 & ~n28930 ;
  assign n28932 = ~n28929 & ~n28930 ;
  assign n28933 = ~n28931 & ~n28932 ;
  assign n28934 = ~n28105 & ~n28118 ;
  assign n28935 = ~n28933 & ~n28934 ;
  assign n28936 = ~n28933 & ~n28935 ;
  assign n28937 = ~n28934 & ~n28935 ;
  assign n28938 = ~n28936 & ~n28937 ;
  assign n28939 = ~n28922 & ~n28938 ;
  assign n28940 = ~n28922 & ~n28939 ;
  assign n28941 = ~n28938 & ~n28939 ;
  assign n28942 = ~n28940 & ~n28941 ;
  assign n28943 = ~n28581 & ~n28942 ;
  assign n28944 = ~n28581 & ~n28943 ;
  assign n28945 = ~n28942 & ~n28943 ;
  assign n28946 = ~n28944 & ~n28945 ;
  assign n28947 = ~n28149 & ~n28152 ;
  assign n28948 = n28946 & n28947 ;
  assign n28949 = ~n28946 & ~n28947 ;
  assign n28950 = ~n28948 & ~n28949 ;
  assign n28951 = ~n28158 & ~n28161 ;
  assign n28952 = n28950 & ~n28951 ;
  assign n28953 = ~n28950 & n28951 ;
  assign n28954 = ~n28952 & ~n28953 ;
  assign n29345 = n28954 & x194 ;
  assign n28955 = ~n28522 & ~n28535 ;
  assign n28956 = ~x127 & n293 ;
  assign n28957 = ~x125 & n373 ;
  assign n28958 = ~x126 & n288 ;
  assign n28959 = ~n28957 & ~n28958 ;
  assign n28960 = ~n28956 & n28959 ;
  assign n28961 = n296 & n26932 ;
  assign n28962 = n28960 & ~n28961 ;
  assign n28963 = ~x5 & ~n28962 ;
  assign n28964 = ~x5 & ~n28963 ;
  assign n28965 = ~n28962 & ~n28963 ;
  assign n28966 = ~n28964 & ~n28965 ;
  assign n28967 = ~n28955 & ~n28966 ;
  assign n28968 = ~n28955 & ~n28967 ;
  assign n28969 = ~n28966 & ~n28967 ;
  assign n28970 = ~n28968 & ~n28969 ;
  assign n28971 = ~x121 & n945 ;
  assign n28972 = ~x119 & n1099 ;
  assign n28973 = ~x120 & n940 ;
  assign n28974 = ~n28972 & ~n28973 ;
  assign n28975 = ~n28971 & n28974 ;
  assign n28976 = n948 & n22229 ;
  assign n28977 = n28975 & ~n28976 ;
  assign n28978 = ~x11 & ~n28977 ;
  assign n28979 = ~x11 & ~n28978 ;
  assign n28980 = ~n28977 & ~n28978 ;
  assign n28981 = ~n28979 & ~n28980 ;
  assign n28982 = ~n28483 & ~n28489 ;
  assign n28983 = n28981 & n28982 ;
  assign n28984 = ~n28981 & ~n28982 ;
  assign n28985 = ~n28983 & ~n28984 ;
  assign n28986 = ~x115 & n2093 ;
  assign n28987 = ~x113 & n2275 ;
  assign n28988 = ~x114 & n2088 ;
  assign n28989 = ~n28987 & ~n28988 ;
  assign n28990 = ~n28986 & n28989 ;
  assign n28991 = n2096 & n17683 ;
  assign n28992 = n28990 & ~n28991 ;
  assign n28993 = ~x17 & ~n28992 ;
  assign n28994 = ~x17 & ~n28993 ;
  assign n28995 = ~n28992 & ~n28993 ;
  assign n28996 = ~n28994 & ~n28995 ;
  assign n28997 = ~n28447 & ~n28451 ;
  assign n28998 = n28996 & n28997 ;
  assign n28999 = ~n28996 & ~n28997 ;
  assign n29000 = ~n28998 & ~n28999 ;
  assign n29001 = ~x112 & n2751 ;
  assign n29002 = ~x110 & n3020 ;
  assign n29003 = ~x111 & n2746 ;
  assign n29004 = ~n29002 & ~n29003 ;
  assign n29005 = ~n29001 & n29004 ;
  assign n29006 = n2754 & n15744 ;
  assign n29007 = n29005 & ~n29006 ;
  assign n29008 = ~x20 & ~n29007 ;
  assign n29009 = ~x20 & ~n29008 ;
  assign n29010 = ~n29007 & ~n29008 ;
  assign n29011 = ~n29009 & ~n29010 ;
  assign n29012 = ~n28438 & ~n28444 ;
  assign n29013 = n29011 & n29012 ;
  assign n29014 = ~n29011 & ~n29012 ;
  assign n29015 = ~n29013 & ~n29014 ;
  assign n29016 = ~x109 & n3589 ;
  assign n29017 = ~x107 & n3878 ;
  assign n29018 = ~x108 & n3584 ;
  assign n29019 = ~n29017 & ~n29018 ;
  assign n29020 = ~n29016 & n29019 ;
  assign n29021 = n3592 & n14177 ;
  assign n29022 = n29020 & ~n29021 ;
  assign n29023 = ~x23 & ~n29022 ;
  assign n29024 = ~x23 & ~n29023 ;
  assign n29025 = ~n29022 & ~n29023 ;
  assign n29026 = ~n29024 & ~n29025 ;
  assign n29027 = ~n28424 & n29026 ;
  assign n29028 = n28424 & ~n29026 ;
  assign n29029 = ~n29027 & ~n29028 ;
  assign n29030 = ~x106 & n4531 ;
  assign n29031 = ~x104 & n4847 ;
  assign n29032 = ~x105 & n4526 ;
  assign n29033 = ~n29031 & ~n29032 ;
  assign n29034 = ~n29030 & n29033 ;
  assign n29035 = n4534 & n12447 ;
  assign n29036 = n29034 & ~n29035 ;
  assign n29037 = ~x26 & ~n29036 ;
  assign n29038 = ~x26 & ~n29037 ;
  assign n29039 = ~n29036 & ~n29037 ;
  assign n29040 = ~n29038 & ~n29039 ;
  assign n29041 = ~n28400 & ~n28406 ;
  assign n29042 = n29040 & n29041 ;
  assign n29043 = ~n29040 & ~n29041 ;
  assign n29044 = ~n29042 & ~n29043 ;
  assign n29045 = ~n28381 & ~n28387 ;
  assign n29046 = ~x103 & n5560 ;
  assign n29047 = ~x101 & n5943 ;
  assign n29048 = ~x102 & n5555 ;
  assign n29049 = ~n29047 & ~n29048 ;
  assign n29050 = ~n29046 & n29049 ;
  assign n29051 = ~n5563 & n29050 ;
  assign n29052 = ~n10833 & n29050 ;
  assign n29053 = ~n29051 & ~n29052 ;
  assign n29054 = ~x29 & ~n29053 ;
  assign n29055 = x29 & n29053 ;
  assign n29056 = ~n29054 & ~n29055 ;
  assign n29057 = ~n29045 & ~n29056 ;
  assign n29058 = n29045 & n29056 ;
  assign n29059 = ~n29057 & ~n29058 ;
  assign n29060 = ~n28238 & ~n28240 ;
  assign n29061 = ~n28199 & ~n28205 ;
  assign n29062 = ~x66 & n27427 ;
  assign n29063 = ~x67 & ~n26217 ;
  assign n29064 = ~n29062 & ~n29063 ;
  assign n29065 = ~x2 & ~n29064 ;
  assign n29066 = x2 & n29064 ;
  assign n29067 = ~n29065 & ~n29066 ;
  assign n29068 = ~x70 & n24612 ;
  assign n29069 = ~x68 & n25390 ;
  assign n29070 = ~x69 & n24607 ;
  assign n29071 = ~n29069 & ~n29070 ;
  assign n29072 = ~n29068 & n29071 ;
  assign n29073 = ~n24615 & n29072 ;
  assign n29074 = ~n529 & n29072 ;
  assign n29075 = ~n29073 & ~n29074 ;
  assign n29076 = ~x62 & ~n29075 ;
  assign n29077 = x62 & n29075 ;
  assign n29078 = ~n29076 & ~n29077 ;
  assign n29079 = n29067 & ~n29078 ;
  assign n29080 = ~n29067 & n29078 ;
  assign n29081 = ~n29079 & ~n29080 ;
  assign n29082 = ~n29061 & n29081 ;
  assign n29083 = n29061 & ~n29081 ;
  assign n29084 = ~n29082 & ~n29083 ;
  assign n29085 = ~x73 & n22325 ;
  assign n29086 = ~x71 & n23066 ;
  assign n29087 = ~x72 & n22320 ;
  assign n29088 = ~n29086 & ~n29087 ;
  assign n29089 = ~n29085 & n29088 ;
  assign n29090 = n903 & n22328 ;
  assign n29091 = n29089 & ~n29090 ;
  assign n29092 = ~x59 & ~n29091 ;
  assign n29093 = ~x59 & ~n29092 ;
  assign n29094 = ~n29091 & ~n29092 ;
  assign n29095 = ~n29093 & ~n29094 ;
  assign n29096 = n29084 & ~n29095 ;
  assign n29097 = n29084 & ~n29096 ;
  assign n29098 = ~n29095 & ~n29096 ;
  assign n29099 = ~n29097 & ~n29098 ;
  assign n29100 = ~n28223 & n29099 ;
  assign n29101 = n28223 & ~n29099 ;
  assign n29102 = ~n29100 & ~n29101 ;
  assign n29103 = ~x76 & n20143 ;
  assign n29104 = ~x74 & n20854 ;
  assign n29105 = ~x75 & n20138 ;
  assign n29106 = ~n29104 & ~n29105 ;
  assign n29107 = ~n29103 & n29106 ;
  assign n29108 = n1390 & n20146 ;
  assign n29109 = n29107 & ~n29108 ;
  assign n29110 = ~x56 & ~n29109 ;
  assign n29111 = ~x56 & ~n29110 ;
  assign n29112 = ~n29109 & ~n29110 ;
  assign n29113 = ~n29111 & ~n29112 ;
  assign n29114 = n29102 & n29113 ;
  assign n29115 = ~n29102 & ~n29113 ;
  assign n29116 = ~n29114 & ~n29115 ;
  assign n29117 = ~n29060 & n29116 ;
  assign n29118 = n29060 & ~n29116 ;
  assign n29119 = ~n29117 & ~n29118 ;
  assign n29120 = ~x79 & n18025 ;
  assign n29121 = ~x77 & n18764 ;
  assign n29122 = ~x78 & n18020 ;
  assign n29123 = ~n29121 & ~n29122 ;
  assign n29124 = ~n29120 & n29123 ;
  assign n29125 = n1921 & n18028 ;
  assign n29126 = n29124 & ~n29125 ;
  assign n29127 = ~x53 & ~n29126 ;
  assign n29128 = ~x53 & ~n29127 ;
  assign n29129 = ~n29126 & ~n29127 ;
  assign n29130 = ~n29128 & ~n29129 ;
  assign n29131 = n29119 & ~n29130 ;
  assign n29132 = n29119 & ~n29131 ;
  assign n29133 = ~n29130 & ~n29131 ;
  assign n29134 = ~n29132 & ~n29133 ;
  assign n29135 = ~n28182 & ~n28257 ;
  assign n29136 = ~n28254 & ~n29135 ;
  assign n29137 = n29134 & n29136 ;
  assign n29138 = ~n29134 & ~n29136 ;
  assign n29139 = ~n29137 & ~n29138 ;
  assign n29140 = ~x82 & n16076 ;
  assign n29141 = ~x80 & n16756 ;
  assign n29142 = ~x81 & n16071 ;
  assign n29143 = ~n29141 & ~n29142 ;
  assign n29144 = ~n29140 & n29143 ;
  assign n29145 = n2697 & n16079 ;
  assign n29146 = n29144 & ~n29145 ;
  assign n29147 = ~x50 & ~n29146 ;
  assign n29148 = ~x50 & ~n29147 ;
  assign n29149 = ~n29146 & ~n29147 ;
  assign n29150 = ~n29148 & ~n29149 ;
  assign n29151 = n29139 & ~n29150 ;
  assign n29152 = n29139 & ~n29151 ;
  assign n29153 = ~n29150 & ~n29151 ;
  assign n29154 = ~n29152 & ~n29153 ;
  assign n29155 = ~n28272 & ~n28276 ;
  assign n29156 = n29154 & n29155 ;
  assign n29157 = ~n29154 & ~n29155 ;
  assign n29158 = ~n29156 & ~n29157 ;
  assign n29159 = ~x85 & n14233 ;
  assign n29160 = ~x83 & n14876 ;
  assign n29161 = ~x84 & n14228 ;
  assign n29162 = ~n29160 & ~n29161 ;
  assign n29163 = ~n29159 & n29162 ;
  assign n29164 = n3521 & n14236 ;
  assign n29165 = n29163 & ~n29164 ;
  assign n29166 = ~x47 & ~n29165 ;
  assign n29167 = ~x47 & ~n29166 ;
  assign n29168 = ~n29165 & ~n29166 ;
  assign n29169 = ~n29167 & ~n29168 ;
  assign n29170 = ~n29158 & n29169 ;
  assign n29171 = n29158 & ~n29169 ;
  assign n29172 = ~n29170 & ~n29171 ;
  assign n29173 = ~n28180 & ~n28292 ;
  assign n29174 = ~n28289 & ~n29173 ;
  assign n29175 = n29172 & ~n29174 ;
  assign n29176 = ~n29172 & n29174 ;
  assign n29177 = ~n29175 & ~n29176 ;
  assign n29178 = ~x88 & n12506 ;
  assign n29179 = ~x86 & n13131 ;
  assign n29180 = ~x87 & n12501 ;
  assign n29181 = ~n29179 & ~n29180 ;
  assign n29182 = ~n29178 & n29181 ;
  assign n29183 = n4457 & n12509 ;
  assign n29184 = n29182 & ~n29183 ;
  assign n29185 = ~x44 & ~n29184 ;
  assign n29186 = ~x44 & ~n29185 ;
  assign n29187 = ~n29184 & ~n29185 ;
  assign n29188 = ~n29186 & ~n29187 ;
  assign n29189 = n29177 & ~n29188 ;
  assign n29190 = n29177 & ~n29189 ;
  assign n29191 = ~n29188 & ~n29189 ;
  assign n29192 = ~n29190 & ~n29191 ;
  assign n29193 = ~n28307 & ~n28311 ;
  assign n29194 = n29192 & n29193 ;
  assign n29195 = ~n29192 & ~n29193 ;
  assign n29196 = ~n29194 & ~n29195 ;
  assign n29197 = ~x91 & n10905 ;
  assign n29198 = ~x89 & n11466 ;
  assign n29199 = ~x90 & n10900 ;
  assign n29200 = ~n29198 & ~n29199 ;
  assign n29201 = ~n29197 & n29200 ;
  assign n29202 = n5507 & n10908 ;
  assign n29203 = n29201 & ~n29202 ;
  assign n29204 = ~x41 & ~n29203 ;
  assign n29205 = ~x41 & ~n29204 ;
  assign n29206 = ~n29203 & ~n29204 ;
  assign n29207 = ~n29205 & ~n29206 ;
  assign n29208 = n29196 & ~n29207 ;
  assign n29209 = n29196 & ~n29208 ;
  assign n29210 = ~n29207 & ~n29208 ;
  assign n29211 = ~n29209 & ~n29210 ;
  assign n29212 = ~n28324 & ~n28330 ;
  assign n29213 = n29211 & n29212 ;
  assign n29214 = ~n29211 & ~n29212 ;
  assign n29215 = ~n29213 & ~n29214 ;
  assign n29216 = ~x94 & n9433 ;
  assign n29217 = ~x92 & n9915 ;
  assign n29218 = ~x93 & n9428 ;
  assign n29219 = ~n29217 & ~n29218 ;
  assign n29220 = ~n29216 & n29219 ;
  assign n29221 = n6671 & n9436 ;
  assign n29222 = n29220 & ~n29221 ;
  assign n29223 = ~x38 & ~n29222 ;
  assign n29224 = ~x38 & ~n29223 ;
  assign n29225 = ~n29222 & ~n29223 ;
  assign n29226 = ~n29224 & ~n29225 ;
  assign n29227 = ~n29215 & n29226 ;
  assign n29228 = n29215 & ~n29226 ;
  assign n29229 = ~n29227 & ~n29228 ;
  assign n29230 = ~n28343 & ~n28349 ;
  assign n29231 = n29229 & ~n29230 ;
  assign n29232 = ~n29229 & n29230 ;
  assign n29233 = ~n29231 & ~n29232 ;
  assign n29234 = ~x97 & n8006 ;
  assign n29235 = ~x95 & n8474 ;
  assign n29236 = ~x96 & n8001 ;
  assign n29237 = ~n29235 & ~n29236 ;
  assign n29238 = ~n29234 & n29237 ;
  assign n29239 = n7949 & n8009 ;
  assign n29240 = n29238 & ~n29239 ;
  assign n29241 = ~x35 & ~n29240 ;
  assign n29242 = ~x35 & ~n29241 ;
  assign n29243 = ~n29240 & ~n29241 ;
  assign n29244 = ~n29242 & ~n29243 ;
  assign n29245 = n29233 & ~n29244 ;
  assign n29246 = n29233 & ~n29245 ;
  assign n29247 = ~n29244 & ~n29245 ;
  assign n29248 = ~n29246 & ~n29247 ;
  assign n29249 = ~x100 & n6725 ;
  assign n29250 = ~x98 & n7129 ;
  assign n29251 = ~x99 & n6720 ;
  assign n29252 = ~n29250 & ~n29251 ;
  assign n29253 = ~n29249 & n29252 ;
  assign n29254 = ~n6728 & n29253 ;
  assign n29255 = ~n9338 & n29253 ;
  assign n29256 = ~n29254 & ~n29255 ;
  assign n29257 = ~x32 & ~n29256 ;
  assign n29258 = x32 & n29256 ;
  assign n29259 = ~n29257 & ~n29258 ;
  assign n29260 = ~n28367 & ~n29259 ;
  assign n29261 = ~n28367 & ~n29260 ;
  assign n29262 = ~n29259 & ~n29260 ;
  assign n29263 = ~n29261 & ~n29262 ;
  assign n29264 = ~n29248 & ~n29263 ;
  assign n29265 = ~n29248 & ~n29264 ;
  assign n29266 = ~n29263 & ~n29264 ;
  assign n29267 = ~n29265 & ~n29266 ;
  assign n29268 = n29059 & ~n29267 ;
  assign n29269 = n29059 & ~n29268 ;
  assign n29270 = ~n29267 & ~n29268 ;
  assign n29271 = ~n29269 & ~n29270 ;
  assign n29272 = n29044 & ~n29271 ;
  assign n29273 = ~n29044 & n29271 ;
  assign n29274 = ~n29029 & ~n29273 ;
  assign n29275 = ~n29272 & n29274 ;
  assign n29276 = ~n29029 & ~n29275 ;
  assign n29277 = ~n29273 & ~n29275 ;
  assign n29278 = ~n29272 & n29277 ;
  assign n29279 = ~n29276 & ~n29278 ;
  assign n29280 = n29015 & ~n29279 ;
  assign n29281 = ~n29015 & n29279 ;
  assign n29282 = n29000 & ~n29281 ;
  assign n29283 = ~n29280 & n29282 ;
  assign n29284 = n29000 & ~n29283 ;
  assign n29285 = ~n29281 & ~n29283 ;
  assign n29286 = ~n29280 & n29285 ;
  assign n29287 = ~n29284 & ~n29286 ;
  assign n29288 = ~n28467 & ~n28469 ;
  assign n29289 = ~x118 & n1434 ;
  assign n29290 = ~x116 & n1646 ;
  assign n29291 = ~x117 & n1429 ;
  assign n29292 = ~n29290 & ~n29291 ;
  assign n29293 = ~n29289 & n29292 ;
  assign n29294 = ~n1437 & n29293 ;
  assign n29295 = ~n19736 & n29293 ;
  assign n29296 = ~n29294 & ~n29295 ;
  assign n29297 = ~x14 & ~n29296 ;
  assign n29298 = x14 & n29296 ;
  assign n29299 = ~n29297 & ~n29298 ;
  assign n29300 = ~n29288 & ~n29299 ;
  assign n29301 = ~n29288 & ~n29300 ;
  assign n29302 = ~n29299 & ~n29300 ;
  assign n29303 = ~n29301 & ~n29302 ;
  assign n29304 = ~n29287 & ~n29303 ;
  assign n29305 = ~n29287 & ~n29304 ;
  assign n29306 = ~n29303 & ~n29304 ;
  assign n29307 = ~n29305 & ~n29306 ;
  assign n29308 = n28985 & ~n29307 ;
  assign n29309 = n28985 & ~n29308 ;
  assign n29310 = ~n29307 & ~n29308 ;
  assign n29311 = ~n29309 & ~n29310 ;
  assign n29312 = ~x124 & n574 ;
  assign n29313 = ~x122 & n673 ;
  assign n29314 = ~x123 & n569 ;
  assign n29315 = ~n29313 & ~n29314 ;
  assign n29316 = ~n29312 & n29315 ;
  assign n29317 = n577 & n24176 ;
  assign n29318 = n29316 & ~n29317 ;
  assign n29319 = ~x8 & ~n29318 ;
  assign n29320 = ~x8 & ~n29319 ;
  assign n29321 = ~n29318 & ~n29319 ;
  assign n29322 = ~n29320 & ~n29321 ;
  assign n29323 = ~n28503 & ~n28516 ;
  assign n29324 = ~n29322 & ~n29323 ;
  assign n29325 = ~n29322 & ~n29324 ;
  assign n29326 = ~n29323 & ~n29324 ;
  assign n29327 = ~n29325 & ~n29326 ;
  assign n29328 = ~n29311 & ~n29327 ;
  assign n29329 = ~n29311 & ~n29328 ;
  assign n29330 = ~n29327 & ~n29328 ;
  assign n29331 = ~n29329 & ~n29330 ;
  assign n29332 = ~n28970 & ~n29331 ;
  assign n29333 = ~n28970 & ~n29332 ;
  assign n29334 = ~n29331 & ~n29332 ;
  assign n29335 = ~n29333 & ~n29334 ;
  assign n29336 = ~n28547 & ~n28550 ;
  assign n29337 = n29335 & n29336 ;
  assign n29338 = ~n29335 & ~n29336 ;
  assign n29339 = ~n29337 & ~n29338 ;
  assign n29340 = ~n28556 & ~n28559 ;
  assign n29341 = n29339 & ~n29340 ;
  assign n29342 = ~n29339 & n29340 ;
  assign n29343 = ~n29341 & ~n29342 ;
  assign n29346 = ~n29343 & ~x194 ;
  assign n29347 = ~n29345 & ~n29346 ;
  assign n29348 = ~n28949 & ~n28952 ;
  assign n29349 = ~n28578 & ~n28943 ;
  assign n29350 = x119 & n1434 ;
  assign n29351 = x117 & n1646 ;
  assign n29352 = x118 & n1429 ;
  assign n29353 = ~n29351 & ~n29352 ;
  assign n29354 = ~n29350 & n29353 ;
  assign n29355 = n1437 & n20423 ;
  assign n29356 = n29354 & ~n29355 ;
  assign n29357 = x14 & ~n29356 ;
  assign n29358 = x14 & ~n29357 ;
  assign n29359 = ~n29356 & ~n29357 ;
  assign n29360 = ~n29358 & ~n29359 ;
  assign n29361 = ~n28610 & ~n28894 ;
  assign n29362 = n29360 & n29361 ;
  assign n29363 = ~n29360 & ~n29361 ;
  assign n29364 = ~n29362 & ~n29363 ;
  assign n29365 = x113 & n2751 ;
  assign n29366 = x111 & n3020 ;
  assign n29367 = x112 & n2746 ;
  assign n29368 = ~n29366 & ~n29367 ;
  assign n29369 = ~n29365 & n29368 ;
  assign n29370 = n2754 & n16361 ;
  assign n29371 = n29369 & ~n29370 ;
  assign n29372 = x20 & ~n29371 ;
  assign n29373 = x20 & ~n29372 ;
  assign n29374 = ~n29371 & ~n29372 ;
  assign n29375 = ~n29373 & ~n29374 ;
  assign n29376 = ~n28026 & ~n28637 ;
  assign n29377 = ~n28886 & ~n29376 ;
  assign n29378 = n29375 & n29377 ;
  assign n29379 = ~n29375 & ~n29377 ;
  assign n29380 = ~n29378 & ~n29379 ;
  assign n29381 = x107 & n4531 ;
  assign n29382 = x105 & n4847 ;
  assign n29383 = x106 & n4526 ;
  assign n29384 = ~n29382 & ~n29383 ;
  assign n29385 = ~n29381 & n29384 ;
  assign n29386 = n4534 & n12749 ;
  assign n29387 = n29385 & ~n29386 ;
  assign n29388 = x26 & ~n29387 ;
  assign n29389 = x26 & ~n29388 ;
  assign n29390 = ~n29387 & ~n29388 ;
  assign n29391 = ~n29389 & ~n29390 ;
  assign n29392 = ~n28668 & ~n28879 ;
  assign n29393 = n29391 & n29392 ;
  assign n29394 = ~n29391 & ~n29392 ;
  assign n29395 = ~n29393 & ~n29394 ;
  assign n29396 = ~n28842 & ~n28856 ;
  assign n29397 = x101 & n6725 ;
  assign n29398 = x99 & n7129 ;
  assign n29399 = x100 & n6720 ;
  assign n29400 = ~n29398 & ~n29399 ;
  assign n29401 = ~n29397 & n29400 ;
  assign n29402 = ~n6728 & n29401 ;
  assign n29403 = ~n9601 & n29401 ;
  assign n29404 = ~n29402 & ~n29403 ;
  assign n29405 = x32 & ~n29404 ;
  assign n29406 = ~x32 & n29404 ;
  assign n29407 = ~n29405 & ~n29406 ;
  assign n29408 = ~n29396 & ~n29407 ;
  assign n29409 = n29396 & n29407 ;
  assign n29410 = ~n29408 & ~n29409 ;
  assign n29411 = x98 & n8006 ;
  assign n29412 = x96 & n8474 ;
  assign n29413 = x97 & n8001 ;
  assign n29414 = ~n29412 & ~n29413 ;
  assign n29415 = ~n29411 & n29414 ;
  assign n29416 = n8009 & n8196 ;
  assign n29417 = n29415 & ~n29416 ;
  assign n29418 = x35 & ~n29417 ;
  assign n29419 = x35 & ~n29418 ;
  assign n29420 = ~n29417 & ~n29418 ;
  assign n29421 = ~n29419 & ~n29420 ;
  assign n29422 = ~n28825 & ~n28839 ;
  assign n29423 = x71 & n24612 ;
  assign n29424 = x69 & n25390 ;
  assign n29425 = x70 & n24607 ;
  assign n29426 = ~n29424 & ~n29425 ;
  assign n29427 = ~n29423 & n29426 ;
  assign n29428 = n558 & n24615 ;
  assign n29429 = n29427 & ~n29428 ;
  assign n29430 = x62 & ~n29429 ;
  assign n29431 = x62 & ~n29430 ;
  assign n29432 = ~n29429 & ~n29430 ;
  assign n29433 = ~n29431 & ~n29432 ;
  assign n29434 = x67 & n27024 ;
  assign n29435 = x68 & ~n26217 ;
  assign n29436 = ~n29434 & ~n29435 ;
  assign n29437 = x2 & ~n29436 ;
  assign n29438 = x2 & ~n29437 ;
  assign n29439 = ~n29436 & ~n29437 ;
  assign n29440 = ~n29438 & ~n29439 ;
  assign n29441 = ~n29433 & ~n29440 ;
  assign n29442 = ~n29433 & ~n29441 ;
  assign n29443 = ~n29440 & ~n29441 ;
  assign n29444 = ~n29442 & ~n29443 ;
  assign n29445 = ~n28676 & ~n28690 ;
  assign n29446 = n29444 & n29445 ;
  assign n29447 = ~n29444 & ~n29445 ;
  assign n29448 = ~n29446 & ~n29447 ;
  assign n29449 = x74 & n22325 ;
  assign n29450 = x72 & n23066 ;
  assign n29451 = x73 & n22320 ;
  assign n29452 = ~n29450 & ~n29451 ;
  assign n29453 = ~n29449 & n29452 ;
  assign n29454 = n994 & n22328 ;
  assign n29455 = n29453 & ~n29454 ;
  assign n29456 = x59 & ~n29455 ;
  assign n29457 = x59 & ~n29456 ;
  assign n29458 = ~n29455 & ~n29456 ;
  assign n29459 = ~n29457 & ~n29458 ;
  assign n29460 = n29448 & ~n29459 ;
  assign n29461 = n29448 & ~n29460 ;
  assign n29462 = ~n29459 & ~n29460 ;
  assign n29463 = ~n29461 & ~n29462 ;
  assign n29464 = ~n28693 & ~n28707 ;
  assign n29465 = n29463 & n29464 ;
  assign n29466 = ~n29463 & ~n29464 ;
  assign n29467 = ~n29465 & ~n29466 ;
  assign n29468 = x77 & n20143 ;
  assign n29469 = x75 & n20854 ;
  assign n29470 = x76 & n20138 ;
  assign n29471 = ~n29469 & ~n29470 ;
  assign n29472 = ~n29468 & n29471 ;
  assign n29473 = n1502 & n20146 ;
  assign n29474 = n29472 & ~n29473 ;
  assign n29475 = x56 & ~n29474 ;
  assign n29476 = x56 & ~n29475 ;
  assign n29477 = ~n29474 & ~n29475 ;
  assign n29478 = ~n29476 & ~n29477 ;
  assign n29479 = ~n29467 & n29478 ;
  assign n29480 = n29467 & ~n29478 ;
  assign n29481 = ~n29479 & ~n29480 ;
  assign n29482 = ~n27825 & ~n28710 ;
  assign n29483 = ~n28726 & ~n29482 ;
  assign n29484 = n29481 & ~n29483 ;
  assign n29485 = ~n29481 & n29483 ;
  assign n29486 = ~n29484 & ~n29485 ;
  assign n29487 = x80 & n18025 ;
  assign n29488 = x78 & n18764 ;
  assign n29489 = x79 & n18020 ;
  assign n29490 = ~n29488 & ~n29489 ;
  assign n29491 = ~n29487 & n29490 ;
  assign n29492 = n2028 & n18028 ;
  assign n29493 = n29491 & ~n29492 ;
  assign n29494 = x53 & ~n29493 ;
  assign n29495 = x53 & ~n29494 ;
  assign n29496 = ~n29493 & ~n29494 ;
  assign n29497 = ~n29495 & ~n29496 ;
  assign n29498 = n29486 & ~n29497 ;
  assign n29499 = n29486 & ~n29498 ;
  assign n29500 = ~n29497 & ~n29498 ;
  assign n29501 = ~n29499 & ~n29500 ;
  assign n29502 = ~n28728 & ~n28742 ;
  assign n29503 = n29501 & n29502 ;
  assign n29504 = ~n29501 & ~n29502 ;
  assign n29505 = ~n29503 & ~n29504 ;
  assign n29506 = x83 & n16076 ;
  assign n29507 = x81 & n16756 ;
  assign n29508 = x82 & n16071 ;
  assign n29509 = ~n29507 & ~n29508 ;
  assign n29510 = ~n29506 & n29509 ;
  assign n29511 = n2843 & n16079 ;
  assign n29512 = n29510 & ~n29511 ;
  assign n29513 = x50 & ~n29512 ;
  assign n29514 = x50 & ~n29513 ;
  assign n29515 = ~n29512 & ~n29513 ;
  assign n29516 = ~n29514 & ~n29515 ;
  assign n29517 = n29505 & ~n29516 ;
  assign n29518 = n29505 & ~n29517 ;
  assign n29519 = ~n29516 & ~n29517 ;
  assign n29520 = ~n29518 & ~n29519 ;
  assign n29521 = ~n28749 & ~n28762 ;
  assign n29522 = n29520 & n29521 ;
  assign n29523 = ~n29520 & ~n29521 ;
  assign n29524 = ~n29522 & ~n29523 ;
  assign n29525 = x86 & n14233 ;
  assign n29526 = x84 & n14876 ;
  assign n29527 = x85 & n14228 ;
  assign n29528 = ~n29526 & ~n29527 ;
  assign n29529 = ~n29525 & n29528 ;
  assign n29530 = n3686 & n14236 ;
  assign n29531 = n29529 & ~n29530 ;
  assign n29532 = x47 & ~n29531 ;
  assign n29533 = x47 & ~n29532 ;
  assign n29534 = ~n29531 & ~n29532 ;
  assign n29535 = ~n29533 & ~n29534 ;
  assign n29536 = n29524 & ~n29535 ;
  assign n29537 = n29524 & ~n29536 ;
  assign n29538 = ~n29535 & ~n29536 ;
  assign n29539 = ~n29537 & ~n29538 ;
  assign n29540 = ~n28768 & ~n28782 ;
  assign n29541 = ~n29539 & ~n29540 ;
  assign n29542 = ~n29539 & ~n29541 ;
  assign n29543 = ~n29540 & ~n29541 ;
  assign n29544 = ~n29542 & ~n29543 ;
  assign n29545 = x89 & n12506 ;
  assign n29546 = x87 & n13131 ;
  assign n29547 = x88 & n12501 ;
  assign n29548 = ~n29546 & ~n29547 ;
  assign n29549 = ~n29545 & n29548 ;
  assign n29550 = n4488 & n12509 ;
  assign n29551 = n29549 & ~n29550 ;
  assign n29552 = x44 & ~n29551 ;
  assign n29553 = x44 & ~n29552 ;
  assign n29554 = ~n29551 & ~n29552 ;
  assign n29555 = ~n29553 & ~n29554 ;
  assign n29556 = ~n29544 & ~n29555 ;
  assign n29557 = ~n29544 & ~n29556 ;
  assign n29558 = ~n29555 & ~n29556 ;
  assign n29559 = ~n29557 & ~n29558 ;
  assign n29560 = ~n28786 & ~n28800 ;
  assign n29561 = n29559 & n29560 ;
  assign n29562 = ~n29559 & ~n29560 ;
  assign n29563 = ~n29561 & ~n29562 ;
  assign n29564 = x92 & n10905 ;
  assign n29565 = x90 & n11466 ;
  assign n29566 = x91 & n10900 ;
  assign n29567 = ~n29565 & ~n29566 ;
  assign n29568 = ~n29564 & n29567 ;
  assign n29569 = n5710 & n10908 ;
  assign n29570 = n29568 & ~n29569 ;
  assign n29571 = x41 & ~n29570 ;
  assign n29572 = x41 & ~n29571 ;
  assign n29573 = ~n29570 & ~n29571 ;
  assign n29574 = ~n29572 & ~n29573 ;
  assign n29575 = n29563 & ~n29574 ;
  assign n29576 = n29563 & ~n29575 ;
  assign n29577 = ~n29574 & ~n29575 ;
  assign n29578 = ~n29576 & ~n29577 ;
  assign n29579 = ~n28806 & ~n28819 ;
  assign n29580 = n29578 & n29579 ;
  assign n29581 = ~n29578 & ~n29579 ;
  assign n29582 = ~n29580 & ~n29581 ;
  assign n29583 = x95 & n9433 ;
  assign n29584 = x93 & n9915 ;
  assign n29585 = x94 & n9428 ;
  assign n29586 = ~n29584 & ~n29585 ;
  assign n29587 = ~n29583 & n29586 ;
  assign n29588 = n6894 & n9436 ;
  assign n29589 = n29587 & ~n29588 ;
  assign n29590 = x38 & ~n29589 ;
  assign n29591 = x38 & ~n29590 ;
  assign n29592 = ~n29589 & ~n29590 ;
  assign n29593 = ~n29591 & ~n29592 ;
  assign n29594 = ~n29582 & n29593 ;
  assign n29595 = n29582 & ~n29593 ;
  assign n29596 = ~n29594 & ~n29595 ;
  assign n29597 = ~n29422 & n29596 ;
  assign n29598 = ~n29422 & ~n29597 ;
  assign n29599 = n29596 & ~n29597 ;
  assign n29600 = ~n29598 & ~n29599 ;
  assign n29601 = ~n29421 & ~n29600 ;
  assign n29602 = ~n29421 & ~n29601 ;
  assign n29603 = ~n29600 & ~n29601 ;
  assign n29604 = ~n29602 & ~n29603 ;
  assign n29605 = ~n29410 & n29604 ;
  assign n29606 = n29410 & ~n29604 ;
  assign n29607 = ~n29605 & ~n29606 ;
  assign n29608 = ~n28871 & ~n28875 ;
  assign n29609 = x104 & n5560 ;
  assign n29610 = x102 & n5943 ;
  assign n29611 = x103 & n5555 ;
  assign n29612 = ~n29610 & ~n29611 ;
  assign n29613 = ~n29609 & n29612 ;
  assign n29614 = ~n5563 & n29613 ;
  assign n29615 = ~n11116 & n29613 ;
  assign n29616 = ~n29614 & ~n29615 ;
  assign n29617 = x29 & ~n29616 ;
  assign n29618 = ~x29 & n29616 ;
  assign n29619 = ~n29617 & ~n29618 ;
  assign n29620 = ~n29608 & ~n29619 ;
  assign n29621 = ~n29608 & ~n29620 ;
  assign n29622 = ~n29619 & ~n29620 ;
  assign n29623 = ~n29621 & ~n29622 ;
  assign n29624 = n29607 & ~n29623 ;
  assign n29625 = n29607 & ~n29624 ;
  assign n29626 = ~n29623 & ~n29624 ;
  assign n29627 = ~n29625 & ~n29626 ;
  assign n29628 = n29395 & ~n29627 ;
  assign n29629 = n29395 & ~n29628 ;
  assign n29630 = ~n29627 & ~n29628 ;
  assign n29631 = ~n29629 & ~n29630 ;
  assign n29632 = x110 & n3589 ;
  assign n29633 = x108 & n3878 ;
  assign n29634 = x109 & n3584 ;
  assign n29635 = ~n29633 & ~n29634 ;
  assign n29636 = ~n29632 & n29635 ;
  assign n29637 = n3592 & n14497 ;
  assign n29638 = n29636 & ~n29637 ;
  assign n29639 = x23 & ~n29638 ;
  assign n29640 = x23 & ~n29639 ;
  assign n29641 = ~n29638 & ~n29639 ;
  assign n29642 = ~n29640 & ~n29641 ;
  assign n29643 = ~n28654 & ~n28883 ;
  assign n29644 = ~n29642 & ~n29643 ;
  assign n29645 = ~n29642 & ~n29644 ;
  assign n29646 = ~n29643 & ~n29644 ;
  assign n29647 = ~n29645 & ~n29646 ;
  assign n29648 = ~n29631 & n29647 ;
  assign n29649 = n29631 & ~n29647 ;
  assign n29650 = ~n29648 & ~n29649 ;
  assign n29651 = n29380 & ~n29650 ;
  assign n29652 = n29380 & ~n29651 ;
  assign n29653 = ~n29650 & ~n29651 ;
  assign n29654 = ~n29652 & ~n29653 ;
  assign n29655 = x116 & n2093 ;
  assign n29656 = x114 & n2275 ;
  assign n29657 = x115 & n2088 ;
  assign n29658 = ~n29656 & ~n29657 ;
  assign n29659 = ~n29655 & n29658 ;
  assign n29660 = n2096 & n18336 ;
  assign n29661 = n29659 & ~n29660 ;
  assign n29662 = x17 & ~n29661 ;
  assign n29663 = x17 & ~n29662 ;
  assign n29664 = ~n29661 & ~n29662 ;
  assign n29665 = ~n29663 & ~n29664 ;
  assign n29666 = ~n28625 & ~n28891 ;
  assign n29667 = ~n29665 & ~n29666 ;
  assign n29668 = ~n29665 & ~n29667 ;
  assign n29669 = ~n29666 & ~n29667 ;
  assign n29670 = ~n29668 & ~n29669 ;
  assign n29671 = ~n29654 & n29670 ;
  assign n29672 = n29654 & ~n29670 ;
  assign n29673 = ~n29671 & ~n29672 ;
  assign n29674 = n29364 & ~n29673 ;
  assign n29675 = n29364 & ~n29674 ;
  assign n29676 = ~n29673 & ~n29674 ;
  assign n29677 = ~n29675 & ~n29676 ;
  assign n29678 = ~n28911 & ~n28915 ;
  assign n29679 = x122 & n945 ;
  assign n29680 = x120 & n1099 ;
  assign n29681 = x121 & n940 ;
  assign n29682 = ~n29680 & ~n29681 ;
  assign n29683 = ~n29679 & n29682 ;
  assign n29684 = ~n948 & n29683 ;
  assign n29685 = ~n22622 & n29683 ;
  assign n29686 = ~n29684 & ~n29685 ;
  assign n29687 = x11 & ~n29686 ;
  assign n29688 = ~x11 & n29686 ;
  assign n29689 = ~n29687 & ~n29688 ;
  assign n29690 = ~n29678 & ~n29689 ;
  assign n29691 = ~n29678 & ~n29690 ;
  assign n29692 = ~n29689 & ~n29690 ;
  assign n29693 = ~n29691 & ~n29692 ;
  assign n29694 = ~n29677 & ~n29693 ;
  assign n29695 = ~n29677 & ~n29694 ;
  assign n29696 = ~n29693 & ~n29694 ;
  assign n29697 = ~n29695 & ~n29696 ;
  assign n29698 = ~n28595 & ~n28919 ;
  assign n29699 = x125 & n574 ;
  assign n29700 = x123 & n673 ;
  assign n29701 = x124 & n569 ;
  assign n29702 = ~n29700 & ~n29701 ;
  assign n29703 = ~n29699 & n29702 ;
  assign n29704 = ~n577 & n29703 ;
  assign n29705 = ~n24935 & n29703 ;
  assign n29706 = ~n29704 & ~n29705 ;
  assign n29707 = x8 & ~n29706 ;
  assign n29708 = ~x8 & n29706 ;
  assign n29709 = ~n29707 & ~n29708 ;
  assign n29710 = ~n29698 & ~n29709 ;
  assign n29711 = ~n29698 & ~n29710 ;
  assign n29712 = ~n29709 & ~n29710 ;
  assign n29713 = ~n29711 & ~n29712 ;
  assign n29714 = ~n29697 & ~n29713 ;
  assign n29715 = ~n29697 & ~n29714 ;
  assign n29716 = ~n29713 & ~n29714 ;
  assign n29717 = ~n29715 & ~n29716 ;
  assign n29718 = ~n28935 & ~n28939 ;
  assign n29719 = x126 & n373 ;
  assign n29720 = x127 & n288 ;
  assign n29721 = ~n29719 & ~n29720 ;
  assign n29722 = ~n296 & n29721 ;
  assign n29723 = n26965 & n29721 ;
  assign n29724 = ~n29722 & ~n29723 ;
  assign n29725 = x5 & ~n29724 ;
  assign n29726 = ~x5 & n29724 ;
  assign n29727 = ~n29725 & ~n29726 ;
  assign n29728 = ~n29718 & ~n29727 ;
  assign n29729 = ~n29718 & ~n29728 ;
  assign n29730 = ~n29727 & ~n29728 ;
  assign n29731 = ~n29729 & ~n29730 ;
  assign n29732 = ~n29717 & ~n29731 ;
  assign n29733 = n29717 & ~n29730 ;
  assign n29734 = ~n29729 & n29733 ;
  assign n29735 = ~n29732 & ~n29734 ;
  assign n29736 = ~n29349 & n29735 ;
  assign n29737 = ~n29349 & ~n29736 ;
  assign n29738 = n29735 & ~n29736 ;
  assign n29739 = ~n29737 & ~n29738 ;
  assign n29740 = ~n29348 & ~n29739 ;
  assign n29741 = n29348 & ~n29738 ;
  assign n29742 = ~n29737 & n29741 ;
  assign n29743 = ~n29740 & ~n29742 ;
  assign n30141 = n29743 & x195 ;
  assign n29744 = ~n29338 & ~n29341 ;
  assign n29745 = ~n28967 & ~n29332 ;
  assign n29746 = ~x119 & n1434 ;
  assign n29747 = ~x117 & n1646 ;
  assign n29748 = ~x118 & n1429 ;
  assign n29749 = ~n29747 & ~n29748 ;
  assign n29750 = ~n29746 & n29749 ;
  assign n29751 = n1437 & n20778 ;
  assign n29752 = n29750 & ~n29751 ;
  assign n29753 = ~x14 & ~n29752 ;
  assign n29754 = ~x14 & ~n29753 ;
  assign n29755 = ~n29752 & ~n29753 ;
  assign n29756 = ~n29754 & ~n29755 ;
  assign n29757 = ~n28999 & ~n29283 ;
  assign n29758 = n29756 & n29757 ;
  assign n29759 = ~n29756 & ~n29757 ;
  assign n29760 = ~n29758 & ~n29759 ;
  assign n29761 = ~x113 & n2751 ;
  assign n29762 = ~x111 & n3020 ;
  assign n29763 = ~x112 & n2746 ;
  assign n29764 = ~n29762 & ~n29763 ;
  assign n29765 = ~n29761 & n29764 ;
  assign n29766 = n2754 & n16684 ;
  assign n29767 = n29765 & ~n29766 ;
  assign n29768 = ~x20 & ~n29767 ;
  assign n29769 = ~x20 & ~n29768 ;
  assign n29770 = ~n29767 & ~n29768 ;
  assign n29771 = ~n29769 & ~n29770 ;
  assign n29772 = ~n28424 & ~n29026 ;
  assign n29773 = ~n29275 & ~n29772 ;
  assign n29774 = n29771 & n29773 ;
  assign n29775 = ~n29771 & ~n29773 ;
  assign n29776 = ~n29774 & ~n29775 ;
  assign n29777 = ~x107 & n4531 ;
  assign n29778 = ~x105 & n4847 ;
  assign n29779 = ~x106 & n4526 ;
  assign n29780 = ~n29778 & ~n29779 ;
  assign n29781 = ~n29777 & n29780 ;
  assign n29782 = n4534 & n13034 ;
  assign n29783 = n29781 & ~n29782 ;
  assign n29784 = ~x26 & ~n29783 ;
  assign n29785 = ~x26 & ~n29784 ;
  assign n29786 = ~n29783 & ~n29784 ;
  assign n29787 = ~n29785 & ~n29786 ;
  assign n29788 = ~n29057 & ~n29268 ;
  assign n29789 = n29787 & n29788 ;
  assign n29790 = ~n29787 & ~n29788 ;
  assign n29791 = ~n29789 & ~n29790 ;
  assign n29792 = ~n29231 & ~n29245 ;
  assign n29793 = ~x101 & n6725 ;
  assign n29794 = ~x99 & n7129 ;
  assign n29795 = ~x100 & n6720 ;
  assign n29796 = ~n29794 & ~n29795 ;
  assign n29797 = ~n29793 & n29796 ;
  assign n29798 = ~n6728 & n29797 ;
  assign n29799 = ~n9844 & n29797 ;
  assign n29800 = ~n29798 & ~n29799 ;
  assign n29801 = ~x32 & ~n29800 ;
  assign n29802 = x32 & n29800 ;
  assign n29803 = ~n29801 & ~n29802 ;
  assign n29804 = ~n29792 & ~n29803 ;
  assign n29805 = n29792 & n29803 ;
  assign n29806 = ~n29804 & ~n29805 ;
  assign n29807 = ~x98 & n8006 ;
  assign n29808 = ~x96 & n8474 ;
  assign n29809 = ~x97 & n8001 ;
  assign n29810 = ~n29808 & ~n29809 ;
  assign n29811 = ~n29807 & n29810 ;
  assign n29812 = n8009 & n8426 ;
  assign n29813 = n29811 & ~n29812 ;
  assign n29814 = ~x35 & ~n29813 ;
  assign n29815 = ~x35 & ~n29814 ;
  assign n29816 = ~n29813 & ~n29814 ;
  assign n29817 = ~n29815 & ~n29816 ;
  assign n29818 = ~n29214 & ~n29228 ;
  assign n29819 = ~x71 & n24612 ;
  assign n29820 = ~x69 & n25390 ;
  assign n29821 = ~x70 & n24607 ;
  assign n29822 = ~n29820 & ~n29821 ;
  assign n29823 = ~n29819 & n29822 ;
  assign n29824 = n622 & n24615 ;
  assign n29825 = n29823 & ~n29824 ;
  assign n29826 = ~x62 & ~n29825 ;
  assign n29827 = ~x62 & ~n29826 ;
  assign n29828 = ~n29825 & ~n29826 ;
  assign n29829 = ~n29827 & ~n29828 ;
  assign n29830 = ~x67 & n27427 ;
  assign n29831 = ~x68 & ~n26217 ;
  assign n29832 = ~n29830 & ~n29831 ;
  assign n29833 = ~x2 & ~n29832 ;
  assign n29834 = ~x2 & ~n29833 ;
  assign n29835 = ~n29832 & ~n29833 ;
  assign n29836 = ~n29834 & ~n29835 ;
  assign n29837 = ~n29829 & ~n29836 ;
  assign n29838 = ~n29829 & ~n29837 ;
  assign n29839 = ~n29836 & ~n29837 ;
  assign n29840 = ~n29838 & ~n29839 ;
  assign n29841 = ~n29065 & ~n29079 ;
  assign n29842 = n29840 & n29841 ;
  assign n29843 = ~n29840 & ~n29841 ;
  assign n29844 = ~n29842 & ~n29843 ;
  assign n29845 = ~x74 & n22325 ;
  assign n29846 = ~x72 & n23066 ;
  assign n29847 = ~x73 & n22320 ;
  assign n29848 = ~n29846 & ~n29847 ;
  assign n29849 = ~n29845 & n29848 ;
  assign n29850 = n1066 & n22328 ;
  assign n29851 = n29849 & ~n29850 ;
  assign n29852 = ~x59 & ~n29851 ;
  assign n29853 = ~x59 & ~n29852 ;
  assign n29854 = ~n29851 & ~n29852 ;
  assign n29855 = ~n29853 & ~n29854 ;
  assign n29856 = n29844 & ~n29855 ;
  assign n29857 = n29844 & ~n29856 ;
  assign n29858 = ~n29855 & ~n29856 ;
  assign n29859 = ~n29857 & ~n29858 ;
  assign n29860 = ~n29082 & ~n29096 ;
  assign n29861 = n29859 & n29860 ;
  assign n29862 = ~n29859 & ~n29860 ;
  assign n29863 = ~n29861 & ~n29862 ;
  assign n29864 = ~x77 & n20143 ;
  assign n29865 = ~x75 & n20854 ;
  assign n29866 = ~x76 & n20138 ;
  assign n29867 = ~n29865 & ~n29866 ;
  assign n29868 = ~n29864 & n29867 ;
  assign n29869 = n1594 & n20146 ;
  assign n29870 = n29868 & ~n29869 ;
  assign n29871 = ~x56 & ~n29870 ;
  assign n29872 = ~x56 & ~n29871 ;
  assign n29873 = ~n29870 & ~n29871 ;
  assign n29874 = ~n29872 & ~n29873 ;
  assign n29875 = ~n29863 & n29874 ;
  assign n29876 = n29863 & ~n29874 ;
  assign n29877 = ~n29875 & ~n29876 ;
  assign n29878 = ~n28223 & ~n29099 ;
  assign n29879 = ~n29115 & ~n29878 ;
  assign n29880 = n29877 & ~n29879 ;
  assign n29881 = ~n29877 & n29879 ;
  assign n29882 = ~n29880 & ~n29881 ;
  assign n29883 = ~x80 & n18025 ;
  assign n29884 = ~x78 & n18764 ;
  assign n29885 = ~x79 & n18020 ;
  assign n29886 = ~n29884 & ~n29885 ;
  assign n29887 = ~n29883 & n29886 ;
  assign n29888 = n2145 & n18028 ;
  assign n29889 = n29887 & ~n29888 ;
  assign n29890 = ~x53 & ~n29889 ;
  assign n29891 = ~x53 & ~n29890 ;
  assign n29892 = ~n29889 & ~n29890 ;
  assign n29893 = ~n29891 & ~n29892 ;
  assign n29894 = n29882 & ~n29893 ;
  assign n29895 = n29882 & ~n29894 ;
  assign n29896 = ~n29893 & ~n29894 ;
  assign n29897 = ~n29895 & ~n29896 ;
  assign n29898 = ~n29117 & ~n29131 ;
  assign n29899 = n29897 & n29898 ;
  assign n29900 = ~n29897 & ~n29898 ;
  assign n29901 = ~n29899 & ~n29900 ;
  assign n29902 = ~x83 & n16076 ;
  assign n29903 = ~x81 & n16756 ;
  assign n29904 = ~x82 & n16071 ;
  assign n29905 = ~n29903 & ~n29904 ;
  assign n29906 = ~n29902 & n29905 ;
  assign n29907 = n2972 & n16079 ;
  assign n29908 = n29906 & ~n29907 ;
  assign n29909 = ~x50 & ~n29908 ;
  assign n29910 = ~x50 & ~n29909 ;
  assign n29911 = ~n29908 & ~n29909 ;
  assign n29912 = ~n29910 & ~n29911 ;
  assign n29913 = n29901 & ~n29912 ;
  assign n29914 = n29901 & ~n29913 ;
  assign n29915 = ~n29912 & ~n29913 ;
  assign n29916 = ~n29914 & ~n29915 ;
  assign n29917 = ~n29138 & ~n29151 ;
  assign n29918 = n29916 & n29917 ;
  assign n29919 = ~n29916 & ~n29917 ;
  assign n29920 = ~n29918 & ~n29919 ;
  assign n29921 = ~x86 & n14233 ;
  assign n29922 = ~x84 & n14876 ;
  assign n29923 = ~x85 & n14228 ;
  assign n29924 = ~n29922 & ~n29923 ;
  assign n29925 = ~n29921 & n29924 ;
  assign n29926 = n3832 & n14236 ;
  assign n29927 = n29925 & ~n29926 ;
  assign n29928 = ~x47 & ~n29927 ;
  assign n29929 = ~x47 & ~n29928 ;
  assign n29930 = ~n29927 & ~n29928 ;
  assign n29931 = ~n29929 & ~n29930 ;
  assign n29932 = n29920 & ~n29931 ;
  assign n29933 = n29920 & ~n29932 ;
  assign n29934 = ~n29931 & ~n29932 ;
  assign n29935 = ~n29933 & ~n29934 ;
  assign n29936 = ~n29157 & ~n29171 ;
  assign n29937 = ~n29935 & ~n29936 ;
  assign n29938 = ~n29935 & ~n29937 ;
  assign n29939 = ~n29936 & ~n29937 ;
  assign n29940 = ~n29938 & ~n29939 ;
  assign n29941 = ~x89 & n12506 ;
  assign n29942 = ~x87 & n13131 ;
  assign n29943 = ~x88 & n12501 ;
  assign n29944 = ~n29942 & ~n29943 ;
  assign n29945 = ~n29941 & n29944 ;
  assign n29946 = n4664 & n12509 ;
  assign n29947 = n29945 & ~n29946 ;
  assign n29948 = ~x44 & ~n29947 ;
  assign n29949 = ~x44 & ~n29948 ;
  assign n29950 = ~n29947 & ~n29948 ;
  assign n29951 = ~n29949 & ~n29950 ;
  assign n29952 = ~n29940 & ~n29951 ;
  assign n29953 = ~n29940 & ~n29952 ;
  assign n29954 = ~n29951 & ~n29952 ;
  assign n29955 = ~n29953 & ~n29954 ;
  assign n29956 = ~n29175 & ~n29189 ;
  assign n29957 = n29955 & n29956 ;
  assign n29958 = ~n29955 & ~n29956 ;
  assign n29959 = ~n29957 & ~n29958 ;
  assign n29960 = ~x92 & n10905 ;
  assign n29961 = ~x90 & n11466 ;
  assign n29962 = ~x91 & n10900 ;
  assign n29963 = ~n29961 & ~n29962 ;
  assign n29964 = ~n29960 & n29963 ;
  assign n29965 = n5896 & n10908 ;
  assign n29966 = n29964 & ~n29965 ;
  assign n29967 = ~x41 & ~n29966 ;
  assign n29968 = ~x41 & ~n29967 ;
  assign n29969 = ~n29966 & ~n29967 ;
  assign n29970 = ~n29968 & ~n29969 ;
  assign n29971 = n29959 & ~n29970 ;
  assign n29972 = n29959 & ~n29971 ;
  assign n29973 = ~n29970 & ~n29971 ;
  assign n29974 = ~n29972 & ~n29973 ;
  assign n29975 = ~n29195 & ~n29208 ;
  assign n29976 = n29974 & n29975 ;
  assign n29977 = ~n29974 & ~n29975 ;
  assign n29978 = ~n29976 & ~n29977 ;
  assign n29979 = ~x95 & n9433 ;
  assign n29980 = ~x93 & n9915 ;
  assign n29981 = ~x94 & n9428 ;
  assign n29982 = ~n29980 & ~n29981 ;
  assign n29983 = ~n29979 & n29982 ;
  assign n29984 = n7100 & n9436 ;
  assign n29985 = n29983 & ~n29984 ;
  assign n29986 = ~x38 & ~n29985 ;
  assign n29987 = ~x38 & ~n29986 ;
  assign n29988 = ~n29985 & ~n29986 ;
  assign n29989 = ~n29987 & ~n29988 ;
  assign n29990 = ~n29978 & n29989 ;
  assign n29991 = n29978 & ~n29989 ;
  assign n29992 = ~n29990 & ~n29991 ;
  assign n29993 = ~n29818 & n29992 ;
  assign n29994 = ~n29818 & ~n29993 ;
  assign n29995 = n29992 & ~n29993 ;
  assign n29996 = ~n29994 & ~n29995 ;
  assign n29997 = ~n29817 & ~n29996 ;
  assign n29998 = ~n29817 & ~n29997 ;
  assign n29999 = ~n29996 & ~n29997 ;
  assign n30000 = ~n29998 & ~n29999 ;
  assign n30001 = ~n29806 & n30000 ;
  assign n30002 = n29806 & ~n30000 ;
  assign n30003 = ~n30001 & ~n30002 ;
  assign n30004 = ~n29260 & ~n29264 ;
  assign n30005 = ~x104 & n5560 ;
  assign n30006 = ~x102 & n5943 ;
  assign n30007 = ~x103 & n5555 ;
  assign n30008 = ~n30006 & ~n30007 ;
  assign n30009 = ~n30005 & n30008 ;
  assign n30010 = ~n5563 & n30009 ;
  assign n30011 = ~n11380 & n30009 ;
  assign n30012 = ~n30010 & ~n30011 ;
  assign n30013 = ~x29 & ~n30012 ;
  assign n30014 = x29 & n30012 ;
  assign n30015 = ~n30013 & ~n30014 ;
  assign n30016 = ~n30004 & ~n30015 ;
  assign n30017 = ~n30004 & ~n30016 ;
  assign n30018 = ~n30015 & ~n30016 ;
  assign n30019 = ~n30017 & ~n30018 ;
  assign n30020 = n30003 & ~n30019 ;
  assign n30021 = n30003 & ~n30020 ;
  assign n30022 = ~n30019 & ~n30020 ;
  assign n30023 = ~n30021 & ~n30022 ;
  assign n30024 = n29791 & ~n30023 ;
  assign n30025 = n29791 & ~n30024 ;
  assign n30026 = ~n30023 & ~n30024 ;
  assign n30027 = ~n30025 & ~n30026 ;
  assign n30028 = ~x110 & n3589 ;
  assign n30029 = ~x108 & n3878 ;
  assign n30030 = ~x109 & n3584 ;
  assign n30031 = ~n30029 & ~n30030 ;
  assign n30032 = ~n30028 & n30031 ;
  assign n30033 = n3592 & n14802 ;
  assign n30034 = n30032 & ~n30033 ;
  assign n30035 = ~x23 & ~n30034 ;
  assign n30036 = ~x23 & ~n30035 ;
  assign n30037 = ~n30034 & ~n30035 ;
  assign n30038 = ~n30036 & ~n30037 ;
  assign n30039 = ~n29043 & ~n29272 ;
  assign n30040 = ~n30038 & ~n30039 ;
  assign n30041 = ~n30038 & ~n30040 ;
  assign n30042 = ~n30039 & ~n30040 ;
  assign n30043 = ~n30041 & ~n30042 ;
  assign n30044 = ~n30027 & n30043 ;
  assign n30045 = n30027 & ~n30043 ;
  assign n30046 = ~n30044 & ~n30045 ;
  assign n30047 = n29776 & ~n30046 ;
  assign n30048 = n29776 & ~n30047 ;
  assign n30049 = ~n30046 & ~n30047 ;
  assign n30050 = ~n30048 & ~n30049 ;
  assign n30051 = ~x116 & n2093 ;
  assign n30052 = ~x114 & n2275 ;
  assign n30053 = ~x115 & n2088 ;
  assign n30054 = ~n30052 & ~n30053 ;
  assign n30055 = ~n30051 & n30054 ;
  assign n30056 = n2096 & n18678 ;
  assign n30057 = n30055 & ~n30056 ;
  assign n30058 = ~x17 & ~n30057 ;
  assign n30059 = ~x17 & ~n30058 ;
  assign n30060 = ~n30057 & ~n30058 ;
  assign n30061 = ~n30059 & ~n30060 ;
  assign n30062 = ~n29014 & ~n29280 ;
  assign n30063 = ~n30061 & ~n30062 ;
  assign n30064 = ~n30061 & ~n30063 ;
  assign n30065 = ~n30062 & ~n30063 ;
  assign n30066 = ~n30064 & ~n30065 ;
  assign n30067 = ~n30050 & n30066 ;
  assign n30068 = n30050 & ~n30066 ;
  assign n30069 = ~n30067 & ~n30068 ;
  assign n30070 = n29760 & ~n30069 ;
  assign n30071 = n29760 & ~n30070 ;
  assign n30072 = ~n30069 & ~n30070 ;
  assign n30073 = ~n30071 & ~n30072 ;
  assign n30074 = ~n29300 & ~n29304 ;
  assign n30075 = ~x122 & n945 ;
  assign n30076 = ~x120 & n1099 ;
  assign n30077 = ~x121 & n940 ;
  assign n30078 = ~n30076 & ~n30077 ;
  assign n30079 = ~n30075 & n30078 ;
  assign n30080 = ~n948 & n30079 ;
  assign n30081 = ~n22998 & n30079 ;
  assign n30082 = ~n30080 & ~n30081 ;
  assign n30083 = ~x11 & ~n30082 ;
  assign n30084 = x11 & n30082 ;
  assign n30085 = ~n30083 & ~n30084 ;
  assign n30086 = ~n30074 & ~n30085 ;
  assign n30087 = ~n30074 & ~n30086 ;
  assign n30088 = ~n30085 & ~n30086 ;
  assign n30089 = ~n30087 & ~n30088 ;
  assign n30090 = ~n30073 & ~n30089 ;
  assign n30091 = ~n30073 & ~n30090 ;
  assign n30092 = ~n30089 & ~n30090 ;
  assign n30093 = ~n30091 & ~n30092 ;
  assign n30094 = ~n28984 & ~n29308 ;
  assign n30095 = ~x125 & n574 ;
  assign n30096 = ~x123 & n673 ;
  assign n30097 = ~x124 & n569 ;
  assign n30098 = ~n30096 & ~n30097 ;
  assign n30099 = ~n30095 & n30098 ;
  assign n30100 = ~n577 & n30099 ;
  assign n30101 = ~n25330 & n30099 ;
  assign n30102 = ~n30100 & ~n30101 ;
  assign n30103 = ~x8 & ~n30102 ;
  assign n30104 = x8 & n30102 ;
  assign n30105 = ~n30103 & ~n30104 ;
  assign n30106 = ~n30094 & ~n30105 ;
  assign n30107 = ~n30094 & ~n30106 ;
  assign n30108 = ~n30105 & ~n30106 ;
  assign n30109 = ~n30107 & ~n30108 ;
  assign n30110 = ~n30093 & ~n30109 ;
  assign n30111 = ~n30093 & ~n30110 ;
  assign n30112 = ~n30109 & ~n30110 ;
  assign n30113 = ~n30111 & ~n30112 ;
  assign n30114 = ~n29324 & ~n29328 ;
  assign n30115 = ~x126 & n373 ;
  assign n30116 = ~x127 & n288 ;
  assign n30117 = ~n30115 & ~n30116 ;
  assign n30118 = ~n296 & n30117 ;
  assign n30119 = n27368 & n30117 ;
  assign n30120 = ~n30118 & ~n30119 ;
  assign n30121 = ~x5 & ~n30120 ;
  assign n30122 = x5 & n30120 ;
  assign n30123 = ~n30121 & ~n30122 ;
  assign n30124 = ~n30114 & ~n30123 ;
  assign n30125 = ~n30114 & ~n30124 ;
  assign n30126 = ~n30123 & ~n30124 ;
  assign n30127 = ~n30125 & ~n30126 ;
  assign n30128 = ~n30113 & ~n30127 ;
  assign n30129 = n30113 & ~n30126 ;
  assign n30130 = ~n30125 & n30129 ;
  assign n30131 = ~n30128 & ~n30130 ;
  assign n30132 = ~n29745 & n30131 ;
  assign n30133 = ~n29745 & ~n30132 ;
  assign n30134 = n30131 & ~n30132 ;
  assign n30135 = ~n30133 & ~n30134 ;
  assign n30136 = ~n29744 & ~n30135 ;
  assign n30137 = n29744 & ~n30134 ;
  assign n30138 = ~n30133 & n30137 ;
  assign n30139 = ~n30136 & ~n30138 ;
  assign n30142 = ~n30139 & ~x195 ;
  assign n30143 = ~n30141 & ~n30142 ;
  assign n30144 = ~n29736 & ~n29740 ;
  assign n30145 = ~n29728 & ~n29732 ;
  assign n30146 = ~n29710 & ~n29714 ;
  assign n30147 = x127 & n373 ;
  assign n30148 = n296 & n26962 ;
  assign n30149 = ~n30147 & ~n30148 ;
  assign n30150 = x5 & ~n30149 ;
  assign n30151 = x5 & ~n30150 ;
  assign n30152 = ~n30149 & ~n30150 ;
  assign n30153 = ~n30151 & ~n30152 ;
  assign n30154 = ~n30146 & ~n30153 ;
  assign n30155 = ~n30146 & ~n30154 ;
  assign n30156 = ~n30153 & ~n30154 ;
  assign n30157 = ~n30155 & ~n30156 ;
  assign n30158 = x123 & n945 ;
  assign n30159 = x121 & n1099 ;
  assign n30160 = x122 & n940 ;
  assign n30161 = ~n30159 & ~n30160 ;
  assign n30162 = ~n30158 & n30161 ;
  assign n30163 = n948 & n23382 ;
  assign n30164 = n30162 & ~n30163 ;
  assign n30165 = x11 & ~n30164 ;
  assign n30166 = x11 & ~n30165 ;
  assign n30167 = ~n30164 & ~n30165 ;
  assign n30168 = ~n30166 & ~n30167 ;
  assign n30169 = ~n29363 & ~n29674 ;
  assign n30170 = n30168 & n30169 ;
  assign n30171 = ~n30168 & ~n30169 ;
  assign n30172 = ~n30170 & ~n30171 ;
  assign n30173 = x120 & n1434 ;
  assign n30174 = x118 & n1646 ;
  assign n30175 = x119 & n1429 ;
  assign n30176 = ~n30174 & ~n30175 ;
  assign n30177 = ~n30173 & n30176 ;
  assign n30178 = n1437 & n21143 ;
  assign n30179 = n30177 & ~n30178 ;
  assign n30180 = x14 & ~n30179 ;
  assign n30181 = x14 & ~n30180 ;
  assign n30182 = ~n30179 & ~n30180 ;
  assign n30183 = ~n30181 & ~n30182 ;
  assign n30184 = ~n29654 & ~n29670 ;
  assign n30185 = ~n29667 & ~n30184 ;
  assign n30186 = ~n30183 & ~n30185 ;
  assign n30187 = ~n30183 & ~n30186 ;
  assign n30188 = ~n30185 & ~n30186 ;
  assign n30189 = ~n30187 & ~n30188 ;
  assign n30190 = ~n29379 & ~n29651 ;
  assign n30191 = x117 & n2093 ;
  assign n30192 = x115 & n2275 ;
  assign n30193 = x116 & n2088 ;
  assign n30194 = ~n30192 & ~n30193 ;
  assign n30195 = ~n30191 & n30194 ;
  assign n30196 = ~n2096 & n30195 ;
  assign n30197 = ~n19026 & n30195 ;
  assign n30198 = ~n30196 & ~n30197 ;
  assign n30199 = x17 & ~n30198 ;
  assign n30200 = ~x17 & n30198 ;
  assign n30201 = ~n30199 & ~n30200 ;
  assign n30202 = ~n30190 & ~n30201 ;
  assign n30203 = n30190 & n30201 ;
  assign n30204 = ~n30202 & ~n30203 ;
  assign n30205 = x114 & n2751 ;
  assign n30206 = x112 & n3020 ;
  assign n30207 = x113 & n2746 ;
  assign n30208 = ~n30206 & ~n30207 ;
  assign n30209 = ~n30205 & n30208 ;
  assign n30210 = n2754 & n17012 ;
  assign n30211 = n30209 & ~n30210 ;
  assign n30212 = x20 & ~n30211 ;
  assign n30213 = x20 & ~n30212 ;
  assign n30214 = ~n30211 & ~n30212 ;
  assign n30215 = ~n30213 & ~n30214 ;
  assign n30216 = ~n29631 & ~n29647 ;
  assign n30217 = ~n29644 & ~n30216 ;
  assign n30218 = ~n30215 & ~n30217 ;
  assign n30219 = ~n30215 & ~n30218 ;
  assign n30220 = ~n30217 & ~n30218 ;
  assign n30221 = ~n30219 & ~n30220 ;
  assign n30222 = x111 & n3589 ;
  assign n30223 = x109 & n3878 ;
  assign n30224 = x110 & n3584 ;
  assign n30225 = ~n30223 & ~n30224 ;
  assign n30226 = ~n30222 & n30225 ;
  assign n30227 = n3592 & n15111 ;
  assign n30228 = n30226 & ~n30227 ;
  assign n30229 = x23 & ~n30228 ;
  assign n30230 = x23 & ~n30229 ;
  assign n30231 = ~n30228 & ~n30229 ;
  assign n30232 = ~n30230 & ~n30231 ;
  assign n30233 = ~n29394 & ~n29628 ;
  assign n30234 = n30232 & n30233 ;
  assign n30235 = ~n30232 & ~n30233 ;
  assign n30236 = ~n30234 & ~n30235 ;
  assign n30237 = x105 & n5560 ;
  assign n30238 = x103 & n5943 ;
  assign n30239 = x104 & n5555 ;
  assign n30240 = ~n30238 & ~n30239 ;
  assign n30241 = ~n30237 & n30240 ;
  assign n30242 = n5563 & n11648 ;
  assign n30243 = n30241 & ~n30242 ;
  assign n30244 = x29 & ~n30243 ;
  assign n30245 = x29 & ~n30244 ;
  assign n30246 = ~n30243 & ~n30244 ;
  assign n30247 = ~n30245 & ~n30246 ;
  assign n30248 = ~n29408 & ~n29606 ;
  assign n30249 = n30247 & n30248 ;
  assign n30250 = ~n30247 & ~n30248 ;
  assign n30251 = ~n30249 & ~n30250 ;
  assign n30252 = x72 & n24612 ;
  assign n30253 = x70 & n25390 ;
  assign n30254 = x71 & n24607 ;
  assign n30255 = ~n30253 & ~n30254 ;
  assign n30256 = ~n30252 & n30255 ;
  assign n30257 = n717 & n24615 ;
  assign n30258 = n30256 & ~n30257 ;
  assign n30259 = x62 & ~n30258 ;
  assign n30260 = x62 & ~n30259 ;
  assign n30261 = ~n30258 & ~n30259 ;
  assign n30262 = ~n30260 & ~n30261 ;
  assign n30263 = x68 & n27024 ;
  assign n30264 = x69 & ~n26217 ;
  assign n30265 = ~n30263 & ~n30264 ;
  assign n30266 = x2 & ~n30265 ;
  assign n30267 = x2 & ~n30266 ;
  assign n30268 = ~n30265 & ~n30266 ;
  assign n30269 = ~n30267 & ~n30268 ;
  assign n30270 = ~n30262 & ~n30269 ;
  assign n30271 = ~n30262 & ~n30270 ;
  assign n30272 = ~n30269 & ~n30270 ;
  assign n30273 = ~n30271 & ~n30272 ;
  assign n30274 = ~n29437 & ~n29441 ;
  assign n30275 = n30273 & n30274 ;
  assign n30276 = ~n30273 & ~n30274 ;
  assign n30277 = ~n30275 & ~n30276 ;
  assign n30278 = x75 & n22325 ;
  assign n30279 = x73 & n23066 ;
  assign n30280 = x74 & n22320 ;
  assign n30281 = ~n30279 & ~n30280 ;
  assign n30282 = ~n30278 & n30281 ;
  assign n30283 = n1150 & n22328 ;
  assign n30284 = n30282 & ~n30283 ;
  assign n30285 = x59 & ~n30284 ;
  assign n30286 = x59 & ~n30285 ;
  assign n30287 = ~n30284 & ~n30285 ;
  assign n30288 = ~n30286 & ~n30287 ;
  assign n30289 = ~n30277 & n30288 ;
  assign n30290 = n30277 & ~n30288 ;
  assign n30291 = ~n30289 & ~n30290 ;
  assign n30292 = ~n29447 & ~n29460 ;
  assign n30293 = n30291 & ~n30292 ;
  assign n30294 = ~n30291 & n30292 ;
  assign n30295 = ~n30293 & ~n30294 ;
  assign n30296 = x78 & n20143 ;
  assign n30297 = x76 & n20854 ;
  assign n30298 = x77 & n20138 ;
  assign n30299 = ~n30297 & ~n30298 ;
  assign n30300 = ~n30296 & n30299 ;
  assign n30301 = n1624 & n20146 ;
  assign n30302 = n30300 & ~n30301 ;
  assign n30303 = x56 & ~n30302 ;
  assign n30304 = x56 & ~n30303 ;
  assign n30305 = ~n30302 & ~n30303 ;
  assign n30306 = ~n30304 & ~n30305 ;
  assign n30307 = n30295 & ~n30306 ;
  assign n30308 = n30295 & ~n30307 ;
  assign n30309 = ~n30306 & ~n30307 ;
  assign n30310 = ~n30308 & ~n30309 ;
  assign n30311 = ~n29466 & ~n29480 ;
  assign n30312 = ~n30310 & ~n30311 ;
  assign n30313 = ~n30310 & ~n30312 ;
  assign n30314 = ~n30311 & ~n30312 ;
  assign n30315 = ~n30313 & ~n30314 ;
  assign n30316 = x81 & n18025 ;
  assign n30317 = x79 & n18764 ;
  assign n30318 = x80 & n18020 ;
  assign n30319 = ~n30317 & ~n30318 ;
  assign n30320 = ~n30316 & n30319 ;
  assign n30321 = n2348 & n18028 ;
  assign n30322 = n30320 & ~n30321 ;
  assign n30323 = x53 & ~n30322 ;
  assign n30324 = x53 & ~n30323 ;
  assign n30325 = ~n30322 & ~n30323 ;
  assign n30326 = ~n30324 & ~n30325 ;
  assign n30327 = ~n30315 & ~n30326 ;
  assign n30328 = ~n30315 & ~n30327 ;
  assign n30329 = ~n30326 & ~n30327 ;
  assign n30330 = ~n30328 & ~n30329 ;
  assign n30331 = ~n29484 & ~n29498 ;
  assign n30332 = n30330 & n30331 ;
  assign n30333 = ~n30330 & ~n30331 ;
  assign n30334 = ~n30332 & ~n30333 ;
  assign n30335 = x84 & n16076 ;
  assign n30336 = x82 & n16756 ;
  assign n30337 = x83 & n16071 ;
  assign n30338 = ~n30336 & ~n30337 ;
  assign n30339 = ~n30335 & n30338 ;
  assign n30340 = n3114 & n16079 ;
  assign n30341 = n30339 & ~n30340 ;
  assign n30342 = x50 & ~n30341 ;
  assign n30343 = x50 & ~n30342 ;
  assign n30344 = ~n30341 & ~n30342 ;
  assign n30345 = ~n30343 & ~n30344 ;
  assign n30346 = ~n30334 & n30345 ;
  assign n30347 = n30334 & ~n30345 ;
  assign n30348 = ~n30346 & ~n30347 ;
  assign n30349 = ~n29504 & ~n29517 ;
  assign n30350 = n30348 & ~n30349 ;
  assign n30351 = ~n30348 & n30349 ;
  assign n30352 = ~n30350 & ~n30351 ;
  assign n30353 = x87 & n14233 ;
  assign n30354 = x85 & n14876 ;
  assign n30355 = x86 & n14228 ;
  assign n30356 = ~n30354 & ~n30355 ;
  assign n30357 = ~n30353 & n30356 ;
  assign n30358 = n3991 & n14236 ;
  assign n30359 = n30357 & ~n30358 ;
  assign n30360 = x47 & ~n30359 ;
  assign n30361 = x47 & ~n30360 ;
  assign n30362 = ~n30359 & ~n30360 ;
  assign n30363 = ~n30361 & ~n30362 ;
  assign n30364 = n30352 & ~n30363 ;
  assign n30365 = n30352 & ~n30364 ;
  assign n30366 = ~n30363 & ~n30364 ;
  assign n30367 = ~n30365 & ~n30366 ;
  assign n30368 = ~n29523 & ~n29536 ;
  assign n30369 = n30367 & n30368 ;
  assign n30370 = ~n30367 & ~n30368 ;
  assign n30371 = ~n30369 & ~n30370 ;
  assign n30372 = x90 & n12506 ;
  assign n30373 = x88 & n13131 ;
  assign n30374 = x89 & n12501 ;
  assign n30375 = ~n30373 & ~n30374 ;
  assign n30376 = ~n30372 & n30375 ;
  assign n30377 = n4986 & n12509 ;
  assign n30378 = n30376 & ~n30377 ;
  assign n30379 = x44 & ~n30378 ;
  assign n30380 = x44 & ~n30379 ;
  assign n30381 = ~n30378 & ~n30379 ;
  assign n30382 = ~n30380 & ~n30381 ;
  assign n30383 = n30371 & ~n30382 ;
  assign n30384 = n30371 & ~n30383 ;
  assign n30385 = ~n30382 & ~n30383 ;
  assign n30386 = ~n30384 & ~n30385 ;
  assign n30387 = ~n29541 & ~n29556 ;
  assign n30388 = n30386 & n30387 ;
  assign n30389 = ~n30386 & ~n30387 ;
  assign n30390 = ~n30388 & ~n30389 ;
  assign n30391 = x93 & n10905 ;
  assign n30392 = x91 & n11466 ;
  assign n30393 = x92 & n10900 ;
  assign n30394 = ~n30392 & ~n30393 ;
  assign n30395 = ~n30391 & n30394 ;
  assign n30396 = n6094 & n10908 ;
  assign n30397 = n30395 & ~n30396 ;
  assign n30398 = x41 & ~n30397 ;
  assign n30399 = x41 & ~n30398 ;
  assign n30400 = ~n30397 & ~n30398 ;
  assign n30401 = ~n30399 & ~n30400 ;
  assign n30402 = n30390 & ~n30401 ;
  assign n30403 = n30390 & ~n30402 ;
  assign n30404 = ~n30401 & ~n30402 ;
  assign n30405 = ~n30403 & ~n30404 ;
  assign n30406 = ~n29562 & ~n29575 ;
  assign n30407 = n30405 & n30406 ;
  assign n30408 = ~n30405 & ~n30406 ;
  assign n30409 = ~n30407 & ~n30408 ;
  assign n30410 = x96 & n9433 ;
  assign n30411 = x94 & n9915 ;
  assign n30412 = x95 & n9428 ;
  assign n30413 = ~n30411 & ~n30412 ;
  assign n30414 = ~n30410 & n30413 ;
  assign n30415 = n7321 & n9436 ;
  assign n30416 = n30414 & ~n30415 ;
  assign n30417 = x38 & ~n30416 ;
  assign n30418 = x38 & ~n30417 ;
  assign n30419 = ~n30416 & ~n30417 ;
  assign n30420 = ~n30418 & ~n30419 ;
  assign n30421 = ~n30409 & n30420 ;
  assign n30422 = n30409 & ~n30420 ;
  assign n30423 = ~n30421 & ~n30422 ;
  assign n30424 = ~n29581 & ~n29595 ;
  assign n30425 = n30423 & ~n30424 ;
  assign n30426 = ~n30423 & n30424 ;
  assign n30427 = ~n30425 & ~n30426 ;
  assign n30428 = x99 & n8006 ;
  assign n30429 = x97 & n8474 ;
  assign n30430 = x98 & n8001 ;
  assign n30431 = ~n30429 & ~n30430 ;
  assign n30432 = ~n30428 & n30431 ;
  assign n30433 = n8009 & n8660 ;
  assign n30434 = n30432 & ~n30433 ;
  assign n30435 = x35 & ~n30434 ;
  assign n30436 = x35 & ~n30435 ;
  assign n30437 = ~n30434 & ~n30435 ;
  assign n30438 = ~n30436 & ~n30437 ;
  assign n30439 = n30427 & ~n30438 ;
  assign n30440 = n30427 & ~n30439 ;
  assign n30441 = ~n30438 & ~n30439 ;
  assign n30442 = ~n30440 & ~n30441 ;
  assign n30443 = ~n29597 & ~n29601 ;
  assign n30444 = x102 & n6725 ;
  assign n30445 = x100 & n7129 ;
  assign n30446 = x101 & n6720 ;
  assign n30447 = ~n30445 & ~n30446 ;
  assign n30448 = ~n30444 & n30447 ;
  assign n30449 = ~n6728 & n30448 ;
  assign n30450 = ~n10092 & n30448 ;
  assign n30451 = ~n30449 & ~n30450 ;
  assign n30452 = x32 & ~n30451 ;
  assign n30453 = ~x32 & n30451 ;
  assign n30454 = ~n30452 & ~n30453 ;
  assign n30455 = ~n30443 & ~n30454 ;
  assign n30456 = n30443 & n30454 ;
  assign n30457 = ~n30455 & ~n30456 ;
  assign n30458 = ~n30442 & n30457 ;
  assign n30459 = ~n30442 & ~n30458 ;
  assign n30460 = n30457 & ~n30458 ;
  assign n30461 = ~n30459 & ~n30460 ;
  assign n30462 = n30251 & ~n30461 ;
  assign n30463 = n30251 & ~n30462 ;
  assign n30464 = ~n30461 & ~n30462 ;
  assign n30465 = ~n30463 & ~n30464 ;
  assign n30466 = ~n29620 & ~n29624 ;
  assign n30467 = x108 & n4531 ;
  assign n30468 = x106 & n4847 ;
  assign n30469 = x107 & n4526 ;
  assign n30470 = ~n30468 & ~n30469 ;
  assign n30471 = ~n30467 & n30470 ;
  assign n30472 = ~n4534 & n30471 ;
  assign n30473 = ~n13323 & n30471 ;
  assign n30474 = ~n30472 & ~n30473 ;
  assign n30475 = x26 & ~n30474 ;
  assign n30476 = ~x26 & n30474 ;
  assign n30477 = ~n30475 & ~n30476 ;
  assign n30478 = ~n30466 & ~n30477 ;
  assign n30479 = ~n30466 & ~n30478 ;
  assign n30480 = ~n30477 & ~n30478 ;
  assign n30481 = ~n30479 & ~n30480 ;
  assign n30482 = ~n30465 & ~n30481 ;
  assign n30483 = ~n30465 & ~n30482 ;
  assign n30484 = ~n30481 & ~n30482 ;
  assign n30485 = ~n30483 & ~n30484 ;
  assign n30486 = n30236 & ~n30485 ;
  assign n30487 = n30236 & ~n30486 ;
  assign n30488 = ~n30485 & ~n30486 ;
  assign n30489 = ~n30487 & ~n30488 ;
  assign n30490 = ~n30221 & n30489 ;
  assign n30491 = n30221 & ~n30489 ;
  assign n30492 = ~n30490 & ~n30491 ;
  assign n30493 = n30204 & ~n30492 ;
  assign n30494 = n30204 & ~n30493 ;
  assign n30495 = ~n30492 & ~n30493 ;
  assign n30496 = ~n30494 & ~n30495 ;
  assign n30497 = ~n30189 & n30496 ;
  assign n30498 = n30189 & ~n30496 ;
  assign n30499 = ~n30497 & ~n30498 ;
  assign n30500 = n30172 & ~n30499 ;
  assign n30501 = n30172 & ~n30500 ;
  assign n30502 = ~n30499 & ~n30500 ;
  assign n30503 = ~n30501 & ~n30502 ;
  assign n30504 = ~n29690 & ~n29694 ;
  assign n30505 = x126 & n574 ;
  assign n30506 = x124 & n673 ;
  assign n30507 = x125 & n569 ;
  assign n30508 = ~n30506 & ~n30507 ;
  assign n30509 = ~n30505 & n30508 ;
  assign n30510 = ~n577 & n30509 ;
  assign n30511 = ~n25735 & n30509 ;
  assign n30512 = ~n30510 & ~n30511 ;
  assign n30513 = x8 & ~n30512 ;
  assign n30514 = ~x8 & n30512 ;
  assign n30515 = ~n30513 & ~n30514 ;
  assign n30516 = ~n30504 & ~n30515 ;
  assign n30517 = ~n30504 & ~n30516 ;
  assign n30518 = ~n30515 & ~n30516 ;
  assign n30519 = ~n30517 & ~n30518 ;
  assign n30520 = ~n30503 & ~n30519 ;
  assign n30521 = n30503 & ~n30518 ;
  assign n30522 = ~n30517 & n30521 ;
  assign n30523 = ~n30520 & ~n30522 ;
  assign n30524 = ~n30157 & n30523 ;
  assign n30525 = n30157 & ~n30523 ;
  assign n30526 = ~n30524 & ~n30525 ;
  assign n30527 = ~n30145 & n30526 ;
  assign n30528 = ~n30145 & ~n30527 ;
  assign n30529 = n30526 & ~n30527 ;
  assign n30530 = ~n30528 & ~n30529 ;
  assign n30531 = ~n30144 & ~n30530 ;
  assign n30532 = n30144 & ~n30529 ;
  assign n30533 = ~n30528 & n30532 ;
  assign n30534 = ~n30531 & ~n30533 ;
  assign n30927 = n30534 & x196 ;
  assign n30535 = ~n30132 & ~n30136 ;
  assign n30536 = ~n30124 & ~n30128 ;
  assign n30537 = ~n30106 & ~n30110 ;
  assign n30538 = ~x127 & n373 ;
  assign n30539 = n296 & n27365 ;
  assign n30540 = ~n30538 & ~n30539 ;
  assign n30541 = ~x5 & ~n30540 ;
  assign n30542 = ~x5 & ~n30541 ;
  assign n30543 = ~n30540 & ~n30541 ;
  assign n30544 = ~n30542 & ~n30543 ;
  assign n30545 = ~n30537 & ~n30544 ;
  assign n30546 = ~n30537 & ~n30545 ;
  assign n30547 = ~n30544 & ~n30545 ;
  assign n30548 = ~n30546 & ~n30547 ;
  assign n30549 = ~x123 & n945 ;
  assign n30550 = ~x121 & n1099 ;
  assign n30551 = ~x122 & n940 ;
  assign n30552 = ~n30550 & ~n30551 ;
  assign n30553 = ~n30549 & n30552 ;
  assign n30554 = n948 & n23760 ;
  assign n30555 = n30553 & ~n30554 ;
  assign n30556 = ~x11 & ~n30555 ;
  assign n30557 = ~x11 & ~n30556 ;
  assign n30558 = ~n30555 & ~n30556 ;
  assign n30559 = ~n30557 & ~n30558 ;
  assign n30560 = ~n29759 & ~n30070 ;
  assign n30561 = n30559 & n30560 ;
  assign n30562 = ~n30559 & ~n30560 ;
  assign n30563 = ~n30561 & ~n30562 ;
  assign n30564 = ~x120 & n1434 ;
  assign n30565 = ~x118 & n1646 ;
  assign n30566 = ~x119 & n1429 ;
  assign n30567 = ~n30565 & ~n30566 ;
  assign n30568 = ~n30564 & n30567 ;
  assign n30569 = n1437 & n21501 ;
  assign n30570 = n30568 & ~n30569 ;
  assign n30571 = ~x14 & ~n30570 ;
  assign n30572 = ~x14 & ~n30571 ;
  assign n30573 = ~n30570 & ~n30571 ;
  assign n30574 = ~n30572 & ~n30573 ;
  assign n30575 = ~n30050 & ~n30066 ;
  assign n30576 = ~n30063 & ~n30575 ;
  assign n30577 = ~n30574 & ~n30576 ;
  assign n30578 = ~n30574 & ~n30577 ;
  assign n30579 = ~n30576 & ~n30577 ;
  assign n30580 = ~n30578 & ~n30579 ;
  assign n30581 = ~n29775 & ~n30047 ;
  assign n30582 = ~x117 & n2093 ;
  assign n30583 = ~x115 & n2275 ;
  assign n30584 = ~x116 & n2088 ;
  assign n30585 = ~n30583 & ~n30584 ;
  assign n30586 = ~n30582 & n30585 ;
  assign n30587 = ~n2096 & n30586 ;
  assign n30588 = ~n19365 & n30586 ;
  assign n30589 = ~n30587 & ~n30588 ;
  assign n30590 = ~x17 & ~n30589 ;
  assign n30591 = x17 & n30589 ;
  assign n30592 = ~n30590 & ~n30591 ;
  assign n30593 = ~n30581 & ~n30592 ;
  assign n30594 = n30581 & n30592 ;
  assign n30595 = ~n30593 & ~n30594 ;
  assign n30596 = ~x114 & n2751 ;
  assign n30597 = ~x112 & n3020 ;
  assign n30598 = ~x113 & n2746 ;
  assign n30599 = ~n30597 & ~n30598 ;
  assign n30600 = ~n30596 & n30599 ;
  assign n30601 = n2754 & n17333 ;
  assign n30602 = n30600 & ~n30601 ;
  assign n30603 = ~x20 & ~n30602 ;
  assign n30604 = ~x20 & ~n30603 ;
  assign n30605 = ~n30602 & ~n30603 ;
  assign n30606 = ~n30604 & ~n30605 ;
  assign n30607 = ~n30027 & ~n30043 ;
  assign n30608 = ~n30040 & ~n30607 ;
  assign n30609 = ~n30606 & ~n30608 ;
  assign n30610 = ~n30606 & ~n30609 ;
  assign n30611 = ~n30608 & ~n30609 ;
  assign n30612 = ~n30610 & ~n30611 ;
  assign n30613 = ~x111 & n3589 ;
  assign n30614 = ~x109 & n3878 ;
  assign n30615 = ~x110 & n3584 ;
  assign n30616 = ~n30614 & ~n30615 ;
  assign n30617 = ~n30613 & n30616 ;
  assign n30618 = n3592 & n15411 ;
  assign n30619 = n30617 & ~n30618 ;
  assign n30620 = ~x23 & ~n30619 ;
  assign n30621 = ~x23 & ~n30620 ;
  assign n30622 = ~n30619 & ~n30620 ;
  assign n30623 = ~n30621 & ~n30622 ;
  assign n30624 = ~n29790 & ~n30024 ;
  assign n30625 = n30623 & n30624 ;
  assign n30626 = ~n30623 & ~n30624 ;
  assign n30627 = ~n30625 & ~n30626 ;
  assign n30628 = ~x105 & n5560 ;
  assign n30629 = ~x103 & n5943 ;
  assign n30630 = ~x104 & n5555 ;
  assign n30631 = ~n30629 & ~n30630 ;
  assign n30632 = ~n30628 & n30631 ;
  assign n30633 = n5563 & n11907 ;
  assign n30634 = n30632 & ~n30633 ;
  assign n30635 = ~x29 & ~n30634 ;
  assign n30636 = ~x29 & ~n30635 ;
  assign n30637 = ~n30634 & ~n30635 ;
  assign n30638 = ~n30636 & ~n30637 ;
  assign n30639 = ~n29804 & ~n30002 ;
  assign n30640 = n30638 & n30639 ;
  assign n30641 = ~n30638 & ~n30639 ;
  assign n30642 = ~n30640 & ~n30641 ;
  assign n30643 = ~x72 & n24612 ;
  assign n30644 = ~x70 & n25390 ;
  assign n30645 = ~x71 & n24607 ;
  assign n30646 = ~n30644 & ~n30645 ;
  assign n30647 = ~n30643 & n30646 ;
  assign n30648 = n773 & n24615 ;
  assign n30649 = n30647 & ~n30648 ;
  assign n30650 = ~x62 & ~n30649 ;
  assign n30651 = ~x62 & ~n30650 ;
  assign n30652 = ~n30649 & ~n30650 ;
  assign n30653 = ~n30651 & ~n30652 ;
  assign n30654 = ~x68 & n27427 ;
  assign n30655 = ~x69 & ~n26217 ;
  assign n30656 = ~n30654 & ~n30655 ;
  assign n30657 = ~x2 & ~n30656 ;
  assign n30658 = ~x2 & ~n30657 ;
  assign n30659 = ~n30656 & ~n30657 ;
  assign n30660 = ~n30658 & ~n30659 ;
  assign n30661 = ~n30653 & ~n30660 ;
  assign n30662 = ~n30653 & ~n30661 ;
  assign n30663 = ~n30660 & ~n30661 ;
  assign n30664 = ~n30662 & ~n30663 ;
  assign n30665 = ~n29833 & ~n29837 ;
  assign n30666 = n30664 & n30665 ;
  assign n30667 = ~n30664 & ~n30665 ;
  assign n30668 = ~n30666 & ~n30667 ;
  assign n30669 = ~x75 & n22325 ;
  assign n30670 = ~x73 & n23066 ;
  assign n30671 = ~x74 & n22320 ;
  assign n30672 = ~n30670 & ~n30671 ;
  assign n30673 = ~n30669 & n30672 ;
  assign n30674 = n1225 & n22328 ;
  assign n30675 = n30673 & ~n30674 ;
  assign n30676 = ~x59 & ~n30675 ;
  assign n30677 = ~x59 & ~n30676 ;
  assign n30678 = ~n30675 & ~n30676 ;
  assign n30679 = ~n30677 & ~n30678 ;
  assign n30680 = ~n30668 & n30679 ;
  assign n30681 = n30668 & ~n30679 ;
  assign n30682 = ~n30680 & ~n30681 ;
  assign n30683 = ~n29843 & ~n29856 ;
  assign n30684 = n30682 & ~n30683 ;
  assign n30685 = ~n30682 & n30683 ;
  assign n30686 = ~n30684 & ~n30685 ;
  assign n30687 = ~x78 & n20143 ;
  assign n30688 = ~x76 & n20854 ;
  assign n30689 = ~x77 & n20138 ;
  assign n30690 = ~n30688 & ~n30689 ;
  assign n30691 = ~n30687 & n30690 ;
  assign n30692 = n1718 & n20146 ;
  assign n30693 = n30691 & ~n30692 ;
  assign n30694 = ~x56 & ~n30693 ;
  assign n30695 = ~x56 & ~n30694 ;
  assign n30696 = ~n30693 & ~n30694 ;
  assign n30697 = ~n30695 & ~n30696 ;
  assign n30698 = n30686 & ~n30697 ;
  assign n30699 = n30686 & ~n30698 ;
  assign n30700 = ~n30697 & ~n30698 ;
  assign n30701 = ~n30699 & ~n30700 ;
  assign n30702 = ~n29862 & ~n29876 ;
  assign n30703 = ~n30701 & ~n30702 ;
  assign n30704 = ~n30701 & ~n30703 ;
  assign n30705 = ~n30702 & ~n30703 ;
  assign n30706 = ~n30704 & ~n30705 ;
  assign n30707 = ~x81 & n18025 ;
  assign n30708 = ~x79 & n18764 ;
  assign n30709 = ~x80 & n18020 ;
  assign n30710 = ~n30708 & ~n30709 ;
  assign n30711 = ~n30707 & n30710 ;
  assign n30712 = n2460 & n18028 ;
  assign n30713 = n30711 & ~n30712 ;
  assign n30714 = ~x53 & ~n30713 ;
  assign n30715 = ~x53 & ~n30714 ;
  assign n30716 = ~n30713 & ~n30714 ;
  assign n30717 = ~n30715 & ~n30716 ;
  assign n30718 = ~n30706 & ~n30717 ;
  assign n30719 = ~n30706 & ~n30718 ;
  assign n30720 = ~n30717 & ~n30718 ;
  assign n30721 = ~n30719 & ~n30720 ;
  assign n30722 = ~n29880 & ~n29894 ;
  assign n30723 = n30721 & n30722 ;
  assign n30724 = ~n30721 & ~n30722 ;
  assign n30725 = ~n30723 & ~n30724 ;
  assign n30726 = ~x84 & n16076 ;
  assign n30727 = ~x82 & n16756 ;
  assign n30728 = ~x83 & n16071 ;
  assign n30729 = ~n30727 & ~n30728 ;
  assign n30730 = ~n30726 & n30729 ;
  assign n30731 = n3247 & n16079 ;
  assign n30732 = n30730 & ~n30731 ;
  assign n30733 = ~x50 & ~n30732 ;
  assign n30734 = ~x50 & ~n30733 ;
  assign n30735 = ~n30732 & ~n30733 ;
  assign n30736 = ~n30734 & ~n30735 ;
  assign n30737 = ~n30725 & n30736 ;
  assign n30738 = n30725 & ~n30736 ;
  assign n30739 = ~n30737 & ~n30738 ;
  assign n30740 = ~n29900 & ~n29913 ;
  assign n30741 = n30739 & ~n30740 ;
  assign n30742 = ~n30739 & n30740 ;
  assign n30743 = ~n30741 & ~n30742 ;
  assign n30744 = ~x87 & n14233 ;
  assign n30745 = ~x85 & n14876 ;
  assign n30746 = ~x86 & n14228 ;
  assign n30747 = ~n30745 & ~n30746 ;
  assign n30748 = ~n30744 & n30747 ;
  assign n30749 = n4143 & n14236 ;
  assign n30750 = n30748 & ~n30749 ;
  assign n30751 = ~x47 & ~n30750 ;
  assign n30752 = ~x47 & ~n30751 ;
  assign n30753 = ~n30750 & ~n30751 ;
  assign n30754 = ~n30752 & ~n30753 ;
  assign n30755 = n30743 & ~n30754 ;
  assign n30756 = n30743 & ~n30755 ;
  assign n30757 = ~n30754 & ~n30755 ;
  assign n30758 = ~n30756 & ~n30757 ;
  assign n30759 = ~n29919 & ~n29932 ;
  assign n30760 = n30758 & n30759 ;
  assign n30761 = ~n30758 & ~n30759 ;
  assign n30762 = ~n30760 & ~n30761 ;
  assign n30763 = ~x90 & n12506 ;
  assign n30764 = ~x88 & n13131 ;
  assign n30765 = ~x89 & n12501 ;
  assign n30766 = ~n30764 & ~n30765 ;
  assign n30767 = ~n30763 & n30766 ;
  assign n30768 = n5155 & n12509 ;
  assign n30769 = n30767 & ~n30768 ;
  assign n30770 = ~x44 & ~n30769 ;
  assign n30771 = ~x44 & ~n30770 ;
  assign n30772 = ~n30769 & ~n30770 ;
  assign n30773 = ~n30771 & ~n30772 ;
  assign n30774 = n30762 & ~n30773 ;
  assign n30775 = n30762 & ~n30774 ;
  assign n30776 = ~n30773 & ~n30774 ;
  assign n30777 = ~n30775 & ~n30776 ;
  assign n30778 = ~n29937 & ~n29952 ;
  assign n30779 = n30777 & n30778 ;
  assign n30780 = ~n30777 & ~n30778 ;
  assign n30781 = ~n30779 & ~n30780 ;
  assign n30782 = ~x93 & n10905 ;
  assign n30783 = ~x91 & n11466 ;
  assign n30784 = ~x92 & n10900 ;
  assign n30785 = ~n30783 & ~n30784 ;
  assign n30786 = ~n30782 & n30785 ;
  assign n30787 = n6285 & n10908 ;
  assign n30788 = n30786 & ~n30787 ;
  assign n30789 = ~x41 & ~n30788 ;
  assign n30790 = ~x41 & ~n30789 ;
  assign n30791 = ~n30788 & ~n30789 ;
  assign n30792 = ~n30790 & ~n30791 ;
  assign n30793 = n30781 & ~n30792 ;
  assign n30794 = n30781 & ~n30793 ;
  assign n30795 = ~n30792 & ~n30793 ;
  assign n30796 = ~n30794 & ~n30795 ;
  assign n30797 = ~n29958 & ~n29971 ;
  assign n30798 = n30796 & n30797 ;
  assign n30799 = ~n30796 & ~n30797 ;
  assign n30800 = ~n30798 & ~n30799 ;
  assign n30801 = ~x96 & n9433 ;
  assign n30802 = ~x94 & n9915 ;
  assign n30803 = ~x95 & n9428 ;
  assign n30804 = ~n30802 & ~n30803 ;
  assign n30805 = ~n30801 & n30804 ;
  assign n30806 = n7531 & n9436 ;
  assign n30807 = n30805 & ~n30806 ;
  assign n30808 = ~x38 & ~n30807 ;
  assign n30809 = ~x38 & ~n30808 ;
  assign n30810 = ~n30807 & ~n30808 ;
  assign n30811 = ~n30809 & ~n30810 ;
  assign n30812 = ~n30800 & n30811 ;
  assign n30813 = n30800 & ~n30811 ;
  assign n30814 = ~n30812 & ~n30813 ;
  assign n30815 = ~n29977 & ~n29991 ;
  assign n30816 = n30814 & ~n30815 ;
  assign n30817 = ~n30814 & n30815 ;
  assign n30818 = ~n30816 & ~n30817 ;
  assign n30819 = ~x99 & n8006 ;
  assign n30820 = ~x97 & n8474 ;
  assign n30821 = ~x98 & n8001 ;
  assign n30822 = ~n30820 & ~n30821 ;
  assign n30823 = ~n30819 & n30822 ;
  assign n30824 = n8009 & n8885 ;
  assign n30825 = n30823 & ~n30824 ;
  assign n30826 = ~x35 & ~n30825 ;
  assign n30827 = ~x35 & ~n30826 ;
  assign n30828 = ~n30825 & ~n30826 ;
  assign n30829 = ~n30827 & ~n30828 ;
  assign n30830 = n30818 & ~n30829 ;
  assign n30831 = n30818 & ~n30830 ;
  assign n30832 = ~n30829 & ~n30830 ;
  assign n30833 = ~n30831 & ~n30832 ;
  assign n30834 = ~n29993 & ~n29997 ;
  assign n30835 = ~x102 & n6725 ;
  assign n30836 = ~x100 & n7129 ;
  assign n30837 = ~x101 & n6720 ;
  assign n30838 = ~n30836 & ~n30837 ;
  assign n30839 = ~n30835 & n30838 ;
  assign n30840 = ~n6728 & n30839 ;
  assign n30841 = ~n10333 & n30839 ;
  assign n30842 = ~n30840 & ~n30841 ;
  assign n30843 = ~x32 & ~n30842 ;
  assign n30844 = x32 & n30842 ;
  assign n30845 = ~n30843 & ~n30844 ;
  assign n30846 = ~n30834 & ~n30845 ;
  assign n30847 = n30834 & n30845 ;
  assign n30848 = ~n30846 & ~n30847 ;
  assign n30849 = ~n30833 & n30848 ;
  assign n30850 = ~n30833 & ~n30849 ;
  assign n30851 = n30848 & ~n30849 ;
  assign n30852 = ~n30850 & ~n30851 ;
  assign n30853 = n30642 & ~n30852 ;
  assign n30854 = n30642 & ~n30853 ;
  assign n30855 = ~n30852 & ~n30853 ;
  assign n30856 = ~n30854 & ~n30855 ;
  assign n30857 = ~n30016 & ~n30020 ;
  assign n30858 = ~x108 & n4531 ;
  assign n30859 = ~x106 & n4847 ;
  assign n30860 = ~x107 & n4526 ;
  assign n30861 = ~n30859 & ~n30860 ;
  assign n30862 = ~n30858 & n30861 ;
  assign n30863 = ~n4534 & n30862 ;
  assign n30864 = ~n13601 & n30862 ;
  assign n30865 = ~n30863 & ~n30864 ;
  assign n30866 = ~x26 & ~n30865 ;
  assign n30867 = x26 & n30865 ;
  assign n30868 = ~n30866 & ~n30867 ;
  assign n30869 = ~n30857 & ~n30868 ;
  assign n30870 = ~n30857 & ~n30869 ;
  assign n30871 = ~n30868 & ~n30869 ;
  assign n30872 = ~n30870 & ~n30871 ;
  assign n30873 = ~n30856 & ~n30872 ;
  assign n30874 = ~n30856 & ~n30873 ;
  assign n30875 = ~n30872 & ~n30873 ;
  assign n30876 = ~n30874 & ~n30875 ;
  assign n30877 = n30627 & ~n30876 ;
  assign n30878 = n30627 & ~n30877 ;
  assign n30879 = ~n30876 & ~n30877 ;
  assign n30880 = ~n30878 & ~n30879 ;
  assign n30881 = ~n30612 & n30880 ;
  assign n30882 = n30612 & ~n30880 ;
  assign n30883 = ~n30881 & ~n30882 ;
  assign n30884 = n30595 & ~n30883 ;
  assign n30885 = n30595 & ~n30884 ;
  assign n30886 = ~n30883 & ~n30884 ;
  assign n30887 = ~n30885 & ~n30886 ;
  assign n30888 = ~n30580 & n30887 ;
  assign n30889 = n30580 & ~n30887 ;
  assign n30890 = ~n30888 & ~n30889 ;
  assign n30891 = n30563 & ~n30890 ;
  assign n30892 = n30563 & ~n30891 ;
  assign n30893 = ~n30890 & ~n30891 ;
  assign n30894 = ~n30892 & ~n30893 ;
  assign n30895 = ~n30086 & ~n30090 ;
  assign n30896 = ~x126 & n574 ;
  assign n30897 = ~x124 & n673 ;
  assign n30898 = ~x125 & n569 ;
  assign n30899 = ~n30897 & ~n30898 ;
  assign n30900 = ~n30896 & n30899 ;
  assign n30901 = ~n577 & n30900 ;
  assign n30902 = ~n26128 & n30900 ;
  assign n30903 = ~n30901 & ~n30902 ;
  assign n30904 = ~x8 & ~n30903 ;
  assign n30905 = x8 & n30903 ;
  assign n30906 = ~n30904 & ~n30905 ;
  assign n30907 = ~n30895 & ~n30906 ;
  assign n30908 = ~n30895 & ~n30907 ;
  assign n30909 = ~n30906 & ~n30907 ;
  assign n30910 = ~n30908 & ~n30909 ;
  assign n30911 = ~n30894 & ~n30910 ;
  assign n30912 = n30894 & ~n30909 ;
  assign n30913 = ~n30908 & n30912 ;
  assign n30914 = ~n30911 & ~n30913 ;
  assign n30915 = ~n30548 & n30914 ;
  assign n30916 = n30548 & ~n30914 ;
  assign n30917 = ~n30915 & ~n30916 ;
  assign n30918 = ~n30536 & n30917 ;
  assign n30919 = ~n30536 & ~n30918 ;
  assign n30920 = n30917 & ~n30918 ;
  assign n30921 = ~n30919 & ~n30920 ;
  assign n30922 = ~n30535 & ~n30921 ;
  assign n30923 = n30535 & ~n30920 ;
  assign n30924 = ~n30919 & n30923 ;
  assign n30925 = ~n30922 & ~n30924 ;
  assign n30928 = ~n30925 & ~x196 ;
  assign n30929 = ~n30927 & ~n30928 ;
  assign n30930 = ~n30527 & ~n30531 ;
  assign n30931 = ~n30154 & ~n30524 ;
  assign n30932 = ~n30516 & ~n30520 ;
  assign n30933 = x127 & n574 ;
  assign n30934 = x125 & n673 ;
  assign n30935 = x126 & n569 ;
  assign n30936 = ~n30934 & ~n30935 ;
  assign n30937 = ~n30933 & n30936 ;
  assign n30938 = n577 & n26533 ;
  assign n30939 = n30937 & ~n30938 ;
  assign n30940 = x8 & ~n30939 ;
  assign n30941 = x8 & ~n30940 ;
  assign n30942 = ~n30939 & ~n30940 ;
  assign n30943 = ~n30941 & ~n30942 ;
  assign n30944 = ~n30932 & ~n30943 ;
  assign n30945 = ~n30932 & ~n30944 ;
  assign n30946 = ~n30943 & ~n30944 ;
  assign n30947 = ~n30945 & ~n30946 ;
  assign n30948 = x124 & n945 ;
  assign n30949 = x122 & n1099 ;
  assign n30950 = x123 & n940 ;
  assign n30951 = ~n30949 & ~n30950 ;
  assign n30952 = ~n30948 & n30951 ;
  assign n30953 = n948 & n23796 ;
  assign n30954 = n30952 & ~n30953 ;
  assign n30955 = x11 & ~n30954 ;
  assign n30956 = x11 & ~n30955 ;
  assign n30957 = ~n30954 & ~n30955 ;
  assign n30958 = ~n30956 & ~n30957 ;
  assign n30959 = ~n30171 & ~n30500 ;
  assign n30960 = n30958 & n30959 ;
  assign n30961 = ~n30958 & ~n30959 ;
  assign n30962 = ~n30960 & ~n30961 ;
  assign n30963 = ~n30202 & ~n30493 ;
  assign n30964 = x118 & n2093 ;
  assign n30965 = x116 & n2275 ;
  assign n30966 = x117 & n2088 ;
  assign n30967 = ~n30965 & ~n30966 ;
  assign n30968 = ~n30964 & n30967 ;
  assign n30969 = n2096 & n19395 ;
  assign n30970 = n30968 & ~n30969 ;
  assign n30971 = x17 & ~n30970 ;
  assign n30972 = x17 & ~n30971 ;
  assign n30973 = ~n30970 & ~n30971 ;
  assign n30974 = ~n30972 & ~n30973 ;
  assign n30975 = ~n30963 & ~n30974 ;
  assign n30976 = ~n30963 & ~n30975 ;
  assign n30977 = ~n30974 & ~n30975 ;
  assign n30978 = ~n30976 & ~n30977 ;
  assign n30979 = x112 & n3589 ;
  assign n30980 = x110 & n3878 ;
  assign n30981 = x111 & n3584 ;
  assign n30982 = ~n30980 & ~n30981 ;
  assign n30983 = ~n30979 & n30982 ;
  assign n30984 = n3592 & n15442 ;
  assign n30985 = n30983 & ~n30984 ;
  assign n30986 = x23 & ~n30985 ;
  assign n30987 = x23 & ~n30986 ;
  assign n30988 = ~n30985 & ~n30986 ;
  assign n30989 = ~n30987 & ~n30988 ;
  assign n30990 = ~n30235 & ~n30486 ;
  assign n30991 = n30989 & n30990 ;
  assign n30992 = ~n30989 & ~n30990 ;
  assign n30993 = ~n30991 & ~n30992 ;
  assign n30994 = ~n30478 & ~n30482 ;
  assign n30995 = x109 & n4531 ;
  assign n30996 = x107 & n4847 ;
  assign n30997 = x108 & n4526 ;
  assign n30998 = ~n30996 & ~n30997 ;
  assign n30999 = ~n30995 & n30998 ;
  assign n31000 = n4534 & n13894 ;
  assign n31001 = n30999 & ~n31000 ;
  assign n31002 = x26 & ~n31001 ;
  assign n31003 = x26 & ~n31002 ;
  assign n31004 = ~n31001 & ~n31002 ;
  assign n31005 = ~n31003 & ~n31004 ;
  assign n31006 = ~n30994 & ~n31005 ;
  assign n31007 = ~n30994 & ~n31006 ;
  assign n31008 = ~n31005 & ~n31006 ;
  assign n31009 = ~n31007 & ~n31008 ;
  assign n31010 = x106 & n5560 ;
  assign n31011 = x104 & n5943 ;
  assign n31012 = x105 & n5555 ;
  assign n31013 = ~n31011 & ~n31012 ;
  assign n31014 = ~n31010 & n31013 ;
  assign n31015 = n5563 & n12181 ;
  assign n31016 = n31014 & ~n31015 ;
  assign n31017 = x29 & ~n31016 ;
  assign n31018 = x29 & ~n31017 ;
  assign n31019 = ~n31016 & ~n31017 ;
  assign n31020 = ~n31018 & ~n31019 ;
  assign n31021 = ~n30250 & ~n30462 ;
  assign n31022 = n31020 & n31021 ;
  assign n31023 = ~n31020 & ~n31021 ;
  assign n31024 = ~n31022 & ~n31023 ;
  assign n31025 = ~n30425 & ~n30439 ;
  assign n31026 = ~n30408 & ~n30422 ;
  assign n31027 = ~n30389 & ~n30402 ;
  assign n31028 = ~n30350 & ~n30364 ;
  assign n31029 = ~n30333 & ~n30347 ;
  assign n31030 = ~n30276 & ~n30290 ;
  assign n31031 = x76 & n22325 ;
  assign n31032 = x74 & n23066 ;
  assign n31033 = x75 & n22320 ;
  assign n31034 = ~n31032 & ~n31033 ;
  assign n31035 = ~n31031 & n31034 ;
  assign n31036 = n1311 & n22328 ;
  assign n31037 = n31035 & ~n31036 ;
  assign n31038 = x59 & ~n31037 ;
  assign n31039 = x59 & ~n31038 ;
  assign n31040 = ~n31037 & ~n31038 ;
  assign n31041 = ~n31039 & ~n31040 ;
  assign n31042 = ~n30266 & ~n30270 ;
  assign n31043 = x69 & n27024 ;
  assign n31044 = x70 & ~n26217 ;
  assign n31045 = ~n31043 & ~n31044 ;
  assign n31046 = x2 & ~x5 ;
  assign n31047 = ~x2 & x5 ;
  assign n31048 = ~n31046 & ~n31047 ;
  assign n31049 = ~n31045 & ~n31048 ;
  assign n31050 = n31045 & n31048 ;
  assign n31051 = ~n31049 & ~n31050 ;
  assign n31052 = n31042 & ~n31051 ;
  assign n31053 = ~n31042 & n31051 ;
  assign n31054 = ~n31052 & ~n31053 ;
  assign n31055 = x73 & n24612 ;
  assign n31056 = x71 & n25390 ;
  assign n31057 = x72 & n24607 ;
  assign n31058 = ~n31056 & ~n31057 ;
  assign n31059 = ~n31055 & n31058 ;
  assign n31060 = n843 & n24615 ;
  assign n31061 = n31059 & ~n31060 ;
  assign n31062 = x62 & ~n31061 ;
  assign n31063 = x62 & ~n31062 ;
  assign n31064 = ~n31061 & ~n31062 ;
  assign n31065 = ~n31063 & ~n31064 ;
  assign n31066 = ~n31054 & n31065 ;
  assign n31067 = n31054 & ~n31065 ;
  assign n31068 = ~n31066 & ~n31067 ;
  assign n31069 = ~n31041 & n31068 ;
  assign n31070 = ~n31041 & ~n31069 ;
  assign n31071 = n31068 & ~n31069 ;
  assign n31072 = ~n31070 & ~n31071 ;
  assign n31073 = ~n31030 & ~n31072 ;
  assign n31074 = ~n31030 & ~n31073 ;
  assign n31075 = ~n31072 & ~n31073 ;
  assign n31076 = ~n31074 & ~n31075 ;
  assign n31077 = x79 & n20143 ;
  assign n31078 = x77 & n20854 ;
  assign n31079 = x78 & n20138 ;
  assign n31080 = ~n31078 & ~n31079 ;
  assign n31081 = ~n31077 & n31080 ;
  assign n31082 = n1817 & n20146 ;
  assign n31083 = n31081 & ~n31082 ;
  assign n31084 = x56 & ~n31083 ;
  assign n31085 = x56 & ~n31084 ;
  assign n31086 = ~n31083 & ~n31084 ;
  assign n31087 = ~n31085 & ~n31086 ;
  assign n31088 = ~n31076 & ~n31087 ;
  assign n31089 = ~n31076 & ~n31088 ;
  assign n31090 = ~n31087 & ~n31088 ;
  assign n31091 = ~n31089 & ~n31090 ;
  assign n31092 = ~n30293 & ~n30307 ;
  assign n31093 = n31091 & n31092 ;
  assign n31094 = ~n31091 & ~n31092 ;
  assign n31095 = ~n31093 & ~n31094 ;
  assign n31096 = x82 & n18025 ;
  assign n31097 = x80 & n18764 ;
  assign n31098 = x81 & n18020 ;
  assign n31099 = ~n31097 & ~n31098 ;
  assign n31100 = ~n31096 & n31099 ;
  assign n31101 = n2584 & n18028 ;
  assign n31102 = n31100 & ~n31101 ;
  assign n31103 = x53 & ~n31102 ;
  assign n31104 = x53 & ~n31103 ;
  assign n31105 = ~n31102 & ~n31103 ;
  assign n31106 = ~n31104 & ~n31105 ;
  assign n31107 = n31095 & ~n31106 ;
  assign n31108 = n31095 & ~n31107 ;
  assign n31109 = ~n31106 & ~n31107 ;
  assign n31110 = ~n31108 & ~n31109 ;
  assign n31111 = ~n30312 & ~n30327 ;
  assign n31112 = n31110 & n31111 ;
  assign n31113 = ~n31110 & ~n31111 ;
  assign n31114 = ~n31112 & ~n31113 ;
  assign n31115 = x85 & n16076 ;
  assign n31116 = x83 & n16756 ;
  assign n31117 = x84 & n16071 ;
  assign n31118 = ~n31116 & ~n31117 ;
  assign n31119 = ~n31115 & n31118 ;
  assign n31120 = n3389 & n16079 ;
  assign n31121 = n31119 & ~n31120 ;
  assign n31122 = x50 & ~n31121 ;
  assign n31123 = x50 & ~n31122 ;
  assign n31124 = ~n31121 & ~n31122 ;
  assign n31125 = ~n31123 & ~n31124 ;
  assign n31126 = n31114 & ~n31125 ;
  assign n31127 = n31114 & ~n31126 ;
  assign n31128 = ~n31125 & ~n31126 ;
  assign n31129 = ~n31127 & ~n31128 ;
  assign n31130 = ~n31029 & n31129 ;
  assign n31131 = n31029 & ~n31129 ;
  assign n31132 = ~n31130 & ~n31131 ;
  assign n31133 = x88 & n14233 ;
  assign n31134 = x86 & n14876 ;
  assign n31135 = x87 & n14228 ;
  assign n31136 = ~n31134 & ~n31135 ;
  assign n31137 = ~n31133 & n31136 ;
  assign n31138 = n4305 & n14236 ;
  assign n31139 = n31137 & ~n31138 ;
  assign n31140 = x47 & ~n31139 ;
  assign n31141 = x47 & ~n31140 ;
  assign n31142 = ~n31139 & ~n31140 ;
  assign n31143 = ~n31141 & ~n31142 ;
  assign n31144 = ~n31132 & ~n31143 ;
  assign n31145 = n31132 & n31143 ;
  assign n31146 = ~n31144 & ~n31145 ;
  assign n31147 = n31028 & ~n31146 ;
  assign n31148 = ~n31028 & n31146 ;
  assign n31149 = ~n31147 & ~n31148 ;
  assign n31150 = x91 & n12506 ;
  assign n31151 = x89 & n13131 ;
  assign n31152 = x90 & n12501 ;
  assign n31153 = ~n31151 & ~n31152 ;
  assign n31154 = ~n31150 & n31153 ;
  assign n31155 = n5336 & n12509 ;
  assign n31156 = n31154 & ~n31155 ;
  assign n31157 = x44 & ~n31156 ;
  assign n31158 = x44 & ~n31157 ;
  assign n31159 = ~n31156 & ~n31157 ;
  assign n31160 = ~n31158 & ~n31159 ;
  assign n31161 = n31149 & ~n31160 ;
  assign n31162 = n31149 & ~n31161 ;
  assign n31163 = ~n31160 & ~n31161 ;
  assign n31164 = ~n31162 & ~n31163 ;
  assign n31165 = ~n30370 & ~n30383 ;
  assign n31166 = n31164 & n31165 ;
  assign n31167 = ~n31164 & ~n31165 ;
  assign n31168 = ~n31166 & ~n31167 ;
  assign n31169 = x94 & n10905 ;
  assign n31170 = x92 & n11466 ;
  assign n31171 = x93 & n10900 ;
  assign n31172 = ~n31170 & ~n31171 ;
  assign n31173 = ~n31169 & n31172 ;
  assign n31174 = n6483 & n10908 ;
  assign n31175 = n31173 & ~n31174 ;
  assign n31176 = x41 & ~n31175 ;
  assign n31177 = x41 & ~n31176 ;
  assign n31178 = ~n31175 & ~n31176 ;
  assign n31179 = ~n31177 & ~n31178 ;
  assign n31180 = n31168 & ~n31179 ;
  assign n31181 = ~n31168 & n31179 ;
  assign n31182 = ~n31027 & ~n31181 ;
  assign n31183 = ~n31180 & n31182 ;
  assign n31184 = ~n31027 & ~n31183 ;
  assign n31185 = ~n31180 & ~n31183 ;
  assign n31186 = ~n31181 & n31185 ;
  assign n31187 = ~n31184 & ~n31186 ;
  assign n31188 = x97 & n9433 ;
  assign n31189 = x95 & n9915 ;
  assign n31190 = x96 & n9428 ;
  assign n31191 = ~n31189 & ~n31190 ;
  assign n31192 = ~n31188 & n31191 ;
  assign n31193 = n7745 & n9436 ;
  assign n31194 = n31192 & ~n31193 ;
  assign n31195 = x38 & ~n31194 ;
  assign n31196 = x38 & ~n31195 ;
  assign n31197 = ~n31194 & ~n31195 ;
  assign n31198 = ~n31196 & ~n31197 ;
  assign n31199 = ~n31187 & ~n31198 ;
  assign n31200 = ~n31187 & ~n31199 ;
  assign n31201 = ~n31198 & ~n31199 ;
  assign n31202 = ~n31200 & ~n31201 ;
  assign n31203 = ~n31026 & n31202 ;
  assign n31204 = n31026 & ~n31202 ;
  assign n31205 = ~n31203 & ~n31204 ;
  assign n31206 = x100 & n8006 ;
  assign n31207 = x98 & n8474 ;
  assign n31208 = x99 & n8001 ;
  assign n31209 = ~n31207 & ~n31208 ;
  assign n31210 = ~n31206 & n31209 ;
  assign n31211 = n8009 & n9115 ;
  assign n31212 = n31210 & ~n31211 ;
  assign n31213 = x35 & ~n31212 ;
  assign n31214 = x35 & ~n31213 ;
  assign n31215 = ~n31212 & ~n31213 ;
  assign n31216 = ~n31214 & ~n31215 ;
  assign n31217 = ~n31205 & ~n31216 ;
  assign n31218 = n31205 & n31216 ;
  assign n31219 = ~n31217 & ~n31218 ;
  assign n31220 = n31025 & ~n31219 ;
  assign n31221 = ~n31025 & n31219 ;
  assign n31222 = ~n31220 & ~n31221 ;
  assign n31223 = x103 & n6725 ;
  assign n31224 = x101 & n7129 ;
  assign n31225 = x102 & n6720 ;
  assign n31226 = ~n31224 & ~n31225 ;
  assign n31227 = ~n31223 & n31226 ;
  assign n31228 = n6728 & n10588 ;
  assign n31229 = n31227 & ~n31228 ;
  assign n31230 = x32 & ~n31229 ;
  assign n31231 = x32 & ~n31230 ;
  assign n31232 = ~n31229 & ~n31230 ;
  assign n31233 = ~n31231 & ~n31232 ;
  assign n31234 = ~n30455 & ~n30458 ;
  assign n31235 = n31233 & n31234 ;
  assign n31236 = ~n31233 & ~n31234 ;
  assign n31237 = ~n31235 & ~n31236 ;
  assign n31238 = n31222 & n31237 ;
  assign n31239 = ~n31222 & ~n31237 ;
  assign n31240 = ~n31238 & ~n31239 ;
  assign n31241 = n31024 & n31240 ;
  assign n31242 = ~n31024 & ~n31240 ;
  assign n31243 = ~n31241 & ~n31242 ;
  assign n31244 = ~n31009 & ~n31243 ;
  assign n31245 = n31009 & n31243 ;
  assign n31246 = ~n31244 & ~n31245 ;
  assign n31247 = n30993 & ~n31246 ;
  assign n31248 = n30993 & ~n31247 ;
  assign n31249 = ~n31246 & ~n31247 ;
  assign n31250 = ~n31248 & ~n31249 ;
  assign n31251 = x115 & n2751 ;
  assign n31252 = x113 & n3020 ;
  assign n31253 = x114 & n2746 ;
  assign n31254 = ~n31252 & ~n31253 ;
  assign n31255 = ~n31251 & n31254 ;
  assign n31256 = n2754 & n17364 ;
  assign n31257 = n31255 & ~n31256 ;
  assign n31258 = x20 & ~n31257 ;
  assign n31259 = x20 & ~n31258 ;
  assign n31260 = ~n31257 & ~n31258 ;
  assign n31261 = ~n31259 & ~n31260 ;
  assign n31262 = ~n30221 & ~n30489 ;
  assign n31263 = ~n30218 & ~n31262 ;
  assign n31264 = ~n31261 & ~n31263 ;
  assign n31265 = n31261 & n31263 ;
  assign n31266 = ~n31264 & ~n31265 ;
  assign n31267 = ~n31250 & n31266 ;
  assign n31268 = ~n31250 & ~n31267 ;
  assign n31269 = n31266 & ~n31267 ;
  assign n31270 = ~n31268 & ~n31269 ;
  assign n31271 = ~n30978 & ~n31270 ;
  assign n31272 = ~n30978 & ~n31271 ;
  assign n31273 = ~n31270 & ~n31271 ;
  assign n31274 = ~n31272 & ~n31273 ;
  assign n31275 = x121 & n1434 ;
  assign n31276 = x119 & n1646 ;
  assign n31277 = x120 & n1429 ;
  assign n31278 = ~n31276 & ~n31277 ;
  assign n31279 = ~n31275 & n31278 ;
  assign n31280 = n1437 & n21870 ;
  assign n31281 = n31279 & ~n31280 ;
  assign n31282 = x14 & ~n31281 ;
  assign n31283 = x14 & ~n31282 ;
  assign n31284 = ~n31281 & ~n31282 ;
  assign n31285 = ~n31283 & ~n31284 ;
  assign n31286 = ~n30189 & ~n30496 ;
  assign n31287 = ~n30186 & ~n31286 ;
  assign n31288 = ~n31285 & ~n31287 ;
  assign n31289 = n31285 & n31287 ;
  assign n31290 = ~n31288 & ~n31289 ;
  assign n31291 = ~n31274 & n31290 ;
  assign n31292 = ~n31274 & ~n31291 ;
  assign n31293 = n31290 & ~n31291 ;
  assign n31294 = ~n31292 & ~n31293 ;
  assign n31295 = n30962 & ~n31294 ;
  assign n31296 = n30962 & ~n31295 ;
  assign n31297 = ~n31294 & ~n31295 ;
  assign n31298 = ~n31296 & ~n31297 ;
  assign n31299 = ~n30947 & n31298 ;
  assign n31300 = n30947 & ~n31298 ;
  assign n31301 = ~n31299 & ~n31300 ;
  assign n31302 = ~n30931 & ~n31301 ;
  assign n31303 = n30931 & n31301 ;
  assign n31304 = ~n31302 & ~n31303 ;
  assign n31305 = ~n30930 & n31304 ;
  assign n31306 = n30930 & ~n31304 ;
  assign n31307 = ~n31305 & ~n31306 ;
  assign n31684 = n31307 & x197 ;
  assign n31308 = ~n30918 & ~n30922 ;
  assign n31309 = ~n30545 & ~n30915 ;
  assign n31310 = ~n30907 & ~n30911 ;
  assign n31311 = ~x127 & n574 ;
  assign n31312 = ~x125 & n673 ;
  assign n31313 = ~x126 & n569 ;
  assign n31314 = ~n31312 & ~n31313 ;
  assign n31315 = ~n31311 & n31314 ;
  assign n31316 = n577 & n26932 ;
  assign n31317 = n31315 & ~n31316 ;
  assign n31318 = ~x8 & ~n31317 ;
  assign n31319 = ~x8 & ~n31318 ;
  assign n31320 = ~n31317 & ~n31318 ;
  assign n31321 = ~n31319 & ~n31320 ;
  assign n31322 = ~n31310 & ~n31321 ;
  assign n31323 = ~n31310 & ~n31322 ;
  assign n31324 = ~n31321 & ~n31322 ;
  assign n31325 = ~n31323 & ~n31324 ;
  assign n31326 = ~x124 & n945 ;
  assign n31327 = ~x122 & n1099 ;
  assign n31328 = ~x123 & n940 ;
  assign n31329 = ~n31327 & ~n31328 ;
  assign n31330 = ~n31326 & n31329 ;
  assign n31331 = n948 & n24176 ;
  assign n31332 = n31330 & ~n31331 ;
  assign n31333 = ~x11 & ~n31332 ;
  assign n31334 = ~x11 & ~n31333 ;
  assign n31335 = ~n31332 & ~n31333 ;
  assign n31336 = ~n31334 & ~n31335 ;
  assign n31337 = ~n30562 & ~n30891 ;
  assign n31338 = n31336 & n31337 ;
  assign n31339 = ~n31336 & ~n31337 ;
  assign n31340 = ~n31338 & ~n31339 ;
  assign n31341 = ~n30593 & ~n30884 ;
  assign n31342 = ~x118 & n2093 ;
  assign n31343 = ~x116 & n2275 ;
  assign n31344 = ~x117 & n2088 ;
  assign n31345 = ~n31343 & ~n31344 ;
  assign n31346 = ~n31342 & n31345 ;
  assign n31347 = n2096 & n19736 ;
  assign n31348 = n31346 & ~n31347 ;
  assign n31349 = ~x17 & ~n31348 ;
  assign n31350 = ~x17 & ~n31349 ;
  assign n31351 = ~n31348 & ~n31349 ;
  assign n31352 = ~n31350 & ~n31351 ;
  assign n31353 = ~n31341 & ~n31352 ;
  assign n31354 = ~n31341 & ~n31353 ;
  assign n31355 = ~n31352 & ~n31353 ;
  assign n31356 = ~n31354 & ~n31355 ;
  assign n31357 = ~x112 & n3589 ;
  assign n31358 = ~x110 & n3878 ;
  assign n31359 = ~x111 & n3584 ;
  assign n31360 = ~n31358 & ~n31359 ;
  assign n31361 = ~n31357 & n31360 ;
  assign n31362 = n3592 & n15744 ;
  assign n31363 = n31361 & ~n31362 ;
  assign n31364 = ~x23 & ~n31363 ;
  assign n31365 = ~x23 & ~n31364 ;
  assign n31366 = ~n31363 & ~n31364 ;
  assign n31367 = ~n31365 & ~n31366 ;
  assign n31368 = ~n30626 & ~n30877 ;
  assign n31369 = n31367 & n31368 ;
  assign n31370 = ~n31367 & ~n31368 ;
  assign n31371 = ~n31369 & ~n31370 ;
  assign n31372 = ~n30869 & ~n30873 ;
  assign n31373 = ~x109 & n4531 ;
  assign n31374 = ~x107 & n4847 ;
  assign n31375 = ~x108 & n4526 ;
  assign n31376 = ~n31374 & ~n31375 ;
  assign n31377 = ~n31373 & n31376 ;
  assign n31378 = n4534 & n14177 ;
  assign n31379 = n31377 & ~n31378 ;
  assign n31380 = ~x26 & ~n31379 ;
  assign n31381 = ~x26 & ~n31380 ;
  assign n31382 = ~n31379 & ~n31380 ;
  assign n31383 = ~n31381 & ~n31382 ;
  assign n31384 = ~n31372 & ~n31383 ;
  assign n31385 = ~n31372 & ~n31384 ;
  assign n31386 = ~n31383 & ~n31384 ;
  assign n31387 = ~n31385 & ~n31386 ;
  assign n31388 = ~x106 & n5560 ;
  assign n31389 = ~x104 & n5943 ;
  assign n31390 = ~x105 & n5555 ;
  assign n31391 = ~n31389 & ~n31390 ;
  assign n31392 = ~n31388 & n31391 ;
  assign n31393 = n5563 & n12447 ;
  assign n31394 = n31392 & ~n31393 ;
  assign n31395 = ~x29 & ~n31394 ;
  assign n31396 = ~x29 & ~n31395 ;
  assign n31397 = ~n31394 & ~n31395 ;
  assign n31398 = ~n31396 & ~n31397 ;
  assign n31399 = ~n30641 & ~n30853 ;
  assign n31400 = n31398 & n31399 ;
  assign n31401 = ~n31398 & ~n31399 ;
  assign n31402 = ~n31400 & ~n31401 ;
  assign n31403 = ~n30816 & ~n30830 ;
  assign n31404 = ~n30799 & ~n30813 ;
  assign n31405 = ~n30780 & ~n30793 ;
  assign n31406 = ~n30741 & ~n30755 ;
  assign n31407 = ~n30724 & ~n30738 ;
  assign n31408 = ~n30667 & ~n30681 ;
  assign n31409 = ~x76 & n22325 ;
  assign n31410 = ~x74 & n23066 ;
  assign n31411 = ~x75 & n22320 ;
  assign n31412 = ~n31410 & ~n31411 ;
  assign n31413 = ~n31409 & n31412 ;
  assign n31414 = n1390 & n22328 ;
  assign n31415 = n31413 & ~n31414 ;
  assign n31416 = ~x59 & ~n31415 ;
  assign n31417 = ~x59 & ~n31416 ;
  assign n31418 = ~n31415 & ~n31416 ;
  assign n31419 = ~n31417 & ~n31418 ;
  assign n31420 = ~n30657 & ~n30661 ;
  assign n31421 = ~x69 & n27427 ;
  assign n31422 = ~x70 & ~n26217 ;
  assign n31423 = ~n31421 & ~n31422 ;
  assign n31424 = ~n31048 & ~n31423 ;
  assign n31425 = n31048 & n31423 ;
  assign n31426 = ~n31424 & ~n31425 ;
  assign n31427 = n31420 & ~n31426 ;
  assign n31428 = ~n31420 & n31426 ;
  assign n31429 = ~n31427 & ~n31428 ;
  assign n31430 = ~x73 & n24612 ;
  assign n31431 = ~x71 & n25390 ;
  assign n31432 = ~x72 & n24607 ;
  assign n31433 = ~n31431 & ~n31432 ;
  assign n31434 = ~n31430 & n31433 ;
  assign n31435 = n903 & n24615 ;
  assign n31436 = n31434 & ~n31435 ;
  assign n31437 = ~x62 & ~n31436 ;
  assign n31438 = ~x62 & ~n31437 ;
  assign n31439 = ~n31436 & ~n31437 ;
  assign n31440 = ~n31438 & ~n31439 ;
  assign n31441 = ~n31429 & n31440 ;
  assign n31442 = n31429 & ~n31440 ;
  assign n31443 = ~n31441 & ~n31442 ;
  assign n31444 = ~n31419 & n31443 ;
  assign n31445 = ~n31419 & ~n31444 ;
  assign n31446 = n31443 & ~n31444 ;
  assign n31447 = ~n31445 & ~n31446 ;
  assign n31448 = ~n31408 & ~n31447 ;
  assign n31449 = ~n31408 & ~n31448 ;
  assign n31450 = ~n31447 & ~n31448 ;
  assign n31451 = ~n31449 & ~n31450 ;
  assign n31452 = ~x79 & n20143 ;
  assign n31453 = ~x77 & n20854 ;
  assign n31454 = ~x78 & n20138 ;
  assign n31455 = ~n31453 & ~n31454 ;
  assign n31456 = ~n31452 & n31455 ;
  assign n31457 = n1921 & n20146 ;
  assign n31458 = n31456 & ~n31457 ;
  assign n31459 = ~x56 & ~n31458 ;
  assign n31460 = ~x56 & ~n31459 ;
  assign n31461 = ~n31458 & ~n31459 ;
  assign n31462 = ~n31460 & ~n31461 ;
  assign n31463 = ~n31451 & ~n31462 ;
  assign n31464 = ~n31451 & ~n31463 ;
  assign n31465 = ~n31462 & ~n31463 ;
  assign n31466 = ~n31464 & ~n31465 ;
  assign n31467 = ~n30684 & ~n30698 ;
  assign n31468 = n31466 & n31467 ;
  assign n31469 = ~n31466 & ~n31467 ;
  assign n31470 = ~n31468 & ~n31469 ;
  assign n31471 = ~x82 & n18025 ;
  assign n31472 = ~x80 & n18764 ;
  assign n31473 = ~x81 & n18020 ;
  assign n31474 = ~n31472 & ~n31473 ;
  assign n31475 = ~n31471 & n31474 ;
  assign n31476 = n2697 & n18028 ;
  assign n31477 = n31475 & ~n31476 ;
  assign n31478 = ~x53 & ~n31477 ;
  assign n31479 = ~x53 & ~n31478 ;
  assign n31480 = ~n31477 & ~n31478 ;
  assign n31481 = ~n31479 & ~n31480 ;
  assign n31482 = n31470 & ~n31481 ;
  assign n31483 = n31470 & ~n31482 ;
  assign n31484 = ~n31481 & ~n31482 ;
  assign n31485 = ~n31483 & ~n31484 ;
  assign n31486 = ~n30703 & ~n30718 ;
  assign n31487 = n31485 & n31486 ;
  assign n31488 = ~n31485 & ~n31486 ;
  assign n31489 = ~n31487 & ~n31488 ;
  assign n31490 = ~x85 & n16076 ;
  assign n31491 = ~x83 & n16756 ;
  assign n31492 = ~x84 & n16071 ;
  assign n31493 = ~n31491 & ~n31492 ;
  assign n31494 = ~n31490 & n31493 ;
  assign n31495 = n3521 & n16079 ;
  assign n31496 = n31494 & ~n31495 ;
  assign n31497 = ~x50 & ~n31496 ;
  assign n31498 = ~x50 & ~n31497 ;
  assign n31499 = ~n31496 & ~n31497 ;
  assign n31500 = ~n31498 & ~n31499 ;
  assign n31501 = n31489 & ~n31500 ;
  assign n31502 = n31489 & ~n31501 ;
  assign n31503 = ~n31500 & ~n31501 ;
  assign n31504 = ~n31502 & ~n31503 ;
  assign n31505 = ~n31407 & n31504 ;
  assign n31506 = n31407 & ~n31504 ;
  assign n31507 = ~n31505 & ~n31506 ;
  assign n31508 = ~x88 & n14233 ;
  assign n31509 = ~x86 & n14876 ;
  assign n31510 = ~x87 & n14228 ;
  assign n31511 = ~n31509 & ~n31510 ;
  assign n31512 = ~n31508 & n31511 ;
  assign n31513 = n4457 & n14236 ;
  assign n31514 = n31512 & ~n31513 ;
  assign n31515 = ~x47 & ~n31514 ;
  assign n31516 = ~x47 & ~n31515 ;
  assign n31517 = ~n31514 & ~n31515 ;
  assign n31518 = ~n31516 & ~n31517 ;
  assign n31519 = ~n31507 & ~n31518 ;
  assign n31520 = n31507 & n31518 ;
  assign n31521 = ~n31519 & ~n31520 ;
  assign n31522 = n31406 & ~n31521 ;
  assign n31523 = ~n31406 & n31521 ;
  assign n31524 = ~n31522 & ~n31523 ;
  assign n31525 = ~x91 & n12506 ;
  assign n31526 = ~x89 & n13131 ;
  assign n31527 = ~x90 & n12501 ;
  assign n31528 = ~n31526 & ~n31527 ;
  assign n31529 = ~n31525 & n31528 ;
  assign n31530 = n5507 & n12509 ;
  assign n31531 = n31529 & ~n31530 ;
  assign n31532 = ~x44 & ~n31531 ;
  assign n31533 = ~x44 & ~n31532 ;
  assign n31534 = ~n31531 & ~n31532 ;
  assign n31535 = ~n31533 & ~n31534 ;
  assign n31536 = n31524 & ~n31535 ;
  assign n31537 = n31524 & ~n31536 ;
  assign n31538 = ~n31535 & ~n31536 ;
  assign n31539 = ~n31537 & ~n31538 ;
  assign n31540 = ~n30761 & ~n30774 ;
  assign n31541 = n31539 & n31540 ;
  assign n31542 = ~n31539 & ~n31540 ;
  assign n31543 = ~n31541 & ~n31542 ;
  assign n31544 = ~x94 & n10905 ;
  assign n31545 = ~x92 & n11466 ;
  assign n31546 = ~x93 & n10900 ;
  assign n31547 = ~n31545 & ~n31546 ;
  assign n31548 = ~n31544 & n31547 ;
  assign n31549 = n6671 & n10908 ;
  assign n31550 = n31548 & ~n31549 ;
  assign n31551 = ~x41 & ~n31550 ;
  assign n31552 = ~x41 & ~n31551 ;
  assign n31553 = ~n31550 & ~n31551 ;
  assign n31554 = ~n31552 & ~n31553 ;
  assign n31555 = n31543 & ~n31554 ;
  assign n31556 = ~n31543 & n31554 ;
  assign n31557 = ~n31405 & ~n31556 ;
  assign n31558 = ~n31555 & n31557 ;
  assign n31559 = ~n31405 & ~n31558 ;
  assign n31560 = ~n31555 & ~n31558 ;
  assign n31561 = ~n31556 & n31560 ;
  assign n31562 = ~n31559 & ~n31561 ;
  assign n31563 = ~x97 & n9433 ;
  assign n31564 = ~x95 & n9915 ;
  assign n31565 = ~x96 & n9428 ;
  assign n31566 = ~n31564 & ~n31565 ;
  assign n31567 = ~n31563 & n31566 ;
  assign n31568 = n7949 & n9436 ;
  assign n31569 = n31567 & ~n31568 ;
  assign n31570 = ~x38 & ~n31569 ;
  assign n31571 = ~x38 & ~n31570 ;
  assign n31572 = ~n31569 & ~n31570 ;
  assign n31573 = ~n31571 & ~n31572 ;
  assign n31574 = ~n31562 & ~n31573 ;
  assign n31575 = ~n31562 & ~n31574 ;
  assign n31576 = ~n31573 & ~n31574 ;
  assign n31577 = ~n31575 & ~n31576 ;
  assign n31578 = ~n31404 & n31577 ;
  assign n31579 = n31404 & ~n31577 ;
  assign n31580 = ~n31578 & ~n31579 ;
  assign n31581 = ~x100 & n8006 ;
  assign n31582 = ~x98 & n8474 ;
  assign n31583 = ~x99 & n8001 ;
  assign n31584 = ~n31582 & ~n31583 ;
  assign n31585 = ~n31581 & n31584 ;
  assign n31586 = n8009 & n9338 ;
  assign n31587 = n31585 & ~n31586 ;
  assign n31588 = ~x35 & ~n31587 ;
  assign n31589 = ~x35 & ~n31588 ;
  assign n31590 = ~n31587 & ~n31588 ;
  assign n31591 = ~n31589 & ~n31590 ;
  assign n31592 = ~n31580 & ~n31591 ;
  assign n31593 = n31580 & n31591 ;
  assign n31594 = ~n31592 & ~n31593 ;
  assign n31595 = n31403 & ~n31594 ;
  assign n31596 = ~n31403 & n31594 ;
  assign n31597 = ~n31595 & ~n31596 ;
  assign n31598 = ~x103 & n6725 ;
  assign n31599 = ~x101 & n7129 ;
  assign n31600 = ~x102 & n6720 ;
  assign n31601 = ~n31599 & ~n31600 ;
  assign n31602 = ~n31598 & n31601 ;
  assign n31603 = n6728 & n10833 ;
  assign n31604 = n31602 & ~n31603 ;
  assign n31605 = ~x32 & ~n31604 ;
  assign n31606 = ~x32 & ~n31605 ;
  assign n31607 = ~n31604 & ~n31605 ;
  assign n31608 = ~n31606 & ~n31607 ;
  assign n31609 = ~n30846 & ~n30849 ;
  assign n31610 = n31608 & n31609 ;
  assign n31611 = ~n31608 & ~n31609 ;
  assign n31612 = ~n31610 & ~n31611 ;
  assign n31613 = n31597 & n31612 ;
  assign n31614 = ~n31597 & ~n31612 ;
  assign n31615 = ~n31613 & ~n31614 ;
  assign n31616 = n31402 & n31615 ;
  assign n31617 = ~n31402 & ~n31615 ;
  assign n31618 = ~n31616 & ~n31617 ;
  assign n31619 = ~n31387 & ~n31618 ;
  assign n31620 = n31387 & n31618 ;
  assign n31621 = ~n31619 & ~n31620 ;
  assign n31622 = n31371 & ~n31621 ;
  assign n31623 = n31371 & ~n31622 ;
  assign n31624 = ~n31621 & ~n31622 ;
  assign n31625 = ~n31623 & ~n31624 ;
  assign n31626 = ~x115 & n2751 ;
  assign n31627 = ~x113 & n3020 ;
  assign n31628 = ~x114 & n2746 ;
  assign n31629 = ~n31627 & ~n31628 ;
  assign n31630 = ~n31626 & n31629 ;
  assign n31631 = n2754 & n17683 ;
  assign n31632 = n31630 & ~n31631 ;
  assign n31633 = ~x20 & ~n31632 ;
  assign n31634 = ~x20 & ~n31633 ;
  assign n31635 = ~n31632 & ~n31633 ;
  assign n31636 = ~n31634 & ~n31635 ;
  assign n31637 = ~n30612 & ~n30880 ;
  assign n31638 = ~n30609 & ~n31637 ;
  assign n31639 = ~n31636 & ~n31638 ;
  assign n31640 = n31636 & n31638 ;
  assign n31641 = ~n31639 & ~n31640 ;
  assign n31642 = ~n31625 & n31641 ;
  assign n31643 = ~n31625 & ~n31642 ;
  assign n31644 = n31641 & ~n31642 ;
  assign n31645 = ~n31643 & ~n31644 ;
  assign n31646 = ~n31356 & ~n31645 ;
  assign n31647 = ~n31356 & ~n31646 ;
  assign n31648 = ~n31645 & ~n31646 ;
  assign n31649 = ~n31647 & ~n31648 ;
  assign n31650 = ~x121 & n1434 ;
  assign n31651 = ~x119 & n1646 ;
  assign n31652 = ~x120 & n1429 ;
  assign n31653 = ~n31651 & ~n31652 ;
  assign n31654 = ~n31650 & n31653 ;
  assign n31655 = n1437 & n22229 ;
  assign n31656 = n31654 & ~n31655 ;
  assign n31657 = ~x14 & ~n31656 ;
  assign n31658 = ~x14 & ~n31657 ;
  assign n31659 = ~n31656 & ~n31657 ;
  assign n31660 = ~n31658 & ~n31659 ;
  assign n31661 = ~n30580 & ~n30887 ;
  assign n31662 = ~n30577 & ~n31661 ;
  assign n31663 = ~n31660 & ~n31662 ;
  assign n31664 = n31660 & n31662 ;
  assign n31665 = ~n31663 & ~n31664 ;
  assign n31666 = ~n31649 & n31665 ;
  assign n31667 = ~n31649 & ~n31666 ;
  assign n31668 = n31665 & ~n31666 ;
  assign n31669 = ~n31667 & ~n31668 ;
  assign n31670 = n31340 & ~n31669 ;
  assign n31671 = n31340 & ~n31670 ;
  assign n31672 = ~n31669 & ~n31670 ;
  assign n31673 = ~n31671 & ~n31672 ;
  assign n31674 = ~n31325 & n31673 ;
  assign n31675 = n31325 & ~n31673 ;
  assign n31676 = ~n31674 & ~n31675 ;
  assign n31677 = ~n31309 & ~n31676 ;
  assign n31678 = n31309 & n31676 ;
  assign n31679 = ~n31677 & ~n31678 ;
  assign n31680 = ~n31308 & n31679 ;
  assign n31681 = n31308 & ~n31679 ;
  assign n31682 = ~n31680 & ~n31681 ;
  assign n31685 = ~n31682 & ~x197 ;
  assign n31686 = ~n31684 & ~n31685 ;
  assign n31687 = ~n30961 & ~n31295 ;
  assign n31688 = x126 & n673 ;
  assign n31689 = x127 & n569 ;
  assign n31690 = ~n31688 & ~n31689 ;
  assign n31691 = ~n577 & n31690 ;
  assign n31692 = n26965 & n31690 ;
  assign n31693 = ~n31691 & ~n31692 ;
  assign n31694 = x8 & ~n31693 ;
  assign n31695 = ~x8 & n31693 ;
  assign n31696 = ~n31694 & ~n31695 ;
  assign n31697 = ~n31687 & ~n31696 ;
  assign n31698 = n31687 & n31696 ;
  assign n31699 = ~n31697 & ~n31698 ;
  assign n31700 = x125 & n945 ;
  assign n31701 = x123 & n1099 ;
  assign n31702 = x124 & n940 ;
  assign n31703 = ~n31701 & ~n31702 ;
  assign n31704 = ~n31700 & n31703 ;
  assign n31705 = n948 & n24935 ;
  assign n31706 = n31704 & ~n31705 ;
  assign n31707 = x11 & ~n31706 ;
  assign n31708 = x11 & ~n31707 ;
  assign n31709 = ~n31706 & ~n31707 ;
  assign n31710 = ~n31708 & ~n31709 ;
  assign n31711 = ~n31288 & ~n31291 ;
  assign n31712 = n31710 & n31711 ;
  assign n31713 = ~n31710 & ~n31711 ;
  assign n31714 = ~n31712 & ~n31713 ;
  assign n31715 = ~n30975 & ~n31271 ;
  assign n31716 = x122 & n1434 ;
  assign n31717 = x120 & n1646 ;
  assign n31718 = x121 & n1429 ;
  assign n31719 = ~n31717 & ~n31718 ;
  assign n31720 = ~n31716 & n31719 ;
  assign n31721 = ~n1437 & n31720 ;
  assign n31722 = ~n22622 & n31720 ;
  assign n31723 = ~n31721 & ~n31722 ;
  assign n31724 = x14 & ~n31723 ;
  assign n31725 = ~x14 & n31723 ;
  assign n31726 = ~n31724 & ~n31725 ;
  assign n31727 = ~n31715 & ~n31726 ;
  assign n31728 = n31715 & n31726 ;
  assign n31729 = ~n31727 & ~n31728 ;
  assign n31730 = x119 & n2093 ;
  assign n31731 = x117 & n2275 ;
  assign n31732 = x118 & n2088 ;
  assign n31733 = ~n31731 & ~n31732 ;
  assign n31734 = ~n31730 & n31733 ;
  assign n31735 = n2096 & n20423 ;
  assign n31736 = n31734 & ~n31735 ;
  assign n31737 = x17 & ~n31736 ;
  assign n31738 = x17 & ~n31737 ;
  assign n31739 = ~n31736 & ~n31737 ;
  assign n31740 = ~n31738 & ~n31739 ;
  assign n31741 = ~n31264 & ~n31267 ;
  assign n31742 = n31740 & n31741 ;
  assign n31743 = ~n31740 & ~n31741 ;
  assign n31744 = ~n31742 & ~n31743 ;
  assign n31745 = x116 & n2751 ;
  assign n31746 = x114 & n3020 ;
  assign n31747 = x115 & n2746 ;
  assign n31748 = ~n31746 & ~n31747 ;
  assign n31749 = ~n31745 & n31748 ;
  assign n31750 = n2754 & n18336 ;
  assign n31751 = n31749 & ~n31750 ;
  assign n31752 = x20 & ~n31751 ;
  assign n31753 = x20 & ~n31752 ;
  assign n31754 = ~n31751 & ~n31752 ;
  assign n31755 = ~n31753 & ~n31754 ;
  assign n31756 = ~n30992 & ~n31247 ;
  assign n31757 = n31755 & n31756 ;
  assign n31758 = ~n31755 & ~n31756 ;
  assign n31759 = ~n31757 & ~n31758 ;
  assign n31760 = x113 & n3589 ;
  assign n31761 = x111 & n3878 ;
  assign n31762 = x112 & n3584 ;
  assign n31763 = ~n31761 & ~n31762 ;
  assign n31764 = ~n31760 & n31763 ;
  assign n31765 = n3592 & n16361 ;
  assign n31766 = n31764 & ~n31765 ;
  assign n31767 = x23 & ~n31766 ;
  assign n31768 = x23 & ~n31767 ;
  assign n31769 = ~n31766 & ~n31767 ;
  assign n31770 = ~n31768 & ~n31769 ;
  assign n31771 = ~n31009 & n31243 ;
  assign n31772 = ~n31006 & ~n31771 ;
  assign n31773 = ~n31770 & ~n31772 ;
  assign n31774 = ~n31770 & ~n31773 ;
  assign n31775 = ~n31772 & ~n31773 ;
  assign n31776 = ~n31774 & ~n31775 ;
  assign n31777 = ~n31023 & ~n31241 ;
  assign n31778 = x110 & n4531 ;
  assign n31779 = x108 & n4847 ;
  assign n31780 = x109 & n4526 ;
  assign n31781 = ~n31779 & ~n31780 ;
  assign n31782 = ~n31778 & n31781 ;
  assign n31783 = ~n4534 & n31782 ;
  assign n31784 = ~n14497 & n31782 ;
  assign n31785 = ~n31783 & ~n31784 ;
  assign n31786 = x26 & ~n31785 ;
  assign n31787 = ~x26 & n31785 ;
  assign n31788 = ~n31786 & ~n31787 ;
  assign n31789 = ~n31777 & ~n31788 ;
  assign n31790 = n31777 & n31788 ;
  assign n31791 = ~n31789 & ~n31790 ;
  assign n31792 = x107 & n5560 ;
  assign n31793 = x105 & n5943 ;
  assign n31794 = x106 & n5555 ;
  assign n31795 = ~n31793 & ~n31794 ;
  assign n31796 = ~n31792 & n31795 ;
  assign n31797 = n5563 & n12749 ;
  assign n31798 = n31796 & ~n31797 ;
  assign n31799 = x29 & ~n31798 ;
  assign n31800 = x29 & ~n31799 ;
  assign n31801 = ~n31798 & ~n31799 ;
  assign n31802 = ~n31800 & ~n31801 ;
  assign n31803 = ~n31236 & ~n31238 ;
  assign n31804 = ~n31802 & ~n31803 ;
  assign n31805 = ~n31802 & ~n31804 ;
  assign n31806 = ~n31803 & ~n31804 ;
  assign n31807 = ~n31805 & ~n31806 ;
  assign n31808 = x104 & n6725 ;
  assign n31809 = x102 & n7129 ;
  assign n31810 = x103 & n6720 ;
  assign n31811 = ~n31809 & ~n31810 ;
  assign n31812 = ~n31808 & n31811 ;
  assign n31813 = n6728 & n11116 ;
  assign n31814 = n31812 & ~n31813 ;
  assign n31815 = x32 & ~n31814 ;
  assign n31816 = x32 & ~n31815 ;
  assign n31817 = ~n31814 & ~n31815 ;
  assign n31818 = ~n31816 & ~n31817 ;
  assign n31819 = ~n31217 & ~n31221 ;
  assign n31820 = n31818 & n31819 ;
  assign n31821 = ~n31818 & ~n31819 ;
  assign n31822 = ~n31820 & ~n31821 ;
  assign n31823 = x101 & n8006 ;
  assign n31824 = x99 & n8474 ;
  assign n31825 = x100 & n8001 ;
  assign n31826 = ~n31824 & ~n31825 ;
  assign n31827 = ~n31823 & n31826 ;
  assign n31828 = n8009 & n9601 ;
  assign n31829 = n31827 & ~n31828 ;
  assign n31830 = x35 & ~n31829 ;
  assign n31831 = x35 & ~n31830 ;
  assign n31832 = ~n31829 & ~n31830 ;
  assign n31833 = ~n31831 & ~n31832 ;
  assign n31834 = ~n31026 & ~n31202 ;
  assign n31835 = ~n31199 & ~n31834 ;
  assign n31836 = x98 & n9433 ;
  assign n31837 = x96 & n9915 ;
  assign n31838 = x97 & n9428 ;
  assign n31839 = ~n31837 & ~n31838 ;
  assign n31840 = ~n31836 & n31839 ;
  assign n31841 = n8196 & n9436 ;
  assign n31842 = n31840 & ~n31841 ;
  assign n31843 = x38 & ~n31842 ;
  assign n31844 = x38 & ~n31843 ;
  assign n31845 = ~n31842 & ~n31843 ;
  assign n31846 = ~n31844 & ~n31845 ;
  assign n31847 = ~n31053 & ~n31067 ;
  assign n31848 = ~x2 & ~x5 ;
  assign n31849 = ~n31049 & ~n31848 ;
  assign n31850 = x70 & n27024 ;
  assign n31851 = x71 & ~n26217 ;
  assign n31852 = ~n31850 & ~n31851 ;
  assign n31853 = ~n31849 & n31852 ;
  assign n31854 = n31849 & ~n31852 ;
  assign n31855 = ~n31853 & ~n31854 ;
  assign n31856 = x74 & n24612 ;
  assign n31857 = x72 & n25390 ;
  assign n31858 = x73 & n24607 ;
  assign n31859 = ~n31857 & ~n31858 ;
  assign n31860 = ~n31856 & n31859 ;
  assign n31861 = ~n24615 & n31860 ;
  assign n31862 = ~n994 & n31860 ;
  assign n31863 = ~n31861 & ~n31862 ;
  assign n31864 = x62 & ~n31863 ;
  assign n31865 = ~x62 & n31863 ;
  assign n31866 = ~n31864 & ~n31865 ;
  assign n31867 = n31855 & ~n31866 ;
  assign n31868 = ~n31855 & n31866 ;
  assign n31869 = ~n31867 & ~n31868 ;
  assign n31870 = ~n31847 & n31869 ;
  assign n31871 = n31847 & ~n31869 ;
  assign n31872 = ~n31870 & ~n31871 ;
  assign n31873 = x77 & n22325 ;
  assign n31874 = x75 & n23066 ;
  assign n31875 = x76 & n22320 ;
  assign n31876 = ~n31874 & ~n31875 ;
  assign n31877 = ~n31873 & n31876 ;
  assign n31878 = n1502 & n22328 ;
  assign n31879 = n31877 & ~n31878 ;
  assign n31880 = x59 & ~n31879 ;
  assign n31881 = x59 & ~n31880 ;
  assign n31882 = ~n31879 & ~n31880 ;
  assign n31883 = ~n31881 & ~n31882 ;
  assign n31884 = n31872 & ~n31883 ;
  assign n31885 = n31872 & ~n31884 ;
  assign n31886 = ~n31883 & ~n31884 ;
  assign n31887 = ~n31885 & ~n31886 ;
  assign n31888 = ~n31069 & ~n31073 ;
  assign n31889 = n31887 & n31888 ;
  assign n31890 = ~n31887 & ~n31888 ;
  assign n31891 = ~n31889 & ~n31890 ;
  assign n31892 = x80 & n20143 ;
  assign n31893 = x78 & n20854 ;
  assign n31894 = x79 & n20138 ;
  assign n31895 = ~n31893 & ~n31894 ;
  assign n31896 = ~n31892 & n31895 ;
  assign n31897 = n2028 & n20146 ;
  assign n31898 = n31896 & ~n31897 ;
  assign n31899 = x56 & ~n31898 ;
  assign n31900 = x56 & ~n31899 ;
  assign n31901 = ~n31898 & ~n31899 ;
  assign n31902 = ~n31900 & ~n31901 ;
  assign n31903 = n31891 & ~n31902 ;
  assign n31904 = n31891 & ~n31903 ;
  assign n31905 = ~n31902 & ~n31903 ;
  assign n31906 = ~n31904 & ~n31905 ;
  assign n31907 = ~n31088 & ~n31094 ;
  assign n31908 = n31906 & n31907 ;
  assign n31909 = ~n31906 & ~n31907 ;
  assign n31910 = ~n31908 & ~n31909 ;
  assign n31911 = x83 & n18025 ;
  assign n31912 = x81 & n18764 ;
  assign n31913 = x82 & n18020 ;
  assign n31914 = ~n31912 & ~n31913 ;
  assign n31915 = ~n31911 & n31914 ;
  assign n31916 = n2843 & n18028 ;
  assign n31917 = n31915 & ~n31916 ;
  assign n31918 = x53 & ~n31917 ;
  assign n31919 = x53 & ~n31918 ;
  assign n31920 = ~n31917 & ~n31918 ;
  assign n31921 = ~n31919 & ~n31920 ;
  assign n31922 = n31910 & ~n31921 ;
  assign n31923 = n31910 & ~n31922 ;
  assign n31924 = ~n31921 & ~n31922 ;
  assign n31925 = ~n31923 & ~n31924 ;
  assign n31926 = ~n31107 & ~n31113 ;
  assign n31927 = n31925 & n31926 ;
  assign n31928 = ~n31925 & ~n31926 ;
  assign n31929 = ~n31927 & ~n31928 ;
  assign n31930 = x86 & n16076 ;
  assign n31931 = x84 & n16756 ;
  assign n31932 = x85 & n16071 ;
  assign n31933 = ~n31931 & ~n31932 ;
  assign n31934 = ~n31930 & n31933 ;
  assign n31935 = n3686 & n16079 ;
  assign n31936 = n31934 & ~n31935 ;
  assign n31937 = x50 & ~n31936 ;
  assign n31938 = x50 & ~n31937 ;
  assign n31939 = ~n31936 & ~n31937 ;
  assign n31940 = ~n31938 & ~n31939 ;
  assign n31941 = n31929 & ~n31940 ;
  assign n31942 = n31929 & ~n31941 ;
  assign n31943 = ~n31940 & ~n31941 ;
  assign n31944 = ~n31942 & ~n31943 ;
  assign n31945 = ~n31029 & ~n31129 ;
  assign n31946 = ~n31126 & ~n31945 ;
  assign n31947 = n31944 & n31946 ;
  assign n31948 = ~n31944 & ~n31946 ;
  assign n31949 = ~n31947 & ~n31948 ;
  assign n31950 = x89 & n14233 ;
  assign n31951 = x87 & n14876 ;
  assign n31952 = x88 & n14228 ;
  assign n31953 = ~n31951 & ~n31952 ;
  assign n31954 = ~n31950 & n31953 ;
  assign n31955 = n4488 & n14236 ;
  assign n31956 = n31954 & ~n31955 ;
  assign n31957 = x47 & ~n31956 ;
  assign n31958 = x47 & ~n31957 ;
  assign n31959 = ~n31956 & ~n31957 ;
  assign n31960 = ~n31958 & ~n31959 ;
  assign n31961 = n31949 & ~n31960 ;
  assign n31962 = n31949 & ~n31961 ;
  assign n31963 = ~n31960 & ~n31961 ;
  assign n31964 = ~n31962 & ~n31963 ;
  assign n31965 = ~n31144 & ~n31148 ;
  assign n31966 = n31964 & n31965 ;
  assign n31967 = ~n31964 & ~n31965 ;
  assign n31968 = ~n31966 & ~n31967 ;
  assign n31969 = x92 & n12506 ;
  assign n31970 = x90 & n13131 ;
  assign n31971 = x91 & n12501 ;
  assign n31972 = ~n31970 & ~n31971 ;
  assign n31973 = ~n31969 & n31972 ;
  assign n31974 = n5710 & n12509 ;
  assign n31975 = n31973 & ~n31974 ;
  assign n31976 = x44 & ~n31975 ;
  assign n31977 = x44 & ~n31976 ;
  assign n31978 = ~n31975 & ~n31976 ;
  assign n31979 = ~n31977 & ~n31978 ;
  assign n31980 = n31968 & ~n31979 ;
  assign n31981 = n31968 & ~n31980 ;
  assign n31982 = ~n31979 & ~n31980 ;
  assign n31983 = ~n31981 & ~n31982 ;
  assign n31984 = ~n31161 & ~n31167 ;
  assign n31985 = n31983 & n31984 ;
  assign n31986 = ~n31983 & ~n31984 ;
  assign n31987 = ~n31985 & ~n31986 ;
  assign n31988 = x95 & n10905 ;
  assign n31989 = x93 & n11466 ;
  assign n31990 = x94 & n10900 ;
  assign n31991 = ~n31989 & ~n31990 ;
  assign n31992 = ~n31988 & n31991 ;
  assign n31993 = n6894 & n10908 ;
  assign n31994 = n31992 & ~n31993 ;
  assign n31995 = x41 & ~n31994 ;
  assign n31996 = x41 & ~n31995 ;
  assign n31997 = ~n31994 & ~n31995 ;
  assign n31998 = ~n31996 & ~n31997 ;
  assign n31999 = ~n31987 & n31998 ;
  assign n32000 = n31987 & ~n31998 ;
  assign n32001 = ~n31999 & ~n32000 ;
  assign n32002 = ~n31185 & n32001 ;
  assign n32003 = n31185 & ~n32001 ;
  assign n32004 = ~n32002 & ~n32003 ;
  assign n32005 = ~n31846 & n32004 ;
  assign n32006 = n31846 & ~n32004 ;
  assign n32007 = ~n32005 & ~n32006 ;
  assign n32008 = ~n31835 & n32007 ;
  assign n32009 = n31835 & ~n32007 ;
  assign n32010 = ~n32008 & ~n32009 ;
  assign n32011 = ~n31833 & n32010 ;
  assign n32012 = ~n31833 & ~n32011 ;
  assign n32013 = n32010 & ~n32011 ;
  assign n32014 = ~n32012 & ~n32013 ;
  assign n32015 = n31822 & ~n32014 ;
  assign n32016 = n31822 & ~n32015 ;
  assign n32017 = ~n32014 & ~n32015 ;
  assign n32018 = ~n32016 & ~n32017 ;
  assign n32019 = ~n31807 & n32018 ;
  assign n32020 = n31807 & ~n32018 ;
  assign n32021 = ~n32019 & ~n32020 ;
  assign n32022 = n31791 & ~n32021 ;
  assign n32023 = n31791 & ~n32022 ;
  assign n32024 = ~n32021 & ~n32022 ;
  assign n32025 = ~n32023 & ~n32024 ;
  assign n32026 = ~n31776 & n32025 ;
  assign n32027 = n31776 & ~n32025 ;
  assign n32028 = ~n32026 & ~n32027 ;
  assign n32029 = n31759 & ~n32028 ;
  assign n32030 = n31759 & ~n32029 ;
  assign n32031 = ~n32028 & ~n32029 ;
  assign n32032 = ~n32030 & ~n32031 ;
  assign n32033 = n31744 & ~n32032 ;
  assign n32034 = ~n31744 & n32032 ;
  assign n32035 = n31729 & ~n32034 ;
  assign n32036 = ~n32033 & n32035 ;
  assign n32037 = n31729 & ~n32036 ;
  assign n32038 = ~n32034 & ~n32036 ;
  assign n32039 = ~n32033 & n32038 ;
  assign n32040 = ~n32037 & ~n32039 ;
  assign n32041 = n31714 & ~n32040 ;
  assign n32042 = ~n31714 & n32040 ;
  assign n32043 = n31699 & ~n32042 ;
  assign n32044 = ~n32041 & n32043 ;
  assign n32045 = n31699 & ~n32044 ;
  assign n32046 = ~n32042 & ~n32044 ;
  assign n32047 = ~n32041 & n32046 ;
  assign n32048 = ~n32045 & ~n32047 ;
  assign n32049 = ~n30947 & ~n31298 ;
  assign n32050 = ~n30944 & ~n32049 ;
  assign n32051 = ~n32048 & ~n32050 ;
  assign n32052 = ~n32048 & ~n32051 ;
  assign n32053 = ~n32050 & ~n32051 ;
  assign n32054 = ~n32052 & ~n32053 ;
  assign n32055 = ~n31302 & ~n31305 ;
  assign n32056 = ~n32054 & ~n32055 ;
  assign n32057 = n32054 & n32055 ;
  assign n32058 = ~n32056 & ~n32057 ;
  assign n32432 = n32058 & x198 ;
  assign n32059 = ~n31339 & ~n31670 ;
  assign n32060 = ~x126 & n673 ;
  assign n32061 = ~x127 & n569 ;
  assign n32062 = ~n32060 & ~n32061 ;
  assign n32063 = ~n577 & n32062 ;
  assign n32064 = n27368 & n32062 ;
  assign n32065 = ~n32063 & ~n32064 ;
  assign n32066 = ~x8 & ~n32065 ;
  assign n32067 = x8 & n32065 ;
  assign n32068 = ~n32066 & ~n32067 ;
  assign n32069 = ~n32059 & ~n32068 ;
  assign n32070 = n32059 & n32068 ;
  assign n32071 = ~n32069 & ~n32070 ;
  assign n32072 = ~x125 & n945 ;
  assign n32073 = ~x123 & n1099 ;
  assign n32074 = ~x124 & n940 ;
  assign n32075 = ~n32073 & ~n32074 ;
  assign n32076 = ~n32072 & n32075 ;
  assign n32077 = n948 & n25330 ;
  assign n32078 = n32076 & ~n32077 ;
  assign n32079 = ~x11 & ~n32078 ;
  assign n32080 = ~x11 & ~n32079 ;
  assign n32081 = ~n32078 & ~n32079 ;
  assign n32082 = ~n32080 & ~n32081 ;
  assign n32083 = ~n31663 & ~n31666 ;
  assign n32084 = n32082 & n32083 ;
  assign n32085 = ~n32082 & ~n32083 ;
  assign n32086 = ~n32084 & ~n32085 ;
  assign n32087 = ~n31353 & ~n31646 ;
  assign n32088 = ~x122 & n1434 ;
  assign n32089 = ~x120 & n1646 ;
  assign n32090 = ~x121 & n1429 ;
  assign n32091 = ~n32089 & ~n32090 ;
  assign n32092 = ~n32088 & n32091 ;
  assign n32093 = ~n1437 & n32092 ;
  assign n32094 = ~n22998 & n32092 ;
  assign n32095 = ~n32093 & ~n32094 ;
  assign n32096 = ~x14 & ~n32095 ;
  assign n32097 = x14 & n32095 ;
  assign n32098 = ~n32096 & ~n32097 ;
  assign n32099 = ~n32087 & ~n32098 ;
  assign n32100 = n32087 & n32098 ;
  assign n32101 = ~n32099 & ~n32100 ;
  assign n32102 = ~x119 & n2093 ;
  assign n32103 = ~x117 & n2275 ;
  assign n32104 = ~x118 & n2088 ;
  assign n32105 = ~n32103 & ~n32104 ;
  assign n32106 = ~n32102 & n32105 ;
  assign n32107 = n2096 & n20778 ;
  assign n32108 = n32106 & ~n32107 ;
  assign n32109 = ~x17 & ~n32108 ;
  assign n32110 = ~x17 & ~n32109 ;
  assign n32111 = ~n32108 & ~n32109 ;
  assign n32112 = ~n32110 & ~n32111 ;
  assign n32113 = ~n31639 & ~n31642 ;
  assign n32114 = n32112 & n32113 ;
  assign n32115 = ~n32112 & ~n32113 ;
  assign n32116 = ~n32114 & ~n32115 ;
  assign n32117 = ~x116 & n2751 ;
  assign n32118 = ~x114 & n3020 ;
  assign n32119 = ~x115 & n2746 ;
  assign n32120 = ~n32118 & ~n32119 ;
  assign n32121 = ~n32117 & n32120 ;
  assign n32122 = n2754 & n18678 ;
  assign n32123 = n32121 & ~n32122 ;
  assign n32124 = ~x20 & ~n32123 ;
  assign n32125 = ~x20 & ~n32124 ;
  assign n32126 = ~n32123 & ~n32124 ;
  assign n32127 = ~n32125 & ~n32126 ;
  assign n32128 = ~n31370 & ~n31622 ;
  assign n32129 = n32127 & n32128 ;
  assign n32130 = ~n32127 & ~n32128 ;
  assign n32131 = ~n32129 & ~n32130 ;
  assign n32132 = ~x113 & n3589 ;
  assign n32133 = ~x111 & n3878 ;
  assign n32134 = ~x112 & n3584 ;
  assign n32135 = ~n32133 & ~n32134 ;
  assign n32136 = ~n32132 & n32135 ;
  assign n32137 = n3592 & n16684 ;
  assign n32138 = n32136 & ~n32137 ;
  assign n32139 = ~x23 & ~n32138 ;
  assign n32140 = ~x23 & ~n32139 ;
  assign n32141 = ~n32138 & ~n32139 ;
  assign n32142 = ~n32140 & ~n32141 ;
  assign n32143 = ~n31387 & n31618 ;
  assign n32144 = ~n31384 & ~n32143 ;
  assign n32145 = ~n32142 & ~n32144 ;
  assign n32146 = ~n32142 & ~n32145 ;
  assign n32147 = ~n32144 & ~n32145 ;
  assign n32148 = ~n32146 & ~n32147 ;
  assign n32149 = ~n31401 & ~n31616 ;
  assign n32150 = ~x110 & n4531 ;
  assign n32151 = ~x108 & n4847 ;
  assign n32152 = ~x109 & n4526 ;
  assign n32153 = ~n32151 & ~n32152 ;
  assign n32154 = ~n32150 & n32153 ;
  assign n32155 = ~n4534 & n32154 ;
  assign n32156 = ~n14802 & n32154 ;
  assign n32157 = ~n32155 & ~n32156 ;
  assign n32158 = ~x26 & ~n32157 ;
  assign n32159 = x26 & n32157 ;
  assign n32160 = ~n32158 & ~n32159 ;
  assign n32161 = ~n32149 & ~n32160 ;
  assign n32162 = n32149 & n32160 ;
  assign n32163 = ~n32161 & ~n32162 ;
  assign n32164 = ~x107 & n5560 ;
  assign n32165 = ~x105 & n5943 ;
  assign n32166 = ~x106 & n5555 ;
  assign n32167 = ~n32165 & ~n32166 ;
  assign n32168 = ~n32164 & n32167 ;
  assign n32169 = n5563 & n13034 ;
  assign n32170 = n32168 & ~n32169 ;
  assign n32171 = ~x29 & ~n32170 ;
  assign n32172 = ~x29 & ~n32171 ;
  assign n32173 = ~n32170 & ~n32171 ;
  assign n32174 = ~n32172 & ~n32173 ;
  assign n32175 = ~n31611 & ~n31613 ;
  assign n32176 = ~n32174 & ~n32175 ;
  assign n32177 = ~n32174 & ~n32176 ;
  assign n32178 = ~n32175 & ~n32176 ;
  assign n32179 = ~n32177 & ~n32178 ;
  assign n32180 = ~x104 & n6725 ;
  assign n32181 = ~x102 & n7129 ;
  assign n32182 = ~x103 & n6720 ;
  assign n32183 = ~n32181 & ~n32182 ;
  assign n32184 = ~n32180 & n32183 ;
  assign n32185 = n6728 & n11380 ;
  assign n32186 = n32184 & ~n32185 ;
  assign n32187 = ~x32 & ~n32186 ;
  assign n32188 = ~x32 & ~n32187 ;
  assign n32189 = ~n32186 & ~n32187 ;
  assign n32190 = ~n32188 & ~n32189 ;
  assign n32191 = ~n31592 & ~n31596 ;
  assign n32192 = n32190 & n32191 ;
  assign n32193 = ~n32190 & ~n32191 ;
  assign n32194 = ~n32192 & ~n32193 ;
  assign n32195 = ~x101 & n8006 ;
  assign n32196 = ~x99 & n8474 ;
  assign n32197 = ~x100 & n8001 ;
  assign n32198 = ~n32196 & ~n32197 ;
  assign n32199 = ~n32195 & n32198 ;
  assign n32200 = n8009 & n9844 ;
  assign n32201 = n32199 & ~n32200 ;
  assign n32202 = ~x35 & ~n32201 ;
  assign n32203 = ~x35 & ~n32202 ;
  assign n32204 = ~n32201 & ~n32202 ;
  assign n32205 = ~n32203 & ~n32204 ;
  assign n32206 = ~n31404 & ~n31577 ;
  assign n32207 = ~n31574 & ~n32206 ;
  assign n32208 = ~x98 & n9433 ;
  assign n32209 = ~x96 & n9915 ;
  assign n32210 = ~x97 & n9428 ;
  assign n32211 = ~n32209 & ~n32210 ;
  assign n32212 = ~n32208 & n32211 ;
  assign n32213 = n8426 & n9436 ;
  assign n32214 = n32212 & ~n32213 ;
  assign n32215 = ~x38 & ~n32214 ;
  assign n32216 = ~x38 & ~n32215 ;
  assign n32217 = ~n32214 & ~n32215 ;
  assign n32218 = ~n32216 & ~n32217 ;
  assign n32219 = ~n31428 & ~n31442 ;
  assign n32220 = x2 & x5 ;
  assign n32221 = ~n31424 & ~n32220 ;
  assign n32222 = ~x70 & n27427 ;
  assign n32223 = ~x71 & ~n26217 ;
  assign n32224 = ~n32222 & ~n32223 ;
  assign n32225 = ~n32221 & n32224 ;
  assign n32226 = n32221 & ~n32224 ;
  assign n32227 = ~n32225 & ~n32226 ;
  assign n32228 = ~x74 & n24612 ;
  assign n32229 = ~x72 & n25390 ;
  assign n32230 = ~x73 & n24607 ;
  assign n32231 = ~n32229 & ~n32230 ;
  assign n32232 = ~n32228 & n32231 ;
  assign n32233 = ~n24615 & n32232 ;
  assign n32234 = ~n1066 & n32232 ;
  assign n32235 = ~n32233 & ~n32234 ;
  assign n32236 = ~x62 & ~n32235 ;
  assign n32237 = x62 & n32235 ;
  assign n32238 = ~n32236 & ~n32237 ;
  assign n32239 = n32227 & ~n32238 ;
  assign n32240 = ~n32227 & n32238 ;
  assign n32241 = ~n32239 & ~n32240 ;
  assign n32242 = ~n32219 & n32241 ;
  assign n32243 = n32219 & ~n32241 ;
  assign n32244 = ~n32242 & ~n32243 ;
  assign n32245 = ~x77 & n22325 ;
  assign n32246 = ~x75 & n23066 ;
  assign n32247 = ~x76 & n22320 ;
  assign n32248 = ~n32246 & ~n32247 ;
  assign n32249 = ~n32245 & n32248 ;
  assign n32250 = n1594 & n22328 ;
  assign n32251 = n32249 & ~n32250 ;
  assign n32252 = ~x59 & ~n32251 ;
  assign n32253 = ~x59 & ~n32252 ;
  assign n32254 = ~n32251 & ~n32252 ;
  assign n32255 = ~n32253 & ~n32254 ;
  assign n32256 = n32244 & ~n32255 ;
  assign n32257 = n32244 & ~n32256 ;
  assign n32258 = ~n32255 & ~n32256 ;
  assign n32259 = ~n32257 & ~n32258 ;
  assign n32260 = ~n31444 & ~n31448 ;
  assign n32261 = n32259 & n32260 ;
  assign n32262 = ~n32259 & ~n32260 ;
  assign n32263 = ~n32261 & ~n32262 ;
  assign n32264 = ~x80 & n20143 ;
  assign n32265 = ~x78 & n20854 ;
  assign n32266 = ~x79 & n20138 ;
  assign n32267 = ~n32265 & ~n32266 ;
  assign n32268 = ~n32264 & n32267 ;
  assign n32269 = n2145 & n20146 ;
  assign n32270 = n32268 & ~n32269 ;
  assign n32271 = ~x56 & ~n32270 ;
  assign n32272 = ~x56 & ~n32271 ;
  assign n32273 = ~n32270 & ~n32271 ;
  assign n32274 = ~n32272 & ~n32273 ;
  assign n32275 = n32263 & ~n32274 ;
  assign n32276 = n32263 & ~n32275 ;
  assign n32277 = ~n32274 & ~n32275 ;
  assign n32278 = ~n32276 & ~n32277 ;
  assign n32279 = ~n31463 & ~n31469 ;
  assign n32280 = n32278 & n32279 ;
  assign n32281 = ~n32278 & ~n32279 ;
  assign n32282 = ~n32280 & ~n32281 ;
  assign n32283 = ~x83 & n18025 ;
  assign n32284 = ~x81 & n18764 ;
  assign n32285 = ~x82 & n18020 ;
  assign n32286 = ~n32284 & ~n32285 ;
  assign n32287 = ~n32283 & n32286 ;
  assign n32288 = n2972 & n18028 ;
  assign n32289 = n32287 & ~n32288 ;
  assign n32290 = ~x53 & ~n32289 ;
  assign n32291 = ~x53 & ~n32290 ;
  assign n32292 = ~n32289 & ~n32290 ;
  assign n32293 = ~n32291 & ~n32292 ;
  assign n32294 = n32282 & ~n32293 ;
  assign n32295 = n32282 & ~n32294 ;
  assign n32296 = ~n32293 & ~n32294 ;
  assign n32297 = ~n32295 & ~n32296 ;
  assign n32298 = ~n31482 & ~n31488 ;
  assign n32299 = n32297 & n32298 ;
  assign n32300 = ~n32297 & ~n32298 ;
  assign n32301 = ~n32299 & ~n32300 ;
  assign n32302 = ~x86 & n16076 ;
  assign n32303 = ~x84 & n16756 ;
  assign n32304 = ~x85 & n16071 ;
  assign n32305 = ~n32303 & ~n32304 ;
  assign n32306 = ~n32302 & n32305 ;
  assign n32307 = n3832 & n16079 ;
  assign n32308 = n32306 & ~n32307 ;
  assign n32309 = ~x50 & ~n32308 ;
  assign n32310 = ~x50 & ~n32309 ;
  assign n32311 = ~n32308 & ~n32309 ;
  assign n32312 = ~n32310 & ~n32311 ;
  assign n32313 = n32301 & ~n32312 ;
  assign n32314 = n32301 & ~n32313 ;
  assign n32315 = ~n32312 & ~n32313 ;
  assign n32316 = ~n32314 & ~n32315 ;
  assign n32317 = ~n31407 & ~n31504 ;
  assign n32318 = ~n31501 & ~n32317 ;
  assign n32319 = n32316 & n32318 ;
  assign n32320 = ~n32316 & ~n32318 ;
  assign n32321 = ~n32319 & ~n32320 ;
  assign n32322 = ~x89 & n14233 ;
  assign n32323 = ~x87 & n14876 ;
  assign n32324 = ~x88 & n14228 ;
  assign n32325 = ~n32323 & ~n32324 ;
  assign n32326 = ~n32322 & n32325 ;
  assign n32327 = n4664 & n14236 ;
  assign n32328 = n32326 & ~n32327 ;
  assign n32329 = ~x47 & ~n32328 ;
  assign n32330 = ~x47 & ~n32329 ;
  assign n32331 = ~n32328 & ~n32329 ;
  assign n32332 = ~n32330 & ~n32331 ;
  assign n32333 = n32321 & ~n32332 ;
  assign n32334 = n32321 & ~n32333 ;
  assign n32335 = ~n32332 & ~n32333 ;
  assign n32336 = ~n32334 & ~n32335 ;
  assign n32337 = ~n31519 & ~n31523 ;
  assign n32338 = n32336 & n32337 ;
  assign n32339 = ~n32336 & ~n32337 ;
  assign n32340 = ~n32338 & ~n32339 ;
  assign n32341 = ~x92 & n12506 ;
  assign n32342 = ~x90 & n13131 ;
  assign n32343 = ~x91 & n12501 ;
  assign n32344 = ~n32342 & ~n32343 ;
  assign n32345 = ~n32341 & n32344 ;
  assign n32346 = n5896 & n12509 ;
  assign n32347 = n32345 & ~n32346 ;
  assign n32348 = ~x44 & ~n32347 ;
  assign n32349 = ~x44 & ~n32348 ;
  assign n32350 = ~n32347 & ~n32348 ;
  assign n32351 = ~n32349 & ~n32350 ;
  assign n32352 = n32340 & ~n32351 ;
  assign n32353 = n32340 & ~n32352 ;
  assign n32354 = ~n32351 & ~n32352 ;
  assign n32355 = ~n32353 & ~n32354 ;
  assign n32356 = ~n31536 & ~n31542 ;
  assign n32357 = n32355 & n32356 ;
  assign n32358 = ~n32355 & ~n32356 ;
  assign n32359 = ~n32357 & ~n32358 ;
  assign n32360 = ~x95 & n10905 ;
  assign n32361 = ~x93 & n11466 ;
  assign n32362 = ~x94 & n10900 ;
  assign n32363 = ~n32361 & ~n32362 ;
  assign n32364 = ~n32360 & n32363 ;
  assign n32365 = n7100 & n10908 ;
  assign n32366 = n32364 & ~n32365 ;
  assign n32367 = ~x41 & ~n32366 ;
  assign n32368 = ~x41 & ~n32367 ;
  assign n32369 = ~n32366 & ~n32367 ;
  assign n32370 = ~n32368 & ~n32369 ;
  assign n32371 = ~n32359 & n32370 ;
  assign n32372 = n32359 & ~n32370 ;
  assign n32373 = ~n32371 & ~n32372 ;
  assign n32374 = ~n31560 & n32373 ;
  assign n32375 = n31560 & ~n32373 ;
  assign n32376 = ~n32374 & ~n32375 ;
  assign n32377 = ~n32218 & n32376 ;
  assign n32378 = n32218 & ~n32376 ;
  assign n32379 = ~n32377 & ~n32378 ;
  assign n32380 = ~n32207 & n32379 ;
  assign n32381 = n32207 & ~n32379 ;
  assign n32382 = ~n32380 & ~n32381 ;
  assign n32383 = ~n32205 & n32382 ;
  assign n32384 = ~n32205 & ~n32383 ;
  assign n32385 = n32382 & ~n32383 ;
  assign n32386 = ~n32384 & ~n32385 ;
  assign n32387 = n32194 & ~n32386 ;
  assign n32388 = n32194 & ~n32387 ;
  assign n32389 = ~n32386 & ~n32387 ;
  assign n32390 = ~n32388 & ~n32389 ;
  assign n32391 = ~n32179 & n32390 ;
  assign n32392 = n32179 & ~n32390 ;
  assign n32393 = ~n32391 & ~n32392 ;
  assign n32394 = n32163 & ~n32393 ;
  assign n32395 = n32163 & ~n32394 ;
  assign n32396 = ~n32393 & ~n32394 ;
  assign n32397 = ~n32395 & ~n32396 ;
  assign n32398 = ~n32148 & n32397 ;
  assign n32399 = n32148 & ~n32397 ;
  assign n32400 = ~n32398 & ~n32399 ;
  assign n32401 = n32131 & ~n32400 ;
  assign n32402 = n32131 & ~n32401 ;
  assign n32403 = ~n32400 & ~n32401 ;
  assign n32404 = ~n32402 & ~n32403 ;
  assign n32405 = n32116 & ~n32404 ;
  assign n32406 = ~n32116 & n32404 ;
  assign n32407 = n32101 & ~n32406 ;
  assign n32408 = ~n32405 & n32407 ;
  assign n32409 = n32101 & ~n32408 ;
  assign n32410 = ~n32406 & ~n32408 ;
  assign n32411 = ~n32405 & n32410 ;
  assign n32412 = ~n32409 & ~n32411 ;
  assign n32413 = n32086 & ~n32412 ;
  assign n32414 = ~n32086 & n32412 ;
  assign n32415 = n32071 & ~n32414 ;
  assign n32416 = ~n32413 & n32415 ;
  assign n32417 = n32071 & ~n32416 ;
  assign n32418 = ~n32414 & ~n32416 ;
  assign n32419 = ~n32413 & n32418 ;
  assign n32420 = ~n32417 & ~n32419 ;
  assign n32421 = ~n31325 & ~n31673 ;
  assign n32422 = ~n31322 & ~n32421 ;
  assign n32423 = ~n32420 & ~n32422 ;
  assign n32424 = ~n32420 & ~n32423 ;
  assign n32425 = ~n32422 & ~n32423 ;
  assign n32426 = ~n32424 & ~n32425 ;
  assign n32427 = ~n31677 & ~n31680 ;
  assign n32428 = ~n32426 & ~n32427 ;
  assign n32429 = n32426 & n32427 ;
  assign n32430 = ~n32428 & ~n32429 ;
  assign n32433 = ~n32430 & ~x198 ;
  assign n32434 = ~n32432 & ~n32433 ;
  assign n32435 = ~n32051 & ~n32056 ;
  assign n32436 = ~n31697 & ~n32044 ;
  assign n32437 = ~n31713 & ~n32041 ;
  assign n32438 = x127 & n673 ;
  assign n32439 = n577 & n26962 ;
  assign n32440 = ~n32438 & ~n32439 ;
  assign n32441 = x8 & ~n32440 ;
  assign n32442 = x8 & ~n32441 ;
  assign n32443 = ~n32440 & ~n32441 ;
  assign n32444 = ~n32442 & ~n32443 ;
  assign n32445 = ~n32437 & ~n32444 ;
  assign n32446 = ~n32437 & ~n32445 ;
  assign n32447 = ~n32444 & ~n32445 ;
  assign n32448 = ~n32446 & ~n32447 ;
  assign n32449 = x120 & n2093 ;
  assign n32450 = x118 & n2275 ;
  assign n32451 = x119 & n2088 ;
  assign n32452 = ~n32450 & ~n32451 ;
  assign n32453 = ~n32449 & n32452 ;
  assign n32454 = n2096 & n21143 ;
  assign n32455 = n32453 & ~n32454 ;
  assign n32456 = x17 & ~n32455 ;
  assign n32457 = x17 & ~n32456 ;
  assign n32458 = ~n32455 & ~n32456 ;
  assign n32459 = ~n32457 & ~n32458 ;
  assign n32460 = ~n31758 & ~n32029 ;
  assign n32461 = n32459 & n32460 ;
  assign n32462 = ~n32459 & ~n32460 ;
  assign n32463 = ~n32461 & ~n32462 ;
  assign n32464 = x114 & n3589 ;
  assign n32465 = x112 & n3878 ;
  assign n32466 = x113 & n3584 ;
  assign n32467 = ~n32465 & ~n32466 ;
  assign n32468 = ~n32464 & n32467 ;
  assign n32469 = n3592 & n17012 ;
  assign n32470 = n32468 & ~n32469 ;
  assign n32471 = x23 & ~n32470 ;
  assign n32472 = x23 & ~n32471 ;
  assign n32473 = ~n32470 & ~n32471 ;
  assign n32474 = ~n32472 & ~n32473 ;
  assign n32475 = ~n31789 & ~n32022 ;
  assign n32476 = n32474 & n32475 ;
  assign n32477 = ~n32474 & ~n32475 ;
  assign n32478 = ~n32476 & ~n32477 ;
  assign n32479 = x111 & n4531 ;
  assign n32480 = x109 & n4847 ;
  assign n32481 = x110 & n4526 ;
  assign n32482 = ~n32480 & ~n32481 ;
  assign n32483 = ~n32479 & n32482 ;
  assign n32484 = n4534 & n15111 ;
  assign n32485 = n32483 & ~n32484 ;
  assign n32486 = x26 & ~n32485 ;
  assign n32487 = x26 & ~n32486 ;
  assign n32488 = ~n32485 & ~n32486 ;
  assign n32489 = ~n32487 & ~n32488 ;
  assign n32490 = ~n31807 & ~n32018 ;
  assign n32491 = ~n31804 & ~n32490 ;
  assign n32492 = ~n32489 & ~n32491 ;
  assign n32493 = ~n32489 & ~n32492 ;
  assign n32494 = ~n32491 & ~n32492 ;
  assign n32495 = ~n32493 & ~n32494 ;
  assign n32496 = x105 & n6725 ;
  assign n32497 = x103 & n7129 ;
  assign n32498 = x104 & n6720 ;
  assign n32499 = ~n32497 & ~n32498 ;
  assign n32500 = ~n32496 & n32499 ;
  assign n32501 = n6728 & n11648 ;
  assign n32502 = n32500 & ~n32501 ;
  assign n32503 = x32 & ~n32502 ;
  assign n32504 = x32 & ~n32503 ;
  assign n32505 = ~n32502 & ~n32503 ;
  assign n32506 = ~n32504 & ~n32505 ;
  assign n32507 = ~n32008 & ~n32011 ;
  assign n32508 = n32506 & n32507 ;
  assign n32509 = ~n32506 & ~n32507 ;
  assign n32510 = ~n32508 & ~n32509 ;
  assign n32511 = ~n31928 & ~n31941 ;
  assign n32512 = x87 & n16076 ;
  assign n32513 = x85 & n16756 ;
  assign n32514 = x86 & n16071 ;
  assign n32515 = ~n32513 & ~n32514 ;
  assign n32516 = ~n32512 & n32515 ;
  assign n32517 = n3991 & n16079 ;
  assign n32518 = n32516 & ~n32517 ;
  assign n32519 = x50 & ~n32518 ;
  assign n32520 = x50 & ~n32519 ;
  assign n32521 = ~n32518 & ~n32519 ;
  assign n32522 = ~n32520 & ~n32521 ;
  assign n32523 = ~n31909 & ~n31922 ;
  assign n32524 = ~n31870 & ~n31884 ;
  assign n32525 = ~n31853 & ~n31867 ;
  assign n32526 = x71 & n27024 ;
  assign n32527 = x72 & ~n26217 ;
  assign n32528 = ~n32526 & ~n32527 ;
  assign n32529 = n31852 & ~n32528 ;
  assign n32530 = ~n31852 & n32528 ;
  assign n32531 = ~n32525 & ~n32530 ;
  assign n32532 = ~n32529 & n32531 ;
  assign n32533 = ~n32525 & ~n32532 ;
  assign n32534 = ~n32530 & ~n32532 ;
  assign n32535 = ~n32529 & n32534 ;
  assign n32536 = ~n32533 & ~n32535 ;
  assign n32537 = x75 & n24612 ;
  assign n32538 = x73 & n25390 ;
  assign n32539 = x74 & n24607 ;
  assign n32540 = ~n32538 & ~n32539 ;
  assign n32541 = ~n32537 & n32540 ;
  assign n32542 = n1150 & n24615 ;
  assign n32543 = n32541 & ~n32542 ;
  assign n32544 = x62 & ~n32543 ;
  assign n32545 = x62 & ~n32544 ;
  assign n32546 = ~n32543 & ~n32544 ;
  assign n32547 = ~n32545 & ~n32546 ;
  assign n32548 = ~n32536 & n32547 ;
  assign n32549 = n32536 & ~n32547 ;
  assign n32550 = ~n32548 & ~n32549 ;
  assign n32551 = x78 & n22325 ;
  assign n32552 = x76 & n23066 ;
  assign n32553 = x77 & n22320 ;
  assign n32554 = ~n32552 & ~n32553 ;
  assign n32555 = ~n32551 & n32554 ;
  assign n32556 = n1624 & n22328 ;
  assign n32557 = n32555 & ~n32556 ;
  assign n32558 = x59 & ~n32557 ;
  assign n32559 = x59 & ~n32558 ;
  assign n32560 = ~n32557 & ~n32558 ;
  assign n32561 = ~n32559 & ~n32560 ;
  assign n32562 = ~n32550 & ~n32561 ;
  assign n32563 = n32550 & n32561 ;
  assign n32564 = ~n32562 & ~n32563 ;
  assign n32565 = n32524 & ~n32564 ;
  assign n32566 = ~n32524 & n32564 ;
  assign n32567 = ~n32565 & ~n32566 ;
  assign n32568 = x81 & n20143 ;
  assign n32569 = x79 & n20854 ;
  assign n32570 = x80 & n20138 ;
  assign n32571 = ~n32569 & ~n32570 ;
  assign n32572 = ~n32568 & n32571 ;
  assign n32573 = n2348 & n20146 ;
  assign n32574 = n32572 & ~n32573 ;
  assign n32575 = x56 & ~n32574 ;
  assign n32576 = x56 & ~n32575 ;
  assign n32577 = ~n32574 & ~n32575 ;
  assign n32578 = ~n32576 & ~n32577 ;
  assign n32579 = n32567 & ~n32578 ;
  assign n32580 = n32567 & ~n32579 ;
  assign n32581 = ~n32578 & ~n32579 ;
  assign n32582 = ~n32580 & ~n32581 ;
  assign n32583 = ~n31890 & ~n31903 ;
  assign n32584 = n32582 & n32583 ;
  assign n32585 = ~n32582 & ~n32583 ;
  assign n32586 = ~n32584 & ~n32585 ;
  assign n32587 = x84 & n18025 ;
  assign n32588 = x82 & n18764 ;
  assign n32589 = x83 & n18020 ;
  assign n32590 = ~n32588 & ~n32589 ;
  assign n32591 = ~n32587 & n32590 ;
  assign n32592 = n3114 & n18028 ;
  assign n32593 = n32591 & ~n32592 ;
  assign n32594 = x53 & ~n32593 ;
  assign n32595 = x53 & ~n32594 ;
  assign n32596 = ~n32593 & ~n32594 ;
  assign n32597 = ~n32595 & ~n32596 ;
  assign n32598 = ~n32586 & n32597 ;
  assign n32599 = n32586 & ~n32597 ;
  assign n32600 = ~n32598 & ~n32599 ;
  assign n32601 = ~n32523 & n32600 ;
  assign n32602 = ~n32523 & ~n32601 ;
  assign n32603 = n32600 & ~n32601 ;
  assign n32604 = ~n32602 & ~n32603 ;
  assign n32605 = ~n32522 & ~n32604 ;
  assign n32606 = n32522 & ~n32603 ;
  assign n32607 = ~n32602 & n32606 ;
  assign n32608 = ~n32605 & ~n32607 ;
  assign n32609 = ~n32511 & n32608 ;
  assign n32610 = n32511 & ~n32608 ;
  assign n32611 = ~n32609 & ~n32610 ;
  assign n32612 = x90 & n14233 ;
  assign n32613 = x88 & n14876 ;
  assign n32614 = x89 & n14228 ;
  assign n32615 = ~n32613 & ~n32614 ;
  assign n32616 = ~n32612 & n32615 ;
  assign n32617 = n4986 & n14236 ;
  assign n32618 = n32616 & ~n32617 ;
  assign n32619 = x47 & ~n32618 ;
  assign n32620 = x47 & ~n32619 ;
  assign n32621 = ~n32618 & ~n32619 ;
  assign n32622 = ~n32620 & ~n32621 ;
  assign n32623 = n32611 & ~n32622 ;
  assign n32624 = n32611 & ~n32623 ;
  assign n32625 = ~n32622 & ~n32623 ;
  assign n32626 = ~n32624 & ~n32625 ;
  assign n32627 = ~n31948 & ~n31961 ;
  assign n32628 = n32626 & n32627 ;
  assign n32629 = ~n32626 & ~n32627 ;
  assign n32630 = ~n32628 & ~n32629 ;
  assign n32631 = x93 & n12506 ;
  assign n32632 = x91 & n13131 ;
  assign n32633 = x92 & n12501 ;
  assign n32634 = ~n32632 & ~n32633 ;
  assign n32635 = ~n32631 & n32634 ;
  assign n32636 = n6094 & n12509 ;
  assign n32637 = n32635 & ~n32636 ;
  assign n32638 = x44 & ~n32637 ;
  assign n32639 = x44 & ~n32638 ;
  assign n32640 = ~n32637 & ~n32638 ;
  assign n32641 = ~n32639 & ~n32640 ;
  assign n32642 = n32630 & ~n32641 ;
  assign n32643 = n32630 & ~n32642 ;
  assign n32644 = ~n32641 & ~n32642 ;
  assign n32645 = ~n32643 & ~n32644 ;
  assign n32646 = ~n31967 & ~n31980 ;
  assign n32647 = n32645 & n32646 ;
  assign n32648 = ~n32645 & ~n32646 ;
  assign n32649 = ~n32647 & ~n32648 ;
  assign n32650 = x96 & n10905 ;
  assign n32651 = x94 & n11466 ;
  assign n32652 = x95 & n10900 ;
  assign n32653 = ~n32651 & ~n32652 ;
  assign n32654 = ~n32650 & n32653 ;
  assign n32655 = n7321 & n10908 ;
  assign n32656 = n32654 & ~n32655 ;
  assign n32657 = x41 & ~n32656 ;
  assign n32658 = x41 & ~n32657 ;
  assign n32659 = ~n32656 & ~n32657 ;
  assign n32660 = ~n32658 & ~n32659 ;
  assign n32661 = ~n32649 & n32660 ;
  assign n32662 = n32649 & ~n32660 ;
  assign n32663 = ~n32661 & ~n32662 ;
  assign n32664 = ~n31986 & ~n32000 ;
  assign n32665 = n32663 & ~n32664 ;
  assign n32666 = ~n32663 & n32664 ;
  assign n32667 = ~n32665 & ~n32666 ;
  assign n32668 = x99 & n9433 ;
  assign n32669 = x97 & n9915 ;
  assign n32670 = x98 & n9428 ;
  assign n32671 = ~n32669 & ~n32670 ;
  assign n32672 = ~n32668 & n32671 ;
  assign n32673 = n8660 & n9436 ;
  assign n32674 = n32672 & ~n32673 ;
  assign n32675 = x38 & ~n32674 ;
  assign n32676 = x38 & ~n32675 ;
  assign n32677 = ~n32674 & ~n32675 ;
  assign n32678 = ~n32676 & ~n32677 ;
  assign n32679 = n32667 & ~n32678 ;
  assign n32680 = n32667 & ~n32679 ;
  assign n32681 = ~n32678 & ~n32679 ;
  assign n32682 = ~n32680 & ~n32681 ;
  assign n32683 = ~n32002 & ~n32005 ;
  assign n32684 = n32682 & n32683 ;
  assign n32685 = ~n32682 & ~n32683 ;
  assign n32686 = ~n32684 & ~n32685 ;
  assign n32687 = x102 & n8006 ;
  assign n32688 = x100 & n8474 ;
  assign n32689 = x101 & n8001 ;
  assign n32690 = ~n32688 & ~n32689 ;
  assign n32691 = ~n32687 & n32690 ;
  assign n32692 = n8009 & n10092 ;
  assign n32693 = n32691 & ~n32692 ;
  assign n32694 = x35 & ~n32693 ;
  assign n32695 = x35 & ~n32694 ;
  assign n32696 = ~n32693 & ~n32694 ;
  assign n32697 = ~n32695 & ~n32696 ;
  assign n32698 = n32686 & ~n32697 ;
  assign n32699 = ~n32686 & n32697 ;
  assign n32700 = n32510 & ~n32699 ;
  assign n32701 = ~n32698 & n32700 ;
  assign n32702 = n32510 & ~n32701 ;
  assign n32703 = ~n32699 & ~n32701 ;
  assign n32704 = ~n32698 & n32703 ;
  assign n32705 = ~n32702 & ~n32704 ;
  assign n32706 = ~n31821 & ~n32015 ;
  assign n32707 = x108 & n5560 ;
  assign n32708 = x106 & n5943 ;
  assign n32709 = x107 & n5555 ;
  assign n32710 = ~n32708 & ~n32709 ;
  assign n32711 = ~n32707 & n32710 ;
  assign n32712 = ~n5563 & n32711 ;
  assign n32713 = ~n13323 & n32711 ;
  assign n32714 = ~n32712 & ~n32713 ;
  assign n32715 = x29 & ~n32714 ;
  assign n32716 = ~x29 & n32714 ;
  assign n32717 = ~n32715 & ~n32716 ;
  assign n32718 = ~n32706 & ~n32717 ;
  assign n32719 = ~n32706 & ~n32718 ;
  assign n32720 = ~n32717 & ~n32718 ;
  assign n32721 = ~n32719 & ~n32720 ;
  assign n32722 = ~n32705 & ~n32721 ;
  assign n32723 = ~n32705 & ~n32722 ;
  assign n32724 = ~n32721 & ~n32722 ;
  assign n32725 = ~n32723 & ~n32724 ;
  assign n32726 = ~n32495 & ~n32725 ;
  assign n32727 = ~n32495 & ~n32726 ;
  assign n32728 = ~n32725 & ~n32726 ;
  assign n32729 = ~n32727 & ~n32728 ;
  assign n32730 = ~n32478 & n32729 ;
  assign n32731 = n32478 & ~n32729 ;
  assign n32732 = ~n32730 & ~n32731 ;
  assign n32733 = ~n31776 & ~n32025 ;
  assign n32734 = ~n31773 & ~n32733 ;
  assign n32735 = x117 & n2751 ;
  assign n32736 = x115 & n3020 ;
  assign n32737 = x116 & n2746 ;
  assign n32738 = ~n32736 & ~n32737 ;
  assign n32739 = ~n32735 & n32738 ;
  assign n32740 = ~n2754 & n32739 ;
  assign n32741 = ~n19026 & n32739 ;
  assign n32742 = ~n32740 & ~n32741 ;
  assign n32743 = x20 & ~n32742 ;
  assign n32744 = ~x20 & n32742 ;
  assign n32745 = ~n32743 & ~n32744 ;
  assign n32746 = ~n32734 & ~n32745 ;
  assign n32747 = ~n32734 & ~n32746 ;
  assign n32748 = ~n32745 & ~n32746 ;
  assign n32749 = ~n32747 & ~n32748 ;
  assign n32750 = n32732 & ~n32749 ;
  assign n32751 = n32732 & ~n32750 ;
  assign n32752 = ~n32749 & ~n32750 ;
  assign n32753 = ~n32751 & ~n32752 ;
  assign n32754 = n32463 & ~n32753 ;
  assign n32755 = n32463 & ~n32754 ;
  assign n32756 = ~n32753 & ~n32754 ;
  assign n32757 = ~n32755 & ~n32756 ;
  assign n32758 = x123 & n1434 ;
  assign n32759 = x121 & n1646 ;
  assign n32760 = x122 & n1429 ;
  assign n32761 = ~n32759 & ~n32760 ;
  assign n32762 = ~n32758 & n32761 ;
  assign n32763 = n1437 & n23382 ;
  assign n32764 = n32762 & ~n32763 ;
  assign n32765 = x14 & ~n32764 ;
  assign n32766 = x14 & ~n32765 ;
  assign n32767 = ~n32764 & ~n32765 ;
  assign n32768 = ~n32766 & ~n32767 ;
  assign n32769 = ~n31743 & ~n32033 ;
  assign n32770 = ~n32768 & ~n32769 ;
  assign n32771 = ~n32768 & ~n32770 ;
  assign n32772 = ~n32769 & ~n32770 ;
  assign n32773 = ~n32771 & ~n32772 ;
  assign n32774 = ~n32757 & n32773 ;
  assign n32775 = n32757 & ~n32773 ;
  assign n32776 = ~n32774 & ~n32775 ;
  assign n32777 = ~n31727 & ~n32036 ;
  assign n32778 = x126 & n945 ;
  assign n32779 = x124 & n1099 ;
  assign n32780 = x125 & n940 ;
  assign n32781 = ~n32779 & ~n32780 ;
  assign n32782 = ~n32778 & n32781 ;
  assign n32783 = ~n948 & n32782 ;
  assign n32784 = ~n25735 & n32782 ;
  assign n32785 = ~n32783 & ~n32784 ;
  assign n32786 = x11 & ~n32785 ;
  assign n32787 = ~x11 & n32785 ;
  assign n32788 = ~n32786 & ~n32787 ;
  assign n32789 = ~n32777 & ~n32788 ;
  assign n32790 = ~n32777 & ~n32789 ;
  assign n32791 = ~n32788 & ~n32789 ;
  assign n32792 = ~n32790 & ~n32791 ;
  assign n32793 = ~n32776 & ~n32792 ;
  assign n32794 = n32776 & ~n32791 ;
  assign n32795 = ~n32790 & n32794 ;
  assign n32796 = ~n32793 & ~n32795 ;
  assign n32797 = ~n32448 & n32796 ;
  assign n32798 = n32448 & ~n32796 ;
  assign n32799 = ~n32797 & ~n32798 ;
  assign n32800 = ~n32436 & n32799 ;
  assign n32801 = ~n32436 & ~n32800 ;
  assign n32802 = n32799 & ~n32800 ;
  assign n32803 = ~n32801 & ~n32802 ;
  assign n32804 = ~n32435 & ~n32803 ;
  assign n32805 = n32435 & ~n32802 ;
  assign n32806 = ~n32801 & n32805 ;
  assign n32807 = ~n32804 & ~n32806 ;
  assign n33182 = n32807 & x199 ;
  assign n32808 = ~n32423 & ~n32428 ;
  assign n32809 = ~n32069 & ~n32416 ;
  assign n32810 = ~n32085 & ~n32413 ;
  assign n32811 = ~x127 & n673 ;
  assign n32812 = n577 & n27365 ;
  assign n32813 = ~n32811 & ~n32812 ;
  assign n32814 = ~x8 & ~n32813 ;
  assign n32815 = ~x8 & ~n32814 ;
  assign n32816 = ~n32813 & ~n32814 ;
  assign n32817 = ~n32815 & ~n32816 ;
  assign n32818 = ~n32810 & ~n32817 ;
  assign n32819 = ~n32810 & ~n32818 ;
  assign n32820 = ~n32817 & ~n32818 ;
  assign n32821 = ~n32819 & ~n32820 ;
  assign n32822 = ~x120 & n2093 ;
  assign n32823 = ~x118 & n2275 ;
  assign n32824 = ~x119 & n2088 ;
  assign n32825 = ~n32823 & ~n32824 ;
  assign n32826 = ~n32822 & n32825 ;
  assign n32827 = n2096 & n21501 ;
  assign n32828 = n32826 & ~n32827 ;
  assign n32829 = ~x17 & ~n32828 ;
  assign n32830 = ~x17 & ~n32829 ;
  assign n32831 = ~n32828 & ~n32829 ;
  assign n32832 = ~n32830 & ~n32831 ;
  assign n32833 = ~n32130 & ~n32401 ;
  assign n32834 = n32832 & n32833 ;
  assign n32835 = ~n32832 & ~n32833 ;
  assign n32836 = ~n32834 & ~n32835 ;
  assign n32837 = ~x114 & n3589 ;
  assign n32838 = ~x112 & n3878 ;
  assign n32839 = ~x113 & n3584 ;
  assign n32840 = ~n32838 & ~n32839 ;
  assign n32841 = ~n32837 & n32840 ;
  assign n32842 = n3592 & n17333 ;
  assign n32843 = n32841 & ~n32842 ;
  assign n32844 = ~x23 & ~n32843 ;
  assign n32845 = ~x23 & ~n32844 ;
  assign n32846 = ~n32843 & ~n32844 ;
  assign n32847 = ~n32845 & ~n32846 ;
  assign n32848 = ~n32161 & ~n32394 ;
  assign n32849 = n32847 & n32848 ;
  assign n32850 = ~n32847 & ~n32848 ;
  assign n32851 = ~n32849 & ~n32850 ;
  assign n32852 = ~x111 & n4531 ;
  assign n32853 = ~x109 & n4847 ;
  assign n32854 = ~x110 & n4526 ;
  assign n32855 = ~n32853 & ~n32854 ;
  assign n32856 = ~n32852 & n32855 ;
  assign n32857 = n4534 & n15411 ;
  assign n32858 = n32856 & ~n32857 ;
  assign n32859 = ~x26 & ~n32858 ;
  assign n32860 = ~x26 & ~n32859 ;
  assign n32861 = ~n32858 & ~n32859 ;
  assign n32862 = ~n32860 & ~n32861 ;
  assign n32863 = ~n32179 & ~n32390 ;
  assign n32864 = ~n32176 & ~n32863 ;
  assign n32865 = ~n32862 & ~n32864 ;
  assign n32866 = ~n32862 & ~n32865 ;
  assign n32867 = ~n32864 & ~n32865 ;
  assign n32868 = ~n32866 & ~n32867 ;
  assign n32869 = ~x105 & n6725 ;
  assign n32870 = ~x103 & n7129 ;
  assign n32871 = ~x104 & n6720 ;
  assign n32872 = ~n32870 & ~n32871 ;
  assign n32873 = ~n32869 & n32872 ;
  assign n32874 = n6728 & n11907 ;
  assign n32875 = n32873 & ~n32874 ;
  assign n32876 = ~x32 & ~n32875 ;
  assign n32877 = ~x32 & ~n32876 ;
  assign n32878 = ~n32875 & ~n32876 ;
  assign n32879 = ~n32877 & ~n32878 ;
  assign n32880 = ~n32380 & ~n32383 ;
  assign n32881 = n32879 & n32880 ;
  assign n32882 = ~n32879 & ~n32880 ;
  assign n32883 = ~n32881 & ~n32882 ;
  assign n32884 = ~n32300 & ~n32313 ;
  assign n32885 = ~x87 & n16076 ;
  assign n32886 = ~x85 & n16756 ;
  assign n32887 = ~x86 & n16071 ;
  assign n32888 = ~n32886 & ~n32887 ;
  assign n32889 = ~n32885 & n32888 ;
  assign n32890 = n4143 & n16079 ;
  assign n32891 = n32889 & ~n32890 ;
  assign n32892 = ~x50 & ~n32891 ;
  assign n32893 = ~x50 & ~n32892 ;
  assign n32894 = ~n32891 & ~n32892 ;
  assign n32895 = ~n32893 & ~n32894 ;
  assign n32896 = ~n32281 & ~n32294 ;
  assign n32897 = ~n32242 & ~n32256 ;
  assign n32898 = ~n32225 & ~n32239 ;
  assign n32899 = ~x71 & n27427 ;
  assign n32900 = ~x72 & ~n26217 ;
  assign n32901 = ~n32899 & ~n32900 ;
  assign n32902 = n32224 & ~n32901 ;
  assign n32903 = ~n32224 & n32901 ;
  assign n32904 = ~n32898 & ~n32903 ;
  assign n32905 = ~n32902 & n32904 ;
  assign n32906 = ~n32898 & ~n32905 ;
  assign n32907 = ~n32903 & ~n32905 ;
  assign n32908 = ~n32902 & n32907 ;
  assign n32909 = ~n32906 & ~n32908 ;
  assign n32910 = ~x75 & n24612 ;
  assign n32911 = ~x73 & n25390 ;
  assign n32912 = ~x74 & n24607 ;
  assign n32913 = ~n32911 & ~n32912 ;
  assign n32914 = ~n32910 & n32913 ;
  assign n32915 = n1225 & n24615 ;
  assign n32916 = n32914 & ~n32915 ;
  assign n32917 = ~x62 & ~n32916 ;
  assign n32918 = ~x62 & ~n32917 ;
  assign n32919 = ~n32916 & ~n32917 ;
  assign n32920 = ~n32918 & ~n32919 ;
  assign n32921 = ~n32909 & n32920 ;
  assign n32922 = n32909 & ~n32920 ;
  assign n32923 = ~n32921 & ~n32922 ;
  assign n32924 = ~x78 & n22325 ;
  assign n32925 = ~x76 & n23066 ;
  assign n32926 = ~x77 & n22320 ;
  assign n32927 = ~n32925 & ~n32926 ;
  assign n32928 = ~n32924 & n32927 ;
  assign n32929 = n1718 & n22328 ;
  assign n32930 = n32928 & ~n32929 ;
  assign n32931 = ~x59 & ~n32930 ;
  assign n32932 = ~x59 & ~n32931 ;
  assign n32933 = ~n32930 & ~n32931 ;
  assign n32934 = ~n32932 & ~n32933 ;
  assign n32935 = ~n32923 & ~n32934 ;
  assign n32936 = n32923 & n32934 ;
  assign n32937 = ~n32935 & ~n32936 ;
  assign n32938 = n32897 & ~n32937 ;
  assign n32939 = ~n32897 & n32937 ;
  assign n32940 = ~n32938 & ~n32939 ;
  assign n32941 = ~x81 & n20143 ;
  assign n32942 = ~x79 & n20854 ;
  assign n32943 = ~x80 & n20138 ;
  assign n32944 = ~n32942 & ~n32943 ;
  assign n32945 = ~n32941 & n32944 ;
  assign n32946 = n2460 & n20146 ;
  assign n32947 = n32945 & ~n32946 ;
  assign n32948 = ~x56 & ~n32947 ;
  assign n32949 = ~x56 & ~n32948 ;
  assign n32950 = ~n32947 & ~n32948 ;
  assign n32951 = ~n32949 & ~n32950 ;
  assign n32952 = n32940 & ~n32951 ;
  assign n32953 = n32940 & ~n32952 ;
  assign n32954 = ~n32951 & ~n32952 ;
  assign n32955 = ~n32953 & ~n32954 ;
  assign n32956 = ~n32262 & ~n32275 ;
  assign n32957 = n32955 & n32956 ;
  assign n32958 = ~n32955 & ~n32956 ;
  assign n32959 = ~n32957 & ~n32958 ;
  assign n32960 = ~x84 & n18025 ;
  assign n32961 = ~x82 & n18764 ;
  assign n32962 = ~x83 & n18020 ;
  assign n32963 = ~n32961 & ~n32962 ;
  assign n32964 = ~n32960 & n32963 ;
  assign n32965 = n3247 & n18028 ;
  assign n32966 = n32964 & ~n32965 ;
  assign n32967 = ~x53 & ~n32966 ;
  assign n32968 = ~x53 & ~n32967 ;
  assign n32969 = ~n32966 & ~n32967 ;
  assign n32970 = ~n32968 & ~n32969 ;
  assign n32971 = ~n32959 & n32970 ;
  assign n32972 = n32959 & ~n32970 ;
  assign n32973 = ~n32971 & ~n32972 ;
  assign n32974 = ~n32896 & n32973 ;
  assign n32975 = ~n32896 & ~n32974 ;
  assign n32976 = n32973 & ~n32974 ;
  assign n32977 = ~n32975 & ~n32976 ;
  assign n32978 = ~n32895 & ~n32977 ;
  assign n32979 = n32895 & ~n32976 ;
  assign n32980 = ~n32975 & n32979 ;
  assign n32981 = ~n32978 & ~n32980 ;
  assign n32982 = ~n32884 & n32981 ;
  assign n32983 = n32884 & ~n32981 ;
  assign n32984 = ~n32982 & ~n32983 ;
  assign n32985 = ~x90 & n14233 ;
  assign n32986 = ~x88 & n14876 ;
  assign n32987 = ~x89 & n14228 ;
  assign n32988 = ~n32986 & ~n32987 ;
  assign n32989 = ~n32985 & n32988 ;
  assign n32990 = n5155 & n14236 ;
  assign n32991 = n32989 & ~n32990 ;
  assign n32992 = ~x47 & ~n32991 ;
  assign n32993 = ~x47 & ~n32992 ;
  assign n32994 = ~n32991 & ~n32992 ;
  assign n32995 = ~n32993 & ~n32994 ;
  assign n32996 = n32984 & ~n32995 ;
  assign n32997 = n32984 & ~n32996 ;
  assign n32998 = ~n32995 & ~n32996 ;
  assign n32999 = ~n32997 & ~n32998 ;
  assign n33000 = ~n32320 & ~n32333 ;
  assign n33001 = n32999 & n33000 ;
  assign n33002 = ~n32999 & ~n33000 ;
  assign n33003 = ~n33001 & ~n33002 ;
  assign n33004 = ~x93 & n12506 ;
  assign n33005 = ~x91 & n13131 ;
  assign n33006 = ~x92 & n12501 ;
  assign n33007 = ~n33005 & ~n33006 ;
  assign n33008 = ~n33004 & n33007 ;
  assign n33009 = n6285 & n12509 ;
  assign n33010 = n33008 & ~n33009 ;
  assign n33011 = ~x44 & ~n33010 ;
  assign n33012 = ~x44 & ~n33011 ;
  assign n33013 = ~n33010 & ~n33011 ;
  assign n33014 = ~n33012 & ~n33013 ;
  assign n33015 = n33003 & ~n33014 ;
  assign n33016 = n33003 & ~n33015 ;
  assign n33017 = ~n33014 & ~n33015 ;
  assign n33018 = ~n33016 & ~n33017 ;
  assign n33019 = ~n32339 & ~n32352 ;
  assign n33020 = n33018 & n33019 ;
  assign n33021 = ~n33018 & ~n33019 ;
  assign n33022 = ~n33020 & ~n33021 ;
  assign n33023 = ~x96 & n10905 ;
  assign n33024 = ~x94 & n11466 ;
  assign n33025 = ~x95 & n10900 ;
  assign n33026 = ~n33024 & ~n33025 ;
  assign n33027 = ~n33023 & n33026 ;
  assign n33028 = n7531 & n10908 ;
  assign n33029 = n33027 & ~n33028 ;
  assign n33030 = ~x41 & ~n33029 ;
  assign n33031 = ~x41 & ~n33030 ;
  assign n33032 = ~n33029 & ~n33030 ;
  assign n33033 = ~n33031 & ~n33032 ;
  assign n33034 = ~n33022 & n33033 ;
  assign n33035 = n33022 & ~n33033 ;
  assign n33036 = ~n33034 & ~n33035 ;
  assign n33037 = ~n32358 & ~n32372 ;
  assign n33038 = n33036 & ~n33037 ;
  assign n33039 = ~n33036 & n33037 ;
  assign n33040 = ~n33038 & ~n33039 ;
  assign n33041 = ~x99 & n9433 ;
  assign n33042 = ~x97 & n9915 ;
  assign n33043 = ~x98 & n9428 ;
  assign n33044 = ~n33042 & ~n33043 ;
  assign n33045 = ~n33041 & n33044 ;
  assign n33046 = n8885 & n9436 ;
  assign n33047 = n33045 & ~n33046 ;
  assign n33048 = ~x38 & ~n33047 ;
  assign n33049 = ~x38 & ~n33048 ;
  assign n33050 = ~n33047 & ~n33048 ;
  assign n33051 = ~n33049 & ~n33050 ;
  assign n33052 = n33040 & ~n33051 ;
  assign n33053 = n33040 & ~n33052 ;
  assign n33054 = ~n33051 & ~n33052 ;
  assign n33055 = ~n33053 & ~n33054 ;
  assign n33056 = ~n32374 & ~n32377 ;
  assign n33057 = n33055 & n33056 ;
  assign n33058 = ~n33055 & ~n33056 ;
  assign n33059 = ~n33057 & ~n33058 ;
  assign n33060 = ~x102 & n8006 ;
  assign n33061 = ~x100 & n8474 ;
  assign n33062 = ~x101 & n8001 ;
  assign n33063 = ~n33061 & ~n33062 ;
  assign n33064 = ~n33060 & n33063 ;
  assign n33065 = n8009 & n10333 ;
  assign n33066 = n33064 & ~n33065 ;
  assign n33067 = ~x35 & ~n33066 ;
  assign n33068 = ~x35 & ~n33067 ;
  assign n33069 = ~n33066 & ~n33067 ;
  assign n33070 = ~n33068 & ~n33069 ;
  assign n33071 = n33059 & ~n33070 ;
  assign n33072 = ~n33059 & n33070 ;
  assign n33073 = n32883 & ~n33072 ;
  assign n33074 = ~n33071 & n33073 ;
  assign n33075 = n32883 & ~n33074 ;
  assign n33076 = ~n33072 & ~n33074 ;
  assign n33077 = ~n33071 & n33076 ;
  assign n33078 = ~n33075 & ~n33077 ;
  assign n33079 = ~n32193 & ~n32387 ;
  assign n33080 = ~x108 & n5560 ;
  assign n33081 = ~x106 & n5943 ;
  assign n33082 = ~x107 & n5555 ;
  assign n33083 = ~n33081 & ~n33082 ;
  assign n33084 = ~n33080 & n33083 ;
  assign n33085 = ~n5563 & n33084 ;
  assign n33086 = ~n13601 & n33084 ;
  assign n33087 = ~n33085 & ~n33086 ;
  assign n33088 = ~x29 & ~n33087 ;
  assign n33089 = x29 & n33087 ;
  assign n33090 = ~n33088 & ~n33089 ;
  assign n33091 = ~n33079 & ~n33090 ;
  assign n33092 = ~n33079 & ~n33091 ;
  assign n33093 = ~n33090 & ~n33091 ;
  assign n33094 = ~n33092 & ~n33093 ;
  assign n33095 = ~n33078 & ~n33094 ;
  assign n33096 = ~n33078 & ~n33095 ;
  assign n33097 = ~n33094 & ~n33095 ;
  assign n33098 = ~n33096 & ~n33097 ;
  assign n33099 = ~n32868 & ~n33098 ;
  assign n33100 = ~n32868 & ~n33099 ;
  assign n33101 = ~n33098 & ~n33099 ;
  assign n33102 = ~n33100 & ~n33101 ;
  assign n33103 = ~n32851 & n33102 ;
  assign n33104 = n32851 & ~n33102 ;
  assign n33105 = ~n33103 & ~n33104 ;
  assign n33106 = ~n32148 & ~n32397 ;
  assign n33107 = ~n32145 & ~n33106 ;
  assign n33108 = ~x117 & n2751 ;
  assign n33109 = ~x115 & n3020 ;
  assign n33110 = ~x116 & n2746 ;
  assign n33111 = ~n33109 & ~n33110 ;
  assign n33112 = ~n33108 & n33111 ;
  assign n33113 = ~n2754 & n33112 ;
  assign n33114 = ~n19365 & n33112 ;
  assign n33115 = ~n33113 & ~n33114 ;
  assign n33116 = ~x20 & ~n33115 ;
  assign n33117 = x20 & n33115 ;
  assign n33118 = ~n33116 & ~n33117 ;
  assign n33119 = ~n33107 & ~n33118 ;
  assign n33120 = ~n33107 & ~n33119 ;
  assign n33121 = ~n33118 & ~n33119 ;
  assign n33122 = ~n33120 & ~n33121 ;
  assign n33123 = n33105 & ~n33122 ;
  assign n33124 = n33105 & ~n33123 ;
  assign n33125 = ~n33122 & ~n33123 ;
  assign n33126 = ~n33124 & ~n33125 ;
  assign n33127 = n32836 & ~n33126 ;
  assign n33128 = n32836 & ~n33127 ;
  assign n33129 = ~n33126 & ~n33127 ;
  assign n33130 = ~n33128 & ~n33129 ;
  assign n33131 = ~x123 & n1434 ;
  assign n33132 = ~x121 & n1646 ;
  assign n33133 = ~x122 & n1429 ;
  assign n33134 = ~n33132 & ~n33133 ;
  assign n33135 = ~n33131 & n33134 ;
  assign n33136 = n1437 & n23760 ;
  assign n33137 = n33135 & ~n33136 ;
  assign n33138 = ~x14 & ~n33137 ;
  assign n33139 = ~x14 & ~n33138 ;
  assign n33140 = ~n33137 & ~n33138 ;
  assign n33141 = ~n33139 & ~n33140 ;
  assign n33142 = ~n32115 & ~n32405 ;
  assign n33143 = ~n33141 & ~n33142 ;
  assign n33144 = ~n33141 & ~n33143 ;
  assign n33145 = ~n33142 & ~n33143 ;
  assign n33146 = ~n33144 & ~n33145 ;
  assign n33147 = ~n33130 & n33146 ;
  assign n33148 = n33130 & ~n33146 ;
  assign n33149 = ~n33147 & ~n33148 ;
  assign n33150 = ~n32099 & ~n32408 ;
  assign n33151 = ~x126 & n945 ;
  assign n33152 = ~x124 & n1099 ;
  assign n33153 = ~x125 & n940 ;
  assign n33154 = ~n33152 & ~n33153 ;
  assign n33155 = ~n33151 & n33154 ;
  assign n33156 = ~n948 & n33155 ;
  assign n33157 = ~n26128 & n33155 ;
  assign n33158 = ~n33156 & ~n33157 ;
  assign n33159 = ~x11 & ~n33158 ;
  assign n33160 = x11 & n33158 ;
  assign n33161 = ~n33159 & ~n33160 ;
  assign n33162 = ~n33150 & ~n33161 ;
  assign n33163 = ~n33150 & ~n33162 ;
  assign n33164 = ~n33161 & ~n33162 ;
  assign n33165 = ~n33163 & ~n33164 ;
  assign n33166 = ~n33149 & ~n33165 ;
  assign n33167 = n33149 & ~n33164 ;
  assign n33168 = ~n33163 & n33167 ;
  assign n33169 = ~n33166 & ~n33168 ;
  assign n33170 = ~n32821 & n33169 ;
  assign n33171 = n32821 & ~n33169 ;
  assign n33172 = ~n33170 & ~n33171 ;
  assign n33173 = ~n32809 & n33172 ;
  assign n33174 = ~n32809 & ~n33173 ;
  assign n33175 = n33172 & ~n33173 ;
  assign n33176 = ~n33174 & ~n33175 ;
  assign n33177 = ~n32808 & ~n33176 ;
  assign n33178 = n32808 & ~n33175 ;
  assign n33179 = ~n33174 & n33178 ;
  assign n33180 = ~n33177 & ~n33179 ;
  assign n33183 = ~n33180 & ~x199 ;
  assign n33184 = ~n33182 & ~n33183 ;
  assign n33185 = ~n32800 & ~n32804 ;
  assign n33186 = ~n32445 & ~n32797 ;
  assign n33187 = ~n32789 & ~n32793 ;
  assign n33188 = x127 & n945 ;
  assign n33189 = x125 & n1099 ;
  assign n33190 = x126 & n940 ;
  assign n33191 = ~n33189 & ~n33190 ;
  assign n33192 = ~n33188 & n33191 ;
  assign n33193 = n948 & n26533 ;
  assign n33194 = n33192 & ~n33193 ;
  assign n33195 = x11 & ~n33194 ;
  assign n33196 = x11 & ~n33195 ;
  assign n33197 = ~n33194 & ~n33195 ;
  assign n33198 = ~n33196 & ~n33197 ;
  assign n33199 = ~n33187 & ~n33198 ;
  assign n33200 = ~n33187 & ~n33199 ;
  assign n33201 = ~n33198 & ~n33199 ;
  assign n33202 = ~n33200 & ~n33201 ;
  assign n33203 = ~n32757 & ~n32773 ;
  assign n33204 = ~n32770 & ~n33203 ;
  assign n33205 = x124 & n1434 ;
  assign n33206 = x122 & n1646 ;
  assign n33207 = x123 & n1429 ;
  assign n33208 = ~n33206 & ~n33207 ;
  assign n33209 = ~n33205 & n33208 ;
  assign n33210 = n1437 & n23796 ;
  assign n33211 = n33209 & ~n33210 ;
  assign n33212 = x14 & ~n33211 ;
  assign n33213 = x14 & ~n33212 ;
  assign n33214 = ~n33211 & ~n33212 ;
  assign n33215 = ~n33213 & ~n33214 ;
  assign n33216 = ~n33204 & n33215 ;
  assign n33217 = n33204 & ~n33215 ;
  assign n33218 = ~n33216 & ~n33217 ;
  assign n33219 = x121 & n2093 ;
  assign n33220 = x119 & n2275 ;
  assign n33221 = x120 & n2088 ;
  assign n33222 = ~n33220 & ~n33221 ;
  assign n33223 = ~n33219 & n33222 ;
  assign n33224 = n2096 & n21870 ;
  assign n33225 = n33223 & ~n33224 ;
  assign n33226 = x17 & ~n33225 ;
  assign n33227 = x17 & ~n33226 ;
  assign n33228 = ~n33225 & ~n33226 ;
  assign n33229 = ~n33227 & ~n33228 ;
  assign n33230 = ~n32462 & ~n32754 ;
  assign n33231 = n33229 & n33230 ;
  assign n33232 = ~n33229 & ~n33230 ;
  assign n33233 = ~n33231 & ~n33232 ;
  assign n33234 = ~n32746 & ~n32750 ;
  assign n33235 = x118 & n2751 ;
  assign n33236 = x116 & n3020 ;
  assign n33237 = x117 & n2746 ;
  assign n33238 = ~n33236 & ~n33237 ;
  assign n33239 = ~n33235 & n33238 ;
  assign n33240 = n2754 & n19395 ;
  assign n33241 = n33239 & ~n33240 ;
  assign n33242 = x20 & ~n33241 ;
  assign n33243 = x20 & ~n33242 ;
  assign n33244 = ~n33241 & ~n33242 ;
  assign n33245 = ~n33243 & ~n33244 ;
  assign n33246 = ~n33234 & ~n33245 ;
  assign n33247 = ~n33234 & ~n33246 ;
  assign n33248 = ~n33245 & ~n33246 ;
  assign n33249 = ~n33247 & ~n33248 ;
  assign n33250 = x112 & n4531 ;
  assign n33251 = x110 & n4847 ;
  assign n33252 = x111 & n4526 ;
  assign n33253 = ~n33251 & ~n33252 ;
  assign n33254 = ~n33250 & n33253 ;
  assign n33255 = n4534 & n15442 ;
  assign n33256 = n33254 & ~n33255 ;
  assign n33257 = x26 & ~n33256 ;
  assign n33258 = x26 & ~n33257 ;
  assign n33259 = ~n33256 & ~n33257 ;
  assign n33260 = ~n33258 & ~n33259 ;
  assign n33261 = ~n32492 & ~n32726 ;
  assign n33262 = n33260 & n33261 ;
  assign n33263 = ~n33260 & ~n33261 ;
  assign n33264 = ~n33262 & ~n33263 ;
  assign n33265 = ~n32718 & ~n32722 ;
  assign n33266 = x109 & n5560 ;
  assign n33267 = x107 & n5943 ;
  assign n33268 = x108 & n5555 ;
  assign n33269 = ~n33267 & ~n33268 ;
  assign n33270 = ~n33266 & n33269 ;
  assign n33271 = n5563 & n13894 ;
  assign n33272 = n33270 & ~n33271 ;
  assign n33273 = x29 & ~n33272 ;
  assign n33274 = x29 & ~n33273 ;
  assign n33275 = ~n33272 & ~n33273 ;
  assign n33276 = ~n33274 & ~n33275 ;
  assign n33277 = ~n33265 & ~n33276 ;
  assign n33278 = ~n33265 & ~n33277 ;
  assign n33279 = ~n33276 & ~n33277 ;
  assign n33280 = ~n33278 & ~n33279 ;
  assign n33281 = ~n32509 & ~n32701 ;
  assign n33282 = x106 & n6725 ;
  assign n33283 = x104 & n7129 ;
  assign n33284 = x105 & n6720 ;
  assign n33285 = ~n33283 & ~n33284 ;
  assign n33286 = ~n33282 & n33285 ;
  assign n33287 = n6728 & n12181 ;
  assign n33288 = n33286 & ~n33287 ;
  assign n33289 = x32 & ~n33288 ;
  assign n33290 = x32 & ~n33289 ;
  assign n33291 = ~n33288 & ~n33289 ;
  assign n33292 = ~n33290 & ~n33291 ;
  assign n33293 = ~n33281 & ~n33292 ;
  assign n33294 = ~n33281 & ~n33293 ;
  assign n33295 = ~n33292 & ~n33293 ;
  assign n33296 = ~n33294 & ~n33295 ;
  assign n33297 = ~n32665 & ~n32679 ;
  assign n33298 = ~n32648 & ~n32662 ;
  assign n33299 = ~n32629 & ~n32642 ;
  assign n33300 = ~n32601 & ~n32605 ;
  assign n33301 = x88 & n16076 ;
  assign n33302 = x86 & n16756 ;
  assign n33303 = x87 & n16071 ;
  assign n33304 = ~n33302 & ~n33303 ;
  assign n33305 = ~n33301 & n33304 ;
  assign n33306 = n4305 & n16079 ;
  assign n33307 = n33305 & ~n33306 ;
  assign n33308 = x50 & ~n33307 ;
  assign n33309 = x50 & ~n33308 ;
  assign n33310 = ~n33307 & ~n33308 ;
  assign n33311 = ~n33309 & ~n33310 ;
  assign n33312 = ~n32536 & ~n32547 ;
  assign n33313 = ~n32562 & ~n33312 ;
  assign n33314 = x76 & n24612 ;
  assign n33315 = x74 & n25390 ;
  assign n33316 = x75 & n24607 ;
  assign n33317 = ~n33315 & ~n33316 ;
  assign n33318 = ~n33314 & n33317 ;
  assign n33319 = n1311 & n24615 ;
  assign n33320 = n33318 & ~n33319 ;
  assign n33321 = x62 & ~n33320 ;
  assign n33322 = x62 & ~n33321 ;
  assign n33323 = ~n33320 & ~n33321 ;
  assign n33324 = ~n33322 & ~n33323 ;
  assign n33325 = x72 & n27024 ;
  assign n33326 = x73 & ~n26217 ;
  assign n33327 = ~n33325 & ~n33326 ;
  assign n33328 = x8 & ~n32528 ;
  assign n33329 = ~x8 & n32528 ;
  assign n33330 = ~n33328 & ~n33329 ;
  assign n33331 = ~n33327 & ~n33330 ;
  assign n33332 = n33327 & n33330 ;
  assign n33333 = ~n33331 & ~n33332 ;
  assign n33334 = ~n32534 & n33333 ;
  assign n33335 = n32534 & ~n33333 ;
  assign n33336 = ~n33334 & ~n33335 ;
  assign n33337 = n33324 & n33336 ;
  assign n33338 = ~n33324 & ~n33336 ;
  assign n33339 = ~n33337 & ~n33338 ;
  assign n33340 = x79 & n22325 ;
  assign n33341 = x77 & n23066 ;
  assign n33342 = x78 & n22320 ;
  assign n33343 = ~n33341 & ~n33342 ;
  assign n33344 = ~n33340 & n33343 ;
  assign n33345 = n1817 & n22328 ;
  assign n33346 = n33344 & ~n33345 ;
  assign n33347 = x59 & ~n33346 ;
  assign n33348 = x59 & ~n33347 ;
  assign n33349 = ~n33346 & ~n33347 ;
  assign n33350 = ~n33348 & ~n33349 ;
  assign n33351 = ~n33339 & ~n33350 ;
  assign n33352 = n33339 & n33350 ;
  assign n33353 = ~n33351 & ~n33352 ;
  assign n33354 = ~n33313 & n33353 ;
  assign n33355 = n33313 & ~n33353 ;
  assign n33356 = ~n33354 & ~n33355 ;
  assign n33357 = x82 & n20143 ;
  assign n33358 = x80 & n20854 ;
  assign n33359 = x81 & n20138 ;
  assign n33360 = ~n33358 & ~n33359 ;
  assign n33361 = ~n33357 & n33360 ;
  assign n33362 = n2584 & n20146 ;
  assign n33363 = n33361 & ~n33362 ;
  assign n33364 = x56 & ~n33363 ;
  assign n33365 = x56 & ~n33364 ;
  assign n33366 = ~n33363 & ~n33364 ;
  assign n33367 = ~n33365 & ~n33366 ;
  assign n33368 = n33356 & ~n33367 ;
  assign n33369 = n33356 & ~n33368 ;
  assign n33370 = ~n33367 & ~n33368 ;
  assign n33371 = ~n33369 & ~n33370 ;
  assign n33372 = ~n32566 & ~n32579 ;
  assign n33373 = n33371 & n33372 ;
  assign n33374 = ~n33371 & ~n33372 ;
  assign n33375 = ~n33373 & ~n33374 ;
  assign n33376 = x85 & n18025 ;
  assign n33377 = x83 & n18764 ;
  assign n33378 = x84 & n18020 ;
  assign n33379 = ~n33377 & ~n33378 ;
  assign n33380 = ~n33376 & n33379 ;
  assign n33381 = n3389 & n18028 ;
  assign n33382 = n33380 & ~n33381 ;
  assign n33383 = x53 & ~n33382 ;
  assign n33384 = x53 & ~n33383 ;
  assign n33385 = ~n33382 & ~n33383 ;
  assign n33386 = ~n33384 & ~n33385 ;
  assign n33387 = n33375 & ~n33386 ;
  assign n33388 = n33375 & ~n33387 ;
  assign n33389 = ~n33386 & ~n33387 ;
  assign n33390 = ~n33388 & ~n33389 ;
  assign n33391 = ~n32585 & ~n32599 ;
  assign n33392 = ~n33390 & ~n33391 ;
  assign n33393 = n33390 & n33391 ;
  assign n33394 = ~n33392 & ~n33393 ;
  assign n33395 = ~n33311 & n33394 ;
  assign n33396 = ~n33311 & ~n33395 ;
  assign n33397 = n33394 & ~n33395 ;
  assign n33398 = ~n33396 & ~n33397 ;
  assign n33399 = ~n33300 & ~n33398 ;
  assign n33400 = ~n33300 & ~n33399 ;
  assign n33401 = ~n33398 & ~n33399 ;
  assign n33402 = ~n33400 & ~n33401 ;
  assign n33403 = x91 & n14233 ;
  assign n33404 = x89 & n14876 ;
  assign n33405 = x90 & n14228 ;
  assign n33406 = ~n33404 & ~n33405 ;
  assign n33407 = ~n33403 & n33406 ;
  assign n33408 = n5336 & n14236 ;
  assign n33409 = n33407 & ~n33408 ;
  assign n33410 = x47 & ~n33409 ;
  assign n33411 = x47 & ~n33410 ;
  assign n33412 = ~n33409 & ~n33410 ;
  assign n33413 = ~n33411 & ~n33412 ;
  assign n33414 = ~n33402 & ~n33413 ;
  assign n33415 = ~n33402 & ~n33414 ;
  assign n33416 = ~n33413 & ~n33414 ;
  assign n33417 = ~n33415 & ~n33416 ;
  assign n33418 = ~n32609 & ~n32623 ;
  assign n33419 = n33417 & n33418 ;
  assign n33420 = ~n33417 & ~n33418 ;
  assign n33421 = ~n33419 & ~n33420 ;
  assign n33422 = x94 & n12506 ;
  assign n33423 = x92 & n13131 ;
  assign n33424 = x93 & n12501 ;
  assign n33425 = ~n33423 & ~n33424 ;
  assign n33426 = ~n33422 & n33425 ;
  assign n33427 = n6483 & n12509 ;
  assign n33428 = n33426 & ~n33427 ;
  assign n33429 = x44 & ~n33428 ;
  assign n33430 = x44 & ~n33429 ;
  assign n33431 = ~n33428 & ~n33429 ;
  assign n33432 = ~n33430 & ~n33431 ;
  assign n33433 = n33421 & ~n33432 ;
  assign n33434 = ~n33421 & n33432 ;
  assign n33435 = ~n33299 & ~n33434 ;
  assign n33436 = ~n33433 & n33435 ;
  assign n33437 = ~n33299 & ~n33436 ;
  assign n33438 = ~n33433 & ~n33436 ;
  assign n33439 = ~n33434 & n33438 ;
  assign n33440 = ~n33437 & ~n33439 ;
  assign n33441 = x97 & n10905 ;
  assign n33442 = x95 & n11466 ;
  assign n33443 = x96 & n10900 ;
  assign n33444 = ~n33442 & ~n33443 ;
  assign n33445 = ~n33441 & n33444 ;
  assign n33446 = n7745 & n10908 ;
  assign n33447 = n33445 & ~n33446 ;
  assign n33448 = x41 & ~n33447 ;
  assign n33449 = x41 & ~n33448 ;
  assign n33450 = ~n33447 & ~n33448 ;
  assign n33451 = ~n33449 & ~n33450 ;
  assign n33452 = ~n33440 & ~n33451 ;
  assign n33453 = ~n33440 & ~n33452 ;
  assign n33454 = ~n33451 & ~n33452 ;
  assign n33455 = ~n33453 & ~n33454 ;
  assign n33456 = ~n33298 & n33455 ;
  assign n33457 = n33298 & ~n33455 ;
  assign n33458 = ~n33456 & ~n33457 ;
  assign n33459 = x100 & n9433 ;
  assign n33460 = x98 & n9915 ;
  assign n33461 = x99 & n9428 ;
  assign n33462 = ~n33460 & ~n33461 ;
  assign n33463 = ~n33459 & n33462 ;
  assign n33464 = n9115 & n9436 ;
  assign n33465 = n33463 & ~n33464 ;
  assign n33466 = x38 & ~n33465 ;
  assign n33467 = x38 & ~n33466 ;
  assign n33468 = ~n33465 & ~n33466 ;
  assign n33469 = ~n33467 & ~n33468 ;
  assign n33470 = ~n33458 & ~n33469 ;
  assign n33471 = n33458 & n33469 ;
  assign n33472 = ~n33470 & ~n33471 ;
  assign n33473 = n33297 & ~n33472 ;
  assign n33474 = ~n33297 & n33472 ;
  assign n33475 = ~n33473 & ~n33474 ;
  assign n33476 = x103 & n8006 ;
  assign n33477 = x101 & n8474 ;
  assign n33478 = x102 & n8001 ;
  assign n33479 = ~n33477 & ~n33478 ;
  assign n33480 = ~n33476 & n33479 ;
  assign n33481 = n8009 & n10588 ;
  assign n33482 = n33480 & ~n33481 ;
  assign n33483 = x35 & ~n33482 ;
  assign n33484 = x35 & ~n33483 ;
  assign n33485 = ~n33482 & ~n33483 ;
  assign n33486 = ~n33484 & ~n33485 ;
  assign n33487 = n33475 & ~n33486 ;
  assign n33488 = n33475 & ~n33487 ;
  assign n33489 = ~n33486 & ~n33487 ;
  assign n33490 = ~n33488 & ~n33489 ;
  assign n33491 = ~n32685 & ~n32698 ;
  assign n33492 = ~n33490 & ~n33491 ;
  assign n33493 = ~n33490 & ~n33492 ;
  assign n33494 = ~n33491 & ~n33492 ;
  assign n33495 = ~n33493 & ~n33494 ;
  assign n33496 = ~n33296 & ~n33495 ;
  assign n33497 = ~n33296 & ~n33496 ;
  assign n33498 = ~n33495 & ~n33496 ;
  assign n33499 = ~n33497 & ~n33498 ;
  assign n33500 = ~n33280 & n33499 ;
  assign n33501 = n33280 & ~n33499 ;
  assign n33502 = ~n33500 & ~n33501 ;
  assign n33503 = n33264 & ~n33502 ;
  assign n33504 = n33264 & ~n33503 ;
  assign n33505 = ~n33502 & ~n33503 ;
  assign n33506 = ~n33504 & ~n33505 ;
  assign n33507 = x115 & n3589 ;
  assign n33508 = x113 & n3878 ;
  assign n33509 = x114 & n3584 ;
  assign n33510 = ~n33508 & ~n33509 ;
  assign n33511 = ~n33507 & n33510 ;
  assign n33512 = n3592 & n17364 ;
  assign n33513 = n33511 & ~n33512 ;
  assign n33514 = x23 & ~n33513 ;
  assign n33515 = x23 & ~n33514 ;
  assign n33516 = ~n33513 & ~n33514 ;
  assign n33517 = ~n33515 & ~n33516 ;
  assign n33518 = ~n32477 & ~n32731 ;
  assign n33519 = ~n33517 & ~n33518 ;
  assign n33520 = n33517 & n33518 ;
  assign n33521 = ~n33519 & ~n33520 ;
  assign n33522 = ~n33506 & n33521 ;
  assign n33523 = ~n33506 & ~n33522 ;
  assign n33524 = n33521 & ~n33522 ;
  assign n33525 = ~n33523 & ~n33524 ;
  assign n33526 = ~n33249 & ~n33525 ;
  assign n33527 = ~n33249 & ~n33526 ;
  assign n33528 = ~n33525 & ~n33526 ;
  assign n33529 = ~n33527 & ~n33528 ;
  assign n33530 = n33233 & ~n33529 ;
  assign n33531 = ~n33233 & n33529 ;
  assign n33532 = ~n33218 & ~n33531 ;
  assign n33533 = ~n33530 & n33532 ;
  assign n33534 = ~n33218 & ~n33533 ;
  assign n33535 = ~n33531 & ~n33533 ;
  assign n33536 = ~n33530 & n33535 ;
  assign n33537 = ~n33534 & ~n33536 ;
  assign n33538 = ~n33202 & n33537 ;
  assign n33539 = n33202 & ~n33537 ;
  assign n33540 = ~n33538 & ~n33539 ;
  assign n33541 = ~n33186 & ~n33540 ;
  assign n33542 = ~n33186 & ~n33541 ;
  assign n33543 = ~n33540 & ~n33541 ;
  assign n33544 = ~n33542 & ~n33543 ;
  assign n33545 = ~n33185 & ~n33544 ;
  assign n33546 = n33185 & ~n33543 ;
  assign n33547 = ~n33542 & n33546 ;
  assign n33548 = ~n33545 & ~n33547 ;
  assign n33914 = n33548 & x200 ;
  assign n33549 = ~n33173 & ~n33177 ;
  assign n33550 = ~n32818 & ~n33170 ;
  assign n33551 = ~n33162 & ~n33166 ;
  assign n33552 = ~x127 & n945 ;
  assign n33553 = ~x125 & n1099 ;
  assign n33554 = ~x126 & n940 ;
  assign n33555 = ~n33553 & ~n33554 ;
  assign n33556 = ~n33552 & n33555 ;
  assign n33557 = n948 & n26932 ;
  assign n33558 = n33556 & ~n33557 ;
  assign n33559 = ~x11 & ~n33558 ;
  assign n33560 = ~x11 & ~n33559 ;
  assign n33561 = ~n33558 & ~n33559 ;
  assign n33562 = ~n33560 & ~n33561 ;
  assign n33563 = ~n33551 & ~n33562 ;
  assign n33564 = ~n33551 & ~n33563 ;
  assign n33565 = ~n33562 & ~n33563 ;
  assign n33566 = ~n33564 & ~n33565 ;
  assign n33567 = ~n33130 & ~n33146 ;
  assign n33568 = ~n33143 & ~n33567 ;
  assign n33569 = ~x124 & n1434 ;
  assign n33570 = ~x122 & n1646 ;
  assign n33571 = ~x123 & n1429 ;
  assign n33572 = ~n33570 & ~n33571 ;
  assign n33573 = ~n33569 & n33572 ;
  assign n33574 = n1437 & n24176 ;
  assign n33575 = n33573 & ~n33574 ;
  assign n33576 = ~x14 & ~n33575 ;
  assign n33577 = ~x14 & ~n33576 ;
  assign n33578 = ~n33575 & ~n33576 ;
  assign n33579 = ~n33577 & ~n33578 ;
  assign n33580 = ~n33568 & n33579 ;
  assign n33581 = n33568 & ~n33579 ;
  assign n33582 = ~n33580 & ~n33581 ;
  assign n33583 = ~x121 & n2093 ;
  assign n33584 = ~x119 & n2275 ;
  assign n33585 = ~x120 & n2088 ;
  assign n33586 = ~n33584 & ~n33585 ;
  assign n33587 = ~n33583 & n33586 ;
  assign n33588 = n2096 & n22229 ;
  assign n33589 = n33587 & ~n33588 ;
  assign n33590 = ~x17 & ~n33589 ;
  assign n33591 = ~x17 & ~n33590 ;
  assign n33592 = ~n33589 & ~n33590 ;
  assign n33593 = ~n33591 & ~n33592 ;
  assign n33594 = ~n32835 & ~n33127 ;
  assign n33595 = n33593 & n33594 ;
  assign n33596 = ~n33593 & ~n33594 ;
  assign n33597 = ~n33595 & ~n33596 ;
  assign n33598 = ~n33119 & ~n33123 ;
  assign n33599 = ~x118 & n2751 ;
  assign n33600 = ~x116 & n3020 ;
  assign n33601 = ~x117 & n2746 ;
  assign n33602 = ~n33600 & ~n33601 ;
  assign n33603 = ~n33599 & n33602 ;
  assign n33604 = n2754 & n19736 ;
  assign n33605 = n33603 & ~n33604 ;
  assign n33606 = ~x20 & ~n33605 ;
  assign n33607 = ~x20 & ~n33606 ;
  assign n33608 = ~n33605 & ~n33606 ;
  assign n33609 = ~n33607 & ~n33608 ;
  assign n33610 = ~n33598 & ~n33609 ;
  assign n33611 = ~n33598 & ~n33610 ;
  assign n33612 = ~n33609 & ~n33610 ;
  assign n33613 = ~n33611 & ~n33612 ;
  assign n33614 = ~x112 & n4531 ;
  assign n33615 = ~x110 & n4847 ;
  assign n33616 = ~x111 & n4526 ;
  assign n33617 = ~n33615 & ~n33616 ;
  assign n33618 = ~n33614 & n33617 ;
  assign n33619 = n4534 & n15744 ;
  assign n33620 = n33618 & ~n33619 ;
  assign n33621 = ~x26 & ~n33620 ;
  assign n33622 = ~x26 & ~n33621 ;
  assign n33623 = ~n33620 & ~n33621 ;
  assign n33624 = ~n33622 & ~n33623 ;
  assign n33625 = ~n32865 & ~n33099 ;
  assign n33626 = n33624 & n33625 ;
  assign n33627 = ~n33624 & ~n33625 ;
  assign n33628 = ~n33626 & ~n33627 ;
  assign n33629 = ~n33091 & ~n33095 ;
  assign n33630 = ~x109 & n5560 ;
  assign n33631 = ~x107 & n5943 ;
  assign n33632 = ~x108 & n5555 ;
  assign n33633 = ~n33631 & ~n33632 ;
  assign n33634 = ~n33630 & n33633 ;
  assign n33635 = n5563 & n14177 ;
  assign n33636 = n33634 & ~n33635 ;
  assign n33637 = ~x29 & ~n33636 ;
  assign n33638 = ~x29 & ~n33637 ;
  assign n33639 = ~n33636 & ~n33637 ;
  assign n33640 = ~n33638 & ~n33639 ;
  assign n33641 = ~n33629 & ~n33640 ;
  assign n33642 = ~n33629 & ~n33641 ;
  assign n33643 = ~n33640 & ~n33641 ;
  assign n33644 = ~n33642 & ~n33643 ;
  assign n33645 = ~n32882 & ~n33074 ;
  assign n33646 = ~x106 & n6725 ;
  assign n33647 = ~x104 & n7129 ;
  assign n33648 = ~x105 & n6720 ;
  assign n33649 = ~n33647 & ~n33648 ;
  assign n33650 = ~n33646 & n33649 ;
  assign n33651 = n6728 & n12447 ;
  assign n33652 = n33650 & ~n33651 ;
  assign n33653 = ~x32 & ~n33652 ;
  assign n33654 = ~x32 & ~n33653 ;
  assign n33655 = ~n33652 & ~n33653 ;
  assign n33656 = ~n33654 & ~n33655 ;
  assign n33657 = ~n33645 & ~n33656 ;
  assign n33658 = ~n33645 & ~n33657 ;
  assign n33659 = ~n33656 & ~n33657 ;
  assign n33660 = ~n33658 & ~n33659 ;
  assign n33661 = ~n33038 & ~n33052 ;
  assign n33662 = ~n33021 & ~n33035 ;
  assign n33663 = ~n33002 & ~n33015 ;
  assign n33664 = ~n32974 & ~n32978 ;
  assign n33665 = ~x88 & n16076 ;
  assign n33666 = ~x86 & n16756 ;
  assign n33667 = ~x87 & n16071 ;
  assign n33668 = ~n33666 & ~n33667 ;
  assign n33669 = ~n33665 & n33668 ;
  assign n33670 = n4457 & n16079 ;
  assign n33671 = n33669 & ~n33670 ;
  assign n33672 = ~x50 & ~n33671 ;
  assign n33673 = ~x50 & ~n33672 ;
  assign n33674 = ~n33671 & ~n33672 ;
  assign n33675 = ~n33673 & ~n33674 ;
  assign n33676 = ~n32909 & ~n32920 ;
  assign n33677 = ~n32935 & ~n33676 ;
  assign n33678 = ~x76 & n24612 ;
  assign n33679 = ~x74 & n25390 ;
  assign n33680 = ~x75 & n24607 ;
  assign n33681 = ~n33679 & ~n33680 ;
  assign n33682 = ~n33678 & n33681 ;
  assign n33683 = n1390 & n24615 ;
  assign n33684 = n33682 & ~n33683 ;
  assign n33685 = ~x62 & ~n33684 ;
  assign n33686 = ~x62 & ~n33685 ;
  assign n33687 = ~n33684 & ~n33685 ;
  assign n33688 = ~n33686 & ~n33687 ;
  assign n33689 = ~x72 & n27427 ;
  assign n33690 = ~x73 & ~n26217 ;
  assign n33691 = ~n33689 & ~n33690 ;
  assign n33692 = ~x8 & ~n32901 ;
  assign n33693 = x8 & n32901 ;
  assign n33694 = ~n33692 & ~n33693 ;
  assign n33695 = ~n33691 & ~n33694 ;
  assign n33696 = n33691 & n33694 ;
  assign n33697 = ~n33695 & ~n33696 ;
  assign n33698 = ~n32907 & n33697 ;
  assign n33699 = n32907 & ~n33697 ;
  assign n33700 = ~n33698 & ~n33699 ;
  assign n33701 = n33688 & n33700 ;
  assign n33702 = ~n33688 & ~n33700 ;
  assign n33703 = ~n33701 & ~n33702 ;
  assign n33704 = ~x79 & n22325 ;
  assign n33705 = ~x77 & n23066 ;
  assign n33706 = ~x78 & n22320 ;
  assign n33707 = ~n33705 & ~n33706 ;
  assign n33708 = ~n33704 & n33707 ;
  assign n33709 = n1921 & n22328 ;
  assign n33710 = n33708 & ~n33709 ;
  assign n33711 = ~x59 & ~n33710 ;
  assign n33712 = ~x59 & ~n33711 ;
  assign n33713 = ~n33710 & ~n33711 ;
  assign n33714 = ~n33712 & ~n33713 ;
  assign n33715 = ~n33703 & ~n33714 ;
  assign n33716 = n33703 & n33714 ;
  assign n33717 = ~n33715 & ~n33716 ;
  assign n33718 = ~n33677 & n33717 ;
  assign n33719 = n33677 & ~n33717 ;
  assign n33720 = ~n33718 & ~n33719 ;
  assign n33721 = ~x82 & n20143 ;
  assign n33722 = ~x80 & n20854 ;
  assign n33723 = ~x81 & n20138 ;
  assign n33724 = ~n33722 & ~n33723 ;
  assign n33725 = ~n33721 & n33724 ;
  assign n33726 = n2697 & n20146 ;
  assign n33727 = n33725 & ~n33726 ;
  assign n33728 = ~x56 & ~n33727 ;
  assign n33729 = ~x56 & ~n33728 ;
  assign n33730 = ~n33727 & ~n33728 ;
  assign n33731 = ~n33729 & ~n33730 ;
  assign n33732 = n33720 & ~n33731 ;
  assign n33733 = n33720 & ~n33732 ;
  assign n33734 = ~n33731 & ~n33732 ;
  assign n33735 = ~n33733 & ~n33734 ;
  assign n33736 = ~n32939 & ~n32952 ;
  assign n33737 = n33735 & n33736 ;
  assign n33738 = ~n33735 & ~n33736 ;
  assign n33739 = ~n33737 & ~n33738 ;
  assign n33740 = ~x85 & n18025 ;
  assign n33741 = ~x83 & n18764 ;
  assign n33742 = ~x84 & n18020 ;
  assign n33743 = ~n33741 & ~n33742 ;
  assign n33744 = ~n33740 & n33743 ;
  assign n33745 = n3521 & n18028 ;
  assign n33746 = n33744 & ~n33745 ;
  assign n33747 = ~x53 & ~n33746 ;
  assign n33748 = ~x53 & ~n33747 ;
  assign n33749 = ~n33746 & ~n33747 ;
  assign n33750 = ~n33748 & ~n33749 ;
  assign n33751 = n33739 & ~n33750 ;
  assign n33752 = n33739 & ~n33751 ;
  assign n33753 = ~n33750 & ~n33751 ;
  assign n33754 = ~n33752 & ~n33753 ;
  assign n33755 = ~n32958 & ~n32972 ;
  assign n33756 = ~n33754 & ~n33755 ;
  assign n33757 = n33754 & n33755 ;
  assign n33758 = ~n33756 & ~n33757 ;
  assign n33759 = ~n33675 & n33758 ;
  assign n33760 = ~n33675 & ~n33759 ;
  assign n33761 = n33758 & ~n33759 ;
  assign n33762 = ~n33760 & ~n33761 ;
  assign n33763 = ~n33664 & ~n33762 ;
  assign n33764 = ~n33664 & ~n33763 ;
  assign n33765 = ~n33762 & ~n33763 ;
  assign n33766 = ~n33764 & ~n33765 ;
  assign n33767 = ~x91 & n14233 ;
  assign n33768 = ~x89 & n14876 ;
  assign n33769 = ~x90 & n14228 ;
  assign n33770 = ~n33768 & ~n33769 ;
  assign n33771 = ~n33767 & n33770 ;
  assign n33772 = n5507 & n14236 ;
  assign n33773 = n33771 & ~n33772 ;
  assign n33774 = ~x47 & ~n33773 ;
  assign n33775 = ~x47 & ~n33774 ;
  assign n33776 = ~n33773 & ~n33774 ;
  assign n33777 = ~n33775 & ~n33776 ;
  assign n33778 = ~n33766 & ~n33777 ;
  assign n33779 = ~n33766 & ~n33778 ;
  assign n33780 = ~n33777 & ~n33778 ;
  assign n33781 = ~n33779 & ~n33780 ;
  assign n33782 = ~n32982 & ~n32996 ;
  assign n33783 = n33781 & n33782 ;
  assign n33784 = ~n33781 & ~n33782 ;
  assign n33785 = ~n33783 & ~n33784 ;
  assign n33786 = ~x94 & n12506 ;
  assign n33787 = ~x92 & n13131 ;
  assign n33788 = ~x93 & n12501 ;
  assign n33789 = ~n33787 & ~n33788 ;
  assign n33790 = ~n33786 & n33789 ;
  assign n33791 = n6671 & n12509 ;
  assign n33792 = n33790 & ~n33791 ;
  assign n33793 = ~x44 & ~n33792 ;
  assign n33794 = ~x44 & ~n33793 ;
  assign n33795 = ~n33792 & ~n33793 ;
  assign n33796 = ~n33794 & ~n33795 ;
  assign n33797 = n33785 & ~n33796 ;
  assign n33798 = ~n33785 & n33796 ;
  assign n33799 = ~n33663 & ~n33798 ;
  assign n33800 = ~n33797 & n33799 ;
  assign n33801 = ~n33663 & ~n33800 ;
  assign n33802 = ~n33797 & ~n33800 ;
  assign n33803 = ~n33798 & n33802 ;
  assign n33804 = ~n33801 & ~n33803 ;
  assign n33805 = ~x97 & n10905 ;
  assign n33806 = ~x95 & n11466 ;
  assign n33807 = ~x96 & n10900 ;
  assign n33808 = ~n33806 & ~n33807 ;
  assign n33809 = ~n33805 & n33808 ;
  assign n33810 = n7949 & n10908 ;
  assign n33811 = n33809 & ~n33810 ;
  assign n33812 = ~x41 & ~n33811 ;
  assign n33813 = ~x41 & ~n33812 ;
  assign n33814 = ~n33811 & ~n33812 ;
  assign n33815 = ~n33813 & ~n33814 ;
  assign n33816 = ~n33804 & ~n33815 ;
  assign n33817 = ~n33804 & ~n33816 ;
  assign n33818 = ~n33815 & ~n33816 ;
  assign n33819 = ~n33817 & ~n33818 ;
  assign n33820 = ~n33662 & n33819 ;
  assign n33821 = n33662 & ~n33819 ;
  assign n33822 = ~n33820 & ~n33821 ;
  assign n33823 = ~x100 & n9433 ;
  assign n33824 = ~x98 & n9915 ;
  assign n33825 = ~x99 & n9428 ;
  assign n33826 = ~n33824 & ~n33825 ;
  assign n33827 = ~n33823 & n33826 ;
  assign n33828 = n9338 & n9436 ;
  assign n33829 = n33827 & ~n33828 ;
  assign n33830 = ~x38 & ~n33829 ;
  assign n33831 = ~x38 & ~n33830 ;
  assign n33832 = ~n33829 & ~n33830 ;
  assign n33833 = ~n33831 & ~n33832 ;
  assign n33834 = ~n33822 & ~n33833 ;
  assign n33835 = n33822 & n33833 ;
  assign n33836 = ~n33834 & ~n33835 ;
  assign n33837 = n33661 & ~n33836 ;
  assign n33838 = ~n33661 & n33836 ;
  assign n33839 = ~n33837 & ~n33838 ;
  assign n33840 = ~x103 & n8006 ;
  assign n33841 = ~x101 & n8474 ;
  assign n33842 = ~x102 & n8001 ;
  assign n33843 = ~n33841 & ~n33842 ;
  assign n33844 = ~n33840 & n33843 ;
  assign n33845 = n8009 & n10833 ;
  assign n33846 = n33844 & ~n33845 ;
  assign n33847 = ~x35 & ~n33846 ;
  assign n33848 = ~x35 & ~n33847 ;
  assign n33849 = ~n33846 & ~n33847 ;
  assign n33850 = ~n33848 & ~n33849 ;
  assign n33851 = n33839 & ~n33850 ;
  assign n33852 = n33839 & ~n33851 ;
  assign n33853 = ~n33850 & ~n33851 ;
  assign n33854 = ~n33852 & ~n33853 ;
  assign n33855 = ~n33058 & ~n33071 ;
  assign n33856 = ~n33854 & ~n33855 ;
  assign n33857 = ~n33854 & ~n33856 ;
  assign n33858 = ~n33855 & ~n33856 ;
  assign n33859 = ~n33857 & ~n33858 ;
  assign n33860 = ~n33660 & ~n33859 ;
  assign n33861 = ~n33660 & ~n33860 ;
  assign n33862 = ~n33859 & ~n33860 ;
  assign n33863 = ~n33861 & ~n33862 ;
  assign n33864 = ~n33644 & n33863 ;
  assign n33865 = n33644 & ~n33863 ;
  assign n33866 = ~n33864 & ~n33865 ;
  assign n33867 = n33628 & ~n33866 ;
  assign n33868 = n33628 & ~n33867 ;
  assign n33869 = ~n33866 & ~n33867 ;
  assign n33870 = ~n33868 & ~n33869 ;
  assign n33871 = ~x115 & n3589 ;
  assign n33872 = ~x113 & n3878 ;
  assign n33873 = ~x114 & n3584 ;
  assign n33874 = ~n33872 & ~n33873 ;
  assign n33875 = ~n33871 & n33874 ;
  assign n33876 = n3592 & n17683 ;
  assign n33877 = n33875 & ~n33876 ;
  assign n33878 = ~x23 & ~n33877 ;
  assign n33879 = ~x23 & ~n33878 ;
  assign n33880 = ~n33877 & ~n33878 ;
  assign n33881 = ~n33879 & ~n33880 ;
  assign n33882 = ~n32850 & ~n33104 ;
  assign n33883 = ~n33881 & ~n33882 ;
  assign n33884 = n33881 & n33882 ;
  assign n33885 = ~n33883 & ~n33884 ;
  assign n33886 = ~n33870 & n33885 ;
  assign n33887 = ~n33870 & ~n33886 ;
  assign n33888 = n33885 & ~n33886 ;
  assign n33889 = ~n33887 & ~n33888 ;
  assign n33890 = ~n33613 & ~n33889 ;
  assign n33891 = ~n33613 & ~n33890 ;
  assign n33892 = ~n33889 & ~n33890 ;
  assign n33893 = ~n33891 & ~n33892 ;
  assign n33894 = n33597 & ~n33893 ;
  assign n33895 = ~n33597 & n33893 ;
  assign n33896 = ~n33582 & ~n33895 ;
  assign n33897 = ~n33894 & n33896 ;
  assign n33898 = ~n33582 & ~n33897 ;
  assign n33899 = ~n33895 & ~n33897 ;
  assign n33900 = ~n33894 & n33899 ;
  assign n33901 = ~n33898 & ~n33900 ;
  assign n33902 = ~n33566 & n33901 ;
  assign n33903 = n33566 & ~n33901 ;
  assign n33904 = ~n33902 & ~n33903 ;
  assign n33905 = ~n33550 & ~n33904 ;
  assign n33906 = ~n33550 & ~n33905 ;
  assign n33907 = ~n33904 & ~n33905 ;
  assign n33908 = ~n33906 & ~n33907 ;
  assign n33909 = ~n33549 & ~n33908 ;
  assign n33910 = n33549 & ~n33907 ;
  assign n33911 = ~n33906 & n33910 ;
  assign n33912 = ~n33909 & ~n33911 ;
  assign n33915 = ~n33912 & ~x200 ;
  assign n33916 = ~n33914 & ~n33915 ;
  assign n33917 = ~n33541 & ~n33545 ;
  assign n33918 = ~n33202 & ~n33537 ;
  assign n33919 = ~n33199 & ~n33918 ;
  assign n33920 = x125 & n1434 ;
  assign n33921 = x123 & n1646 ;
  assign n33922 = x124 & n1429 ;
  assign n33923 = ~n33921 & ~n33922 ;
  assign n33924 = ~n33920 & n33923 ;
  assign n33925 = n1437 & n24935 ;
  assign n33926 = n33924 & ~n33925 ;
  assign n33927 = x14 & ~n33926 ;
  assign n33928 = x14 & ~n33927 ;
  assign n33929 = ~n33926 & ~n33927 ;
  assign n33930 = ~n33928 & ~n33929 ;
  assign n33931 = ~n33232 & ~n33530 ;
  assign n33932 = ~n33930 & ~n33931 ;
  assign n33933 = ~n33930 & ~n33932 ;
  assign n33934 = ~n33931 & ~n33932 ;
  assign n33935 = ~n33933 & ~n33934 ;
  assign n33936 = x119 & n2751 ;
  assign n33937 = x117 & n3020 ;
  assign n33938 = x118 & n2746 ;
  assign n33939 = ~n33937 & ~n33938 ;
  assign n33940 = ~n33936 & n33939 ;
  assign n33941 = n2754 & n20423 ;
  assign n33942 = n33940 & ~n33941 ;
  assign n33943 = x20 & ~n33942 ;
  assign n33944 = x20 & ~n33943 ;
  assign n33945 = ~n33942 & ~n33943 ;
  assign n33946 = ~n33944 & ~n33945 ;
  assign n33947 = ~n33519 & ~n33522 ;
  assign n33948 = n33946 & n33947 ;
  assign n33949 = ~n33946 & ~n33947 ;
  assign n33950 = ~n33948 & ~n33949 ;
  assign n33951 = x116 & n3589 ;
  assign n33952 = x114 & n3878 ;
  assign n33953 = x115 & n3584 ;
  assign n33954 = ~n33952 & ~n33953 ;
  assign n33955 = ~n33951 & n33954 ;
  assign n33956 = n3592 & n18336 ;
  assign n33957 = n33955 & ~n33956 ;
  assign n33958 = x23 & ~n33957 ;
  assign n33959 = x23 & ~n33958 ;
  assign n33960 = ~n33957 & ~n33958 ;
  assign n33961 = ~n33959 & ~n33960 ;
  assign n33962 = ~n33263 & ~n33503 ;
  assign n33963 = n33961 & n33962 ;
  assign n33964 = ~n33961 & ~n33962 ;
  assign n33965 = ~n33963 & ~n33964 ;
  assign n33966 = x113 & n4531 ;
  assign n33967 = x111 & n4847 ;
  assign n33968 = x112 & n4526 ;
  assign n33969 = ~n33967 & ~n33968 ;
  assign n33970 = ~n33966 & n33969 ;
  assign n33971 = n4534 & n16361 ;
  assign n33972 = n33970 & ~n33971 ;
  assign n33973 = x26 & ~n33972 ;
  assign n33974 = x26 & ~n33973 ;
  assign n33975 = ~n33972 & ~n33973 ;
  assign n33976 = ~n33974 & ~n33975 ;
  assign n33977 = ~n33280 & ~n33499 ;
  assign n33978 = ~n33277 & ~n33977 ;
  assign n33979 = ~n33976 & ~n33978 ;
  assign n33980 = ~n33976 & ~n33979 ;
  assign n33981 = ~n33978 & ~n33979 ;
  assign n33982 = ~n33980 & ~n33981 ;
  assign n33983 = x107 & n6725 ;
  assign n33984 = x105 & n7129 ;
  assign n33985 = x106 & n6720 ;
  assign n33986 = ~n33984 & ~n33985 ;
  assign n33987 = ~n33983 & n33986 ;
  assign n33988 = n6728 & n12749 ;
  assign n33989 = n33987 & ~n33988 ;
  assign n33990 = x32 & ~n33989 ;
  assign n33991 = x32 & ~n33990 ;
  assign n33992 = ~n33989 & ~n33990 ;
  assign n33993 = ~n33991 & ~n33992 ;
  assign n33994 = ~n33487 & ~n33492 ;
  assign n33995 = n33993 & n33994 ;
  assign n33996 = ~n33993 & ~n33994 ;
  assign n33997 = ~n33995 & ~n33996 ;
  assign n33998 = x104 & n8006 ;
  assign n33999 = x102 & n8474 ;
  assign n34000 = x103 & n8001 ;
  assign n34001 = ~n33999 & ~n34000 ;
  assign n34002 = ~n33998 & n34001 ;
  assign n34003 = n8009 & n11116 ;
  assign n34004 = n34002 & ~n34003 ;
  assign n34005 = x35 & ~n34004 ;
  assign n34006 = x35 & ~n34005 ;
  assign n34007 = ~n34004 & ~n34005 ;
  assign n34008 = ~n34006 & ~n34007 ;
  assign n34009 = ~n33470 & ~n33474 ;
  assign n34010 = x101 & n9433 ;
  assign n34011 = x99 & n9915 ;
  assign n34012 = x100 & n9428 ;
  assign n34013 = ~n34011 & ~n34012 ;
  assign n34014 = ~n34010 & n34013 ;
  assign n34015 = n9436 & n9601 ;
  assign n34016 = n34014 & ~n34015 ;
  assign n34017 = x38 & ~n34016 ;
  assign n34018 = x38 & ~n34017 ;
  assign n34019 = ~n34016 & ~n34017 ;
  assign n34020 = ~n34018 & ~n34019 ;
  assign n34021 = ~n33298 & ~n33455 ;
  assign n34022 = ~n33452 & ~n34021 ;
  assign n34023 = x98 & n10905 ;
  assign n34024 = x96 & n11466 ;
  assign n34025 = x97 & n10900 ;
  assign n34026 = ~n34024 & ~n34025 ;
  assign n34027 = ~n34023 & n34026 ;
  assign n34028 = n8196 & n10908 ;
  assign n34029 = n34027 & ~n34028 ;
  assign n34030 = x41 & ~n34029 ;
  assign n34031 = x41 & ~n34030 ;
  assign n34032 = ~n34029 & ~n34030 ;
  assign n34033 = ~n34031 & ~n34032 ;
  assign n34034 = x77 & n24612 ;
  assign n34035 = x75 & n25390 ;
  assign n34036 = x76 & n24607 ;
  assign n34037 = ~n34035 & ~n34036 ;
  assign n34038 = ~n34034 & n34037 ;
  assign n34039 = n1502 & n24615 ;
  assign n34040 = n34038 & ~n34039 ;
  assign n34041 = x62 & ~n34040 ;
  assign n34042 = x62 & ~n34041 ;
  assign n34043 = ~n34040 & ~n34041 ;
  assign n34044 = ~n34042 & ~n34043 ;
  assign n34045 = x73 & n27024 ;
  assign n34046 = x74 & ~n26217 ;
  assign n34047 = ~n34045 & ~n34046 ;
  assign n34048 = ~x8 & ~n32528 ;
  assign n34049 = ~n33331 & ~n34048 ;
  assign n34050 = n34047 & ~n34049 ;
  assign n34051 = n34047 & ~n34050 ;
  assign n34052 = ~n34049 & ~n34050 ;
  assign n34053 = ~n34051 & ~n34052 ;
  assign n34054 = ~n34044 & ~n34053 ;
  assign n34055 = ~n34044 & ~n34054 ;
  assign n34056 = ~n34053 & ~n34054 ;
  assign n34057 = ~n34055 & ~n34056 ;
  assign n34058 = ~n33324 & n33336 ;
  assign n34059 = ~n33334 & ~n34058 ;
  assign n34060 = ~n34057 & ~n34059 ;
  assign n34061 = ~n34057 & ~n34060 ;
  assign n34062 = ~n34059 & ~n34060 ;
  assign n34063 = ~n34061 & ~n34062 ;
  assign n34064 = x80 & n22325 ;
  assign n34065 = x78 & n23066 ;
  assign n34066 = x79 & n22320 ;
  assign n34067 = ~n34065 & ~n34066 ;
  assign n34068 = ~n34064 & n34067 ;
  assign n34069 = n2028 & n22328 ;
  assign n34070 = n34068 & ~n34069 ;
  assign n34071 = x59 & ~n34070 ;
  assign n34072 = x59 & ~n34071 ;
  assign n34073 = ~n34070 & ~n34071 ;
  assign n34074 = ~n34072 & ~n34073 ;
  assign n34075 = ~n34063 & ~n34074 ;
  assign n34076 = ~n34063 & ~n34075 ;
  assign n34077 = ~n34074 & ~n34075 ;
  assign n34078 = ~n34076 & ~n34077 ;
  assign n34079 = ~n33351 & ~n33354 ;
  assign n34080 = n34078 & n34079 ;
  assign n34081 = ~n34078 & ~n34079 ;
  assign n34082 = ~n34080 & ~n34081 ;
  assign n34083 = x83 & n20143 ;
  assign n34084 = x81 & n20854 ;
  assign n34085 = x82 & n20138 ;
  assign n34086 = ~n34084 & ~n34085 ;
  assign n34087 = ~n34083 & n34086 ;
  assign n34088 = n2843 & n20146 ;
  assign n34089 = n34087 & ~n34088 ;
  assign n34090 = x56 & ~n34089 ;
  assign n34091 = x56 & ~n34090 ;
  assign n34092 = ~n34089 & ~n34090 ;
  assign n34093 = ~n34091 & ~n34092 ;
  assign n34094 = n34082 & ~n34093 ;
  assign n34095 = n34082 & ~n34094 ;
  assign n34096 = ~n34093 & ~n34094 ;
  assign n34097 = ~n34095 & ~n34096 ;
  assign n34098 = ~n33368 & ~n33374 ;
  assign n34099 = n34097 & n34098 ;
  assign n34100 = ~n34097 & ~n34098 ;
  assign n34101 = ~n34099 & ~n34100 ;
  assign n34102 = x86 & n18025 ;
  assign n34103 = x84 & n18764 ;
  assign n34104 = x85 & n18020 ;
  assign n34105 = ~n34103 & ~n34104 ;
  assign n34106 = ~n34102 & n34105 ;
  assign n34107 = n3686 & n18028 ;
  assign n34108 = n34106 & ~n34107 ;
  assign n34109 = x53 & ~n34108 ;
  assign n34110 = x53 & ~n34109 ;
  assign n34111 = ~n34108 & ~n34109 ;
  assign n34112 = ~n34110 & ~n34111 ;
  assign n34113 = n34101 & ~n34112 ;
  assign n34114 = n34101 & ~n34113 ;
  assign n34115 = ~n34112 & ~n34113 ;
  assign n34116 = ~n34114 & ~n34115 ;
  assign n34117 = ~n33387 & ~n33392 ;
  assign n34118 = n34116 & n34117 ;
  assign n34119 = ~n34116 & ~n34117 ;
  assign n34120 = ~n34118 & ~n34119 ;
  assign n34121 = x89 & n16076 ;
  assign n34122 = x87 & n16756 ;
  assign n34123 = x88 & n16071 ;
  assign n34124 = ~n34122 & ~n34123 ;
  assign n34125 = ~n34121 & n34124 ;
  assign n34126 = n4488 & n16079 ;
  assign n34127 = n34125 & ~n34126 ;
  assign n34128 = x50 & ~n34127 ;
  assign n34129 = x50 & ~n34128 ;
  assign n34130 = ~n34127 & ~n34128 ;
  assign n34131 = ~n34129 & ~n34130 ;
  assign n34132 = n34120 & ~n34131 ;
  assign n34133 = n34120 & ~n34132 ;
  assign n34134 = ~n34131 & ~n34132 ;
  assign n34135 = ~n34133 & ~n34134 ;
  assign n34136 = ~n33395 & ~n33399 ;
  assign n34137 = n34135 & n34136 ;
  assign n34138 = ~n34135 & ~n34136 ;
  assign n34139 = ~n34137 & ~n34138 ;
  assign n34140 = x92 & n14233 ;
  assign n34141 = x90 & n14876 ;
  assign n34142 = x91 & n14228 ;
  assign n34143 = ~n34141 & ~n34142 ;
  assign n34144 = ~n34140 & n34143 ;
  assign n34145 = n5710 & n14236 ;
  assign n34146 = n34144 & ~n34145 ;
  assign n34147 = x47 & ~n34146 ;
  assign n34148 = x47 & ~n34147 ;
  assign n34149 = ~n34146 & ~n34147 ;
  assign n34150 = ~n34148 & ~n34149 ;
  assign n34151 = n34139 & ~n34150 ;
  assign n34152 = n34139 & ~n34151 ;
  assign n34153 = ~n34150 & ~n34151 ;
  assign n34154 = ~n34152 & ~n34153 ;
  assign n34155 = ~n33414 & ~n33420 ;
  assign n34156 = n34154 & n34155 ;
  assign n34157 = ~n34154 & ~n34155 ;
  assign n34158 = ~n34156 & ~n34157 ;
  assign n34159 = x95 & n12506 ;
  assign n34160 = x93 & n13131 ;
  assign n34161 = x94 & n12501 ;
  assign n34162 = ~n34160 & ~n34161 ;
  assign n34163 = ~n34159 & n34162 ;
  assign n34164 = n6894 & n12509 ;
  assign n34165 = n34163 & ~n34164 ;
  assign n34166 = x44 & ~n34165 ;
  assign n34167 = x44 & ~n34166 ;
  assign n34168 = ~n34165 & ~n34166 ;
  assign n34169 = ~n34167 & ~n34168 ;
  assign n34170 = ~n34158 & n34169 ;
  assign n34171 = n34158 & ~n34169 ;
  assign n34172 = ~n34170 & ~n34171 ;
  assign n34173 = ~n33438 & n34172 ;
  assign n34174 = n33438 & ~n34172 ;
  assign n34175 = ~n34173 & ~n34174 ;
  assign n34176 = ~n34033 & n34175 ;
  assign n34177 = n34033 & ~n34175 ;
  assign n34178 = ~n34176 & ~n34177 ;
  assign n34179 = ~n34022 & n34178 ;
  assign n34180 = ~n34022 & ~n34179 ;
  assign n34181 = n34178 & ~n34179 ;
  assign n34182 = ~n34180 & ~n34181 ;
  assign n34183 = ~n34020 & ~n34182 ;
  assign n34184 = n34020 & ~n34181 ;
  assign n34185 = ~n34180 & n34184 ;
  assign n34186 = ~n34183 & ~n34185 ;
  assign n34187 = ~n34009 & n34186 ;
  assign n34188 = ~n34009 & ~n34187 ;
  assign n34189 = n34186 & ~n34187 ;
  assign n34190 = ~n34188 & ~n34189 ;
  assign n34191 = ~n34008 & ~n34190 ;
  assign n34192 = ~n34008 & ~n34191 ;
  assign n34193 = ~n34190 & ~n34191 ;
  assign n34194 = ~n34192 & ~n34193 ;
  assign n34195 = n33997 & ~n34194 ;
  assign n34196 = n33997 & ~n34195 ;
  assign n34197 = ~n34194 & ~n34195 ;
  assign n34198 = ~n34196 & ~n34197 ;
  assign n34199 = ~n33293 & ~n33496 ;
  assign n34200 = x110 & n5560 ;
  assign n34201 = x108 & n5943 ;
  assign n34202 = x109 & n5555 ;
  assign n34203 = ~n34201 & ~n34202 ;
  assign n34204 = ~n34200 & n34203 ;
  assign n34205 = ~n5563 & n34204 ;
  assign n34206 = ~n14497 & n34204 ;
  assign n34207 = ~n34205 & ~n34206 ;
  assign n34208 = x29 & ~n34207 ;
  assign n34209 = ~x29 & n34207 ;
  assign n34210 = ~n34208 & ~n34209 ;
  assign n34211 = ~n34199 & ~n34210 ;
  assign n34212 = ~n34199 & ~n34211 ;
  assign n34213 = ~n34210 & ~n34211 ;
  assign n34214 = ~n34212 & ~n34213 ;
  assign n34215 = ~n34198 & ~n34214 ;
  assign n34216 = ~n34198 & ~n34215 ;
  assign n34217 = ~n34214 & ~n34215 ;
  assign n34218 = ~n34216 & ~n34217 ;
  assign n34219 = ~n33982 & ~n34218 ;
  assign n34220 = ~n33982 & ~n34219 ;
  assign n34221 = ~n34218 & ~n34219 ;
  assign n34222 = ~n34220 & ~n34221 ;
  assign n34223 = n33965 & ~n34222 ;
  assign n34224 = ~n33965 & n34222 ;
  assign n34225 = n33950 & ~n34224 ;
  assign n34226 = ~n34223 & n34225 ;
  assign n34227 = n33950 & ~n34226 ;
  assign n34228 = ~n34224 & ~n34226 ;
  assign n34229 = ~n34223 & n34228 ;
  assign n34230 = ~n34227 & ~n34229 ;
  assign n34231 = ~n33246 & ~n33526 ;
  assign n34232 = x122 & n2093 ;
  assign n34233 = x120 & n2275 ;
  assign n34234 = x121 & n2088 ;
  assign n34235 = ~n34233 & ~n34234 ;
  assign n34236 = ~n34232 & n34235 ;
  assign n34237 = ~n2096 & n34236 ;
  assign n34238 = ~n22622 & n34236 ;
  assign n34239 = ~n34237 & ~n34238 ;
  assign n34240 = x17 & ~n34239 ;
  assign n34241 = ~x17 & n34239 ;
  assign n34242 = ~n34240 & ~n34241 ;
  assign n34243 = ~n34231 & ~n34242 ;
  assign n34244 = ~n34231 & ~n34243 ;
  assign n34245 = ~n34242 & ~n34243 ;
  assign n34246 = ~n34244 & ~n34245 ;
  assign n34247 = ~n34230 & ~n34246 ;
  assign n34248 = ~n34230 & ~n34247 ;
  assign n34249 = ~n34246 & ~n34247 ;
  assign n34250 = ~n34248 & ~n34249 ;
  assign n34251 = ~n33935 & ~n34250 ;
  assign n34252 = ~n33935 & ~n34251 ;
  assign n34253 = ~n34250 & ~n34251 ;
  assign n34254 = ~n34252 & ~n34253 ;
  assign n34255 = ~n33204 & ~n33215 ;
  assign n34256 = ~n33533 & ~n34255 ;
  assign n34257 = x126 & n1099 ;
  assign n34258 = x127 & n940 ;
  assign n34259 = ~n34257 & ~n34258 ;
  assign n34260 = ~n948 & n34259 ;
  assign n34261 = n26965 & n34259 ;
  assign n34262 = ~n34260 & ~n34261 ;
  assign n34263 = x11 & ~n34262 ;
  assign n34264 = ~x11 & n34262 ;
  assign n34265 = ~n34263 & ~n34264 ;
  assign n34266 = ~n34256 & ~n34265 ;
  assign n34267 = ~n34256 & ~n34266 ;
  assign n34268 = ~n34265 & ~n34266 ;
  assign n34269 = ~n34267 & ~n34268 ;
  assign n34270 = ~n34254 & ~n34269 ;
  assign n34271 = n34254 & ~n34268 ;
  assign n34272 = ~n34267 & n34271 ;
  assign n34273 = ~n34270 & ~n34272 ;
  assign n34274 = ~n33919 & n34273 ;
  assign n34275 = ~n33919 & ~n34274 ;
  assign n34276 = n34273 & ~n34274 ;
  assign n34277 = ~n34275 & ~n34276 ;
  assign n34278 = ~n33917 & ~n34277 ;
  assign n34279 = n33917 & ~n34276 ;
  assign n34280 = ~n34275 & n34279 ;
  assign n34281 = ~n34278 & ~n34280 ;
  assign n34648 = n34281 & x201 ;
  assign n34282 = ~n33905 & ~n33909 ;
  assign n34283 = ~n33566 & ~n33901 ;
  assign n34284 = ~n33563 & ~n34283 ;
  assign n34285 = ~x125 & n1434 ;
  assign n34286 = ~x123 & n1646 ;
  assign n34287 = ~x124 & n1429 ;
  assign n34288 = ~n34286 & ~n34287 ;
  assign n34289 = ~n34285 & n34288 ;
  assign n34290 = n1437 & n25330 ;
  assign n34291 = n34289 & ~n34290 ;
  assign n34292 = ~x14 & ~n34291 ;
  assign n34293 = ~x14 & ~n34292 ;
  assign n34294 = ~n34291 & ~n34292 ;
  assign n34295 = ~n34293 & ~n34294 ;
  assign n34296 = ~n33596 & ~n33894 ;
  assign n34297 = ~n34295 & ~n34296 ;
  assign n34298 = ~n34295 & ~n34297 ;
  assign n34299 = ~n34296 & ~n34297 ;
  assign n34300 = ~n34298 & ~n34299 ;
  assign n34301 = ~x119 & n2751 ;
  assign n34302 = ~x117 & n3020 ;
  assign n34303 = ~x118 & n2746 ;
  assign n34304 = ~n34302 & ~n34303 ;
  assign n34305 = ~n34301 & n34304 ;
  assign n34306 = n2754 & n20778 ;
  assign n34307 = n34305 & ~n34306 ;
  assign n34308 = ~x20 & ~n34307 ;
  assign n34309 = ~x20 & ~n34308 ;
  assign n34310 = ~n34307 & ~n34308 ;
  assign n34311 = ~n34309 & ~n34310 ;
  assign n34312 = ~n33883 & ~n33886 ;
  assign n34313 = n34311 & n34312 ;
  assign n34314 = ~n34311 & ~n34312 ;
  assign n34315 = ~n34313 & ~n34314 ;
  assign n34316 = ~x116 & n3589 ;
  assign n34317 = ~x114 & n3878 ;
  assign n34318 = ~x115 & n3584 ;
  assign n34319 = ~n34317 & ~n34318 ;
  assign n34320 = ~n34316 & n34319 ;
  assign n34321 = n3592 & n18678 ;
  assign n34322 = n34320 & ~n34321 ;
  assign n34323 = ~x23 & ~n34322 ;
  assign n34324 = ~x23 & ~n34323 ;
  assign n34325 = ~n34322 & ~n34323 ;
  assign n34326 = ~n34324 & ~n34325 ;
  assign n34327 = ~n33627 & ~n33867 ;
  assign n34328 = n34326 & n34327 ;
  assign n34329 = ~n34326 & ~n34327 ;
  assign n34330 = ~n34328 & ~n34329 ;
  assign n34331 = ~x113 & n4531 ;
  assign n34332 = ~x111 & n4847 ;
  assign n34333 = ~x112 & n4526 ;
  assign n34334 = ~n34332 & ~n34333 ;
  assign n34335 = ~n34331 & n34334 ;
  assign n34336 = n4534 & n16684 ;
  assign n34337 = n34335 & ~n34336 ;
  assign n34338 = ~x26 & ~n34337 ;
  assign n34339 = ~x26 & ~n34338 ;
  assign n34340 = ~n34337 & ~n34338 ;
  assign n34341 = ~n34339 & ~n34340 ;
  assign n34342 = ~n33644 & ~n33863 ;
  assign n34343 = ~n33641 & ~n34342 ;
  assign n34344 = ~n34341 & ~n34343 ;
  assign n34345 = ~n34341 & ~n34344 ;
  assign n34346 = ~n34343 & ~n34344 ;
  assign n34347 = ~n34345 & ~n34346 ;
  assign n34348 = ~x107 & n6725 ;
  assign n34349 = ~x105 & n7129 ;
  assign n34350 = ~x106 & n6720 ;
  assign n34351 = ~n34349 & ~n34350 ;
  assign n34352 = ~n34348 & n34351 ;
  assign n34353 = n6728 & n13034 ;
  assign n34354 = n34352 & ~n34353 ;
  assign n34355 = ~x32 & ~n34354 ;
  assign n34356 = ~x32 & ~n34355 ;
  assign n34357 = ~n34354 & ~n34355 ;
  assign n34358 = ~n34356 & ~n34357 ;
  assign n34359 = ~n33851 & ~n33856 ;
  assign n34360 = n34358 & n34359 ;
  assign n34361 = ~n34358 & ~n34359 ;
  assign n34362 = ~n34360 & ~n34361 ;
  assign n34363 = ~x104 & n8006 ;
  assign n34364 = ~x102 & n8474 ;
  assign n34365 = ~x103 & n8001 ;
  assign n34366 = ~n34364 & ~n34365 ;
  assign n34367 = ~n34363 & n34366 ;
  assign n34368 = n8009 & n11380 ;
  assign n34369 = n34367 & ~n34368 ;
  assign n34370 = ~x35 & ~n34369 ;
  assign n34371 = ~x35 & ~n34370 ;
  assign n34372 = ~n34369 & ~n34370 ;
  assign n34373 = ~n34371 & ~n34372 ;
  assign n34374 = ~n33834 & ~n33838 ;
  assign n34375 = ~x101 & n9433 ;
  assign n34376 = ~x99 & n9915 ;
  assign n34377 = ~x100 & n9428 ;
  assign n34378 = ~n34376 & ~n34377 ;
  assign n34379 = ~n34375 & n34378 ;
  assign n34380 = n9436 & n9844 ;
  assign n34381 = n34379 & ~n34380 ;
  assign n34382 = ~x38 & ~n34381 ;
  assign n34383 = ~x38 & ~n34382 ;
  assign n34384 = ~n34381 & ~n34382 ;
  assign n34385 = ~n34383 & ~n34384 ;
  assign n34386 = ~n33662 & ~n33819 ;
  assign n34387 = ~n33816 & ~n34386 ;
  assign n34388 = ~x98 & n10905 ;
  assign n34389 = ~x96 & n11466 ;
  assign n34390 = ~x97 & n10900 ;
  assign n34391 = ~n34389 & ~n34390 ;
  assign n34392 = ~n34388 & n34391 ;
  assign n34393 = n8426 & n10908 ;
  assign n34394 = n34392 & ~n34393 ;
  assign n34395 = ~x41 & ~n34394 ;
  assign n34396 = ~x41 & ~n34395 ;
  assign n34397 = ~n34394 & ~n34395 ;
  assign n34398 = ~n34396 & ~n34397 ;
  assign n34399 = ~x77 & n24612 ;
  assign n34400 = ~x75 & n25390 ;
  assign n34401 = ~x76 & n24607 ;
  assign n34402 = ~n34400 & ~n34401 ;
  assign n34403 = ~n34399 & n34402 ;
  assign n34404 = n1594 & n24615 ;
  assign n34405 = n34403 & ~n34404 ;
  assign n34406 = ~x62 & ~n34405 ;
  assign n34407 = ~x62 & ~n34406 ;
  assign n34408 = ~n34405 & ~n34406 ;
  assign n34409 = ~n34407 & ~n34408 ;
  assign n34410 = ~x73 & n27427 ;
  assign n34411 = ~x74 & ~n26217 ;
  assign n34412 = ~n34410 & ~n34411 ;
  assign n34413 = x8 & ~n32901 ;
  assign n34414 = ~n33695 & ~n34413 ;
  assign n34415 = n34412 & ~n34414 ;
  assign n34416 = n34412 & ~n34415 ;
  assign n34417 = ~n34414 & ~n34415 ;
  assign n34418 = ~n34416 & ~n34417 ;
  assign n34419 = ~n34409 & ~n34418 ;
  assign n34420 = ~n34409 & ~n34419 ;
  assign n34421 = ~n34418 & ~n34419 ;
  assign n34422 = ~n34420 & ~n34421 ;
  assign n34423 = ~n33688 & n33700 ;
  assign n34424 = ~n33698 & ~n34423 ;
  assign n34425 = ~n34422 & ~n34424 ;
  assign n34426 = ~n34422 & ~n34425 ;
  assign n34427 = ~n34424 & ~n34425 ;
  assign n34428 = ~n34426 & ~n34427 ;
  assign n34429 = ~x80 & n22325 ;
  assign n34430 = ~x78 & n23066 ;
  assign n34431 = ~x79 & n22320 ;
  assign n34432 = ~n34430 & ~n34431 ;
  assign n34433 = ~n34429 & n34432 ;
  assign n34434 = n2145 & n22328 ;
  assign n34435 = n34433 & ~n34434 ;
  assign n34436 = ~x59 & ~n34435 ;
  assign n34437 = ~x59 & ~n34436 ;
  assign n34438 = ~n34435 & ~n34436 ;
  assign n34439 = ~n34437 & ~n34438 ;
  assign n34440 = ~n34428 & ~n34439 ;
  assign n34441 = ~n34428 & ~n34440 ;
  assign n34442 = ~n34439 & ~n34440 ;
  assign n34443 = ~n34441 & ~n34442 ;
  assign n34444 = ~n33715 & ~n33718 ;
  assign n34445 = n34443 & n34444 ;
  assign n34446 = ~n34443 & ~n34444 ;
  assign n34447 = ~n34445 & ~n34446 ;
  assign n34448 = ~x83 & n20143 ;
  assign n34449 = ~x81 & n20854 ;
  assign n34450 = ~x82 & n20138 ;
  assign n34451 = ~n34449 & ~n34450 ;
  assign n34452 = ~n34448 & n34451 ;
  assign n34453 = n2972 & n20146 ;
  assign n34454 = n34452 & ~n34453 ;
  assign n34455 = ~x56 & ~n34454 ;
  assign n34456 = ~x56 & ~n34455 ;
  assign n34457 = ~n34454 & ~n34455 ;
  assign n34458 = ~n34456 & ~n34457 ;
  assign n34459 = n34447 & ~n34458 ;
  assign n34460 = n34447 & ~n34459 ;
  assign n34461 = ~n34458 & ~n34459 ;
  assign n34462 = ~n34460 & ~n34461 ;
  assign n34463 = ~n33732 & ~n33738 ;
  assign n34464 = n34462 & n34463 ;
  assign n34465 = ~n34462 & ~n34463 ;
  assign n34466 = ~n34464 & ~n34465 ;
  assign n34467 = ~x86 & n18025 ;
  assign n34468 = ~x84 & n18764 ;
  assign n34469 = ~x85 & n18020 ;
  assign n34470 = ~n34468 & ~n34469 ;
  assign n34471 = ~n34467 & n34470 ;
  assign n34472 = n3832 & n18028 ;
  assign n34473 = n34471 & ~n34472 ;
  assign n34474 = ~x53 & ~n34473 ;
  assign n34475 = ~x53 & ~n34474 ;
  assign n34476 = ~n34473 & ~n34474 ;
  assign n34477 = ~n34475 & ~n34476 ;
  assign n34478 = n34466 & ~n34477 ;
  assign n34479 = n34466 & ~n34478 ;
  assign n34480 = ~n34477 & ~n34478 ;
  assign n34481 = ~n34479 & ~n34480 ;
  assign n34482 = ~n33751 & ~n33756 ;
  assign n34483 = n34481 & n34482 ;
  assign n34484 = ~n34481 & ~n34482 ;
  assign n34485 = ~n34483 & ~n34484 ;
  assign n34486 = ~x89 & n16076 ;
  assign n34487 = ~x87 & n16756 ;
  assign n34488 = ~x88 & n16071 ;
  assign n34489 = ~n34487 & ~n34488 ;
  assign n34490 = ~n34486 & n34489 ;
  assign n34491 = n4664 & n16079 ;
  assign n34492 = n34490 & ~n34491 ;
  assign n34493 = ~x50 & ~n34492 ;
  assign n34494 = ~x50 & ~n34493 ;
  assign n34495 = ~n34492 & ~n34493 ;
  assign n34496 = ~n34494 & ~n34495 ;
  assign n34497 = n34485 & ~n34496 ;
  assign n34498 = n34485 & ~n34497 ;
  assign n34499 = ~n34496 & ~n34497 ;
  assign n34500 = ~n34498 & ~n34499 ;
  assign n34501 = ~n33759 & ~n33763 ;
  assign n34502 = n34500 & n34501 ;
  assign n34503 = ~n34500 & ~n34501 ;
  assign n34504 = ~n34502 & ~n34503 ;
  assign n34505 = ~x92 & n14233 ;
  assign n34506 = ~x90 & n14876 ;
  assign n34507 = ~x91 & n14228 ;
  assign n34508 = ~n34506 & ~n34507 ;
  assign n34509 = ~n34505 & n34508 ;
  assign n34510 = n5896 & n14236 ;
  assign n34511 = n34509 & ~n34510 ;
  assign n34512 = ~x47 & ~n34511 ;
  assign n34513 = ~x47 & ~n34512 ;
  assign n34514 = ~n34511 & ~n34512 ;
  assign n34515 = ~n34513 & ~n34514 ;
  assign n34516 = n34504 & ~n34515 ;
  assign n34517 = n34504 & ~n34516 ;
  assign n34518 = ~n34515 & ~n34516 ;
  assign n34519 = ~n34517 & ~n34518 ;
  assign n34520 = ~n33778 & ~n33784 ;
  assign n34521 = n34519 & n34520 ;
  assign n34522 = ~n34519 & ~n34520 ;
  assign n34523 = ~n34521 & ~n34522 ;
  assign n34524 = ~x95 & n12506 ;
  assign n34525 = ~x93 & n13131 ;
  assign n34526 = ~x94 & n12501 ;
  assign n34527 = ~n34525 & ~n34526 ;
  assign n34528 = ~n34524 & n34527 ;
  assign n34529 = n7100 & n12509 ;
  assign n34530 = n34528 & ~n34529 ;
  assign n34531 = ~x44 & ~n34530 ;
  assign n34532 = ~x44 & ~n34531 ;
  assign n34533 = ~n34530 & ~n34531 ;
  assign n34534 = ~n34532 & ~n34533 ;
  assign n34535 = ~n34523 & n34534 ;
  assign n34536 = n34523 & ~n34534 ;
  assign n34537 = ~n34535 & ~n34536 ;
  assign n34538 = ~n33802 & n34537 ;
  assign n34539 = n33802 & ~n34537 ;
  assign n34540 = ~n34538 & ~n34539 ;
  assign n34541 = ~n34398 & n34540 ;
  assign n34542 = n34398 & ~n34540 ;
  assign n34543 = ~n34541 & ~n34542 ;
  assign n34544 = ~n34387 & n34543 ;
  assign n34545 = ~n34387 & ~n34544 ;
  assign n34546 = n34543 & ~n34544 ;
  assign n34547 = ~n34545 & ~n34546 ;
  assign n34548 = ~n34385 & ~n34547 ;
  assign n34549 = n34385 & ~n34546 ;
  assign n34550 = ~n34545 & n34549 ;
  assign n34551 = ~n34548 & ~n34550 ;
  assign n34552 = ~n34374 & n34551 ;
  assign n34553 = ~n34374 & ~n34552 ;
  assign n34554 = n34551 & ~n34552 ;
  assign n34555 = ~n34553 & ~n34554 ;
  assign n34556 = ~n34373 & ~n34555 ;
  assign n34557 = ~n34373 & ~n34556 ;
  assign n34558 = ~n34555 & ~n34556 ;
  assign n34559 = ~n34557 & ~n34558 ;
  assign n34560 = n34362 & ~n34559 ;
  assign n34561 = n34362 & ~n34560 ;
  assign n34562 = ~n34559 & ~n34560 ;
  assign n34563 = ~n34561 & ~n34562 ;
  assign n34564 = ~n33657 & ~n33860 ;
  assign n34565 = ~x110 & n5560 ;
  assign n34566 = ~x108 & n5943 ;
  assign n34567 = ~x109 & n5555 ;
  assign n34568 = ~n34566 & ~n34567 ;
  assign n34569 = ~n34565 & n34568 ;
  assign n34570 = ~n5563 & n34569 ;
  assign n34571 = ~n14802 & n34569 ;
  assign n34572 = ~n34570 & ~n34571 ;
  assign n34573 = ~x29 & ~n34572 ;
  assign n34574 = x29 & n34572 ;
  assign n34575 = ~n34573 & ~n34574 ;
  assign n34576 = ~n34564 & ~n34575 ;
  assign n34577 = ~n34564 & ~n34576 ;
  assign n34578 = ~n34575 & ~n34576 ;
  assign n34579 = ~n34577 & ~n34578 ;
  assign n34580 = ~n34563 & ~n34579 ;
  assign n34581 = ~n34563 & ~n34580 ;
  assign n34582 = ~n34579 & ~n34580 ;
  assign n34583 = ~n34581 & ~n34582 ;
  assign n34584 = ~n34347 & ~n34583 ;
  assign n34585 = ~n34347 & ~n34584 ;
  assign n34586 = ~n34583 & ~n34584 ;
  assign n34587 = ~n34585 & ~n34586 ;
  assign n34588 = n34330 & ~n34587 ;
  assign n34589 = ~n34330 & n34587 ;
  assign n34590 = n34315 & ~n34589 ;
  assign n34591 = ~n34588 & n34590 ;
  assign n34592 = n34315 & ~n34591 ;
  assign n34593 = ~n34589 & ~n34591 ;
  assign n34594 = ~n34588 & n34593 ;
  assign n34595 = ~n34592 & ~n34594 ;
  assign n34596 = ~n33610 & ~n33890 ;
  assign n34597 = ~x122 & n2093 ;
  assign n34598 = ~x120 & n2275 ;
  assign n34599 = ~x121 & n2088 ;
  assign n34600 = ~n34598 & ~n34599 ;
  assign n34601 = ~n34597 & n34600 ;
  assign n34602 = ~n2096 & n34601 ;
  assign n34603 = ~n22998 & n34601 ;
  assign n34604 = ~n34602 & ~n34603 ;
  assign n34605 = ~x17 & ~n34604 ;
  assign n34606 = x17 & n34604 ;
  assign n34607 = ~n34605 & ~n34606 ;
  assign n34608 = ~n34596 & ~n34607 ;
  assign n34609 = ~n34596 & ~n34608 ;
  assign n34610 = ~n34607 & ~n34608 ;
  assign n34611 = ~n34609 & ~n34610 ;
  assign n34612 = ~n34595 & ~n34611 ;
  assign n34613 = ~n34595 & ~n34612 ;
  assign n34614 = ~n34611 & ~n34612 ;
  assign n34615 = ~n34613 & ~n34614 ;
  assign n34616 = ~n34300 & ~n34615 ;
  assign n34617 = ~n34300 & ~n34616 ;
  assign n34618 = ~n34615 & ~n34616 ;
  assign n34619 = ~n34617 & ~n34618 ;
  assign n34620 = ~n33568 & ~n33579 ;
  assign n34621 = ~n33897 & ~n34620 ;
  assign n34622 = ~x126 & n1099 ;
  assign n34623 = ~x127 & n940 ;
  assign n34624 = ~n34622 & ~n34623 ;
  assign n34625 = ~n948 & n34624 ;
  assign n34626 = n27368 & n34624 ;
  assign n34627 = ~n34625 & ~n34626 ;
  assign n34628 = ~x11 & ~n34627 ;
  assign n34629 = x11 & n34627 ;
  assign n34630 = ~n34628 & ~n34629 ;
  assign n34631 = ~n34621 & ~n34630 ;
  assign n34632 = ~n34621 & ~n34631 ;
  assign n34633 = ~n34630 & ~n34631 ;
  assign n34634 = ~n34632 & ~n34633 ;
  assign n34635 = ~n34619 & ~n34634 ;
  assign n34636 = n34619 & ~n34633 ;
  assign n34637 = ~n34632 & n34636 ;
  assign n34638 = ~n34635 & ~n34637 ;
  assign n34639 = ~n34284 & n34638 ;
  assign n34640 = ~n34284 & ~n34639 ;
  assign n34641 = n34638 & ~n34639 ;
  assign n34642 = ~n34640 & ~n34641 ;
  assign n34643 = ~n34282 & ~n34642 ;
  assign n34644 = n34282 & ~n34641 ;
  assign n34645 = ~n34640 & n34644 ;
  assign n34646 = ~n34643 & ~n34645 ;
  assign n34649 = ~n34646 & ~x201 ;
  assign n34650 = ~n34648 & ~n34649 ;
  assign n34651 = ~n34274 & ~n34278 ;
  assign n34652 = ~n34266 & ~n34270 ;
  assign n34653 = ~n33932 & ~n34251 ;
  assign n34654 = x127 & n1099 ;
  assign n34655 = n948 & n26962 ;
  assign n34656 = ~n34654 & ~n34655 ;
  assign n34657 = x11 & ~n34656 ;
  assign n34658 = x11 & ~n34657 ;
  assign n34659 = ~n34656 & ~n34657 ;
  assign n34660 = ~n34658 & ~n34659 ;
  assign n34661 = ~n34653 & ~n34660 ;
  assign n34662 = ~n34653 & ~n34661 ;
  assign n34663 = ~n34660 & ~n34661 ;
  assign n34664 = ~n34662 & ~n34663 ;
  assign n34665 = ~n34243 & ~n34247 ;
  assign n34666 = x126 & n1434 ;
  assign n34667 = x124 & n1646 ;
  assign n34668 = x125 & n1429 ;
  assign n34669 = ~n34667 & ~n34668 ;
  assign n34670 = ~n34666 & n34669 ;
  assign n34671 = ~n1437 & n34670 ;
  assign n34672 = ~n25735 & n34670 ;
  assign n34673 = ~n34671 & ~n34672 ;
  assign n34674 = x14 & ~n34673 ;
  assign n34675 = ~x14 & n34673 ;
  assign n34676 = ~n34674 & ~n34675 ;
  assign n34677 = ~n34665 & ~n34676 ;
  assign n34678 = n34665 & n34676 ;
  assign n34679 = ~n34677 & ~n34678 ;
  assign n34680 = x123 & n2093 ;
  assign n34681 = x121 & n2275 ;
  assign n34682 = x122 & n2088 ;
  assign n34683 = ~n34681 & ~n34682 ;
  assign n34684 = ~n34680 & n34683 ;
  assign n34685 = n2096 & n23382 ;
  assign n34686 = n34684 & ~n34685 ;
  assign n34687 = x17 & ~n34686 ;
  assign n34688 = x17 & ~n34687 ;
  assign n34689 = ~n34686 & ~n34687 ;
  assign n34690 = ~n34688 & ~n34689 ;
  assign n34691 = ~n33949 & ~n34226 ;
  assign n34692 = n34690 & n34691 ;
  assign n34693 = ~n34690 & ~n34691 ;
  assign n34694 = ~n34692 & ~n34693 ;
  assign n34695 = x120 & n2751 ;
  assign n34696 = x118 & n3020 ;
  assign n34697 = x119 & n2746 ;
  assign n34698 = ~n34696 & ~n34697 ;
  assign n34699 = ~n34695 & n34698 ;
  assign n34700 = n2754 & n21143 ;
  assign n34701 = n34699 & ~n34700 ;
  assign n34702 = x20 & ~n34701 ;
  assign n34703 = x20 & ~n34702 ;
  assign n34704 = ~n34701 & ~n34702 ;
  assign n34705 = ~n34703 & ~n34704 ;
  assign n34706 = ~n33964 & ~n34223 ;
  assign n34707 = ~n34705 & ~n34706 ;
  assign n34708 = ~n34705 & ~n34707 ;
  assign n34709 = ~n34706 & ~n34707 ;
  assign n34710 = ~n34708 & ~n34709 ;
  assign n34711 = ~n34211 & ~n34215 ;
  assign n34712 = x114 & n4531 ;
  assign n34713 = x112 & n4847 ;
  assign n34714 = x113 & n4526 ;
  assign n34715 = ~n34713 & ~n34714 ;
  assign n34716 = ~n34712 & n34715 ;
  assign n34717 = ~n4534 & n34716 ;
  assign n34718 = ~n17012 & n34716 ;
  assign n34719 = ~n34717 & ~n34718 ;
  assign n34720 = x26 & ~n34719 ;
  assign n34721 = ~x26 & n34719 ;
  assign n34722 = ~n34720 & ~n34721 ;
  assign n34723 = ~n34711 & ~n34722 ;
  assign n34724 = n34711 & n34722 ;
  assign n34725 = ~n34723 & ~n34724 ;
  assign n34726 = x111 & n5560 ;
  assign n34727 = x109 & n5943 ;
  assign n34728 = x110 & n5555 ;
  assign n34729 = ~n34727 & ~n34728 ;
  assign n34730 = ~n34726 & n34729 ;
  assign n34731 = n5563 & n15111 ;
  assign n34732 = n34730 & ~n34731 ;
  assign n34733 = x29 & ~n34732 ;
  assign n34734 = x29 & ~n34733 ;
  assign n34735 = ~n34732 & ~n34733 ;
  assign n34736 = ~n34734 & ~n34735 ;
  assign n34737 = ~n33996 & ~n34195 ;
  assign n34738 = n34736 & n34737 ;
  assign n34739 = ~n34736 & ~n34737 ;
  assign n34740 = ~n34738 & ~n34739 ;
  assign n34741 = ~n34187 & ~n34191 ;
  assign n34742 = x108 & n6725 ;
  assign n34743 = x106 & n7129 ;
  assign n34744 = x107 & n6720 ;
  assign n34745 = ~n34743 & ~n34744 ;
  assign n34746 = ~n34742 & n34745 ;
  assign n34747 = ~n6728 & n34746 ;
  assign n34748 = ~n13323 & n34746 ;
  assign n34749 = ~n34747 & ~n34748 ;
  assign n34750 = x32 & ~n34749 ;
  assign n34751 = ~x32 & n34749 ;
  assign n34752 = ~n34750 & ~n34751 ;
  assign n34753 = ~n34741 & ~n34752 ;
  assign n34754 = n34741 & n34752 ;
  assign n34755 = ~n34753 & ~n34754 ;
  assign n34756 = x105 & n8006 ;
  assign n34757 = x103 & n8474 ;
  assign n34758 = x104 & n8001 ;
  assign n34759 = ~n34757 & ~n34758 ;
  assign n34760 = ~n34756 & n34759 ;
  assign n34761 = n8009 & n11648 ;
  assign n34762 = n34760 & ~n34761 ;
  assign n34763 = x35 & ~n34762 ;
  assign n34764 = x35 & ~n34763 ;
  assign n34765 = ~n34762 & ~n34763 ;
  assign n34766 = ~n34764 & ~n34765 ;
  assign n34767 = ~n34179 & ~n34183 ;
  assign n34768 = ~n34119 & ~n34132 ;
  assign n34769 = x90 & n16076 ;
  assign n34770 = x88 & n16756 ;
  assign n34771 = x89 & n16071 ;
  assign n34772 = ~n34770 & ~n34771 ;
  assign n34773 = ~n34769 & n34772 ;
  assign n34774 = n4986 & n16079 ;
  assign n34775 = n34773 & ~n34774 ;
  assign n34776 = x50 & ~n34775 ;
  assign n34777 = x50 & ~n34776 ;
  assign n34778 = ~n34775 & ~n34776 ;
  assign n34779 = ~n34777 & ~n34778 ;
  assign n34780 = ~n34100 & ~n34113 ;
  assign n34781 = x87 & n18025 ;
  assign n34782 = x85 & n18764 ;
  assign n34783 = x86 & n18020 ;
  assign n34784 = ~n34782 & ~n34783 ;
  assign n34785 = ~n34781 & n34784 ;
  assign n34786 = n3991 & n18028 ;
  assign n34787 = n34785 & ~n34786 ;
  assign n34788 = x53 & ~n34787 ;
  assign n34789 = x53 & ~n34788 ;
  assign n34790 = ~n34787 & ~n34788 ;
  assign n34791 = ~n34789 & ~n34790 ;
  assign n34792 = ~n34081 & ~n34094 ;
  assign n34793 = ~n34050 & ~n34054 ;
  assign n34794 = x74 & n27024 ;
  assign n34795 = x75 & ~n26217 ;
  assign n34796 = ~n34794 & ~n34795 ;
  assign n34797 = n34047 & ~n34796 ;
  assign n34798 = n34047 & ~n34797 ;
  assign n34799 = ~n34796 & ~n34797 ;
  assign n34800 = ~n34798 & ~n34799 ;
  assign n34801 = ~n34793 & ~n34800 ;
  assign n34802 = ~n34793 & ~n34801 ;
  assign n34803 = ~n34800 & ~n34801 ;
  assign n34804 = ~n34802 & ~n34803 ;
  assign n34805 = x78 & n24612 ;
  assign n34806 = x76 & n25390 ;
  assign n34807 = x77 & n24607 ;
  assign n34808 = ~n34806 & ~n34807 ;
  assign n34809 = ~n34805 & n34808 ;
  assign n34810 = n1624 & n24615 ;
  assign n34811 = n34809 & ~n34810 ;
  assign n34812 = x62 & ~n34811 ;
  assign n34813 = x62 & ~n34812 ;
  assign n34814 = ~n34811 & ~n34812 ;
  assign n34815 = ~n34813 & ~n34814 ;
  assign n34816 = ~n34804 & ~n34815 ;
  assign n34817 = ~n34804 & ~n34816 ;
  assign n34818 = ~n34815 & ~n34816 ;
  assign n34819 = ~n34817 & ~n34818 ;
  assign n34820 = x81 & n22325 ;
  assign n34821 = x79 & n23066 ;
  assign n34822 = x80 & n22320 ;
  assign n34823 = ~n34821 & ~n34822 ;
  assign n34824 = ~n34820 & n34823 ;
  assign n34825 = n2348 & n22328 ;
  assign n34826 = n34824 & ~n34825 ;
  assign n34827 = x59 & ~n34826 ;
  assign n34828 = x59 & ~n34827 ;
  assign n34829 = ~n34826 & ~n34827 ;
  assign n34830 = ~n34828 & ~n34829 ;
  assign n34831 = ~n34819 & ~n34830 ;
  assign n34832 = ~n34819 & ~n34831 ;
  assign n34833 = ~n34830 & ~n34831 ;
  assign n34834 = ~n34832 & ~n34833 ;
  assign n34835 = ~n34060 & ~n34075 ;
  assign n34836 = n34834 & n34835 ;
  assign n34837 = ~n34834 & ~n34835 ;
  assign n34838 = ~n34836 & ~n34837 ;
  assign n34839 = x84 & n20143 ;
  assign n34840 = x82 & n20854 ;
  assign n34841 = x83 & n20138 ;
  assign n34842 = ~n34840 & ~n34841 ;
  assign n34843 = ~n34839 & n34842 ;
  assign n34844 = n3114 & n20146 ;
  assign n34845 = n34843 & ~n34844 ;
  assign n34846 = x56 & ~n34845 ;
  assign n34847 = x56 & ~n34846 ;
  assign n34848 = ~n34845 & ~n34846 ;
  assign n34849 = ~n34847 & ~n34848 ;
  assign n34850 = ~n34838 & n34849 ;
  assign n34851 = n34838 & ~n34849 ;
  assign n34852 = ~n34850 & ~n34851 ;
  assign n34853 = ~n34792 & n34852 ;
  assign n34854 = ~n34792 & ~n34853 ;
  assign n34855 = n34852 & ~n34853 ;
  assign n34856 = ~n34854 & ~n34855 ;
  assign n34857 = ~n34791 & ~n34856 ;
  assign n34858 = n34791 & ~n34855 ;
  assign n34859 = ~n34854 & n34858 ;
  assign n34860 = ~n34857 & ~n34859 ;
  assign n34861 = ~n34780 & n34860 ;
  assign n34862 = n34780 & ~n34860 ;
  assign n34863 = ~n34861 & ~n34862 ;
  assign n34864 = ~n34779 & n34863 ;
  assign n34865 = n34779 & ~n34863 ;
  assign n34866 = ~n34864 & ~n34865 ;
  assign n34867 = ~n34768 & n34866 ;
  assign n34868 = n34768 & ~n34866 ;
  assign n34869 = ~n34867 & ~n34868 ;
  assign n34870 = x93 & n14233 ;
  assign n34871 = x91 & n14876 ;
  assign n34872 = x92 & n14228 ;
  assign n34873 = ~n34871 & ~n34872 ;
  assign n34874 = ~n34870 & n34873 ;
  assign n34875 = n6094 & n14236 ;
  assign n34876 = n34874 & ~n34875 ;
  assign n34877 = x47 & ~n34876 ;
  assign n34878 = x47 & ~n34877 ;
  assign n34879 = ~n34876 & ~n34877 ;
  assign n34880 = ~n34878 & ~n34879 ;
  assign n34881 = n34869 & ~n34880 ;
  assign n34882 = n34869 & ~n34881 ;
  assign n34883 = ~n34880 & ~n34881 ;
  assign n34884 = ~n34882 & ~n34883 ;
  assign n34885 = ~n34138 & ~n34151 ;
  assign n34886 = n34884 & n34885 ;
  assign n34887 = ~n34884 & ~n34885 ;
  assign n34888 = ~n34886 & ~n34887 ;
  assign n34889 = x96 & n12506 ;
  assign n34890 = x94 & n13131 ;
  assign n34891 = x95 & n12501 ;
  assign n34892 = ~n34890 & ~n34891 ;
  assign n34893 = ~n34889 & n34892 ;
  assign n34894 = n7321 & n12509 ;
  assign n34895 = n34893 & ~n34894 ;
  assign n34896 = x44 & ~n34895 ;
  assign n34897 = x44 & ~n34896 ;
  assign n34898 = ~n34895 & ~n34896 ;
  assign n34899 = ~n34897 & ~n34898 ;
  assign n34900 = ~n34888 & n34899 ;
  assign n34901 = n34888 & ~n34899 ;
  assign n34902 = ~n34900 & ~n34901 ;
  assign n34903 = ~n34157 & ~n34171 ;
  assign n34904 = n34902 & ~n34903 ;
  assign n34905 = ~n34902 & n34903 ;
  assign n34906 = ~n34904 & ~n34905 ;
  assign n34907 = x99 & n10905 ;
  assign n34908 = x97 & n11466 ;
  assign n34909 = x98 & n10900 ;
  assign n34910 = ~n34908 & ~n34909 ;
  assign n34911 = ~n34907 & n34910 ;
  assign n34912 = n8660 & n10908 ;
  assign n34913 = n34911 & ~n34912 ;
  assign n34914 = x41 & ~n34913 ;
  assign n34915 = x41 & ~n34914 ;
  assign n34916 = ~n34913 & ~n34914 ;
  assign n34917 = ~n34915 & ~n34916 ;
  assign n34918 = n34906 & ~n34917 ;
  assign n34919 = n34906 & ~n34918 ;
  assign n34920 = ~n34917 & ~n34918 ;
  assign n34921 = ~n34919 & ~n34920 ;
  assign n34922 = ~n34173 & ~n34176 ;
  assign n34923 = n34921 & n34922 ;
  assign n34924 = ~n34921 & ~n34922 ;
  assign n34925 = ~n34923 & ~n34924 ;
  assign n34926 = x102 & n9433 ;
  assign n34927 = x100 & n9915 ;
  assign n34928 = x101 & n9428 ;
  assign n34929 = ~n34927 & ~n34928 ;
  assign n34930 = ~n34926 & n34929 ;
  assign n34931 = n9436 & n10092 ;
  assign n34932 = n34930 & ~n34931 ;
  assign n34933 = x38 & ~n34932 ;
  assign n34934 = x38 & ~n34933 ;
  assign n34935 = ~n34932 & ~n34933 ;
  assign n34936 = ~n34934 & ~n34935 ;
  assign n34937 = ~n34925 & n34936 ;
  assign n34938 = n34925 & ~n34936 ;
  assign n34939 = ~n34937 & ~n34938 ;
  assign n34940 = ~n34767 & n34939 ;
  assign n34941 = n34767 & ~n34939 ;
  assign n34942 = ~n34940 & ~n34941 ;
  assign n34943 = ~n34766 & n34942 ;
  assign n34944 = ~n34766 & ~n34943 ;
  assign n34945 = n34942 & ~n34943 ;
  assign n34946 = ~n34944 & ~n34945 ;
  assign n34947 = n34755 & ~n34946 ;
  assign n34948 = n34755 & ~n34947 ;
  assign n34949 = ~n34946 & ~n34947 ;
  assign n34950 = ~n34948 & ~n34949 ;
  assign n34951 = n34740 & ~n34950 ;
  assign n34952 = ~n34740 & n34950 ;
  assign n34953 = n34725 & ~n34952 ;
  assign n34954 = ~n34951 & n34953 ;
  assign n34955 = n34725 & ~n34954 ;
  assign n34956 = ~n34952 & ~n34954 ;
  assign n34957 = ~n34951 & n34956 ;
  assign n34958 = ~n34955 & ~n34957 ;
  assign n34959 = ~n33979 & ~n34219 ;
  assign n34960 = x117 & n3589 ;
  assign n34961 = x115 & n3878 ;
  assign n34962 = x116 & n3584 ;
  assign n34963 = ~n34961 & ~n34962 ;
  assign n34964 = ~n34960 & n34963 ;
  assign n34965 = ~n3592 & n34964 ;
  assign n34966 = ~n19026 & n34964 ;
  assign n34967 = ~n34965 & ~n34966 ;
  assign n34968 = x23 & ~n34967 ;
  assign n34969 = ~x23 & n34967 ;
  assign n34970 = ~n34968 & ~n34969 ;
  assign n34971 = ~n34959 & ~n34970 ;
  assign n34972 = ~n34959 & ~n34971 ;
  assign n34973 = ~n34970 & ~n34971 ;
  assign n34974 = ~n34972 & ~n34973 ;
  assign n34975 = ~n34958 & ~n34974 ;
  assign n34976 = ~n34958 & ~n34975 ;
  assign n34977 = ~n34974 & ~n34975 ;
  assign n34978 = ~n34976 & ~n34977 ;
  assign n34979 = ~n34710 & ~n34978 ;
  assign n34980 = ~n34710 & ~n34979 ;
  assign n34981 = ~n34978 & ~n34979 ;
  assign n34982 = ~n34980 & ~n34981 ;
  assign n34983 = n34694 & ~n34982 ;
  assign n34984 = ~n34694 & n34982 ;
  assign n34985 = n34679 & ~n34984 ;
  assign n34986 = ~n34983 & n34985 ;
  assign n34987 = n34679 & ~n34986 ;
  assign n34988 = ~n34984 & ~n34986 ;
  assign n34989 = ~n34983 & n34988 ;
  assign n34990 = ~n34987 & ~n34989 ;
  assign n34991 = ~n34664 & n34990 ;
  assign n34992 = n34664 & ~n34990 ;
  assign n34993 = ~n34991 & ~n34992 ;
  assign n34994 = ~n34652 & ~n34993 ;
  assign n34995 = ~n34652 & ~n34994 ;
  assign n34996 = ~n34993 & ~n34994 ;
  assign n34997 = ~n34995 & ~n34996 ;
  assign n34998 = ~n34651 & ~n34997 ;
  assign n34999 = n34651 & ~n34996 ;
  assign n35000 = ~n34995 & n34999 ;
  assign n35001 = ~n34998 & ~n35000 ;
  assign n35354 = n35001 & x202 ;
  assign n35002 = ~n34639 & ~n34643 ;
  assign n35003 = ~n34631 & ~n34635 ;
  assign n35004 = ~n34297 & ~n34616 ;
  assign n35005 = ~x127 & n1099 ;
  assign n35006 = n948 & n27365 ;
  assign n35007 = ~n35005 & ~n35006 ;
  assign n35008 = ~x11 & ~n35007 ;
  assign n35009 = ~x11 & ~n35008 ;
  assign n35010 = ~n35007 & ~n35008 ;
  assign n35011 = ~n35009 & ~n35010 ;
  assign n35012 = ~n35004 & ~n35011 ;
  assign n35013 = ~n35004 & ~n35012 ;
  assign n35014 = ~n35011 & ~n35012 ;
  assign n35015 = ~n35013 & ~n35014 ;
  assign n35016 = ~n34608 & ~n34612 ;
  assign n35017 = ~x126 & n1434 ;
  assign n35018 = ~x124 & n1646 ;
  assign n35019 = ~x125 & n1429 ;
  assign n35020 = ~n35018 & ~n35019 ;
  assign n35021 = ~n35017 & n35020 ;
  assign n35022 = ~n1437 & n35021 ;
  assign n35023 = ~n26128 & n35021 ;
  assign n35024 = ~n35022 & ~n35023 ;
  assign n35025 = ~x14 & ~n35024 ;
  assign n35026 = x14 & n35024 ;
  assign n35027 = ~n35025 & ~n35026 ;
  assign n35028 = ~n35016 & ~n35027 ;
  assign n35029 = n35016 & n35027 ;
  assign n35030 = ~n35028 & ~n35029 ;
  assign n35031 = ~x123 & n2093 ;
  assign n35032 = ~x121 & n2275 ;
  assign n35033 = ~x122 & n2088 ;
  assign n35034 = ~n35032 & ~n35033 ;
  assign n35035 = ~n35031 & n35034 ;
  assign n35036 = n2096 & n23760 ;
  assign n35037 = n35035 & ~n35036 ;
  assign n35038 = ~x17 & ~n35037 ;
  assign n35039 = ~x17 & ~n35038 ;
  assign n35040 = ~n35037 & ~n35038 ;
  assign n35041 = ~n35039 & ~n35040 ;
  assign n35042 = ~n34314 & ~n34591 ;
  assign n35043 = n35041 & n35042 ;
  assign n35044 = ~n35041 & ~n35042 ;
  assign n35045 = ~n35043 & ~n35044 ;
  assign n35046 = ~x120 & n2751 ;
  assign n35047 = ~x118 & n3020 ;
  assign n35048 = ~x119 & n2746 ;
  assign n35049 = ~n35047 & ~n35048 ;
  assign n35050 = ~n35046 & n35049 ;
  assign n35051 = n2754 & n21501 ;
  assign n35052 = n35050 & ~n35051 ;
  assign n35053 = ~x20 & ~n35052 ;
  assign n35054 = ~x20 & ~n35053 ;
  assign n35055 = ~n35052 & ~n35053 ;
  assign n35056 = ~n35054 & ~n35055 ;
  assign n35057 = ~n34329 & ~n34588 ;
  assign n35058 = ~n35056 & ~n35057 ;
  assign n35059 = ~n35056 & ~n35058 ;
  assign n35060 = ~n35057 & ~n35058 ;
  assign n35061 = ~n35059 & ~n35060 ;
  assign n35062 = ~n34576 & ~n34580 ;
  assign n35063 = ~x114 & n4531 ;
  assign n35064 = ~x112 & n4847 ;
  assign n35065 = ~x113 & n4526 ;
  assign n35066 = ~n35064 & ~n35065 ;
  assign n35067 = ~n35063 & n35066 ;
  assign n35068 = ~n4534 & n35067 ;
  assign n35069 = ~n17333 & n35067 ;
  assign n35070 = ~n35068 & ~n35069 ;
  assign n35071 = ~x26 & ~n35070 ;
  assign n35072 = x26 & n35070 ;
  assign n35073 = ~n35071 & ~n35072 ;
  assign n35074 = ~n35062 & ~n35073 ;
  assign n35075 = n35062 & n35073 ;
  assign n35076 = ~n35074 & ~n35075 ;
  assign n35077 = ~x111 & n5560 ;
  assign n35078 = ~x109 & n5943 ;
  assign n35079 = ~x110 & n5555 ;
  assign n35080 = ~n35078 & ~n35079 ;
  assign n35081 = ~n35077 & n35080 ;
  assign n35082 = n5563 & n15411 ;
  assign n35083 = n35081 & ~n35082 ;
  assign n35084 = ~x29 & ~n35083 ;
  assign n35085 = ~x29 & ~n35084 ;
  assign n35086 = ~n35083 & ~n35084 ;
  assign n35087 = ~n35085 & ~n35086 ;
  assign n35088 = ~n34361 & ~n34560 ;
  assign n35089 = n35087 & n35088 ;
  assign n35090 = ~n35087 & ~n35088 ;
  assign n35091 = ~n35089 & ~n35090 ;
  assign n35092 = ~n34552 & ~n34556 ;
  assign n35093 = ~x108 & n6725 ;
  assign n35094 = ~x106 & n7129 ;
  assign n35095 = ~x107 & n6720 ;
  assign n35096 = ~n35094 & ~n35095 ;
  assign n35097 = ~n35093 & n35096 ;
  assign n35098 = ~n6728 & n35097 ;
  assign n35099 = ~n13601 & n35097 ;
  assign n35100 = ~n35098 & ~n35099 ;
  assign n35101 = ~x32 & ~n35100 ;
  assign n35102 = x32 & n35100 ;
  assign n35103 = ~n35101 & ~n35102 ;
  assign n35104 = ~n35092 & ~n35103 ;
  assign n35105 = n35092 & n35103 ;
  assign n35106 = ~n35104 & ~n35105 ;
  assign n35107 = ~x105 & n8006 ;
  assign n35108 = ~x103 & n8474 ;
  assign n35109 = ~x104 & n8001 ;
  assign n35110 = ~n35108 & ~n35109 ;
  assign n35111 = ~n35107 & n35110 ;
  assign n35112 = n8009 & n11907 ;
  assign n35113 = n35111 & ~n35112 ;
  assign n35114 = ~x35 & ~n35113 ;
  assign n35115 = ~x35 & ~n35114 ;
  assign n35116 = ~n35113 & ~n35114 ;
  assign n35117 = ~n35115 & ~n35116 ;
  assign n35118 = ~n34544 & ~n34548 ;
  assign n35119 = ~n34484 & ~n34497 ;
  assign n35120 = ~x90 & n16076 ;
  assign n35121 = ~x88 & n16756 ;
  assign n35122 = ~x89 & n16071 ;
  assign n35123 = ~n35121 & ~n35122 ;
  assign n35124 = ~n35120 & n35123 ;
  assign n35125 = n5155 & n16079 ;
  assign n35126 = n35124 & ~n35125 ;
  assign n35127 = ~x50 & ~n35126 ;
  assign n35128 = ~x50 & ~n35127 ;
  assign n35129 = ~n35126 & ~n35127 ;
  assign n35130 = ~n35128 & ~n35129 ;
  assign n35131 = ~n34465 & ~n34478 ;
  assign n35132 = ~x87 & n18025 ;
  assign n35133 = ~x85 & n18764 ;
  assign n35134 = ~x86 & n18020 ;
  assign n35135 = ~n35133 & ~n35134 ;
  assign n35136 = ~n35132 & n35135 ;
  assign n35137 = n4143 & n18028 ;
  assign n35138 = n35136 & ~n35137 ;
  assign n35139 = ~x53 & ~n35138 ;
  assign n35140 = ~x53 & ~n35139 ;
  assign n35141 = ~n35138 & ~n35139 ;
  assign n35142 = ~n35140 & ~n35141 ;
  assign n35143 = ~n34446 & ~n34459 ;
  assign n35144 = ~n34415 & ~n34419 ;
  assign n35145 = ~x74 & n27427 ;
  assign n35146 = ~x75 & ~n26217 ;
  assign n35147 = ~n35145 & ~n35146 ;
  assign n35148 = n34412 & ~n35147 ;
  assign n35149 = n34412 & ~n35148 ;
  assign n35150 = ~n35147 & ~n35148 ;
  assign n35151 = ~n35149 & ~n35150 ;
  assign n35152 = ~n35144 & ~n35151 ;
  assign n35153 = ~n35144 & ~n35152 ;
  assign n35154 = ~n35151 & ~n35152 ;
  assign n35155 = ~n35153 & ~n35154 ;
  assign n35156 = ~x78 & n24612 ;
  assign n35157 = ~x76 & n25390 ;
  assign n35158 = ~x77 & n24607 ;
  assign n35159 = ~n35157 & ~n35158 ;
  assign n35160 = ~n35156 & n35159 ;
  assign n35161 = n1718 & n24615 ;
  assign n35162 = n35160 & ~n35161 ;
  assign n35163 = ~x62 & ~n35162 ;
  assign n35164 = ~x62 & ~n35163 ;
  assign n35165 = ~n35162 & ~n35163 ;
  assign n35166 = ~n35164 & ~n35165 ;
  assign n35167 = ~n35155 & ~n35166 ;
  assign n35168 = ~n35155 & ~n35167 ;
  assign n35169 = ~n35166 & ~n35167 ;
  assign n35170 = ~n35168 & ~n35169 ;
  assign n35171 = ~x81 & n22325 ;
  assign n35172 = ~x79 & n23066 ;
  assign n35173 = ~x80 & n22320 ;
  assign n35174 = ~n35172 & ~n35173 ;
  assign n35175 = ~n35171 & n35174 ;
  assign n35176 = n2460 & n22328 ;
  assign n35177 = n35175 & ~n35176 ;
  assign n35178 = ~x59 & ~n35177 ;
  assign n35179 = ~x59 & ~n35178 ;
  assign n35180 = ~n35177 & ~n35178 ;
  assign n35181 = ~n35179 & ~n35180 ;
  assign n35182 = ~n35170 & ~n35181 ;
  assign n35183 = ~n35170 & ~n35182 ;
  assign n35184 = ~n35181 & ~n35182 ;
  assign n35185 = ~n35183 & ~n35184 ;
  assign n35186 = ~n34425 & ~n34440 ;
  assign n35187 = n35185 & n35186 ;
  assign n35188 = ~n35185 & ~n35186 ;
  assign n35189 = ~n35187 & ~n35188 ;
  assign n35190 = ~x84 & n20143 ;
  assign n35191 = ~x82 & n20854 ;
  assign n35192 = ~x83 & n20138 ;
  assign n35193 = ~n35191 & ~n35192 ;
  assign n35194 = ~n35190 & n35193 ;
  assign n35195 = n3247 & n20146 ;
  assign n35196 = n35194 & ~n35195 ;
  assign n35197 = ~x56 & ~n35196 ;
  assign n35198 = ~x56 & ~n35197 ;
  assign n35199 = ~n35196 & ~n35197 ;
  assign n35200 = ~n35198 & ~n35199 ;
  assign n35201 = ~n35189 & n35200 ;
  assign n35202 = n35189 & ~n35200 ;
  assign n35203 = ~n35201 & ~n35202 ;
  assign n35204 = ~n35143 & n35203 ;
  assign n35205 = ~n35143 & ~n35204 ;
  assign n35206 = n35203 & ~n35204 ;
  assign n35207 = ~n35205 & ~n35206 ;
  assign n35208 = ~n35142 & ~n35207 ;
  assign n35209 = n35142 & ~n35206 ;
  assign n35210 = ~n35205 & n35209 ;
  assign n35211 = ~n35208 & ~n35210 ;
  assign n35212 = ~n35131 & n35211 ;
  assign n35213 = n35131 & ~n35211 ;
  assign n35214 = ~n35212 & ~n35213 ;
  assign n35215 = ~n35130 & n35214 ;
  assign n35216 = n35130 & ~n35214 ;
  assign n35217 = ~n35215 & ~n35216 ;
  assign n35218 = ~n35119 & n35217 ;
  assign n35219 = n35119 & ~n35217 ;
  assign n35220 = ~n35218 & ~n35219 ;
  assign n35221 = ~x93 & n14233 ;
  assign n35222 = ~x91 & n14876 ;
  assign n35223 = ~x92 & n14228 ;
  assign n35224 = ~n35222 & ~n35223 ;
  assign n35225 = ~n35221 & n35224 ;
  assign n35226 = n6285 & n14236 ;
  assign n35227 = n35225 & ~n35226 ;
  assign n35228 = ~x47 & ~n35227 ;
  assign n35229 = ~x47 & ~n35228 ;
  assign n35230 = ~n35227 & ~n35228 ;
  assign n35231 = ~n35229 & ~n35230 ;
  assign n35232 = n35220 & ~n35231 ;
  assign n35233 = n35220 & ~n35232 ;
  assign n35234 = ~n35231 & ~n35232 ;
  assign n35235 = ~n35233 & ~n35234 ;
  assign n35236 = ~n34503 & ~n34516 ;
  assign n35237 = n35235 & n35236 ;
  assign n35238 = ~n35235 & ~n35236 ;
  assign n35239 = ~n35237 & ~n35238 ;
  assign n35240 = ~x96 & n12506 ;
  assign n35241 = ~x94 & n13131 ;
  assign n35242 = ~x95 & n12501 ;
  assign n35243 = ~n35241 & ~n35242 ;
  assign n35244 = ~n35240 & n35243 ;
  assign n35245 = n7531 & n12509 ;
  assign n35246 = n35244 & ~n35245 ;
  assign n35247 = ~x44 & ~n35246 ;
  assign n35248 = ~x44 & ~n35247 ;
  assign n35249 = ~n35246 & ~n35247 ;
  assign n35250 = ~n35248 & ~n35249 ;
  assign n35251 = ~n35239 & n35250 ;
  assign n35252 = n35239 & ~n35250 ;
  assign n35253 = ~n35251 & ~n35252 ;
  assign n35254 = ~n34522 & ~n34536 ;
  assign n35255 = n35253 & ~n35254 ;
  assign n35256 = ~n35253 & n35254 ;
  assign n35257 = ~n35255 & ~n35256 ;
  assign n35258 = ~x99 & n10905 ;
  assign n35259 = ~x97 & n11466 ;
  assign n35260 = ~x98 & n10900 ;
  assign n35261 = ~n35259 & ~n35260 ;
  assign n35262 = ~n35258 & n35261 ;
  assign n35263 = n8885 & n10908 ;
  assign n35264 = n35262 & ~n35263 ;
  assign n35265 = ~x41 & ~n35264 ;
  assign n35266 = ~x41 & ~n35265 ;
  assign n35267 = ~n35264 & ~n35265 ;
  assign n35268 = ~n35266 & ~n35267 ;
  assign n35269 = n35257 & ~n35268 ;
  assign n35270 = n35257 & ~n35269 ;
  assign n35271 = ~n35268 & ~n35269 ;
  assign n35272 = ~n35270 & ~n35271 ;
  assign n35273 = ~n34538 & ~n34541 ;
  assign n35274 = n35272 & n35273 ;
  assign n35275 = ~n35272 & ~n35273 ;
  assign n35276 = ~n35274 & ~n35275 ;
  assign n35277 = ~x102 & n9433 ;
  assign n35278 = ~x100 & n9915 ;
  assign n35279 = ~x101 & n9428 ;
  assign n35280 = ~n35278 & ~n35279 ;
  assign n35281 = ~n35277 & n35280 ;
  assign n35282 = n9436 & n10333 ;
  assign n35283 = n35281 & ~n35282 ;
  assign n35284 = ~x38 & ~n35283 ;
  assign n35285 = ~x38 & ~n35284 ;
  assign n35286 = ~n35283 & ~n35284 ;
  assign n35287 = ~n35285 & ~n35286 ;
  assign n35288 = ~n35276 & n35287 ;
  assign n35289 = n35276 & ~n35287 ;
  assign n35290 = ~n35288 & ~n35289 ;
  assign n35291 = ~n35118 & n35290 ;
  assign n35292 = n35118 & ~n35290 ;
  assign n35293 = ~n35291 & ~n35292 ;
  assign n35294 = ~n35117 & n35293 ;
  assign n35295 = ~n35117 & ~n35294 ;
  assign n35296 = n35293 & ~n35294 ;
  assign n35297 = ~n35295 & ~n35296 ;
  assign n35298 = n35106 & ~n35297 ;
  assign n35299 = n35106 & ~n35298 ;
  assign n35300 = ~n35297 & ~n35298 ;
  assign n35301 = ~n35299 & ~n35300 ;
  assign n35302 = n35091 & ~n35301 ;
  assign n35303 = ~n35091 & n35301 ;
  assign n35304 = n35076 & ~n35303 ;
  assign n35305 = ~n35302 & n35304 ;
  assign n35306 = n35076 & ~n35305 ;
  assign n35307 = ~n35303 & ~n35305 ;
  assign n35308 = ~n35302 & n35307 ;
  assign n35309 = ~n35306 & ~n35308 ;
  assign n35310 = ~n34344 & ~n34584 ;
  assign n35311 = ~x117 & n3589 ;
  assign n35312 = ~x115 & n3878 ;
  assign n35313 = ~x116 & n3584 ;
  assign n35314 = ~n35312 & ~n35313 ;
  assign n35315 = ~n35311 & n35314 ;
  assign n35316 = ~n3592 & n35315 ;
  assign n35317 = ~n19365 & n35315 ;
  assign n35318 = ~n35316 & ~n35317 ;
  assign n35319 = ~x23 & ~n35318 ;
  assign n35320 = x23 & n35318 ;
  assign n35321 = ~n35319 & ~n35320 ;
  assign n35322 = ~n35310 & ~n35321 ;
  assign n35323 = ~n35310 & ~n35322 ;
  assign n35324 = ~n35321 & ~n35322 ;
  assign n35325 = ~n35323 & ~n35324 ;
  assign n35326 = ~n35309 & ~n35325 ;
  assign n35327 = ~n35309 & ~n35326 ;
  assign n35328 = ~n35325 & ~n35326 ;
  assign n35329 = ~n35327 & ~n35328 ;
  assign n35330 = ~n35061 & ~n35329 ;
  assign n35331 = ~n35061 & ~n35330 ;
  assign n35332 = ~n35329 & ~n35330 ;
  assign n35333 = ~n35331 & ~n35332 ;
  assign n35334 = n35045 & ~n35333 ;
  assign n35335 = ~n35045 & n35333 ;
  assign n35336 = n35030 & ~n35335 ;
  assign n35337 = ~n35334 & n35336 ;
  assign n35338 = n35030 & ~n35337 ;
  assign n35339 = ~n35335 & ~n35337 ;
  assign n35340 = ~n35334 & n35339 ;
  assign n35341 = ~n35338 & ~n35340 ;
  assign n35342 = ~n35015 & n35341 ;
  assign n35343 = n35015 & ~n35341 ;
  assign n35344 = ~n35342 & ~n35343 ;
  assign n35345 = ~n35003 & ~n35344 ;
  assign n35346 = ~n35003 & ~n35345 ;
  assign n35347 = ~n35344 & ~n35345 ;
  assign n35348 = ~n35346 & ~n35347 ;
  assign n35349 = ~n35002 & ~n35348 ;
  assign n35350 = n35002 & ~n35347 ;
  assign n35351 = ~n35346 & n35350 ;
  assign n35352 = ~n35349 & ~n35351 ;
  assign n35355 = ~n35352 & ~x202 ;
  assign n35356 = ~n35354 & ~n35355 ;
  assign n35357 = ~n34994 & ~n34998 ;
  assign n35358 = ~n34664 & ~n34990 ;
  assign n35359 = ~n34661 & ~n35358 ;
  assign n35360 = ~n34677 & ~n34986 ;
  assign n35361 = x127 & n1434 ;
  assign n35362 = x125 & n1646 ;
  assign n35363 = x126 & n1429 ;
  assign n35364 = ~n35362 & ~n35363 ;
  assign n35365 = ~n35361 & n35364 ;
  assign n35366 = n1437 & n26533 ;
  assign n35367 = n35365 & ~n35366 ;
  assign n35368 = x14 & ~n35367 ;
  assign n35369 = x14 & ~n35368 ;
  assign n35370 = ~n35367 & ~n35368 ;
  assign n35371 = ~n35369 & ~n35370 ;
  assign n35372 = ~n35360 & ~n35371 ;
  assign n35373 = ~n35360 & ~n35372 ;
  assign n35374 = ~n35371 & ~n35372 ;
  assign n35375 = ~n35373 & ~n35374 ;
  assign n35376 = ~n34693 & ~n34983 ;
  assign n35377 = x124 & n2093 ;
  assign n35378 = x122 & n2275 ;
  assign n35379 = x123 & n2088 ;
  assign n35380 = ~n35378 & ~n35379 ;
  assign n35381 = ~n35377 & n35380 ;
  assign n35382 = n2096 & n23796 ;
  assign n35383 = n35381 & ~n35382 ;
  assign n35384 = x17 & ~n35383 ;
  assign n35385 = x17 & ~n35384 ;
  assign n35386 = ~n35383 & ~n35384 ;
  assign n35387 = ~n35385 & ~n35386 ;
  assign n35388 = ~n35376 & n35387 ;
  assign n35389 = n35376 & ~n35387 ;
  assign n35390 = ~n35388 & ~n35389 ;
  assign n35391 = x121 & n2751 ;
  assign n35392 = x119 & n3020 ;
  assign n35393 = x120 & n2746 ;
  assign n35394 = ~n35392 & ~n35393 ;
  assign n35395 = ~n35391 & n35394 ;
  assign n35396 = n2754 & n21870 ;
  assign n35397 = n35395 & ~n35396 ;
  assign n35398 = x20 & ~n35397 ;
  assign n35399 = x20 & ~n35398 ;
  assign n35400 = ~n35397 & ~n35398 ;
  assign n35401 = ~n35399 & ~n35400 ;
  assign n35402 = ~n34707 & ~n34979 ;
  assign n35403 = n35401 & n35402 ;
  assign n35404 = ~n35401 & ~n35402 ;
  assign n35405 = ~n35403 & ~n35404 ;
  assign n35406 = ~n34971 & ~n34975 ;
  assign n35407 = x118 & n3589 ;
  assign n35408 = x116 & n3878 ;
  assign n35409 = x117 & n3584 ;
  assign n35410 = ~n35408 & ~n35409 ;
  assign n35411 = ~n35407 & n35410 ;
  assign n35412 = n3592 & n19395 ;
  assign n35413 = n35411 & ~n35412 ;
  assign n35414 = x23 & ~n35413 ;
  assign n35415 = x23 & ~n35414 ;
  assign n35416 = ~n35413 & ~n35414 ;
  assign n35417 = ~n35415 & ~n35416 ;
  assign n35418 = ~n35406 & ~n35417 ;
  assign n35419 = ~n35406 & ~n35418 ;
  assign n35420 = ~n35417 & ~n35418 ;
  assign n35421 = ~n35419 & ~n35420 ;
  assign n35422 = x115 & n4531 ;
  assign n35423 = x113 & n4847 ;
  assign n35424 = x114 & n4526 ;
  assign n35425 = ~n35423 & ~n35424 ;
  assign n35426 = ~n35422 & n35425 ;
  assign n35427 = n4534 & n17364 ;
  assign n35428 = n35426 & ~n35427 ;
  assign n35429 = x26 & ~n35428 ;
  assign n35430 = x26 & ~n35429 ;
  assign n35431 = ~n35428 & ~n35429 ;
  assign n35432 = ~n35430 & ~n35431 ;
  assign n35433 = ~n34723 & ~n34954 ;
  assign n35434 = n35432 & n35433 ;
  assign n35435 = ~n35432 & ~n35433 ;
  assign n35436 = ~n35434 & ~n35435 ;
  assign n35437 = ~n34739 & ~n34951 ;
  assign n35438 = x112 & n5560 ;
  assign n35439 = x110 & n5943 ;
  assign n35440 = x111 & n5555 ;
  assign n35441 = ~n35439 & ~n35440 ;
  assign n35442 = ~n35438 & n35441 ;
  assign n35443 = n5563 & n15442 ;
  assign n35444 = n35442 & ~n35443 ;
  assign n35445 = x29 & ~n35444 ;
  assign n35446 = x29 & ~n35445 ;
  assign n35447 = ~n35444 & ~n35445 ;
  assign n35448 = ~n35446 & ~n35447 ;
  assign n35449 = ~n35437 & n35448 ;
  assign n35450 = n35437 & ~n35448 ;
  assign n35451 = ~n35449 & ~n35450 ;
  assign n35452 = ~n34940 & ~n34943 ;
  assign n35453 = ~n34924 & ~n34938 ;
  assign n35454 = ~n34904 & ~n34918 ;
  assign n35455 = ~n34887 & ~n34901 ;
  assign n35456 = ~n34867 & ~n34881 ;
  assign n35457 = ~n34853 & ~n34857 ;
  assign n35458 = x88 & n18025 ;
  assign n35459 = x86 & n18764 ;
  assign n35460 = x87 & n18020 ;
  assign n35461 = ~n35459 & ~n35460 ;
  assign n35462 = ~n35458 & n35461 ;
  assign n35463 = n4305 & n18028 ;
  assign n35464 = n35462 & ~n35463 ;
  assign n35465 = x53 & ~n35464 ;
  assign n35466 = x53 & ~n35465 ;
  assign n35467 = ~n35464 & ~n35465 ;
  assign n35468 = ~n35466 & ~n35467 ;
  assign n35469 = ~n34797 & ~n34801 ;
  assign n35470 = x79 & n24612 ;
  assign n35471 = x77 & n25390 ;
  assign n35472 = x78 & n24607 ;
  assign n35473 = ~n35471 & ~n35472 ;
  assign n35474 = ~n35470 & n35473 ;
  assign n35475 = n1817 & n24615 ;
  assign n35476 = n35474 & ~n35475 ;
  assign n35477 = x62 & ~n35476 ;
  assign n35478 = x62 & ~n35477 ;
  assign n35479 = ~n35476 & ~n35477 ;
  assign n35480 = ~n35478 & ~n35479 ;
  assign n35481 = x75 & n27024 ;
  assign n35482 = x76 & ~n26217 ;
  assign n35483 = ~n35481 & ~n35482 ;
  assign n35484 = x11 & ~n34047 ;
  assign n35485 = ~x11 & n34047 ;
  assign n35486 = ~n35484 & ~n35485 ;
  assign n35487 = ~n35483 & ~n35486 ;
  assign n35488 = n35483 & n35486 ;
  assign n35489 = ~n35487 & ~n35488 ;
  assign n35490 = ~n35480 & n35489 ;
  assign n35491 = ~n35480 & ~n35490 ;
  assign n35492 = n35489 & ~n35490 ;
  assign n35493 = ~n35491 & ~n35492 ;
  assign n35494 = ~n35469 & ~n35493 ;
  assign n35495 = ~n35469 & ~n35494 ;
  assign n35496 = ~n35493 & ~n35494 ;
  assign n35497 = ~n35495 & ~n35496 ;
  assign n35498 = x82 & n22325 ;
  assign n35499 = x80 & n23066 ;
  assign n35500 = x81 & n22320 ;
  assign n35501 = ~n35499 & ~n35500 ;
  assign n35502 = ~n35498 & n35501 ;
  assign n35503 = n2584 & n22328 ;
  assign n35504 = n35502 & ~n35503 ;
  assign n35505 = x59 & ~n35504 ;
  assign n35506 = x59 & ~n35505 ;
  assign n35507 = ~n35504 & ~n35505 ;
  assign n35508 = ~n35506 & ~n35507 ;
  assign n35509 = ~n35497 & ~n35508 ;
  assign n35510 = ~n35497 & ~n35509 ;
  assign n35511 = ~n35508 & ~n35509 ;
  assign n35512 = ~n35510 & ~n35511 ;
  assign n35513 = ~n34816 & ~n34831 ;
  assign n35514 = n35512 & n35513 ;
  assign n35515 = ~n35512 & ~n35513 ;
  assign n35516 = ~n35514 & ~n35515 ;
  assign n35517 = x85 & n20143 ;
  assign n35518 = x83 & n20854 ;
  assign n35519 = x84 & n20138 ;
  assign n35520 = ~n35518 & ~n35519 ;
  assign n35521 = ~n35517 & n35520 ;
  assign n35522 = n3389 & n20146 ;
  assign n35523 = n35521 & ~n35522 ;
  assign n35524 = x56 & ~n35523 ;
  assign n35525 = x56 & ~n35524 ;
  assign n35526 = ~n35523 & ~n35524 ;
  assign n35527 = ~n35525 & ~n35526 ;
  assign n35528 = n35516 & ~n35527 ;
  assign n35529 = n35516 & ~n35528 ;
  assign n35530 = ~n35527 & ~n35528 ;
  assign n35531 = ~n35529 & ~n35530 ;
  assign n35532 = ~n34837 & ~n34851 ;
  assign n35533 = ~n35531 & ~n35532 ;
  assign n35534 = n35531 & n35532 ;
  assign n35535 = ~n35533 & ~n35534 ;
  assign n35536 = ~n35468 & n35535 ;
  assign n35537 = ~n35468 & ~n35536 ;
  assign n35538 = n35535 & ~n35536 ;
  assign n35539 = ~n35537 & ~n35538 ;
  assign n35540 = ~n35457 & ~n35539 ;
  assign n35541 = ~n35457 & ~n35540 ;
  assign n35542 = ~n35539 & ~n35540 ;
  assign n35543 = ~n35541 & ~n35542 ;
  assign n35544 = x91 & n16076 ;
  assign n35545 = x89 & n16756 ;
  assign n35546 = x90 & n16071 ;
  assign n35547 = ~n35545 & ~n35546 ;
  assign n35548 = ~n35544 & n35547 ;
  assign n35549 = n5336 & n16079 ;
  assign n35550 = n35548 & ~n35549 ;
  assign n35551 = x50 & ~n35550 ;
  assign n35552 = x50 & ~n35551 ;
  assign n35553 = ~n35550 & ~n35551 ;
  assign n35554 = ~n35552 & ~n35553 ;
  assign n35555 = ~n35543 & ~n35554 ;
  assign n35556 = ~n35543 & ~n35555 ;
  assign n35557 = ~n35554 & ~n35555 ;
  assign n35558 = ~n35556 & ~n35557 ;
  assign n35559 = ~n34861 & ~n34864 ;
  assign n35560 = n35558 & n35559 ;
  assign n35561 = ~n35558 & ~n35559 ;
  assign n35562 = ~n35560 & ~n35561 ;
  assign n35563 = x94 & n14233 ;
  assign n35564 = x92 & n14876 ;
  assign n35565 = x93 & n14228 ;
  assign n35566 = ~n35564 & ~n35565 ;
  assign n35567 = ~n35563 & n35566 ;
  assign n35568 = n6483 & n14236 ;
  assign n35569 = n35567 & ~n35568 ;
  assign n35570 = x47 & ~n35569 ;
  assign n35571 = x47 & ~n35570 ;
  assign n35572 = ~n35569 & ~n35570 ;
  assign n35573 = ~n35571 & ~n35572 ;
  assign n35574 = n35562 & ~n35573 ;
  assign n35575 = ~n35562 & n35573 ;
  assign n35576 = ~n35456 & ~n35575 ;
  assign n35577 = ~n35574 & n35576 ;
  assign n35578 = ~n35456 & ~n35577 ;
  assign n35579 = ~n35574 & ~n35577 ;
  assign n35580 = ~n35575 & n35579 ;
  assign n35581 = ~n35578 & ~n35580 ;
  assign n35582 = x97 & n12506 ;
  assign n35583 = x95 & n13131 ;
  assign n35584 = x96 & n12501 ;
  assign n35585 = ~n35583 & ~n35584 ;
  assign n35586 = ~n35582 & n35585 ;
  assign n35587 = n7745 & n12509 ;
  assign n35588 = n35586 & ~n35587 ;
  assign n35589 = x44 & ~n35588 ;
  assign n35590 = x44 & ~n35589 ;
  assign n35591 = ~n35588 & ~n35589 ;
  assign n35592 = ~n35590 & ~n35591 ;
  assign n35593 = ~n35581 & ~n35592 ;
  assign n35594 = ~n35581 & ~n35593 ;
  assign n35595 = ~n35592 & ~n35593 ;
  assign n35596 = ~n35594 & ~n35595 ;
  assign n35597 = ~n35455 & n35596 ;
  assign n35598 = n35455 & ~n35596 ;
  assign n35599 = ~n35597 & ~n35598 ;
  assign n35600 = x100 & n10905 ;
  assign n35601 = x98 & n11466 ;
  assign n35602 = x99 & n10900 ;
  assign n35603 = ~n35601 & ~n35602 ;
  assign n35604 = ~n35600 & n35603 ;
  assign n35605 = n9115 & n10908 ;
  assign n35606 = n35604 & ~n35605 ;
  assign n35607 = x41 & ~n35606 ;
  assign n35608 = x41 & ~n35607 ;
  assign n35609 = ~n35606 & ~n35607 ;
  assign n35610 = ~n35608 & ~n35609 ;
  assign n35611 = ~n35599 & ~n35610 ;
  assign n35612 = n35599 & n35610 ;
  assign n35613 = ~n35611 & ~n35612 ;
  assign n35614 = n35454 & ~n35613 ;
  assign n35615 = ~n35454 & n35613 ;
  assign n35616 = ~n35614 & ~n35615 ;
  assign n35617 = x103 & n9433 ;
  assign n35618 = x101 & n9915 ;
  assign n35619 = x102 & n9428 ;
  assign n35620 = ~n35618 & ~n35619 ;
  assign n35621 = ~n35617 & n35620 ;
  assign n35622 = n9436 & n10588 ;
  assign n35623 = n35621 & ~n35622 ;
  assign n35624 = x38 & ~n35623 ;
  assign n35625 = x38 & ~n35624 ;
  assign n35626 = ~n35623 & ~n35624 ;
  assign n35627 = ~n35625 & ~n35626 ;
  assign n35628 = n35616 & ~n35627 ;
  assign n35629 = n35616 & ~n35628 ;
  assign n35630 = ~n35627 & ~n35628 ;
  assign n35631 = ~n35629 & ~n35630 ;
  assign n35632 = ~n35453 & n35631 ;
  assign n35633 = n35453 & ~n35631 ;
  assign n35634 = ~n35632 & ~n35633 ;
  assign n35635 = x106 & n8006 ;
  assign n35636 = x104 & n8474 ;
  assign n35637 = x105 & n8001 ;
  assign n35638 = ~n35636 & ~n35637 ;
  assign n35639 = ~n35635 & n35638 ;
  assign n35640 = n8009 & n12181 ;
  assign n35641 = n35639 & ~n35640 ;
  assign n35642 = x35 & ~n35641 ;
  assign n35643 = x35 & ~n35642 ;
  assign n35644 = ~n35641 & ~n35642 ;
  assign n35645 = ~n35643 & ~n35644 ;
  assign n35646 = ~n35634 & ~n35645 ;
  assign n35647 = n35634 & n35645 ;
  assign n35648 = ~n35646 & ~n35647 ;
  assign n35649 = n35452 & ~n35648 ;
  assign n35650 = ~n35452 & n35648 ;
  assign n35651 = ~n35649 & ~n35650 ;
  assign n35652 = ~n34753 & ~n34947 ;
  assign n35653 = x109 & n6725 ;
  assign n35654 = x107 & n7129 ;
  assign n35655 = x108 & n6720 ;
  assign n35656 = ~n35654 & ~n35655 ;
  assign n35657 = ~n35653 & n35656 ;
  assign n35658 = n6728 & n13894 ;
  assign n35659 = n35657 & ~n35658 ;
  assign n35660 = x32 & ~n35659 ;
  assign n35661 = x32 & ~n35660 ;
  assign n35662 = ~n35659 & ~n35660 ;
  assign n35663 = ~n35661 & ~n35662 ;
  assign n35664 = ~n35652 & ~n35663 ;
  assign n35665 = ~n35652 & ~n35664 ;
  assign n35666 = ~n35663 & ~n35664 ;
  assign n35667 = ~n35665 & ~n35666 ;
  assign n35668 = n35651 & ~n35667 ;
  assign n35669 = ~n35651 & n35667 ;
  assign n35670 = ~n35451 & ~n35669 ;
  assign n35671 = ~n35668 & n35670 ;
  assign n35672 = ~n35451 & ~n35671 ;
  assign n35673 = ~n35669 & ~n35671 ;
  assign n35674 = ~n35668 & n35673 ;
  assign n35675 = ~n35672 & ~n35674 ;
  assign n35676 = n35436 & ~n35675 ;
  assign n35677 = ~n35436 & n35675 ;
  assign n35678 = ~n35421 & ~n35677 ;
  assign n35679 = ~n35676 & n35678 ;
  assign n35680 = ~n35421 & ~n35679 ;
  assign n35681 = ~n35677 & ~n35679 ;
  assign n35682 = ~n35676 & n35681 ;
  assign n35683 = ~n35680 & ~n35682 ;
  assign n35684 = n35405 & ~n35683 ;
  assign n35685 = ~n35405 & n35683 ;
  assign n35686 = ~n35390 & ~n35685 ;
  assign n35687 = ~n35684 & n35686 ;
  assign n35688 = ~n35390 & ~n35687 ;
  assign n35689 = ~n35685 & ~n35687 ;
  assign n35690 = ~n35684 & n35689 ;
  assign n35691 = ~n35688 & ~n35690 ;
  assign n35692 = ~n35375 & n35691 ;
  assign n35693 = n35375 & ~n35691 ;
  assign n35694 = ~n35692 & ~n35693 ;
  assign n35695 = ~n35359 & ~n35694 ;
  assign n35696 = ~n35359 & ~n35695 ;
  assign n35697 = ~n35694 & ~n35695 ;
  assign n35698 = ~n35696 & ~n35697 ;
  assign n35699 = ~n35357 & ~n35698 ;
  assign n35700 = n35357 & ~n35697 ;
  assign n35701 = ~n35696 & n35700 ;
  assign n35702 = ~n35699 & ~n35701 ;
  assign n36050 = n35702 & x203 ;
  assign n35703 = ~n35345 & ~n35349 ;
  assign n35704 = ~n35015 & ~n35341 ;
  assign n35705 = ~n35012 & ~n35704 ;
  assign n35706 = ~n35028 & ~n35337 ;
  assign n35707 = ~x127 & n1434 ;
  assign n35708 = ~x125 & n1646 ;
  assign n35709 = ~x126 & n1429 ;
  assign n35710 = ~n35708 & ~n35709 ;
  assign n35711 = ~n35707 & n35710 ;
  assign n35712 = n1437 & n26932 ;
  assign n35713 = n35711 & ~n35712 ;
  assign n35714 = ~x14 & ~n35713 ;
  assign n35715 = ~x14 & ~n35714 ;
  assign n35716 = ~n35713 & ~n35714 ;
  assign n35717 = ~n35715 & ~n35716 ;
  assign n35718 = ~n35706 & ~n35717 ;
  assign n35719 = ~n35706 & ~n35718 ;
  assign n35720 = ~n35717 & ~n35718 ;
  assign n35721 = ~n35719 & ~n35720 ;
  assign n35722 = ~n35044 & ~n35334 ;
  assign n35723 = ~x124 & n2093 ;
  assign n35724 = ~x122 & n2275 ;
  assign n35725 = ~x123 & n2088 ;
  assign n35726 = ~n35724 & ~n35725 ;
  assign n35727 = ~n35723 & n35726 ;
  assign n35728 = n2096 & n24176 ;
  assign n35729 = n35727 & ~n35728 ;
  assign n35730 = ~x17 & ~n35729 ;
  assign n35731 = ~x17 & ~n35730 ;
  assign n35732 = ~n35729 & ~n35730 ;
  assign n35733 = ~n35731 & ~n35732 ;
  assign n35734 = ~n35722 & n35733 ;
  assign n35735 = n35722 & ~n35733 ;
  assign n35736 = ~n35734 & ~n35735 ;
  assign n35737 = ~x121 & n2751 ;
  assign n35738 = ~x119 & n3020 ;
  assign n35739 = ~x120 & n2746 ;
  assign n35740 = ~n35738 & ~n35739 ;
  assign n35741 = ~n35737 & n35740 ;
  assign n35742 = n2754 & n22229 ;
  assign n35743 = n35741 & ~n35742 ;
  assign n35744 = ~x20 & ~n35743 ;
  assign n35745 = ~x20 & ~n35744 ;
  assign n35746 = ~n35743 & ~n35744 ;
  assign n35747 = ~n35745 & ~n35746 ;
  assign n35748 = ~n35058 & ~n35330 ;
  assign n35749 = n35747 & n35748 ;
  assign n35750 = ~n35747 & ~n35748 ;
  assign n35751 = ~n35749 & ~n35750 ;
  assign n35752 = ~n35322 & ~n35326 ;
  assign n35753 = ~x118 & n3589 ;
  assign n35754 = ~x116 & n3878 ;
  assign n35755 = ~x117 & n3584 ;
  assign n35756 = ~n35754 & ~n35755 ;
  assign n35757 = ~n35753 & n35756 ;
  assign n35758 = n3592 & n19736 ;
  assign n35759 = n35757 & ~n35758 ;
  assign n35760 = ~x23 & ~n35759 ;
  assign n35761 = ~x23 & ~n35760 ;
  assign n35762 = ~n35759 & ~n35760 ;
  assign n35763 = ~n35761 & ~n35762 ;
  assign n35764 = ~n35752 & ~n35763 ;
  assign n35765 = ~n35752 & ~n35764 ;
  assign n35766 = ~n35763 & ~n35764 ;
  assign n35767 = ~n35765 & ~n35766 ;
  assign n35768 = ~x115 & n4531 ;
  assign n35769 = ~x113 & n4847 ;
  assign n35770 = ~x114 & n4526 ;
  assign n35771 = ~n35769 & ~n35770 ;
  assign n35772 = ~n35768 & n35771 ;
  assign n35773 = n4534 & n17683 ;
  assign n35774 = n35772 & ~n35773 ;
  assign n35775 = ~x26 & ~n35774 ;
  assign n35776 = ~x26 & ~n35775 ;
  assign n35777 = ~n35774 & ~n35775 ;
  assign n35778 = ~n35776 & ~n35777 ;
  assign n35779 = ~n35074 & ~n35305 ;
  assign n35780 = n35778 & n35779 ;
  assign n35781 = ~n35778 & ~n35779 ;
  assign n35782 = ~n35780 & ~n35781 ;
  assign n35783 = ~n35090 & ~n35302 ;
  assign n35784 = ~x112 & n5560 ;
  assign n35785 = ~x110 & n5943 ;
  assign n35786 = ~x111 & n5555 ;
  assign n35787 = ~n35785 & ~n35786 ;
  assign n35788 = ~n35784 & n35787 ;
  assign n35789 = n5563 & n15744 ;
  assign n35790 = n35788 & ~n35789 ;
  assign n35791 = ~x29 & ~n35790 ;
  assign n35792 = ~x29 & ~n35791 ;
  assign n35793 = ~n35790 & ~n35791 ;
  assign n35794 = ~n35792 & ~n35793 ;
  assign n35795 = ~n35783 & n35794 ;
  assign n35796 = n35783 & ~n35794 ;
  assign n35797 = ~n35795 & ~n35796 ;
  assign n35798 = ~n35291 & ~n35294 ;
  assign n35799 = ~n35275 & ~n35289 ;
  assign n35800 = ~n35255 & ~n35269 ;
  assign n35801 = ~n35238 & ~n35252 ;
  assign n35802 = ~n35218 & ~n35232 ;
  assign n35803 = ~n35204 & ~n35208 ;
  assign n35804 = ~x88 & n18025 ;
  assign n35805 = ~x86 & n18764 ;
  assign n35806 = ~x87 & n18020 ;
  assign n35807 = ~n35805 & ~n35806 ;
  assign n35808 = ~n35804 & n35807 ;
  assign n35809 = n4457 & n18028 ;
  assign n35810 = n35808 & ~n35809 ;
  assign n35811 = ~x53 & ~n35810 ;
  assign n35812 = ~x53 & ~n35811 ;
  assign n35813 = ~n35810 & ~n35811 ;
  assign n35814 = ~n35812 & ~n35813 ;
  assign n35815 = ~n35148 & ~n35152 ;
  assign n35816 = ~x79 & n24612 ;
  assign n35817 = ~x77 & n25390 ;
  assign n35818 = ~x78 & n24607 ;
  assign n35819 = ~n35817 & ~n35818 ;
  assign n35820 = ~n35816 & n35819 ;
  assign n35821 = n1921 & n24615 ;
  assign n35822 = n35820 & ~n35821 ;
  assign n35823 = ~x62 & ~n35822 ;
  assign n35824 = ~x62 & ~n35823 ;
  assign n35825 = ~n35822 & ~n35823 ;
  assign n35826 = ~n35824 & ~n35825 ;
  assign n35827 = ~x75 & n27427 ;
  assign n35828 = ~x76 & ~n26217 ;
  assign n35829 = ~n35827 & ~n35828 ;
  assign n35830 = ~x11 & ~n34412 ;
  assign n35831 = x11 & n34412 ;
  assign n35832 = ~n35830 & ~n35831 ;
  assign n35833 = ~n35829 & ~n35832 ;
  assign n35834 = n35829 & n35832 ;
  assign n35835 = ~n35833 & ~n35834 ;
  assign n35836 = ~n35826 & n35835 ;
  assign n35837 = ~n35826 & ~n35836 ;
  assign n35838 = n35835 & ~n35836 ;
  assign n35839 = ~n35837 & ~n35838 ;
  assign n35840 = ~n35815 & ~n35839 ;
  assign n35841 = ~n35815 & ~n35840 ;
  assign n35842 = ~n35839 & ~n35840 ;
  assign n35843 = ~n35841 & ~n35842 ;
  assign n35844 = ~x82 & n22325 ;
  assign n35845 = ~x80 & n23066 ;
  assign n35846 = ~x81 & n22320 ;
  assign n35847 = ~n35845 & ~n35846 ;
  assign n35848 = ~n35844 & n35847 ;
  assign n35849 = n2697 & n22328 ;
  assign n35850 = n35848 & ~n35849 ;
  assign n35851 = ~x59 & ~n35850 ;
  assign n35852 = ~x59 & ~n35851 ;
  assign n35853 = ~n35850 & ~n35851 ;
  assign n35854 = ~n35852 & ~n35853 ;
  assign n35855 = ~n35843 & ~n35854 ;
  assign n35856 = ~n35843 & ~n35855 ;
  assign n35857 = ~n35854 & ~n35855 ;
  assign n35858 = ~n35856 & ~n35857 ;
  assign n35859 = ~n35167 & ~n35182 ;
  assign n35860 = n35858 & n35859 ;
  assign n35861 = ~n35858 & ~n35859 ;
  assign n35862 = ~n35860 & ~n35861 ;
  assign n35863 = ~x85 & n20143 ;
  assign n35864 = ~x83 & n20854 ;
  assign n35865 = ~x84 & n20138 ;
  assign n35866 = ~n35864 & ~n35865 ;
  assign n35867 = ~n35863 & n35866 ;
  assign n35868 = n3521 & n20146 ;
  assign n35869 = n35867 & ~n35868 ;
  assign n35870 = ~x56 & ~n35869 ;
  assign n35871 = ~x56 & ~n35870 ;
  assign n35872 = ~n35869 & ~n35870 ;
  assign n35873 = ~n35871 & ~n35872 ;
  assign n35874 = n35862 & ~n35873 ;
  assign n35875 = n35862 & ~n35874 ;
  assign n35876 = ~n35873 & ~n35874 ;
  assign n35877 = ~n35875 & ~n35876 ;
  assign n35878 = ~n35188 & ~n35202 ;
  assign n35879 = ~n35877 & ~n35878 ;
  assign n35880 = n35877 & n35878 ;
  assign n35881 = ~n35879 & ~n35880 ;
  assign n35882 = ~n35814 & n35881 ;
  assign n35883 = ~n35814 & ~n35882 ;
  assign n35884 = n35881 & ~n35882 ;
  assign n35885 = ~n35883 & ~n35884 ;
  assign n35886 = ~n35803 & ~n35885 ;
  assign n35887 = ~n35803 & ~n35886 ;
  assign n35888 = ~n35885 & ~n35886 ;
  assign n35889 = ~n35887 & ~n35888 ;
  assign n35890 = ~x91 & n16076 ;
  assign n35891 = ~x89 & n16756 ;
  assign n35892 = ~x90 & n16071 ;
  assign n35893 = ~n35891 & ~n35892 ;
  assign n35894 = ~n35890 & n35893 ;
  assign n35895 = n5507 & n16079 ;
  assign n35896 = n35894 & ~n35895 ;
  assign n35897 = ~x50 & ~n35896 ;
  assign n35898 = ~x50 & ~n35897 ;
  assign n35899 = ~n35896 & ~n35897 ;
  assign n35900 = ~n35898 & ~n35899 ;
  assign n35901 = ~n35889 & ~n35900 ;
  assign n35902 = ~n35889 & ~n35901 ;
  assign n35903 = ~n35900 & ~n35901 ;
  assign n35904 = ~n35902 & ~n35903 ;
  assign n35905 = ~n35212 & ~n35215 ;
  assign n35906 = n35904 & n35905 ;
  assign n35907 = ~n35904 & ~n35905 ;
  assign n35908 = ~n35906 & ~n35907 ;
  assign n35909 = ~x94 & n14233 ;
  assign n35910 = ~x92 & n14876 ;
  assign n35911 = ~x93 & n14228 ;
  assign n35912 = ~n35910 & ~n35911 ;
  assign n35913 = ~n35909 & n35912 ;
  assign n35914 = n6671 & n14236 ;
  assign n35915 = n35913 & ~n35914 ;
  assign n35916 = ~x47 & ~n35915 ;
  assign n35917 = ~x47 & ~n35916 ;
  assign n35918 = ~n35915 & ~n35916 ;
  assign n35919 = ~n35917 & ~n35918 ;
  assign n35920 = n35908 & ~n35919 ;
  assign n35921 = ~n35908 & n35919 ;
  assign n35922 = ~n35802 & ~n35921 ;
  assign n35923 = ~n35920 & n35922 ;
  assign n35924 = ~n35802 & ~n35923 ;
  assign n35925 = ~n35920 & ~n35923 ;
  assign n35926 = ~n35921 & n35925 ;
  assign n35927 = ~n35924 & ~n35926 ;
  assign n35928 = ~x97 & n12506 ;
  assign n35929 = ~x95 & n13131 ;
  assign n35930 = ~x96 & n12501 ;
  assign n35931 = ~n35929 & ~n35930 ;
  assign n35932 = ~n35928 & n35931 ;
  assign n35933 = n7949 & n12509 ;
  assign n35934 = n35932 & ~n35933 ;
  assign n35935 = ~x44 & ~n35934 ;
  assign n35936 = ~x44 & ~n35935 ;
  assign n35937 = ~n35934 & ~n35935 ;
  assign n35938 = ~n35936 & ~n35937 ;
  assign n35939 = ~n35927 & ~n35938 ;
  assign n35940 = ~n35927 & ~n35939 ;
  assign n35941 = ~n35938 & ~n35939 ;
  assign n35942 = ~n35940 & ~n35941 ;
  assign n35943 = ~n35801 & n35942 ;
  assign n35944 = n35801 & ~n35942 ;
  assign n35945 = ~n35943 & ~n35944 ;
  assign n35946 = ~x100 & n10905 ;
  assign n35947 = ~x98 & n11466 ;
  assign n35948 = ~x99 & n10900 ;
  assign n35949 = ~n35947 & ~n35948 ;
  assign n35950 = ~n35946 & n35949 ;
  assign n35951 = n9338 & n10908 ;
  assign n35952 = n35950 & ~n35951 ;
  assign n35953 = ~x41 & ~n35952 ;
  assign n35954 = ~x41 & ~n35953 ;
  assign n35955 = ~n35952 & ~n35953 ;
  assign n35956 = ~n35954 & ~n35955 ;
  assign n35957 = ~n35945 & ~n35956 ;
  assign n35958 = n35945 & n35956 ;
  assign n35959 = ~n35957 & ~n35958 ;
  assign n35960 = n35800 & ~n35959 ;
  assign n35961 = ~n35800 & n35959 ;
  assign n35962 = ~n35960 & ~n35961 ;
  assign n35963 = ~x103 & n9433 ;
  assign n35964 = ~x101 & n9915 ;
  assign n35965 = ~x102 & n9428 ;
  assign n35966 = ~n35964 & ~n35965 ;
  assign n35967 = ~n35963 & n35966 ;
  assign n35968 = n9436 & n10833 ;
  assign n35969 = n35967 & ~n35968 ;
  assign n35970 = ~x38 & ~n35969 ;
  assign n35971 = ~x38 & ~n35970 ;
  assign n35972 = ~n35969 & ~n35970 ;
  assign n35973 = ~n35971 & ~n35972 ;
  assign n35974 = n35962 & ~n35973 ;
  assign n35975 = n35962 & ~n35974 ;
  assign n35976 = ~n35973 & ~n35974 ;
  assign n35977 = ~n35975 & ~n35976 ;
  assign n35978 = ~n35799 & n35977 ;
  assign n35979 = n35799 & ~n35977 ;
  assign n35980 = ~n35978 & ~n35979 ;
  assign n35981 = ~x106 & n8006 ;
  assign n35982 = ~x104 & n8474 ;
  assign n35983 = ~x105 & n8001 ;
  assign n35984 = ~n35982 & ~n35983 ;
  assign n35985 = ~n35981 & n35984 ;
  assign n35986 = n8009 & n12447 ;
  assign n35987 = n35985 & ~n35986 ;
  assign n35988 = ~x35 & ~n35987 ;
  assign n35989 = ~x35 & ~n35988 ;
  assign n35990 = ~n35987 & ~n35988 ;
  assign n35991 = ~n35989 & ~n35990 ;
  assign n35992 = ~n35980 & ~n35991 ;
  assign n35993 = n35980 & n35991 ;
  assign n35994 = ~n35992 & ~n35993 ;
  assign n35995 = n35798 & ~n35994 ;
  assign n35996 = ~n35798 & n35994 ;
  assign n35997 = ~n35995 & ~n35996 ;
  assign n35998 = ~n35104 & ~n35298 ;
  assign n35999 = ~x109 & n6725 ;
  assign n36000 = ~x107 & n7129 ;
  assign n36001 = ~x108 & n6720 ;
  assign n36002 = ~n36000 & ~n36001 ;
  assign n36003 = ~n35999 & n36002 ;
  assign n36004 = n6728 & n14177 ;
  assign n36005 = n36003 & ~n36004 ;
  assign n36006 = ~x32 & ~n36005 ;
  assign n36007 = ~x32 & ~n36006 ;
  assign n36008 = ~n36005 & ~n36006 ;
  assign n36009 = ~n36007 & ~n36008 ;
  assign n36010 = ~n35998 & ~n36009 ;
  assign n36011 = ~n35998 & ~n36010 ;
  assign n36012 = ~n36009 & ~n36010 ;
  assign n36013 = ~n36011 & ~n36012 ;
  assign n36014 = n35997 & ~n36013 ;
  assign n36015 = ~n35997 & n36013 ;
  assign n36016 = ~n35797 & ~n36015 ;
  assign n36017 = ~n36014 & n36016 ;
  assign n36018 = ~n35797 & ~n36017 ;
  assign n36019 = ~n36015 & ~n36017 ;
  assign n36020 = ~n36014 & n36019 ;
  assign n36021 = ~n36018 & ~n36020 ;
  assign n36022 = n35782 & ~n36021 ;
  assign n36023 = ~n35782 & n36021 ;
  assign n36024 = ~n35767 & ~n36023 ;
  assign n36025 = ~n36022 & n36024 ;
  assign n36026 = ~n35767 & ~n36025 ;
  assign n36027 = ~n36023 & ~n36025 ;
  assign n36028 = ~n36022 & n36027 ;
  assign n36029 = ~n36026 & ~n36028 ;
  assign n36030 = n35751 & ~n36029 ;
  assign n36031 = ~n35751 & n36029 ;
  assign n36032 = ~n35736 & ~n36031 ;
  assign n36033 = ~n36030 & n36032 ;
  assign n36034 = ~n35736 & ~n36033 ;
  assign n36035 = ~n36031 & ~n36033 ;
  assign n36036 = ~n36030 & n36035 ;
  assign n36037 = ~n36034 & ~n36036 ;
  assign n36038 = ~n35721 & n36037 ;
  assign n36039 = n35721 & ~n36037 ;
  assign n36040 = ~n36038 & ~n36039 ;
  assign n36041 = ~n35705 & ~n36040 ;
  assign n36042 = ~n35705 & ~n36041 ;
  assign n36043 = ~n36040 & ~n36041 ;
  assign n36044 = ~n36042 & ~n36043 ;
  assign n36045 = ~n35703 & ~n36044 ;
  assign n36046 = n35703 & ~n36043 ;
  assign n36047 = ~n36042 & n36046 ;
  assign n36048 = ~n36045 & ~n36047 ;
  assign n36051 = ~n36048 & ~x203 ;
  assign n36052 = ~n36050 & ~n36051 ;
  assign n36053 = ~n35695 & ~n35699 ;
  assign n36054 = ~n35375 & ~n35691 ;
  assign n36055 = ~n35372 & ~n36054 ;
  assign n36056 = x125 & n2093 ;
  assign n36057 = x123 & n2275 ;
  assign n36058 = x124 & n2088 ;
  assign n36059 = ~n36057 & ~n36058 ;
  assign n36060 = ~n36056 & n36059 ;
  assign n36061 = n2096 & n24935 ;
  assign n36062 = n36060 & ~n36061 ;
  assign n36063 = x17 & ~n36062 ;
  assign n36064 = x17 & ~n36063 ;
  assign n36065 = ~n36062 & ~n36063 ;
  assign n36066 = ~n36064 & ~n36065 ;
  assign n36067 = ~n35404 & ~n35684 ;
  assign n36068 = ~n36066 & ~n36067 ;
  assign n36069 = ~n36066 & ~n36068 ;
  assign n36070 = ~n36067 & ~n36068 ;
  assign n36071 = ~n36069 & ~n36070 ;
  assign n36072 = x119 & n3589 ;
  assign n36073 = x117 & n3878 ;
  assign n36074 = x118 & n3584 ;
  assign n36075 = ~n36073 & ~n36074 ;
  assign n36076 = ~n36072 & n36075 ;
  assign n36077 = n3592 & n20423 ;
  assign n36078 = n36076 & ~n36077 ;
  assign n36079 = x23 & ~n36078 ;
  assign n36080 = x23 & ~n36079 ;
  assign n36081 = ~n36078 & ~n36079 ;
  assign n36082 = ~n36080 & ~n36081 ;
  assign n36083 = ~n35435 & ~n35676 ;
  assign n36084 = ~n36082 & ~n36083 ;
  assign n36085 = ~n36082 & ~n36084 ;
  assign n36086 = ~n36083 & ~n36084 ;
  assign n36087 = ~n36085 & ~n36086 ;
  assign n36088 = x113 & n5560 ;
  assign n36089 = x111 & n5943 ;
  assign n36090 = x112 & n5555 ;
  assign n36091 = ~n36089 & ~n36090 ;
  assign n36092 = ~n36088 & n36091 ;
  assign n36093 = n5563 & n16361 ;
  assign n36094 = n36092 & ~n36093 ;
  assign n36095 = x29 & ~n36094 ;
  assign n36096 = x29 & ~n36095 ;
  assign n36097 = ~n36094 & ~n36095 ;
  assign n36098 = ~n36096 & ~n36097 ;
  assign n36099 = ~n35664 & ~n35668 ;
  assign n36100 = ~n36098 & ~n36099 ;
  assign n36101 = ~n36098 & ~n36100 ;
  assign n36102 = ~n36099 & ~n36100 ;
  assign n36103 = ~n36101 & ~n36102 ;
  assign n36104 = ~n35453 & ~n35631 ;
  assign n36105 = ~n35628 & ~n36104 ;
  assign n36106 = x104 & n9433 ;
  assign n36107 = x102 & n9915 ;
  assign n36108 = x103 & n9428 ;
  assign n36109 = ~n36107 & ~n36108 ;
  assign n36110 = ~n36106 & n36109 ;
  assign n36111 = n9436 & n11116 ;
  assign n36112 = n36110 & ~n36111 ;
  assign n36113 = x38 & ~n36112 ;
  assign n36114 = x38 & ~n36113 ;
  assign n36115 = ~n36112 & ~n36113 ;
  assign n36116 = ~n36114 & ~n36115 ;
  assign n36117 = ~n35611 & ~n35615 ;
  assign n36118 = x101 & n10905 ;
  assign n36119 = x99 & n11466 ;
  assign n36120 = x100 & n10900 ;
  assign n36121 = ~n36119 & ~n36120 ;
  assign n36122 = ~n36118 & n36121 ;
  assign n36123 = n9601 & n10908 ;
  assign n36124 = n36122 & ~n36123 ;
  assign n36125 = x41 & ~n36124 ;
  assign n36126 = x41 & ~n36125 ;
  assign n36127 = ~n36124 & ~n36125 ;
  assign n36128 = ~n36126 & ~n36127 ;
  assign n36129 = ~n35455 & ~n35596 ;
  assign n36130 = ~n35593 & ~n36129 ;
  assign n36131 = x98 & n12506 ;
  assign n36132 = x96 & n13131 ;
  assign n36133 = x97 & n12501 ;
  assign n36134 = ~n36132 & ~n36133 ;
  assign n36135 = ~n36131 & n36134 ;
  assign n36136 = n8196 & n12509 ;
  assign n36137 = n36135 & ~n36136 ;
  assign n36138 = x44 & ~n36137 ;
  assign n36139 = x44 & ~n36138 ;
  assign n36140 = ~n36137 & ~n36138 ;
  assign n36141 = ~n36139 & ~n36140 ;
  assign n36142 = x95 & n14233 ;
  assign n36143 = x93 & n14876 ;
  assign n36144 = x94 & n14228 ;
  assign n36145 = ~n36143 & ~n36144 ;
  assign n36146 = ~n36142 & n36145 ;
  assign n36147 = n6894 & n14236 ;
  assign n36148 = n36146 & ~n36147 ;
  assign n36149 = x47 & ~n36148 ;
  assign n36150 = x47 & ~n36149 ;
  assign n36151 = ~n36148 & ~n36149 ;
  assign n36152 = ~n36150 & ~n36151 ;
  assign n36153 = ~n35555 & ~n35561 ;
  assign n36154 = x76 & n27024 ;
  assign n36155 = x77 & ~n26217 ;
  assign n36156 = ~n36154 & ~n36155 ;
  assign n36157 = ~x11 & ~n34047 ;
  assign n36158 = ~n35487 & ~n36157 ;
  assign n36159 = n36156 & ~n36158 ;
  assign n36160 = n36156 & ~n36159 ;
  assign n36161 = ~n36158 & ~n36159 ;
  assign n36162 = ~n36160 & ~n36161 ;
  assign n36163 = x80 & n24612 ;
  assign n36164 = x78 & n25390 ;
  assign n36165 = x79 & n24607 ;
  assign n36166 = ~n36164 & ~n36165 ;
  assign n36167 = ~n36163 & n36166 ;
  assign n36168 = n2028 & n24615 ;
  assign n36169 = n36167 & ~n36168 ;
  assign n36170 = x62 & ~n36169 ;
  assign n36171 = x62 & ~n36170 ;
  assign n36172 = ~n36169 & ~n36170 ;
  assign n36173 = ~n36171 & ~n36172 ;
  assign n36174 = ~n36162 & n36173 ;
  assign n36175 = n36162 & ~n36173 ;
  assign n36176 = ~n36174 & ~n36175 ;
  assign n36177 = ~n35490 & ~n35494 ;
  assign n36178 = n36176 & n36177 ;
  assign n36179 = ~n36176 & ~n36177 ;
  assign n36180 = ~n36178 & ~n36179 ;
  assign n36181 = x83 & n22325 ;
  assign n36182 = x81 & n23066 ;
  assign n36183 = x82 & n22320 ;
  assign n36184 = ~n36182 & ~n36183 ;
  assign n36185 = ~n36181 & n36184 ;
  assign n36186 = n2843 & n22328 ;
  assign n36187 = n36185 & ~n36186 ;
  assign n36188 = x59 & ~n36187 ;
  assign n36189 = x59 & ~n36188 ;
  assign n36190 = ~n36187 & ~n36188 ;
  assign n36191 = ~n36189 & ~n36190 ;
  assign n36192 = n36180 & ~n36191 ;
  assign n36193 = n36180 & ~n36192 ;
  assign n36194 = ~n36191 & ~n36192 ;
  assign n36195 = ~n36193 & ~n36194 ;
  assign n36196 = ~n35509 & ~n35515 ;
  assign n36197 = n36195 & n36196 ;
  assign n36198 = ~n36195 & ~n36196 ;
  assign n36199 = ~n36197 & ~n36198 ;
  assign n36200 = x86 & n20143 ;
  assign n36201 = x84 & n20854 ;
  assign n36202 = x85 & n20138 ;
  assign n36203 = ~n36201 & ~n36202 ;
  assign n36204 = ~n36200 & n36203 ;
  assign n36205 = n3686 & n20146 ;
  assign n36206 = n36204 & ~n36205 ;
  assign n36207 = x56 & ~n36206 ;
  assign n36208 = x56 & ~n36207 ;
  assign n36209 = ~n36206 & ~n36207 ;
  assign n36210 = ~n36208 & ~n36209 ;
  assign n36211 = n36199 & ~n36210 ;
  assign n36212 = n36199 & ~n36211 ;
  assign n36213 = ~n36210 & ~n36211 ;
  assign n36214 = ~n36212 & ~n36213 ;
  assign n36215 = ~n35528 & ~n35533 ;
  assign n36216 = n36214 & n36215 ;
  assign n36217 = ~n36214 & ~n36215 ;
  assign n36218 = ~n36216 & ~n36217 ;
  assign n36219 = x89 & n18025 ;
  assign n36220 = x87 & n18764 ;
  assign n36221 = x88 & n18020 ;
  assign n36222 = ~n36220 & ~n36221 ;
  assign n36223 = ~n36219 & n36222 ;
  assign n36224 = n4488 & n18028 ;
  assign n36225 = n36223 & ~n36224 ;
  assign n36226 = x53 & ~n36225 ;
  assign n36227 = x53 & ~n36226 ;
  assign n36228 = ~n36225 & ~n36226 ;
  assign n36229 = ~n36227 & ~n36228 ;
  assign n36230 = n36218 & ~n36229 ;
  assign n36231 = n36218 & ~n36230 ;
  assign n36232 = ~n36229 & ~n36230 ;
  assign n36233 = ~n36231 & ~n36232 ;
  assign n36234 = ~n35536 & ~n35540 ;
  assign n36235 = n36233 & n36234 ;
  assign n36236 = ~n36233 & ~n36234 ;
  assign n36237 = ~n36235 & ~n36236 ;
  assign n36238 = x92 & n16076 ;
  assign n36239 = x90 & n16756 ;
  assign n36240 = x91 & n16071 ;
  assign n36241 = ~n36239 & ~n36240 ;
  assign n36242 = ~n36238 & n36241 ;
  assign n36243 = n5710 & n16079 ;
  assign n36244 = n36242 & ~n36243 ;
  assign n36245 = x50 & ~n36244 ;
  assign n36246 = x50 & ~n36245 ;
  assign n36247 = ~n36244 & ~n36245 ;
  assign n36248 = ~n36246 & ~n36247 ;
  assign n36249 = ~n36237 & n36248 ;
  assign n36250 = n36237 & ~n36248 ;
  assign n36251 = ~n36249 & ~n36250 ;
  assign n36252 = ~n36153 & n36251 ;
  assign n36253 = ~n36153 & ~n36252 ;
  assign n36254 = n36251 & ~n36252 ;
  assign n36255 = ~n36253 & ~n36254 ;
  assign n36256 = ~n36152 & ~n36255 ;
  assign n36257 = n36152 & ~n36254 ;
  assign n36258 = ~n36253 & n36257 ;
  assign n36259 = ~n36256 & ~n36258 ;
  assign n36260 = ~n35579 & n36259 ;
  assign n36261 = n35579 & ~n36259 ;
  assign n36262 = ~n36260 & ~n36261 ;
  assign n36263 = ~n36141 & n36262 ;
  assign n36264 = n36141 & ~n36262 ;
  assign n36265 = ~n36263 & ~n36264 ;
  assign n36266 = ~n36130 & n36265 ;
  assign n36267 = ~n36130 & ~n36266 ;
  assign n36268 = n36265 & ~n36266 ;
  assign n36269 = ~n36267 & ~n36268 ;
  assign n36270 = ~n36128 & ~n36269 ;
  assign n36271 = n36128 & ~n36268 ;
  assign n36272 = ~n36267 & n36271 ;
  assign n36273 = ~n36270 & ~n36272 ;
  assign n36274 = ~n36117 & n36273 ;
  assign n36275 = ~n36117 & ~n36274 ;
  assign n36276 = n36273 & ~n36274 ;
  assign n36277 = ~n36275 & ~n36276 ;
  assign n36278 = ~n36116 & ~n36277 ;
  assign n36279 = n36116 & ~n36276 ;
  assign n36280 = ~n36275 & n36279 ;
  assign n36281 = ~n36278 & ~n36280 ;
  assign n36282 = ~n36105 & n36281 ;
  assign n36283 = n36105 & ~n36281 ;
  assign n36284 = ~n36282 & ~n36283 ;
  assign n36285 = x107 & n8006 ;
  assign n36286 = x105 & n8474 ;
  assign n36287 = x106 & n8001 ;
  assign n36288 = ~n36286 & ~n36287 ;
  assign n36289 = ~n36285 & n36288 ;
  assign n36290 = n8009 & n12749 ;
  assign n36291 = n36289 & ~n36290 ;
  assign n36292 = x35 & ~n36291 ;
  assign n36293 = x35 & ~n36292 ;
  assign n36294 = ~n36291 & ~n36292 ;
  assign n36295 = ~n36293 & ~n36294 ;
  assign n36296 = n36284 & ~n36295 ;
  assign n36297 = n36284 & ~n36296 ;
  assign n36298 = ~n36295 & ~n36296 ;
  assign n36299 = ~n36297 & ~n36298 ;
  assign n36300 = ~n35646 & ~n35650 ;
  assign n36301 = x110 & n6725 ;
  assign n36302 = x108 & n7129 ;
  assign n36303 = x109 & n6720 ;
  assign n36304 = ~n36302 & ~n36303 ;
  assign n36305 = ~n36301 & n36304 ;
  assign n36306 = ~n6728 & n36305 ;
  assign n36307 = ~n14497 & n36305 ;
  assign n36308 = ~n36306 & ~n36307 ;
  assign n36309 = x32 & ~n36308 ;
  assign n36310 = ~x32 & n36308 ;
  assign n36311 = ~n36309 & ~n36310 ;
  assign n36312 = ~n36300 & ~n36311 ;
  assign n36313 = ~n36300 & ~n36312 ;
  assign n36314 = ~n36311 & ~n36312 ;
  assign n36315 = ~n36313 & ~n36314 ;
  assign n36316 = ~n36299 & ~n36315 ;
  assign n36317 = ~n36299 & ~n36316 ;
  assign n36318 = ~n36315 & ~n36316 ;
  assign n36319 = ~n36317 & ~n36318 ;
  assign n36320 = ~n36103 & ~n36319 ;
  assign n36321 = ~n36103 & ~n36320 ;
  assign n36322 = ~n36319 & ~n36320 ;
  assign n36323 = ~n36321 & ~n36322 ;
  assign n36324 = ~n35437 & ~n35448 ;
  assign n36325 = ~n35671 & ~n36324 ;
  assign n36326 = x116 & n4531 ;
  assign n36327 = x114 & n4847 ;
  assign n36328 = x115 & n4526 ;
  assign n36329 = ~n36327 & ~n36328 ;
  assign n36330 = ~n36326 & n36329 ;
  assign n36331 = ~n4534 & n36330 ;
  assign n36332 = ~n18336 & n36330 ;
  assign n36333 = ~n36331 & ~n36332 ;
  assign n36334 = x26 & ~n36333 ;
  assign n36335 = ~x26 & n36333 ;
  assign n36336 = ~n36334 & ~n36335 ;
  assign n36337 = ~n36325 & ~n36336 ;
  assign n36338 = n36325 & n36336 ;
  assign n36339 = ~n36337 & ~n36338 ;
  assign n36340 = ~n36323 & n36339 ;
  assign n36341 = ~n36323 & ~n36340 ;
  assign n36342 = n36339 & ~n36340 ;
  assign n36343 = ~n36341 & ~n36342 ;
  assign n36344 = ~n36087 & ~n36343 ;
  assign n36345 = ~n36087 & ~n36344 ;
  assign n36346 = ~n36343 & ~n36344 ;
  assign n36347 = ~n36345 & ~n36346 ;
  assign n36348 = ~n35418 & ~n35679 ;
  assign n36349 = x122 & n2751 ;
  assign n36350 = x120 & n3020 ;
  assign n36351 = x121 & n2746 ;
  assign n36352 = ~n36350 & ~n36351 ;
  assign n36353 = ~n36349 & n36352 ;
  assign n36354 = ~n2754 & n36353 ;
  assign n36355 = ~n22622 & n36353 ;
  assign n36356 = ~n36354 & ~n36355 ;
  assign n36357 = x20 & ~n36356 ;
  assign n36358 = ~x20 & n36356 ;
  assign n36359 = ~n36357 & ~n36358 ;
  assign n36360 = ~n36348 & ~n36359 ;
  assign n36361 = ~n36348 & ~n36360 ;
  assign n36362 = ~n36359 & ~n36360 ;
  assign n36363 = ~n36361 & ~n36362 ;
  assign n36364 = ~n36347 & ~n36363 ;
  assign n36365 = ~n36347 & ~n36364 ;
  assign n36366 = ~n36363 & ~n36364 ;
  assign n36367 = ~n36365 & ~n36366 ;
  assign n36368 = ~n36071 & ~n36367 ;
  assign n36369 = ~n36071 & ~n36368 ;
  assign n36370 = ~n36367 & ~n36368 ;
  assign n36371 = ~n36369 & ~n36370 ;
  assign n36372 = ~n35376 & ~n35387 ;
  assign n36373 = ~n35687 & ~n36372 ;
  assign n36374 = x126 & n1646 ;
  assign n36375 = x127 & n1429 ;
  assign n36376 = ~n36374 & ~n36375 ;
  assign n36377 = ~n1437 & n36376 ;
  assign n36378 = n26965 & n36376 ;
  assign n36379 = ~n36377 & ~n36378 ;
  assign n36380 = x14 & ~n36379 ;
  assign n36381 = ~x14 & n36379 ;
  assign n36382 = ~n36380 & ~n36381 ;
  assign n36383 = ~n36373 & ~n36382 ;
  assign n36384 = ~n36373 & ~n36383 ;
  assign n36385 = ~n36382 & ~n36383 ;
  assign n36386 = ~n36384 & ~n36385 ;
  assign n36387 = ~n36371 & ~n36386 ;
  assign n36388 = n36371 & ~n36385 ;
  assign n36389 = ~n36384 & n36388 ;
  assign n36390 = ~n36387 & ~n36389 ;
  assign n36391 = ~n36055 & n36390 ;
  assign n36392 = ~n36055 & ~n36391 ;
  assign n36393 = n36390 & ~n36391 ;
  assign n36394 = ~n36392 & ~n36393 ;
  assign n36395 = ~n36053 & ~n36394 ;
  assign n36396 = n36053 & ~n36393 ;
  assign n36397 = ~n36392 & n36396 ;
  assign n36398 = ~n36395 & ~n36397 ;
  assign n36746 = n36398 & x204 ;
  assign n36399 = ~n36041 & ~n36045 ;
  assign n36400 = ~n35721 & ~n36037 ;
  assign n36401 = ~n35718 & ~n36400 ;
  assign n36402 = ~x125 & n2093 ;
  assign n36403 = ~x123 & n2275 ;
  assign n36404 = ~x124 & n2088 ;
  assign n36405 = ~n36403 & ~n36404 ;
  assign n36406 = ~n36402 & n36405 ;
  assign n36407 = n2096 & n25330 ;
  assign n36408 = n36406 & ~n36407 ;
  assign n36409 = ~x17 & ~n36408 ;
  assign n36410 = ~x17 & ~n36409 ;
  assign n36411 = ~n36408 & ~n36409 ;
  assign n36412 = ~n36410 & ~n36411 ;
  assign n36413 = ~n35750 & ~n36030 ;
  assign n36414 = ~n36412 & ~n36413 ;
  assign n36415 = ~n36412 & ~n36414 ;
  assign n36416 = ~n36413 & ~n36414 ;
  assign n36417 = ~n36415 & ~n36416 ;
  assign n36418 = ~x119 & n3589 ;
  assign n36419 = ~x117 & n3878 ;
  assign n36420 = ~x118 & n3584 ;
  assign n36421 = ~n36419 & ~n36420 ;
  assign n36422 = ~n36418 & n36421 ;
  assign n36423 = n3592 & n20778 ;
  assign n36424 = n36422 & ~n36423 ;
  assign n36425 = ~x23 & ~n36424 ;
  assign n36426 = ~x23 & ~n36425 ;
  assign n36427 = ~n36424 & ~n36425 ;
  assign n36428 = ~n36426 & ~n36427 ;
  assign n36429 = ~n35781 & ~n36022 ;
  assign n36430 = ~n36428 & ~n36429 ;
  assign n36431 = ~n36428 & ~n36430 ;
  assign n36432 = ~n36429 & ~n36430 ;
  assign n36433 = ~n36431 & ~n36432 ;
  assign n36434 = ~x113 & n5560 ;
  assign n36435 = ~x111 & n5943 ;
  assign n36436 = ~x112 & n5555 ;
  assign n36437 = ~n36435 & ~n36436 ;
  assign n36438 = ~n36434 & n36437 ;
  assign n36439 = n5563 & n16684 ;
  assign n36440 = n36438 & ~n36439 ;
  assign n36441 = ~x29 & ~n36440 ;
  assign n36442 = ~x29 & ~n36441 ;
  assign n36443 = ~n36440 & ~n36441 ;
  assign n36444 = ~n36442 & ~n36443 ;
  assign n36445 = ~n36010 & ~n36014 ;
  assign n36446 = ~n36444 & ~n36445 ;
  assign n36447 = ~n36444 & ~n36446 ;
  assign n36448 = ~n36445 & ~n36446 ;
  assign n36449 = ~n36447 & ~n36448 ;
  assign n36450 = ~n35799 & ~n35977 ;
  assign n36451 = ~n35974 & ~n36450 ;
  assign n36452 = ~x104 & n9433 ;
  assign n36453 = ~x102 & n9915 ;
  assign n36454 = ~x103 & n9428 ;
  assign n36455 = ~n36453 & ~n36454 ;
  assign n36456 = ~n36452 & n36455 ;
  assign n36457 = n9436 & n11380 ;
  assign n36458 = n36456 & ~n36457 ;
  assign n36459 = ~x38 & ~n36458 ;
  assign n36460 = ~x38 & ~n36459 ;
  assign n36461 = ~n36458 & ~n36459 ;
  assign n36462 = ~n36460 & ~n36461 ;
  assign n36463 = ~n35957 & ~n35961 ;
  assign n36464 = ~x101 & n10905 ;
  assign n36465 = ~x99 & n11466 ;
  assign n36466 = ~x100 & n10900 ;
  assign n36467 = ~n36465 & ~n36466 ;
  assign n36468 = ~n36464 & n36467 ;
  assign n36469 = n9844 & n10908 ;
  assign n36470 = n36468 & ~n36469 ;
  assign n36471 = ~x41 & ~n36470 ;
  assign n36472 = ~x41 & ~n36471 ;
  assign n36473 = ~n36470 & ~n36471 ;
  assign n36474 = ~n36472 & ~n36473 ;
  assign n36475 = ~n35801 & ~n35942 ;
  assign n36476 = ~n35939 & ~n36475 ;
  assign n36477 = ~x98 & n12506 ;
  assign n36478 = ~x96 & n13131 ;
  assign n36479 = ~x97 & n12501 ;
  assign n36480 = ~n36478 & ~n36479 ;
  assign n36481 = ~n36477 & n36480 ;
  assign n36482 = n8426 & n12509 ;
  assign n36483 = n36481 & ~n36482 ;
  assign n36484 = ~x44 & ~n36483 ;
  assign n36485 = ~x44 & ~n36484 ;
  assign n36486 = ~n36483 & ~n36484 ;
  assign n36487 = ~n36485 & ~n36486 ;
  assign n36488 = ~x95 & n14233 ;
  assign n36489 = ~x93 & n14876 ;
  assign n36490 = ~x94 & n14228 ;
  assign n36491 = ~n36489 & ~n36490 ;
  assign n36492 = ~n36488 & n36491 ;
  assign n36493 = n7100 & n14236 ;
  assign n36494 = n36492 & ~n36493 ;
  assign n36495 = ~x47 & ~n36494 ;
  assign n36496 = ~x47 & ~n36495 ;
  assign n36497 = ~n36494 & ~n36495 ;
  assign n36498 = ~n36496 & ~n36497 ;
  assign n36499 = ~n35901 & ~n35907 ;
  assign n36500 = ~x76 & n27427 ;
  assign n36501 = ~x77 & ~n26217 ;
  assign n36502 = ~n36500 & ~n36501 ;
  assign n36503 = x11 & ~n34412 ;
  assign n36504 = ~n35833 & ~n36503 ;
  assign n36505 = n36502 & ~n36504 ;
  assign n36506 = n36502 & ~n36505 ;
  assign n36507 = ~n36504 & ~n36505 ;
  assign n36508 = ~n36506 & ~n36507 ;
  assign n36509 = ~x80 & n24612 ;
  assign n36510 = ~x78 & n25390 ;
  assign n36511 = ~x79 & n24607 ;
  assign n36512 = ~n36510 & ~n36511 ;
  assign n36513 = ~n36509 & n36512 ;
  assign n36514 = n2145 & n24615 ;
  assign n36515 = n36513 & ~n36514 ;
  assign n36516 = ~x62 & ~n36515 ;
  assign n36517 = ~x62 & ~n36516 ;
  assign n36518 = ~n36515 & ~n36516 ;
  assign n36519 = ~n36517 & ~n36518 ;
  assign n36520 = ~n36508 & n36519 ;
  assign n36521 = n36508 & ~n36519 ;
  assign n36522 = ~n36520 & ~n36521 ;
  assign n36523 = ~n35836 & ~n35840 ;
  assign n36524 = n36522 & n36523 ;
  assign n36525 = ~n36522 & ~n36523 ;
  assign n36526 = ~n36524 & ~n36525 ;
  assign n36527 = ~x83 & n22325 ;
  assign n36528 = ~x81 & n23066 ;
  assign n36529 = ~x82 & n22320 ;
  assign n36530 = ~n36528 & ~n36529 ;
  assign n36531 = ~n36527 & n36530 ;
  assign n36532 = n2972 & n22328 ;
  assign n36533 = n36531 & ~n36532 ;
  assign n36534 = ~x59 & ~n36533 ;
  assign n36535 = ~x59 & ~n36534 ;
  assign n36536 = ~n36533 & ~n36534 ;
  assign n36537 = ~n36535 & ~n36536 ;
  assign n36538 = n36526 & ~n36537 ;
  assign n36539 = n36526 & ~n36538 ;
  assign n36540 = ~n36537 & ~n36538 ;
  assign n36541 = ~n36539 & ~n36540 ;
  assign n36542 = ~n35855 & ~n35861 ;
  assign n36543 = n36541 & n36542 ;
  assign n36544 = ~n36541 & ~n36542 ;
  assign n36545 = ~n36543 & ~n36544 ;
  assign n36546 = ~x86 & n20143 ;
  assign n36547 = ~x84 & n20854 ;
  assign n36548 = ~x85 & n20138 ;
  assign n36549 = ~n36547 & ~n36548 ;
  assign n36550 = ~n36546 & n36549 ;
  assign n36551 = n3832 & n20146 ;
  assign n36552 = n36550 & ~n36551 ;
  assign n36553 = ~x56 & ~n36552 ;
  assign n36554 = ~x56 & ~n36553 ;
  assign n36555 = ~n36552 & ~n36553 ;
  assign n36556 = ~n36554 & ~n36555 ;
  assign n36557 = n36545 & ~n36556 ;
  assign n36558 = n36545 & ~n36557 ;
  assign n36559 = ~n36556 & ~n36557 ;
  assign n36560 = ~n36558 & ~n36559 ;
  assign n36561 = ~n35874 & ~n35879 ;
  assign n36562 = n36560 & n36561 ;
  assign n36563 = ~n36560 & ~n36561 ;
  assign n36564 = ~n36562 & ~n36563 ;
  assign n36565 = ~x89 & n18025 ;
  assign n36566 = ~x87 & n18764 ;
  assign n36567 = ~x88 & n18020 ;
  assign n36568 = ~n36566 & ~n36567 ;
  assign n36569 = ~n36565 & n36568 ;
  assign n36570 = n4664 & n18028 ;
  assign n36571 = n36569 & ~n36570 ;
  assign n36572 = ~x53 & ~n36571 ;
  assign n36573 = ~x53 & ~n36572 ;
  assign n36574 = ~n36571 & ~n36572 ;
  assign n36575 = ~n36573 & ~n36574 ;
  assign n36576 = n36564 & ~n36575 ;
  assign n36577 = n36564 & ~n36576 ;
  assign n36578 = ~n36575 & ~n36576 ;
  assign n36579 = ~n36577 & ~n36578 ;
  assign n36580 = ~n35882 & ~n35886 ;
  assign n36581 = n36579 & n36580 ;
  assign n36582 = ~n36579 & ~n36580 ;
  assign n36583 = ~n36581 & ~n36582 ;
  assign n36584 = ~x92 & n16076 ;
  assign n36585 = ~x90 & n16756 ;
  assign n36586 = ~x91 & n16071 ;
  assign n36587 = ~n36585 & ~n36586 ;
  assign n36588 = ~n36584 & n36587 ;
  assign n36589 = n5896 & n16079 ;
  assign n36590 = n36588 & ~n36589 ;
  assign n36591 = ~x50 & ~n36590 ;
  assign n36592 = ~x50 & ~n36591 ;
  assign n36593 = ~n36590 & ~n36591 ;
  assign n36594 = ~n36592 & ~n36593 ;
  assign n36595 = ~n36583 & n36594 ;
  assign n36596 = n36583 & ~n36594 ;
  assign n36597 = ~n36595 & ~n36596 ;
  assign n36598 = ~n36499 & n36597 ;
  assign n36599 = ~n36499 & ~n36598 ;
  assign n36600 = n36597 & ~n36598 ;
  assign n36601 = ~n36599 & ~n36600 ;
  assign n36602 = ~n36498 & ~n36601 ;
  assign n36603 = n36498 & ~n36600 ;
  assign n36604 = ~n36599 & n36603 ;
  assign n36605 = ~n36602 & ~n36604 ;
  assign n36606 = ~n35925 & n36605 ;
  assign n36607 = n35925 & ~n36605 ;
  assign n36608 = ~n36606 & ~n36607 ;
  assign n36609 = ~n36487 & n36608 ;
  assign n36610 = n36487 & ~n36608 ;
  assign n36611 = ~n36609 & ~n36610 ;
  assign n36612 = ~n36476 & n36611 ;
  assign n36613 = ~n36476 & ~n36612 ;
  assign n36614 = n36611 & ~n36612 ;
  assign n36615 = ~n36613 & ~n36614 ;
  assign n36616 = ~n36474 & ~n36615 ;
  assign n36617 = n36474 & ~n36614 ;
  assign n36618 = ~n36613 & n36617 ;
  assign n36619 = ~n36616 & ~n36618 ;
  assign n36620 = ~n36463 & n36619 ;
  assign n36621 = ~n36463 & ~n36620 ;
  assign n36622 = n36619 & ~n36620 ;
  assign n36623 = ~n36621 & ~n36622 ;
  assign n36624 = ~n36462 & ~n36623 ;
  assign n36625 = n36462 & ~n36622 ;
  assign n36626 = ~n36621 & n36625 ;
  assign n36627 = ~n36624 & ~n36626 ;
  assign n36628 = ~n36451 & n36627 ;
  assign n36629 = n36451 & ~n36627 ;
  assign n36630 = ~n36628 & ~n36629 ;
  assign n36631 = ~x107 & n8006 ;
  assign n36632 = ~x105 & n8474 ;
  assign n36633 = ~x106 & n8001 ;
  assign n36634 = ~n36632 & ~n36633 ;
  assign n36635 = ~n36631 & n36634 ;
  assign n36636 = n8009 & n13034 ;
  assign n36637 = n36635 & ~n36636 ;
  assign n36638 = ~x35 & ~n36637 ;
  assign n36639 = ~x35 & ~n36638 ;
  assign n36640 = ~n36637 & ~n36638 ;
  assign n36641 = ~n36639 & ~n36640 ;
  assign n36642 = n36630 & ~n36641 ;
  assign n36643 = n36630 & ~n36642 ;
  assign n36644 = ~n36641 & ~n36642 ;
  assign n36645 = ~n36643 & ~n36644 ;
  assign n36646 = ~n35992 & ~n35996 ;
  assign n36647 = ~x110 & n6725 ;
  assign n36648 = ~x108 & n7129 ;
  assign n36649 = ~x109 & n6720 ;
  assign n36650 = ~n36648 & ~n36649 ;
  assign n36651 = ~n36647 & n36650 ;
  assign n36652 = ~n6728 & n36651 ;
  assign n36653 = ~n14802 & n36651 ;
  assign n36654 = ~n36652 & ~n36653 ;
  assign n36655 = ~x32 & ~n36654 ;
  assign n36656 = x32 & n36654 ;
  assign n36657 = ~n36655 & ~n36656 ;
  assign n36658 = ~n36646 & ~n36657 ;
  assign n36659 = ~n36646 & ~n36658 ;
  assign n36660 = ~n36657 & ~n36658 ;
  assign n36661 = ~n36659 & ~n36660 ;
  assign n36662 = ~n36645 & ~n36661 ;
  assign n36663 = ~n36645 & ~n36662 ;
  assign n36664 = ~n36661 & ~n36662 ;
  assign n36665 = ~n36663 & ~n36664 ;
  assign n36666 = ~n36449 & ~n36665 ;
  assign n36667 = ~n36449 & ~n36666 ;
  assign n36668 = ~n36665 & ~n36666 ;
  assign n36669 = ~n36667 & ~n36668 ;
  assign n36670 = ~n35783 & ~n35794 ;
  assign n36671 = ~n36017 & ~n36670 ;
  assign n36672 = ~x116 & n4531 ;
  assign n36673 = ~x114 & n4847 ;
  assign n36674 = ~x115 & n4526 ;
  assign n36675 = ~n36673 & ~n36674 ;
  assign n36676 = ~n36672 & n36675 ;
  assign n36677 = ~n4534 & n36676 ;
  assign n36678 = ~n18678 & n36676 ;
  assign n36679 = ~n36677 & ~n36678 ;
  assign n36680 = ~x26 & ~n36679 ;
  assign n36681 = x26 & n36679 ;
  assign n36682 = ~n36680 & ~n36681 ;
  assign n36683 = ~n36671 & ~n36682 ;
  assign n36684 = n36671 & n36682 ;
  assign n36685 = ~n36683 & ~n36684 ;
  assign n36686 = ~n36669 & n36685 ;
  assign n36687 = ~n36669 & ~n36686 ;
  assign n36688 = n36685 & ~n36686 ;
  assign n36689 = ~n36687 & ~n36688 ;
  assign n36690 = ~n36433 & ~n36689 ;
  assign n36691 = ~n36433 & ~n36690 ;
  assign n36692 = ~n36689 & ~n36690 ;
  assign n36693 = ~n36691 & ~n36692 ;
  assign n36694 = ~n35764 & ~n36025 ;
  assign n36695 = ~x122 & n2751 ;
  assign n36696 = ~x120 & n3020 ;
  assign n36697 = ~x121 & n2746 ;
  assign n36698 = ~n36696 & ~n36697 ;
  assign n36699 = ~n36695 & n36698 ;
  assign n36700 = ~n2754 & n36699 ;
  assign n36701 = ~n22998 & n36699 ;
  assign n36702 = ~n36700 & ~n36701 ;
  assign n36703 = ~x20 & ~n36702 ;
  assign n36704 = x20 & n36702 ;
  assign n36705 = ~n36703 & ~n36704 ;
  assign n36706 = ~n36694 & ~n36705 ;
  assign n36707 = ~n36694 & ~n36706 ;
  assign n36708 = ~n36705 & ~n36706 ;
  assign n36709 = ~n36707 & ~n36708 ;
  assign n36710 = ~n36693 & ~n36709 ;
  assign n36711 = ~n36693 & ~n36710 ;
  assign n36712 = ~n36709 & ~n36710 ;
  assign n36713 = ~n36711 & ~n36712 ;
  assign n36714 = ~n36417 & ~n36713 ;
  assign n36715 = ~n36417 & ~n36714 ;
  assign n36716 = ~n36713 & ~n36714 ;
  assign n36717 = ~n36715 & ~n36716 ;
  assign n36718 = ~n35722 & ~n35733 ;
  assign n36719 = ~n36033 & ~n36718 ;
  assign n36720 = ~x126 & n1646 ;
  assign n36721 = ~x127 & n1429 ;
  assign n36722 = ~n36720 & ~n36721 ;
  assign n36723 = ~n1437 & n36722 ;
  assign n36724 = n27368 & n36722 ;
  assign n36725 = ~n36723 & ~n36724 ;
  assign n36726 = ~x14 & ~n36725 ;
  assign n36727 = x14 & n36725 ;
  assign n36728 = ~n36726 & ~n36727 ;
  assign n36729 = ~n36719 & ~n36728 ;
  assign n36730 = ~n36719 & ~n36729 ;
  assign n36731 = ~n36728 & ~n36729 ;
  assign n36732 = ~n36730 & ~n36731 ;
  assign n36733 = ~n36717 & ~n36732 ;
  assign n36734 = n36717 & ~n36731 ;
  assign n36735 = ~n36730 & n36734 ;
  assign n36736 = ~n36733 & ~n36735 ;
  assign n36737 = ~n36401 & n36736 ;
  assign n36738 = ~n36401 & ~n36737 ;
  assign n36739 = n36736 & ~n36737 ;
  assign n36740 = ~n36738 & ~n36739 ;
  assign n36741 = ~n36399 & ~n36740 ;
  assign n36742 = n36399 & ~n36739 ;
  assign n36743 = ~n36738 & n36742 ;
  assign n36744 = ~n36741 & ~n36743 ;
  assign n36747 = ~n36744 & ~x204 ;
  assign n36748 = ~n36746 & ~n36747 ;
  assign n36749 = ~n36391 & ~n36395 ;
  assign n36750 = ~n36383 & ~n36387 ;
  assign n36751 = ~n36068 & ~n36368 ;
  assign n36752 = x127 & n1646 ;
  assign n36753 = n1437 & n26962 ;
  assign n36754 = ~n36752 & ~n36753 ;
  assign n36755 = x14 & ~n36754 ;
  assign n36756 = x14 & ~n36755 ;
  assign n36757 = ~n36754 & ~n36755 ;
  assign n36758 = ~n36756 & ~n36757 ;
  assign n36759 = ~n36751 & ~n36758 ;
  assign n36760 = ~n36751 & ~n36759 ;
  assign n36761 = ~n36758 & ~n36759 ;
  assign n36762 = ~n36760 & ~n36761 ;
  assign n36763 = x123 & n2751 ;
  assign n36764 = x121 & n3020 ;
  assign n36765 = x122 & n2746 ;
  assign n36766 = ~n36764 & ~n36765 ;
  assign n36767 = ~n36763 & n36766 ;
  assign n36768 = n2754 & n23382 ;
  assign n36769 = n36767 & ~n36768 ;
  assign n36770 = x20 & ~n36769 ;
  assign n36771 = x20 & ~n36770 ;
  assign n36772 = ~n36769 & ~n36770 ;
  assign n36773 = ~n36771 & ~n36772 ;
  assign n36774 = ~n36084 & ~n36344 ;
  assign n36775 = n36773 & n36774 ;
  assign n36776 = ~n36773 & ~n36774 ;
  assign n36777 = ~n36775 & ~n36776 ;
  assign n36778 = x120 & n3589 ;
  assign n36779 = x118 & n3878 ;
  assign n36780 = x119 & n3584 ;
  assign n36781 = ~n36779 & ~n36780 ;
  assign n36782 = ~n36778 & n36781 ;
  assign n36783 = n3592 & n21143 ;
  assign n36784 = n36782 & ~n36783 ;
  assign n36785 = x23 & ~n36784 ;
  assign n36786 = x23 & ~n36785 ;
  assign n36787 = ~n36784 & ~n36785 ;
  assign n36788 = ~n36786 & ~n36787 ;
  assign n36789 = ~n36337 & ~n36340 ;
  assign n36790 = n36788 & n36789 ;
  assign n36791 = ~n36788 & ~n36789 ;
  assign n36792 = ~n36790 & ~n36791 ;
  assign n36793 = x117 & n4531 ;
  assign n36794 = x115 & n4847 ;
  assign n36795 = x116 & n4526 ;
  assign n36796 = ~n36794 & ~n36795 ;
  assign n36797 = ~n36793 & n36796 ;
  assign n36798 = n4534 & n19026 ;
  assign n36799 = n36797 & ~n36798 ;
  assign n36800 = x26 & ~n36799 ;
  assign n36801 = x26 & ~n36800 ;
  assign n36802 = ~n36799 & ~n36800 ;
  assign n36803 = ~n36801 & ~n36802 ;
  assign n36804 = ~n36100 & ~n36320 ;
  assign n36805 = n36803 & n36804 ;
  assign n36806 = ~n36803 & ~n36804 ;
  assign n36807 = ~n36805 & ~n36806 ;
  assign n36808 = ~n36282 & ~n36296 ;
  assign n36809 = x111 & n6725 ;
  assign n36810 = x109 & n7129 ;
  assign n36811 = x110 & n6720 ;
  assign n36812 = ~n36810 & ~n36811 ;
  assign n36813 = ~n36809 & n36812 ;
  assign n36814 = ~n6728 & n36813 ;
  assign n36815 = ~n15111 & n36813 ;
  assign n36816 = ~n36814 & ~n36815 ;
  assign n36817 = x32 & ~n36816 ;
  assign n36818 = ~x32 & n36816 ;
  assign n36819 = ~n36817 & ~n36818 ;
  assign n36820 = ~n36808 & ~n36819 ;
  assign n36821 = n36808 & n36819 ;
  assign n36822 = ~n36820 & ~n36821 ;
  assign n36823 = x108 & n8006 ;
  assign n36824 = x106 & n8474 ;
  assign n36825 = x107 & n8001 ;
  assign n36826 = ~n36824 & ~n36825 ;
  assign n36827 = ~n36823 & n36826 ;
  assign n36828 = n8009 & n13323 ;
  assign n36829 = n36827 & ~n36828 ;
  assign n36830 = x35 & ~n36829 ;
  assign n36831 = x35 & ~n36830 ;
  assign n36832 = ~n36829 & ~n36830 ;
  assign n36833 = ~n36831 & ~n36832 ;
  assign n36834 = ~n36274 & ~n36278 ;
  assign n36835 = x105 & n9433 ;
  assign n36836 = x103 & n9915 ;
  assign n36837 = x104 & n9428 ;
  assign n36838 = ~n36836 & ~n36837 ;
  assign n36839 = ~n36835 & n36838 ;
  assign n36840 = n9436 & n11648 ;
  assign n36841 = n36839 & ~n36840 ;
  assign n36842 = x38 & ~n36841 ;
  assign n36843 = x38 & ~n36842 ;
  assign n36844 = ~n36841 & ~n36842 ;
  assign n36845 = ~n36843 & ~n36844 ;
  assign n36846 = ~n36266 & ~n36270 ;
  assign n36847 = ~n36252 & ~n36256 ;
  assign n36848 = ~n36217 & ~n36230 ;
  assign n36849 = x90 & n18025 ;
  assign n36850 = x88 & n18764 ;
  assign n36851 = x89 & n18020 ;
  assign n36852 = ~n36850 & ~n36851 ;
  assign n36853 = ~n36849 & n36852 ;
  assign n36854 = n4986 & n18028 ;
  assign n36855 = n36853 & ~n36854 ;
  assign n36856 = x53 & ~n36855 ;
  assign n36857 = x53 & ~n36856 ;
  assign n36858 = ~n36855 & ~n36856 ;
  assign n36859 = ~n36857 & ~n36858 ;
  assign n36860 = ~n36198 & ~n36211 ;
  assign n36861 = ~n36162 & ~n36173 ;
  assign n36862 = ~n36159 & ~n36861 ;
  assign n36863 = x77 & n27024 ;
  assign n36864 = x78 & ~n26217 ;
  assign n36865 = ~n36863 & ~n36864 ;
  assign n36866 = n36156 & ~n36865 ;
  assign n36867 = ~n36156 & n36865 ;
  assign n36868 = ~n36866 & ~n36867 ;
  assign n36869 = x81 & n24612 ;
  assign n36870 = x79 & n25390 ;
  assign n36871 = x80 & n24607 ;
  assign n36872 = ~n36870 & ~n36871 ;
  assign n36873 = ~n36869 & n36872 ;
  assign n36874 = ~n24615 & n36873 ;
  assign n36875 = ~n2348 & n36873 ;
  assign n36876 = ~n36874 & ~n36875 ;
  assign n36877 = x62 & ~n36876 ;
  assign n36878 = ~x62 & n36876 ;
  assign n36879 = ~n36877 & ~n36878 ;
  assign n36880 = n36868 & ~n36879 ;
  assign n36881 = ~n36868 & n36879 ;
  assign n36882 = ~n36880 & ~n36881 ;
  assign n36883 = ~n36862 & n36882 ;
  assign n36884 = n36862 & ~n36882 ;
  assign n36885 = ~n36883 & ~n36884 ;
  assign n36886 = x84 & n22325 ;
  assign n36887 = x82 & n23066 ;
  assign n36888 = x83 & n22320 ;
  assign n36889 = ~n36887 & ~n36888 ;
  assign n36890 = ~n36886 & n36889 ;
  assign n36891 = n3114 & n22328 ;
  assign n36892 = n36890 & ~n36891 ;
  assign n36893 = x59 & ~n36892 ;
  assign n36894 = x59 & ~n36893 ;
  assign n36895 = ~n36892 & ~n36893 ;
  assign n36896 = ~n36894 & ~n36895 ;
  assign n36897 = n36885 & ~n36896 ;
  assign n36898 = n36885 & ~n36897 ;
  assign n36899 = ~n36896 & ~n36897 ;
  assign n36900 = ~n36898 & ~n36899 ;
  assign n36901 = ~n36179 & ~n36192 ;
  assign n36902 = n36900 & n36901 ;
  assign n36903 = ~n36900 & ~n36901 ;
  assign n36904 = ~n36902 & ~n36903 ;
  assign n36905 = x87 & n20143 ;
  assign n36906 = x85 & n20854 ;
  assign n36907 = x86 & n20138 ;
  assign n36908 = ~n36906 & ~n36907 ;
  assign n36909 = ~n36905 & n36908 ;
  assign n36910 = n3991 & n20146 ;
  assign n36911 = n36909 & ~n36910 ;
  assign n36912 = x56 & ~n36911 ;
  assign n36913 = x56 & ~n36912 ;
  assign n36914 = ~n36911 & ~n36912 ;
  assign n36915 = ~n36913 & ~n36914 ;
  assign n36916 = ~n36904 & n36915 ;
  assign n36917 = n36904 & ~n36915 ;
  assign n36918 = ~n36916 & ~n36917 ;
  assign n36919 = ~n36860 & n36918 ;
  assign n36920 = n36860 & ~n36918 ;
  assign n36921 = ~n36919 & ~n36920 ;
  assign n36922 = ~n36859 & n36921 ;
  assign n36923 = n36859 & ~n36921 ;
  assign n36924 = ~n36922 & ~n36923 ;
  assign n36925 = ~n36848 & n36924 ;
  assign n36926 = n36848 & ~n36924 ;
  assign n36927 = ~n36925 & ~n36926 ;
  assign n36928 = x93 & n16076 ;
  assign n36929 = x91 & n16756 ;
  assign n36930 = x92 & n16071 ;
  assign n36931 = ~n36929 & ~n36930 ;
  assign n36932 = ~n36928 & n36931 ;
  assign n36933 = n6094 & n16079 ;
  assign n36934 = n36932 & ~n36933 ;
  assign n36935 = x50 & ~n36934 ;
  assign n36936 = x50 & ~n36935 ;
  assign n36937 = ~n36934 & ~n36935 ;
  assign n36938 = ~n36936 & ~n36937 ;
  assign n36939 = n36927 & ~n36938 ;
  assign n36940 = n36927 & ~n36939 ;
  assign n36941 = ~n36938 & ~n36939 ;
  assign n36942 = ~n36940 & ~n36941 ;
  assign n36943 = ~n36236 & ~n36250 ;
  assign n36944 = ~n36942 & ~n36943 ;
  assign n36945 = ~n36942 & ~n36944 ;
  assign n36946 = ~n36943 & ~n36944 ;
  assign n36947 = ~n36945 & ~n36946 ;
  assign n36948 = x96 & n14233 ;
  assign n36949 = x94 & n14876 ;
  assign n36950 = x95 & n14228 ;
  assign n36951 = ~n36949 & ~n36950 ;
  assign n36952 = ~n36948 & n36951 ;
  assign n36953 = n7321 & n14236 ;
  assign n36954 = n36952 & ~n36953 ;
  assign n36955 = x47 & ~n36954 ;
  assign n36956 = x47 & ~n36955 ;
  assign n36957 = ~n36954 & ~n36955 ;
  assign n36958 = ~n36956 & ~n36957 ;
  assign n36959 = ~n36947 & n36958 ;
  assign n36960 = n36947 & ~n36958 ;
  assign n36961 = ~n36959 & ~n36960 ;
  assign n36962 = n36847 & n36961 ;
  assign n36963 = ~n36847 & ~n36961 ;
  assign n36964 = ~n36962 & ~n36963 ;
  assign n36965 = x99 & n12506 ;
  assign n36966 = x97 & n13131 ;
  assign n36967 = x98 & n12501 ;
  assign n36968 = ~n36966 & ~n36967 ;
  assign n36969 = ~n36965 & n36968 ;
  assign n36970 = n8660 & n12509 ;
  assign n36971 = n36969 & ~n36970 ;
  assign n36972 = x44 & ~n36971 ;
  assign n36973 = x44 & ~n36972 ;
  assign n36974 = ~n36971 & ~n36972 ;
  assign n36975 = ~n36973 & ~n36974 ;
  assign n36976 = n36964 & ~n36975 ;
  assign n36977 = n36964 & ~n36976 ;
  assign n36978 = ~n36975 & ~n36976 ;
  assign n36979 = ~n36977 & ~n36978 ;
  assign n36980 = ~n36260 & ~n36263 ;
  assign n36981 = n36979 & n36980 ;
  assign n36982 = ~n36979 & ~n36980 ;
  assign n36983 = ~n36981 & ~n36982 ;
  assign n36984 = x102 & n10905 ;
  assign n36985 = x100 & n11466 ;
  assign n36986 = x101 & n10900 ;
  assign n36987 = ~n36985 & ~n36986 ;
  assign n36988 = ~n36984 & n36987 ;
  assign n36989 = n10092 & n10908 ;
  assign n36990 = n36988 & ~n36989 ;
  assign n36991 = x41 & ~n36990 ;
  assign n36992 = x41 & ~n36991 ;
  assign n36993 = ~n36990 & ~n36991 ;
  assign n36994 = ~n36992 & ~n36993 ;
  assign n36995 = ~n36983 & n36994 ;
  assign n36996 = n36983 & ~n36994 ;
  assign n36997 = ~n36995 & ~n36996 ;
  assign n36998 = ~n36846 & n36997 ;
  assign n36999 = n36846 & ~n36997 ;
  assign n37000 = ~n36998 & ~n36999 ;
  assign n37001 = ~n36845 & n37000 ;
  assign n37002 = n36845 & ~n37000 ;
  assign n37003 = ~n37001 & ~n37002 ;
  assign n37004 = ~n36834 & n37003 ;
  assign n37005 = n36834 & ~n37003 ;
  assign n37006 = ~n37004 & ~n37005 ;
  assign n37007 = ~n36833 & n37006 ;
  assign n37008 = ~n36833 & ~n37007 ;
  assign n37009 = n37006 & ~n37007 ;
  assign n37010 = ~n37008 & ~n37009 ;
  assign n37011 = n36822 & ~n37010 ;
  assign n37012 = n36822 & ~n37011 ;
  assign n37013 = ~n37010 & ~n37011 ;
  assign n37014 = ~n37012 & ~n37013 ;
  assign n37015 = ~n36312 & ~n36316 ;
  assign n37016 = x114 & n5560 ;
  assign n37017 = x112 & n5943 ;
  assign n37018 = x113 & n5555 ;
  assign n37019 = ~n37017 & ~n37018 ;
  assign n37020 = ~n37016 & n37019 ;
  assign n37021 = ~n5563 & n37020 ;
  assign n37022 = ~n17012 & n37020 ;
  assign n37023 = ~n37021 & ~n37022 ;
  assign n37024 = x29 & ~n37023 ;
  assign n37025 = ~x29 & n37023 ;
  assign n37026 = ~n37024 & ~n37025 ;
  assign n37027 = ~n37015 & ~n37026 ;
  assign n37028 = n37015 & n37026 ;
  assign n37029 = ~n37027 & ~n37028 ;
  assign n37030 = ~n37014 & n37029 ;
  assign n37031 = ~n37014 & ~n37030 ;
  assign n37032 = n37029 & ~n37030 ;
  assign n37033 = ~n37031 & ~n37032 ;
  assign n37034 = n36807 & ~n37033 ;
  assign n37035 = n36807 & ~n37034 ;
  assign n37036 = ~n37033 & ~n37034 ;
  assign n37037 = ~n37035 & ~n37036 ;
  assign n37038 = n36792 & ~n37037 ;
  assign n37039 = ~n36792 & n37037 ;
  assign n37040 = n36777 & ~n37039 ;
  assign n37041 = ~n37038 & n37040 ;
  assign n37042 = n36777 & ~n37041 ;
  assign n37043 = ~n37039 & ~n37041 ;
  assign n37044 = ~n37038 & n37043 ;
  assign n37045 = ~n37042 & ~n37044 ;
  assign n37046 = ~n36360 & ~n36364 ;
  assign n37047 = x126 & n2093 ;
  assign n37048 = x124 & n2275 ;
  assign n37049 = x125 & n2088 ;
  assign n37050 = ~n37048 & ~n37049 ;
  assign n37051 = ~n37047 & n37050 ;
  assign n37052 = ~n2096 & n37051 ;
  assign n37053 = ~n25735 & n37051 ;
  assign n37054 = ~n37052 & ~n37053 ;
  assign n37055 = x17 & ~n37054 ;
  assign n37056 = ~x17 & n37054 ;
  assign n37057 = ~n37055 & ~n37056 ;
  assign n37058 = ~n37046 & ~n37057 ;
  assign n37059 = ~n37046 & ~n37058 ;
  assign n37060 = ~n37057 & ~n37058 ;
  assign n37061 = ~n37059 & ~n37060 ;
  assign n37062 = ~n37045 & ~n37061 ;
  assign n37063 = n37045 & ~n37060 ;
  assign n37064 = ~n37059 & n37063 ;
  assign n37065 = ~n37062 & ~n37064 ;
  assign n37066 = ~n36762 & n37065 ;
  assign n37067 = n36762 & ~n37065 ;
  assign n37068 = ~n37066 & ~n37067 ;
  assign n37069 = ~n36750 & n37068 ;
  assign n37070 = n36750 & ~n37068 ;
  assign n37071 = ~n37069 & ~n37070 ;
  assign n37072 = ~n36749 & n37071 ;
  assign n37073 = n36749 & ~n37071 ;
  assign n37074 = ~n37072 & ~n37073 ;
  assign n37402 = n37074 & x205 ;
  assign n37075 = ~n36737 & ~n36741 ;
  assign n37076 = ~n36729 & ~n36733 ;
  assign n37077 = ~n36414 & ~n36714 ;
  assign n37078 = ~x127 & n1646 ;
  assign n37079 = n1437 & n27365 ;
  assign n37080 = ~n37078 & ~n37079 ;
  assign n37081 = ~x14 & ~n37080 ;
  assign n37082 = ~x14 & ~n37081 ;
  assign n37083 = ~n37080 & ~n37081 ;
  assign n37084 = ~n37082 & ~n37083 ;
  assign n37085 = ~n37077 & ~n37084 ;
  assign n37086 = ~n37077 & ~n37085 ;
  assign n37087 = ~n37084 & ~n37085 ;
  assign n37088 = ~n37086 & ~n37087 ;
  assign n37089 = ~x123 & n2751 ;
  assign n37090 = ~x121 & n3020 ;
  assign n37091 = ~x122 & n2746 ;
  assign n37092 = ~n37090 & ~n37091 ;
  assign n37093 = ~n37089 & n37092 ;
  assign n37094 = n2754 & n23760 ;
  assign n37095 = n37093 & ~n37094 ;
  assign n37096 = ~x20 & ~n37095 ;
  assign n37097 = ~x20 & ~n37096 ;
  assign n37098 = ~n37095 & ~n37096 ;
  assign n37099 = ~n37097 & ~n37098 ;
  assign n37100 = ~n36430 & ~n36690 ;
  assign n37101 = n37099 & n37100 ;
  assign n37102 = ~n37099 & ~n37100 ;
  assign n37103 = ~n37101 & ~n37102 ;
  assign n37104 = ~x120 & n3589 ;
  assign n37105 = ~x118 & n3878 ;
  assign n37106 = ~x119 & n3584 ;
  assign n37107 = ~n37105 & ~n37106 ;
  assign n37108 = ~n37104 & n37107 ;
  assign n37109 = n3592 & n21501 ;
  assign n37110 = n37108 & ~n37109 ;
  assign n37111 = ~x23 & ~n37110 ;
  assign n37112 = ~x23 & ~n37111 ;
  assign n37113 = ~n37110 & ~n37111 ;
  assign n37114 = ~n37112 & ~n37113 ;
  assign n37115 = ~n36683 & ~n36686 ;
  assign n37116 = n37114 & n37115 ;
  assign n37117 = ~n37114 & ~n37115 ;
  assign n37118 = ~n37116 & ~n37117 ;
  assign n37119 = ~x117 & n4531 ;
  assign n37120 = ~x115 & n4847 ;
  assign n37121 = ~x116 & n4526 ;
  assign n37122 = ~n37120 & ~n37121 ;
  assign n37123 = ~n37119 & n37122 ;
  assign n37124 = n4534 & n19365 ;
  assign n37125 = n37123 & ~n37124 ;
  assign n37126 = ~x26 & ~n37125 ;
  assign n37127 = ~x26 & ~n37126 ;
  assign n37128 = ~n37125 & ~n37126 ;
  assign n37129 = ~n37127 & ~n37128 ;
  assign n37130 = ~n36446 & ~n36666 ;
  assign n37131 = n37129 & n37130 ;
  assign n37132 = ~n37129 & ~n37130 ;
  assign n37133 = ~n37131 & ~n37132 ;
  assign n37134 = ~n36628 & ~n36642 ;
  assign n37135 = ~x111 & n6725 ;
  assign n37136 = ~x109 & n7129 ;
  assign n37137 = ~x110 & n6720 ;
  assign n37138 = ~n37136 & ~n37137 ;
  assign n37139 = ~n37135 & n37138 ;
  assign n37140 = ~n6728 & n37139 ;
  assign n37141 = ~n15411 & n37139 ;
  assign n37142 = ~n37140 & ~n37141 ;
  assign n37143 = ~x32 & ~n37142 ;
  assign n37144 = x32 & n37142 ;
  assign n37145 = ~n37143 & ~n37144 ;
  assign n37146 = ~n37134 & ~n37145 ;
  assign n37147 = n37134 & n37145 ;
  assign n37148 = ~n37146 & ~n37147 ;
  assign n37149 = ~x108 & n8006 ;
  assign n37150 = ~x106 & n8474 ;
  assign n37151 = ~x107 & n8001 ;
  assign n37152 = ~n37150 & ~n37151 ;
  assign n37153 = ~n37149 & n37152 ;
  assign n37154 = n8009 & n13601 ;
  assign n37155 = n37153 & ~n37154 ;
  assign n37156 = ~x35 & ~n37155 ;
  assign n37157 = ~x35 & ~n37156 ;
  assign n37158 = ~n37155 & ~n37156 ;
  assign n37159 = ~n37157 & ~n37158 ;
  assign n37160 = ~n36620 & ~n36624 ;
  assign n37161 = ~x105 & n9433 ;
  assign n37162 = ~x103 & n9915 ;
  assign n37163 = ~x104 & n9428 ;
  assign n37164 = ~n37162 & ~n37163 ;
  assign n37165 = ~n37161 & n37164 ;
  assign n37166 = n9436 & n11907 ;
  assign n37167 = n37165 & ~n37166 ;
  assign n37168 = ~x38 & ~n37167 ;
  assign n37169 = ~x38 & ~n37168 ;
  assign n37170 = ~n37167 & ~n37168 ;
  assign n37171 = ~n37169 & ~n37170 ;
  assign n37172 = ~n36612 & ~n36616 ;
  assign n37173 = ~n36598 & ~n36602 ;
  assign n37174 = ~n36563 & ~n36576 ;
  assign n37175 = ~x90 & n18025 ;
  assign n37176 = ~x88 & n18764 ;
  assign n37177 = ~x89 & n18020 ;
  assign n37178 = ~n37176 & ~n37177 ;
  assign n37179 = ~n37175 & n37178 ;
  assign n37180 = n5155 & n18028 ;
  assign n37181 = n37179 & ~n37180 ;
  assign n37182 = ~x53 & ~n37181 ;
  assign n37183 = ~x53 & ~n37182 ;
  assign n37184 = ~n37181 & ~n37182 ;
  assign n37185 = ~n37183 & ~n37184 ;
  assign n37186 = ~n36544 & ~n36557 ;
  assign n37187 = ~n36508 & ~n36519 ;
  assign n37188 = ~n36505 & ~n37187 ;
  assign n37189 = ~x77 & n27427 ;
  assign n37190 = ~x78 & ~n26217 ;
  assign n37191 = ~n37189 & ~n37190 ;
  assign n37192 = n36502 & ~n37191 ;
  assign n37193 = ~n36502 & n37191 ;
  assign n37194 = ~n37192 & ~n37193 ;
  assign n37195 = ~x81 & n24612 ;
  assign n37196 = ~x79 & n25390 ;
  assign n37197 = ~x80 & n24607 ;
  assign n37198 = ~n37196 & ~n37197 ;
  assign n37199 = ~n37195 & n37198 ;
  assign n37200 = ~n24615 & n37199 ;
  assign n37201 = ~n2460 & n37199 ;
  assign n37202 = ~n37200 & ~n37201 ;
  assign n37203 = ~x62 & ~n37202 ;
  assign n37204 = x62 & n37202 ;
  assign n37205 = ~n37203 & ~n37204 ;
  assign n37206 = n37194 & ~n37205 ;
  assign n37207 = ~n37194 & n37205 ;
  assign n37208 = ~n37206 & ~n37207 ;
  assign n37209 = ~n37188 & n37208 ;
  assign n37210 = n37188 & ~n37208 ;
  assign n37211 = ~n37209 & ~n37210 ;
  assign n37212 = ~x84 & n22325 ;
  assign n37213 = ~x82 & n23066 ;
  assign n37214 = ~x83 & n22320 ;
  assign n37215 = ~n37213 & ~n37214 ;
  assign n37216 = ~n37212 & n37215 ;
  assign n37217 = n3247 & n22328 ;
  assign n37218 = n37216 & ~n37217 ;
  assign n37219 = ~x59 & ~n37218 ;
  assign n37220 = ~x59 & ~n37219 ;
  assign n37221 = ~n37218 & ~n37219 ;
  assign n37222 = ~n37220 & ~n37221 ;
  assign n37223 = n37211 & ~n37222 ;
  assign n37224 = n37211 & ~n37223 ;
  assign n37225 = ~n37222 & ~n37223 ;
  assign n37226 = ~n37224 & ~n37225 ;
  assign n37227 = ~n36525 & ~n36538 ;
  assign n37228 = n37226 & n37227 ;
  assign n37229 = ~n37226 & ~n37227 ;
  assign n37230 = ~n37228 & ~n37229 ;
  assign n37231 = ~x87 & n20143 ;
  assign n37232 = ~x85 & n20854 ;
  assign n37233 = ~x86 & n20138 ;
  assign n37234 = ~n37232 & ~n37233 ;
  assign n37235 = ~n37231 & n37234 ;
  assign n37236 = n4143 & n20146 ;
  assign n37237 = n37235 & ~n37236 ;
  assign n37238 = ~x56 & ~n37237 ;
  assign n37239 = ~x56 & ~n37238 ;
  assign n37240 = ~n37237 & ~n37238 ;
  assign n37241 = ~n37239 & ~n37240 ;
  assign n37242 = ~n37230 & n37241 ;
  assign n37243 = n37230 & ~n37241 ;
  assign n37244 = ~n37242 & ~n37243 ;
  assign n37245 = ~n37186 & n37244 ;
  assign n37246 = n37186 & ~n37244 ;
  assign n37247 = ~n37245 & ~n37246 ;
  assign n37248 = ~n37185 & n37247 ;
  assign n37249 = n37185 & ~n37247 ;
  assign n37250 = ~n37248 & ~n37249 ;
  assign n37251 = ~n37174 & n37250 ;
  assign n37252 = n37174 & ~n37250 ;
  assign n37253 = ~n37251 & ~n37252 ;
  assign n37254 = ~x93 & n16076 ;
  assign n37255 = ~x91 & n16756 ;
  assign n37256 = ~x92 & n16071 ;
  assign n37257 = ~n37255 & ~n37256 ;
  assign n37258 = ~n37254 & n37257 ;
  assign n37259 = n6285 & n16079 ;
  assign n37260 = n37258 & ~n37259 ;
  assign n37261 = ~x50 & ~n37260 ;
  assign n37262 = ~x50 & ~n37261 ;
  assign n37263 = ~n37260 & ~n37261 ;
  assign n37264 = ~n37262 & ~n37263 ;
  assign n37265 = n37253 & ~n37264 ;
  assign n37266 = n37253 & ~n37265 ;
  assign n37267 = ~n37264 & ~n37265 ;
  assign n37268 = ~n37266 & ~n37267 ;
  assign n37269 = ~n36582 & ~n36596 ;
  assign n37270 = ~n37268 & ~n37269 ;
  assign n37271 = ~n37268 & ~n37270 ;
  assign n37272 = ~n37269 & ~n37270 ;
  assign n37273 = ~n37271 & ~n37272 ;
  assign n37274 = ~x96 & n14233 ;
  assign n37275 = ~x94 & n14876 ;
  assign n37276 = ~x95 & n14228 ;
  assign n37277 = ~n37275 & ~n37276 ;
  assign n37278 = ~n37274 & n37277 ;
  assign n37279 = n7531 & n14236 ;
  assign n37280 = n37278 & ~n37279 ;
  assign n37281 = ~x47 & ~n37280 ;
  assign n37282 = ~x47 & ~n37281 ;
  assign n37283 = ~n37280 & ~n37281 ;
  assign n37284 = ~n37282 & ~n37283 ;
  assign n37285 = ~n37273 & n37284 ;
  assign n37286 = n37273 & ~n37284 ;
  assign n37287 = ~n37285 & ~n37286 ;
  assign n37288 = n37173 & n37287 ;
  assign n37289 = ~n37173 & ~n37287 ;
  assign n37290 = ~n37288 & ~n37289 ;
  assign n37291 = ~x99 & n12506 ;
  assign n37292 = ~x97 & n13131 ;
  assign n37293 = ~x98 & n12501 ;
  assign n37294 = ~n37292 & ~n37293 ;
  assign n37295 = ~n37291 & n37294 ;
  assign n37296 = n8885 & n12509 ;
  assign n37297 = n37295 & ~n37296 ;
  assign n37298 = ~x44 & ~n37297 ;
  assign n37299 = ~x44 & ~n37298 ;
  assign n37300 = ~n37297 & ~n37298 ;
  assign n37301 = ~n37299 & ~n37300 ;
  assign n37302 = n37290 & ~n37301 ;
  assign n37303 = n37290 & ~n37302 ;
  assign n37304 = ~n37301 & ~n37302 ;
  assign n37305 = ~n37303 & ~n37304 ;
  assign n37306 = ~n36606 & ~n36609 ;
  assign n37307 = n37305 & n37306 ;
  assign n37308 = ~n37305 & ~n37306 ;
  assign n37309 = ~n37307 & ~n37308 ;
  assign n37310 = ~x102 & n10905 ;
  assign n37311 = ~x100 & n11466 ;
  assign n37312 = ~x101 & n10900 ;
  assign n37313 = ~n37311 & ~n37312 ;
  assign n37314 = ~n37310 & n37313 ;
  assign n37315 = n10333 & n10908 ;
  assign n37316 = n37314 & ~n37315 ;
  assign n37317 = ~x41 & ~n37316 ;
  assign n37318 = ~x41 & ~n37317 ;
  assign n37319 = ~n37316 & ~n37317 ;
  assign n37320 = ~n37318 & ~n37319 ;
  assign n37321 = ~n37309 & n37320 ;
  assign n37322 = n37309 & ~n37320 ;
  assign n37323 = ~n37321 & ~n37322 ;
  assign n37324 = ~n37172 & n37323 ;
  assign n37325 = n37172 & ~n37323 ;
  assign n37326 = ~n37324 & ~n37325 ;
  assign n37327 = ~n37171 & n37326 ;
  assign n37328 = n37171 & ~n37326 ;
  assign n37329 = ~n37327 & ~n37328 ;
  assign n37330 = ~n37160 & n37329 ;
  assign n37331 = n37160 & ~n37329 ;
  assign n37332 = ~n37330 & ~n37331 ;
  assign n37333 = ~n37159 & n37332 ;
  assign n37334 = ~n37159 & ~n37333 ;
  assign n37335 = n37332 & ~n37333 ;
  assign n37336 = ~n37334 & ~n37335 ;
  assign n37337 = n37148 & ~n37336 ;
  assign n37338 = n37148 & ~n37337 ;
  assign n37339 = ~n37336 & ~n37337 ;
  assign n37340 = ~n37338 & ~n37339 ;
  assign n37341 = ~n36658 & ~n36662 ;
  assign n37342 = ~x114 & n5560 ;
  assign n37343 = ~x112 & n5943 ;
  assign n37344 = ~x113 & n5555 ;
  assign n37345 = ~n37343 & ~n37344 ;
  assign n37346 = ~n37342 & n37345 ;
  assign n37347 = ~n5563 & n37346 ;
  assign n37348 = ~n17333 & n37346 ;
  assign n37349 = ~n37347 & ~n37348 ;
  assign n37350 = ~x29 & ~n37349 ;
  assign n37351 = x29 & n37349 ;
  assign n37352 = ~n37350 & ~n37351 ;
  assign n37353 = ~n37341 & ~n37352 ;
  assign n37354 = n37341 & n37352 ;
  assign n37355 = ~n37353 & ~n37354 ;
  assign n37356 = ~n37340 & n37355 ;
  assign n37357 = ~n37340 & ~n37356 ;
  assign n37358 = n37355 & ~n37356 ;
  assign n37359 = ~n37357 & ~n37358 ;
  assign n37360 = n37133 & ~n37359 ;
  assign n37361 = n37133 & ~n37360 ;
  assign n37362 = ~n37359 & ~n37360 ;
  assign n37363 = ~n37361 & ~n37362 ;
  assign n37364 = n37118 & ~n37363 ;
  assign n37365 = ~n37118 & n37363 ;
  assign n37366 = n37103 & ~n37365 ;
  assign n37367 = ~n37364 & n37366 ;
  assign n37368 = n37103 & ~n37367 ;
  assign n37369 = ~n37365 & ~n37367 ;
  assign n37370 = ~n37364 & n37369 ;
  assign n37371 = ~n37368 & ~n37370 ;
  assign n37372 = ~n36706 & ~n36710 ;
  assign n37373 = ~x126 & n2093 ;
  assign n37374 = ~x124 & n2275 ;
  assign n37375 = ~x125 & n2088 ;
  assign n37376 = ~n37374 & ~n37375 ;
  assign n37377 = ~n37373 & n37376 ;
  assign n37378 = ~n2096 & n37377 ;
  assign n37379 = ~n26128 & n37377 ;
  assign n37380 = ~n37378 & ~n37379 ;
  assign n37381 = ~x17 & ~n37380 ;
  assign n37382 = x17 & n37380 ;
  assign n37383 = ~n37381 & ~n37382 ;
  assign n37384 = ~n37372 & ~n37383 ;
  assign n37385 = ~n37372 & ~n37384 ;
  assign n37386 = ~n37383 & ~n37384 ;
  assign n37387 = ~n37385 & ~n37386 ;
  assign n37388 = ~n37371 & ~n37387 ;
  assign n37389 = n37371 & ~n37386 ;
  assign n37390 = ~n37385 & n37389 ;
  assign n37391 = ~n37388 & ~n37390 ;
  assign n37392 = ~n37088 & n37391 ;
  assign n37393 = n37088 & ~n37391 ;
  assign n37394 = ~n37392 & ~n37393 ;
  assign n37395 = ~n37076 & n37394 ;
  assign n37396 = n37076 & ~n37394 ;
  assign n37397 = ~n37395 & ~n37396 ;
  assign n37398 = ~n37075 & n37397 ;
  assign n37399 = n37075 & ~n37397 ;
  assign n37400 = ~n37398 & ~n37399 ;
  assign n37403 = ~n37400 & ~x205 ;
  assign n37404 = ~n37402 & ~n37403 ;
  assign n37405 = ~n37058 & ~n37062 ;
  assign n37406 = x127 & n2093 ;
  assign n37407 = x125 & n2275 ;
  assign n37408 = x126 & n2088 ;
  assign n37409 = ~n37407 & ~n37408 ;
  assign n37410 = ~n37406 & n37409 ;
  assign n37411 = n2096 & n26533 ;
  assign n37412 = n37410 & ~n37411 ;
  assign n37413 = x17 & ~n37412 ;
  assign n37414 = x17 & ~n37413 ;
  assign n37415 = ~n37412 & ~n37413 ;
  assign n37416 = ~n37414 & ~n37415 ;
  assign n37417 = ~n37405 & ~n37416 ;
  assign n37418 = ~n37405 & ~n37417 ;
  assign n37419 = ~n37416 & ~n37417 ;
  assign n37420 = ~n37418 & ~n37419 ;
  assign n37421 = x124 & n2751 ;
  assign n37422 = x122 & n3020 ;
  assign n37423 = x123 & n2746 ;
  assign n37424 = ~n37422 & ~n37423 ;
  assign n37425 = ~n37421 & n37424 ;
  assign n37426 = n2754 & n23796 ;
  assign n37427 = n37425 & ~n37426 ;
  assign n37428 = x20 & ~n37427 ;
  assign n37429 = x20 & ~n37428 ;
  assign n37430 = ~n37427 & ~n37428 ;
  assign n37431 = ~n37429 & ~n37430 ;
  assign n37432 = ~n36776 & ~n37041 ;
  assign n37433 = n37431 & n37432 ;
  assign n37434 = ~n37431 & ~n37432 ;
  assign n37435 = ~n37433 & ~n37434 ;
  assign n37436 = ~n36791 & ~n37038 ;
  assign n37437 = x121 & n3589 ;
  assign n37438 = x119 & n3878 ;
  assign n37439 = x120 & n3584 ;
  assign n37440 = ~n37438 & ~n37439 ;
  assign n37441 = ~n37437 & n37440 ;
  assign n37442 = n3592 & n21870 ;
  assign n37443 = n37441 & ~n37442 ;
  assign n37444 = x23 & ~n37443 ;
  assign n37445 = x23 & ~n37444 ;
  assign n37446 = ~n37443 & ~n37444 ;
  assign n37447 = ~n37445 & ~n37446 ;
  assign n37448 = ~n37436 & n37447 ;
  assign n37449 = n37436 & ~n37447 ;
  assign n37450 = ~n37448 & ~n37449 ;
  assign n37451 = x118 & n4531 ;
  assign n37452 = x116 & n4847 ;
  assign n37453 = x117 & n4526 ;
  assign n37454 = ~n37452 & ~n37453 ;
  assign n37455 = ~n37451 & n37454 ;
  assign n37456 = n4534 & n19395 ;
  assign n37457 = n37455 & ~n37456 ;
  assign n37458 = x26 & ~n37457 ;
  assign n37459 = x26 & ~n37458 ;
  assign n37460 = ~n37457 & ~n37458 ;
  assign n37461 = ~n37459 & ~n37460 ;
  assign n37462 = ~n36806 & ~n37034 ;
  assign n37463 = n37461 & n37462 ;
  assign n37464 = ~n37461 & ~n37462 ;
  assign n37465 = ~n37463 & ~n37464 ;
  assign n37466 = x115 & n5560 ;
  assign n37467 = x113 & n5943 ;
  assign n37468 = x114 & n5555 ;
  assign n37469 = ~n37467 & ~n37468 ;
  assign n37470 = ~n37466 & n37469 ;
  assign n37471 = n5563 & n17364 ;
  assign n37472 = n37470 & ~n37471 ;
  assign n37473 = x29 & ~n37472 ;
  assign n37474 = x29 & ~n37473 ;
  assign n37475 = ~n37472 & ~n37473 ;
  assign n37476 = ~n37474 & ~n37475 ;
  assign n37477 = ~n37027 & ~n37030 ;
  assign n37478 = n37476 & n37477 ;
  assign n37479 = ~n37476 & ~n37477 ;
  assign n37480 = ~n37478 & ~n37479 ;
  assign n37481 = ~n36998 & ~n37001 ;
  assign n37482 = ~n36982 & ~n36996 ;
  assign n37483 = ~n36963 & ~n36976 ;
  assign n37484 = ~n36947 & ~n36958 ;
  assign n37485 = ~n36944 & ~n37484 ;
  assign n37486 = ~n36903 & ~n36917 ;
  assign n37487 = x78 & n27024 ;
  assign n37488 = x79 & ~n26217 ;
  assign n37489 = ~n37487 & ~n37488 ;
  assign n37490 = ~x14 & ~n37489 ;
  assign n37491 = ~x14 & ~n37490 ;
  assign n37492 = ~n37489 & ~n37490 ;
  assign n37493 = ~n37491 & ~n37492 ;
  assign n37494 = ~n36156 & ~n37493 ;
  assign n37495 = ~n36156 & ~n37494 ;
  assign n37496 = ~n37493 & ~n37494 ;
  assign n37497 = ~n37495 & ~n37496 ;
  assign n37498 = x82 & n24612 ;
  assign n37499 = x80 & n25390 ;
  assign n37500 = x81 & n24607 ;
  assign n37501 = ~n37499 & ~n37500 ;
  assign n37502 = ~n37498 & n37501 ;
  assign n37503 = n2584 & n24615 ;
  assign n37504 = n37502 & ~n37503 ;
  assign n37505 = x62 & ~n37504 ;
  assign n37506 = x62 & ~n37505 ;
  assign n37507 = ~n37504 & ~n37505 ;
  assign n37508 = ~n37506 & ~n37507 ;
  assign n37509 = ~n37497 & ~n37508 ;
  assign n37510 = ~n37497 & ~n37509 ;
  assign n37511 = ~n37508 & ~n37509 ;
  assign n37512 = ~n37510 & ~n37511 ;
  assign n37513 = ~n36866 & ~n36880 ;
  assign n37514 = n37512 & n37513 ;
  assign n37515 = ~n37512 & ~n37513 ;
  assign n37516 = ~n37514 & ~n37515 ;
  assign n37517 = x85 & n22325 ;
  assign n37518 = x83 & n23066 ;
  assign n37519 = x84 & n22320 ;
  assign n37520 = ~n37518 & ~n37519 ;
  assign n37521 = ~n37517 & n37520 ;
  assign n37522 = n3389 & n22328 ;
  assign n37523 = n37521 & ~n37522 ;
  assign n37524 = x59 & ~n37523 ;
  assign n37525 = x59 & ~n37524 ;
  assign n37526 = ~n37523 & ~n37524 ;
  assign n37527 = ~n37525 & ~n37526 ;
  assign n37528 = n37516 & ~n37527 ;
  assign n37529 = n37516 & ~n37528 ;
  assign n37530 = ~n37527 & ~n37528 ;
  assign n37531 = ~n37529 & ~n37530 ;
  assign n37532 = ~n36883 & ~n36897 ;
  assign n37533 = n37531 & n37532 ;
  assign n37534 = ~n37531 & ~n37532 ;
  assign n37535 = ~n37533 & ~n37534 ;
  assign n37536 = x88 & n20143 ;
  assign n37537 = x86 & n20854 ;
  assign n37538 = x87 & n20138 ;
  assign n37539 = ~n37537 & ~n37538 ;
  assign n37540 = ~n37536 & n37539 ;
  assign n37541 = n4305 & n20146 ;
  assign n37542 = n37540 & ~n37541 ;
  assign n37543 = x56 & ~n37542 ;
  assign n37544 = x56 & ~n37543 ;
  assign n37545 = ~n37542 & ~n37543 ;
  assign n37546 = ~n37544 & ~n37545 ;
  assign n37547 = n37535 & ~n37546 ;
  assign n37548 = ~n37535 & n37546 ;
  assign n37549 = ~n37486 & ~n37548 ;
  assign n37550 = ~n37547 & n37549 ;
  assign n37551 = ~n37486 & ~n37550 ;
  assign n37552 = ~n37547 & ~n37550 ;
  assign n37553 = ~n37548 & n37552 ;
  assign n37554 = ~n37551 & ~n37553 ;
  assign n37555 = x91 & n18025 ;
  assign n37556 = x89 & n18764 ;
  assign n37557 = x90 & n18020 ;
  assign n37558 = ~n37556 & ~n37557 ;
  assign n37559 = ~n37555 & n37558 ;
  assign n37560 = n5336 & n18028 ;
  assign n37561 = n37559 & ~n37560 ;
  assign n37562 = x53 & ~n37561 ;
  assign n37563 = x53 & ~n37562 ;
  assign n37564 = ~n37561 & ~n37562 ;
  assign n37565 = ~n37563 & ~n37564 ;
  assign n37566 = ~n37554 & ~n37565 ;
  assign n37567 = ~n37554 & ~n37566 ;
  assign n37568 = ~n37565 & ~n37566 ;
  assign n37569 = ~n37567 & ~n37568 ;
  assign n37570 = ~n36919 & ~n36922 ;
  assign n37571 = n37569 & n37570 ;
  assign n37572 = ~n37569 & ~n37570 ;
  assign n37573 = ~n37571 & ~n37572 ;
  assign n37574 = x94 & n16076 ;
  assign n37575 = x92 & n16756 ;
  assign n37576 = x93 & n16071 ;
  assign n37577 = ~n37575 & ~n37576 ;
  assign n37578 = ~n37574 & n37577 ;
  assign n37579 = n6483 & n16079 ;
  assign n37580 = n37578 & ~n37579 ;
  assign n37581 = x50 & ~n37580 ;
  assign n37582 = x50 & ~n37581 ;
  assign n37583 = ~n37580 & ~n37581 ;
  assign n37584 = ~n37582 & ~n37583 ;
  assign n37585 = n37573 & ~n37584 ;
  assign n37586 = n37573 & ~n37585 ;
  assign n37587 = ~n37584 & ~n37585 ;
  assign n37588 = ~n37586 & ~n37587 ;
  assign n37589 = ~n36925 & ~n36939 ;
  assign n37590 = n37588 & n37589 ;
  assign n37591 = ~n37588 & ~n37589 ;
  assign n37592 = ~n37590 & ~n37591 ;
  assign n37593 = x97 & n14233 ;
  assign n37594 = x95 & n14876 ;
  assign n37595 = x96 & n14228 ;
  assign n37596 = ~n37594 & ~n37595 ;
  assign n37597 = ~n37593 & n37596 ;
  assign n37598 = n7745 & n14236 ;
  assign n37599 = n37597 & ~n37598 ;
  assign n37600 = x47 & ~n37599 ;
  assign n37601 = x47 & ~n37600 ;
  assign n37602 = ~n37599 & ~n37600 ;
  assign n37603 = ~n37601 & ~n37602 ;
  assign n37604 = n37592 & ~n37603 ;
  assign n37605 = n37592 & ~n37604 ;
  assign n37606 = ~n37603 & ~n37604 ;
  assign n37607 = ~n37605 & ~n37606 ;
  assign n37608 = ~n37485 & n37607 ;
  assign n37609 = n37485 & ~n37607 ;
  assign n37610 = ~n37608 & ~n37609 ;
  assign n37611 = x100 & n12506 ;
  assign n37612 = x98 & n13131 ;
  assign n37613 = x99 & n12501 ;
  assign n37614 = ~n37612 & ~n37613 ;
  assign n37615 = ~n37611 & n37614 ;
  assign n37616 = n9115 & n12509 ;
  assign n37617 = n37615 & ~n37616 ;
  assign n37618 = x44 & ~n37617 ;
  assign n37619 = x44 & ~n37618 ;
  assign n37620 = ~n37617 & ~n37618 ;
  assign n37621 = ~n37619 & ~n37620 ;
  assign n37622 = ~n37610 & ~n37621 ;
  assign n37623 = n37610 & n37621 ;
  assign n37624 = ~n37622 & ~n37623 ;
  assign n37625 = n37483 & ~n37624 ;
  assign n37626 = ~n37483 & n37624 ;
  assign n37627 = ~n37625 & ~n37626 ;
  assign n37628 = x103 & n10905 ;
  assign n37629 = x101 & n11466 ;
  assign n37630 = x102 & n10900 ;
  assign n37631 = ~n37629 & ~n37630 ;
  assign n37632 = ~n37628 & n37631 ;
  assign n37633 = n10588 & n10908 ;
  assign n37634 = n37632 & ~n37633 ;
  assign n37635 = x41 & ~n37634 ;
  assign n37636 = x41 & ~n37635 ;
  assign n37637 = ~n37634 & ~n37635 ;
  assign n37638 = ~n37636 & ~n37637 ;
  assign n37639 = n37627 & ~n37638 ;
  assign n37640 = n37627 & ~n37639 ;
  assign n37641 = ~n37638 & ~n37639 ;
  assign n37642 = ~n37640 & ~n37641 ;
  assign n37643 = ~n37482 & n37642 ;
  assign n37644 = n37482 & ~n37642 ;
  assign n37645 = ~n37643 & ~n37644 ;
  assign n37646 = x106 & n9433 ;
  assign n37647 = x104 & n9915 ;
  assign n37648 = x105 & n9428 ;
  assign n37649 = ~n37647 & ~n37648 ;
  assign n37650 = ~n37646 & n37649 ;
  assign n37651 = n9436 & n12181 ;
  assign n37652 = n37650 & ~n37651 ;
  assign n37653 = x38 & ~n37652 ;
  assign n37654 = x38 & ~n37653 ;
  assign n37655 = ~n37652 & ~n37653 ;
  assign n37656 = ~n37654 & ~n37655 ;
  assign n37657 = ~n37645 & ~n37656 ;
  assign n37658 = n37645 & n37656 ;
  assign n37659 = ~n37657 & ~n37658 ;
  assign n37660 = n37481 & ~n37659 ;
  assign n37661 = ~n37481 & n37659 ;
  assign n37662 = ~n37660 & ~n37661 ;
  assign n37663 = x109 & n8006 ;
  assign n37664 = x107 & n8474 ;
  assign n37665 = x108 & n8001 ;
  assign n37666 = ~n37664 & ~n37665 ;
  assign n37667 = ~n37663 & n37666 ;
  assign n37668 = n8009 & n13894 ;
  assign n37669 = n37667 & ~n37668 ;
  assign n37670 = x35 & ~n37669 ;
  assign n37671 = x35 & ~n37670 ;
  assign n37672 = ~n37669 & ~n37670 ;
  assign n37673 = ~n37671 & ~n37672 ;
  assign n37674 = n37662 & ~n37673 ;
  assign n37675 = n37662 & ~n37674 ;
  assign n37676 = ~n37673 & ~n37674 ;
  assign n37677 = ~n37675 & ~n37676 ;
  assign n37678 = ~n37004 & ~n37007 ;
  assign n37679 = n37677 & n37678 ;
  assign n37680 = ~n37677 & ~n37678 ;
  assign n37681 = ~n37679 & ~n37680 ;
  assign n37682 = ~n36820 & ~n37011 ;
  assign n37683 = x112 & n6725 ;
  assign n37684 = x110 & n7129 ;
  assign n37685 = x111 & n6720 ;
  assign n37686 = ~n37684 & ~n37685 ;
  assign n37687 = ~n37683 & n37686 ;
  assign n37688 = n6728 & n15442 ;
  assign n37689 = n37687 & ~n37688 ;
  assign n37690 = x32 & ~n37689 ;
  assign n37691 = x32 & ~n37690 ;
  assign n37692 = ~n37689 & ~n37690 ;
  assign n37693 = ~n37691 & ~n37692 ;
  assign n37694 = ~n37682 & ~n37693 ;
  assign n37695 = ~n37682 & ~n37694 ;
  assign n37696 = ~n37693 & ~n37694 ;
  assign n37697 = ~n37695 & ~n37696 ;
  assign n37698 = n37681 & ~n37697 ;
  assign n37699 = ~n37681 & n37697 ;
  assign n37700 = n37480 & ~n37699 ;
  assign n37701 = ~n37698 & n37700 ;
  assign n37702 = n37480 & ~n37701 ;
  assign n37703 = ~n37699 & ~n37701 ;
  assign n37704 = ~n37698 & n37703 ;
  assign n37705 = ~n37702 & ~n37704 ;
  assign n37706 = n37465 & ~n37705 ;
  assign n37707 = ~n37465 & n37705 ;
  assign n37708 = ~n37450 & ~n37707 ;
  assign n37709 = ~n37706 & n37708 ;
  assign n37710 = ~n37450 & ~n37709 ;
  assign n37711 = ~n37707 & ~n37709 ;
  assign n37712 = ~n37706 & n37711 ;
  assign n37713 = ~n37710 & ~n37712 ;
  assign n37714 = n37435 & ~n37713 ;
  assign n37715 = ~n37435 & n37713 ;
  assign n37716 = ~n37420 & ~n37715 ;
  assign n37717 = ~n37714 & n37716 ;
  assign n37718 = ~n37420 & ~n37717 ;
  assign n37719 = ~n37715 & ~n37717 ;
  assign n37720 = ~n37714 & n37719 ;
  assign n37721 = ~n37718 & ~n37720 ;
  assign n37722 = ~n36759 & ~n37066 ;
  assign n37723 = n37721 & n37722 ;
  assign n37724 = ~n37721 & ~n37722 ;
  assign n37725 = ~n37723 & ~n37724 ;
  assign n37726 = ~n37069 & ~n37072 ;
  assign n37727 = n37725 & ~n37726 ;
  assign n37728 = ~n37725 & n37726 ;
  assign n37729 = ~n37727 & ~n37728 ;
  assign n38056 = n37729 & x206 ;
  assign n37730 = ~n37384 & ~n37388 ;
  assign n37731 = ~x127 & n2093 ;
  assign n37732 = ~x125 & n2275 ;
  assign n37733 = ~x126 & n2088 ;
  assign n37734 = ~n37732 & ~n37733 ;
  assign n37735 = ~n37731 & n37734 ;
  assign n37736 = n2096 & n26932 ;
  assign n37737 = n37735 & ~n37736 ;
  assign n37738 = ~x17 & ~n37737 ;
  assign n37739 = ~x17 & ~n37738 ;
  assign n37740 = ~n37737 & ~n37738 ;
  assign n37741 = ~n37739 & ~n37740 ;
  assign n37742 = ~n37730 & ~n37741 ;
  assign n37743 = ~n37730 & ~n37742 ;
  assign n37744 = ~n37741 & ~n37742 ;
  assign n37745 = ~n37743 & ~n37744 ;
  assign n37746 = ~x124 & n2751 ;
  assign n37747 = ~x122 & n3020 ;
  assign n37748 = ~x123 & n2746 ;
  assign n37749 = ~n37747 & ~n37748 ;
  assign n37750 = ~n37746 & n37749 ;
  assign n37751 = n2754 & n24176 ;
  assign n37752 = n37750 & ~n37751 ;
  assign n37753 = ~x20 & ~n37752 ;
  assign n37754 = ~x20 & ~n37753 ;
  assign n37755 = ~n37752 & ~n37753 ;
  assign n37756 = ~n37754 & ~n37755 ;
  assign n37757 = ~n37102 & ~n37367 ;
  assign n37758 = n37756 & n37757 ;
  assign n37759 = ~n37756 & ~n37757 ;
  assign n37760 = ~n37758 & ~n37759 ;
  assign n37761 = ~n37117 & ~n37364 ;
  assign n37762 = ~x121 & n3589 ;
  assign n37763 = ~x119 & n3878 ;
  assign n37764 = ~x120 & n3584 ;
  assign n37765 = ~n37763 & ~n37764 ;
  assign n37766 = ~n37762 & n37765 ;
  assign n37767 = n3592 & n22229 ;
  assign n37768 = n37766 & ~n37767 ;
  assign n37769 = ~x23 & ~n37768 ;
  assign n37770 = ~x23 & ~n37769 ;
  assign n37771 = ~n37768 & ~n37769 ;
  assign n37772 = ~n37770 & ~n37771 ;
  assign n37773 = ~n37761 & n37772 ;
  assign n37774 = n37761 & ~n37772 ;
  assign n37775 = ~n37773 & ~n37774 ;
  assign n37776 = ~x118 & n4531 ;
  assign n37777 = ~x116 & n4847 ;
  assign n37778 = ~x117 & n4526 ;
  assign n37779 = ~n37777 & ~n37778 ;
  assign n37780 = ~n37776 & n37779 ;
  assign n37781 = n4534 & n19736 ;
  assign n37782 = n37780 & ~n37781 ;
  assign n37783 = ~x26 & ~n37782 ;
  assign n37784 = ~x26 & ~n37783 ;
  assign n37785 = ~n37782 & ~n37783 ;
  assign n37786 = ~n37784 & ~n37785 ;
  assign n37787 = ~n37132 & ~n37360 ;
  assign n37788 = n37786 & n37787 ;
  assign n37789 = ~n37786 & ~n37787 ;
  assign n37790 = ~n37788 & ~n37789 ;
  assign n37791 = ~x115 & n5560 ;
  assign n37792 = ~x113 & n5943 ;
  assign n37793 = ~x114 & n5555 ;
  assign n37794 = ~n37792 & ~n37793 ;
  assign n37795 = ~n37791 & n37794 ;
  assign n37796 = n5563 & n17683 ;
  assign n37797 = n37795 & ~n37796 ;
  assign n37798 = ~x29 & ~n37797 ;
  assign n37799 = ~x29 & ~n37798 ;
  assign n37800 = ~n37797 & ~n37798 ;
  assign n37801 = ~n37799 & ~n37800 ;
  assign n37802 = ~n37353 & ~n37356 ;
  assign n37803 = n37801 & n37802 ;
  assign n37804 = ~n37801 & ~n37802 ;
  assign n37805 = ~n37803 & ~n37804 ;
  assign n37806 = ~n37324 & ~n37327 ;
  assign n37807 = ~n37308 & ~n37322 ;
  assign n37808 = ~n37289 & ~n37302 ;
  assign n37809 = ~n37273 & ~n37284 ;
  assign n37810 = ~n37270 & ~n37809 ;
  assign n37811 = ~n37229 & ~n37243 ;
  assign n37812 = ~x78 & n27427 ;
  assign n37813 = ~x79 & ~n26217 ;
  assign n37814 = ~n37812 & ~n37813 ;
  assign n37815 = x14 & ~n37814 ;
  assign n37816 = x14 & ~n37815 ;
  assign n37817 = ~n37814 & ~n37815 ;
  assign n37818 = ~n37816 & ~n37817 ;
  assign n37819 = ~n36502 & ~n37818 ;
  assign n37820 = ~n36502 & ~n37819 ;
  assign n37821 = ~n37818 & ~n37819 ;
  assign n37822 = ~n37820 & ~n37821 ;
  assign n37823 = ~x82 & n24612 ;
  assign n37824 = ~x80 & n25390 ;
  assign n37825 = ~x81 & n24607 ;
  assign n37826 = ~n37824 & ~n37825 ;
  assign n37827 = ~n37823 & n37826 ;
  assign n37828 = n2697 & n24615 ;
  assign n37829 = n37827 & ~n37828 ;
  assign n37830 = ~x62 & ~n37829 ;
  assign n37831 = ~x62 & ~n37830 ;
  assign n37832 = ~n37829 & ~n37830 ;
  assign n37833 = ~n37831 & ~n37832 ;
  assign n37834 = ~n37822 & ~n37833 ;
  assign n37835 = ~n37822 & ~n37834 ;
  assign n37836 = ~n37833 & ~n37834 ;
  assign n37837 = ~n37835 & ~n37836 ;
  assign n37838 = ~n37192 & ~n37206 ;
  assign n37839 = n37837 & n37838 ;
  assign n37840 = ~n37837 & ~n37838 ;
  assign n37841 = ~n37839 & ~n37840 ;
  assign n37842 = ~x85 & n22325 ;
  assign n37843 = ~x83 & n23066 ;
  assign n37844 = ~x84 & n22320 ;
  assign n37845 = ~n37843 & ~n37844 ;
  assign n37846 = ~n37842 & n37845 ;
  assign n37847 = n3521 & n22328 ;
  assign n37848 = n37846 & ~n37847 ;
  assign n37849 = ~x59 & ~n37848 ;
  assign n37850 = ~x59 & ~n37849 ;
  assign n37851 = ~n37848 & ~n37849 ;
  assign n37852 = ~n37850 & ~n37851 ;
  assign n37853 = n37841 & ~n37852 ;
  assign n37854 = n37841 & ~n37853 ;
  assign n37855 = ~n37852 & ~n37853 ;
  assign n37856 = ~n37854 & ~n37855 ;
  assign n37857 = ~n37209 & ~n37223 ;
  assign n37858 = n37856 & n37857 ;
  assign n37859 = ~n37856 & ~n37857 ;
  assign n37860 = ~n37858 & ~n37859 ;
  assign n37861 = ~x88 & n20143 ;
  assign n37862 = ~x86 & n20854 ;
  assign n37863 = ~x87 & n20138 ;
  assign n37864 = ~n37862 & ~n37863 ;
  assign n37865 = ~n37861 & n37864 ;
  assign n37866 = n4457 & n20146 ;
  assign n37867 = n37865 & ~n37866 ;
  assign n37868 = ~x56 & ~n37867 ;
  assign n37869 = ~x56 & ~n37868 ;
  assign n37870 = ~n37867 & ~n37868 ;
  assign n37871 = ~n37869 & ~n37870 ;
  assign n37872 = n37860 & ~n37871 ;
  assign n37873 = ~n37860 & n37871 ;
  assign n37874 = ~n37811 & ~n37873 ;
  assign n37875 = ~n37872 & n37874 ;
  assign n37876 = ~n37811 & ~n37875 ;
  assign n37877 = ~n37872 & ~n37875 ;
  assign n37878 = ~n37873 & n37877 ;
  assign n37879 = ~n37876 & ~n37878 ;
  assign n37880 = ~x91 & n18025 ;
  assign n37881 = ~x89 & n18764 ;
  assign n37882 = ~x90 & n18020 ;
  assign n37883 = ~n37881 & ~n37882 ;
  assign n37884 = ~n37880 & n37883 ;
  assign n37885 = n5507 & n18028 ;
  assign n37886 = n37884 & ~n37885 ;
  assign n37887 = ~x53 & ~n37886 ;
  assign n37888 = ~x53 & ~n37887 ;
  assign n37889 = ~n37886 & ~n37887 ;
  assign n37890 = ~n37888 & ~n37889 ;
  assign n37891 = ~n37879 & ~n37890 ;
  assign n37892 = ~n37879 & ~n37891 ;
  assign n37893 = ~n37890 & ~n37891 ;
  assign n37894 = ~n37892 & ~n37893 ;
  assign n37895 = ~n37245 & ~n37248 ;
  assign n37896 = n37894 & n37895 ;
  assign n37897 = ~n37894 & ~n37895 ;
  assign n37898 = ~n37896 & ~n37897 ;
  assign n37899 = ~x94 & n16076 ;
  assign n37900 = ~x92 & n16756 ;
  assign n37901 = ~x93 & n16071 ;
  assign n37902 = ~n37900 & ~n37901 ;
  assign n37903 = ~n37899 & n37902 ;
  assign n37904 = n6671 & n16079 ;
  assign n37905 = n37903 & ~n37904 ;
  assign n37906 = ~x50 & ~n37905 ;
  assign n37907 = ~x50 & ~n37906 ;
  assign n37908 = ~n37905 & ~n37906 ;
  assign n37909 = ~n37907 & ~n37908 ;
  assign n37910 = n37898 & ~n37909 ;
  assign n37911 = n37898 & ~n37910 ;
  assign n37912 = ~n37909 & ~n37910 ;
  assign n37913 = ~n37911 & ~n37912 ;
  assign n37914 = ~n37251 & ~n37265 ;
  assign n37915 = n37913 & n37914 ;
  assign n37916 = ~n37913 & ~n37914 ;
  assign n37917 = ~n37915 & ~n37916 ;
  assign n37918 = ~x97 & n14233 ;
  assign n37919 = ~x95 & n14876 ;
  assign n37920 = ~x96 & n14228 ;
  assign n37921 = ~n37919 & ~n37920 ;
  assign n37922 = ~n37918 & n37921 ;
  assign n37923 = n7949 & n14236 ;
  assign n37924 = n37922 & ~n37923 ;
  assign n37925 = ~x47 & ~n37924 ;
  assign n37926 = ~x47 & ~n37925 ;
  assign n37927 = ~n37924 & ~n37925 ;
  assign n37928 = ~n37926 & ~n37927 ;
  assign n37929 = n37917 & ~n37928 ;
  assign n37930 = n37917 & ~n37929 ;
  assign n37931 = ~n37928 & ~n37929 ;
  assign n37932 = ~n37930 & ~n37931 ;
  assign n37933 = ~n37810 & n37932 ;
  assign n37934 = n37810 & ~n37932 ;
  assign n37935 = ~n37933 & ~n37934 ;
  assign n37936 = ~x100 & n12506 ;
  assign n37937 = ~x98 & n13131 ;
  assign n37938 = ~x99 & n12501 ;
  assign n37939 = ~n37937 & ~n37938 ;
  assign n37940 = ~n37936 & n37939 ;
  assign n37941 = n9338 & n12509 ;
  assign n37942 = n37940 & ~n37941 ;
  assign n37943 = ~x44 & ~n37942 ;
  assign n37944 = ~x44 & ~n37943 ;
  assign n37945 = ~n37942 & ~n37943 ;
  assign n37946 = ~n37944 & ~n37945 ;
  assign n37947 = ~n37935 & ~n37946 ;
  assign n37948 = n37935 & n37946 ;
  assign n37949 = ~n37947 & ~n37948 ;
  assign n37950 = n37808 & ~n37949 ;
  assign n37951 = ~n37808 & n37949 ;
  assign n37952 = ~n37950 & ~n37951 ;
  assign n37953 = ~x103 & n10905 ;
  assign n37954 = ~x101 & n11466 ;
  assign n37955 = ~x102 & n10900 ;
  assign n37956 = ~n37954 & ~n37955 ;
  assign n37957 = ~n37953 & n37956 ;
  assign n37958 = n10833 & n10908 ;
  assign n37959 = n37957 & ~n37958 ;
  assign n37960 = ~x41 & ~n37959 ;
  assign n37961 = ~x41 & ~n37960 ;
  assign n37962 = ~n37959 & ~n37960 ;
  assign n37963 = ~n37961 & ~n37962 ;
  assign n37964 = n37952 & ~n37963 ;
  assign n37965 = n37952 & ~n37964 ;
  assign n37966 = ~n37963 & ~n37964 ;
  assign n37967 = ~n37965 & ~n37966 ;
  assign n37968 = ~n37807 & n37967 ;
  assign n37969 = n37807 & ~n37967 ;
  assign n37970 = ~n37968 & ~n37969 ;
  assign n37971 = ~x106 & n9433 ;
  assign n37972 = ~x104 & n9915 ;
  assign n37973 = ~x105 & n9428 ;
  assign n37974 = ~n37972 & ~n37973 ;
  assign n37975 = ~n37971 & n37974 ;
  assign n37976 = n9436 & n12447 ;
  assign n37977 = n37975 & ~n37976 ;
  assign n37978 = ~x38 & ~n37977 ;
  assign n37979 = ~x38 & ~n37978 ;
  assign n37980 = ~n37977 & ~n37978 ;
  assign n37981 = ~n37979 & ~n37980 ;
  assign n37982 = ~n37970 & ~n37981 ;
  assign n37983 = n37970 & n37981 ;
  assign n37984 = ~n37982 & ~n37983 ;
  assign n37985 = n37806 & ~n37984 ;
  assign n37986 = ~n37806 & n37984 ;
  assign n37987 = ~n37985 & ~n37986 ;
  assign n37988 = ~x109 & n8006 ;
  assign n37989 = ~x107 & n8474 ;
  assign n37990 = ~x108 & n8001 ;
  assign n37991 = ~n37989 & ~n37990 ;
  assign n37992 = ~n37988 & n37991 ;
  assign n37993 = n8009 & n14177 ;
  assign n37994 = n37992 & ~n37993 ;
  assign n37995 = ~x35 & ~n37994 ;
  assign n37996 = ~x35 & ~n37995 ;
  assign n37997 = ~n37994 & ~n37995 ;
  assign n37998 = ~n37996 & ~n37997 ;
  assign n37999 = n37987 & ~n37998 ;
  assign n38000 = n37987 & ~n37999 ;
  assign n38001 = ~n37998 & ~n37999 ;
  assign n38002 = ~n38000 & ~n38001 ;
  assign n38003 = ~n37330 & ~n37333 ;
  assign n38004 = n38002 & n38003 ;
  assign n38005 = ~n38002 & ~n38003 ;
  assign n38006 = ~n38004 & ~n38005 ;
  assign n38007 = ~n37146 & ~n37337 ;
  assign n38008 = ~x112 & n6725 ;
  assign n38009 = ~x110 & n7129 ;
  assign n38010 = ~x111 & n6720 ;
  assign n38011 = ~n38009 & ~n38010 ;
  assign n38012 = ~n38008 & n38011 ;
  assign n38013 = n6728 & n15744 ;
  assign n38014 = n38012 & ~n38013 ;
  assign n38015 = ~x32 & ~n38014 ;
  assign n38016 = ~x32 & ~n38015 ;
  assign n38017 = ~n38014 & ~n38015 ;
  assign n38018 = ~n38016 & ~n38017 ;
  assign n38019 = ~n38007 & ~n38018 ;
  assign n38020 = ~n38007 & ~n38019 ;
  assign n38021 = ~n38018 & ~n38019 ;
  assign n38022 = ~n38020 & ~n38021 ;
  assign n38023 = n38006 & ~n38022 ;
  assign n38024 = ~n38006 & n38022 ;
  assign n38025 = n37805 & ~n38024 ;
  assign n38026 = ~n38023 & n38025 ;
  assign n38027 = n37805 & ~n38026 ;
  assign n38028 = ~n38024 & ~n38026 ;
  assign n38029 = ~n38023 & n38028 ;
  assign n38030 = ~n38027 & ~n38029 ;
  assign n38031 = n37790 & ~n38030 ;
  assign n38032 = ~n37790 & n38030 ;
  assign n38033 = ~n37775 & ~n38032 ;
  assign n38034 = ~n38031 & n38033 ;
  assign n38035 = ~n37775 & ~n38034 ;
  assign n38036 = ~n38032 & ~n38034 ;
  assign n38037 = ~n38031 & n38036 ;
  assign n38038 = ~n38035 & ~n38037 ;
  assign n38039 = n37760 & ~n38038 ;
  assign n38040 = ~n37760 & n38038 ;
  assign n38041 = ~n37745 & ~n38040 ;
  assign n38042 = ~n38039 & n38041 ;
  assign n38043 = ~n37745 & ~n38042 ;
  assign n38044 = ~n38040 & ~n38042 ;
  assign n38045 = ~n38039 & n38044 ;
  assign n38046 = ~n38043 & ~n38045 ;
  assign n38047 = ~n37085 & ~n37392 ;
  assign n38048 = n38046 & n38047 ;
  assign n38049 = ~n38046 & ~n38047 ;
  assign n38050 = ~n38048 & ~n38049 ;
  assign n38051 = ~n37395 & ~n37398 ;
  assign n38052 = n38050 & ~n38051 ;
  assign n38053 = ~n38050 & n38051 ;
  assign n38054 = ~n38052 & ~n38053 ;
  assign n38057 = ~n38054 & ~x206 ;
  assign n38058 = ~n38056 & ~n38057 ;
  assign n38059 = ~n37434 & ~n37714 ;
  assign n38060 = x126 & n2275 ;
  assign n38061 = x127 & n2088 ;
  assign n38062 = ~n38060 & ~n38061 ;
  assign n38063 = ~n2096 & n38062 ;
  assign n38064 = n26965 & n38062 ;
  assign n38065 = ~n38063 & ~n38064 ;
  assign n38066 = x17 & ~n38065 ;
  assign n38067 = ~x17 & n38065 ;
  assign n38068 = ~n38066 & ~n38067 ;
  assign n38069 = ~n38059 & ~n38068 ;
  assign n38070 = n38059 & n38068 ;
  assign n38071 = ~n38069 & ~n38070 ;
  assign n38072 = x125 & n2751 ;
  assign n38073 = x123 & n3020 ;
  assign n38074 = x124 & n2746 ;
  assign n38075 = ~n38073 & ~n38074 ;
  assign n38076 = ~n38072 & n38075 ;
  assign n38077 = n2754 & n24935 ;
  assign n38078 = n38076 & ~n38077 ;
  assign n38079 = x20 & ~n38078 ;
  assign n38080 = x20 & ~n38079 ;
  assign n38081 = ~n38078 & ~n38079 ;
  assign n38082 = ~n38080 & ~n38081 ;
  assign n38083 = ~n37436 & ~n37447 ;
  assign n38084 = ~n37709 & ~n38083 ;
  assign n38085 = n38082 & n38084 ;
  assign n38086 = ~n38082 & ~n38084 ;
  assign n38087 = ~n38085 & ~n38086 ;
  assign n38088 = ~n37464 & ~n37706 ;
  assign n38089 = x122 & n3589 ;
  assign n38090 = x120 & n3878 ;
  assign n38091 = x121 & n3584 ;
  assign n38092 = ~n38090 & ~n38091 ;
  assign n38093 = ~n38089 & n38092 ;
  assign n38094 = ~n3592 & n38093 ;
  assign n38095 = ~n22622 & n38093 ;
  assign n38096 = ~n38094 & ~n38095 ;
  assign n38097 = x23 & ~n38096 ;
  assign n38098 = ~x23 & n38096 ;
  assign n38099 = ~n38097 & ~n38098 ;
  assign n38100 = ~n38088 & ~n38099 ;
  assign n38101 = n38088 & n38099 ;
  assign n38102 = ~n38100 & ~n38101 ;
  assign n38103 = x119 & n4531 ;
  assign n38104 = x117 & n4847 ;
  assign n38105 = x118 & n4526 ;
  assign n38106 = ~n38104 & ~n38105 ;
  assign n38107 = ~n38103 & n38106 ;
  assign n38108 = n4534 & n20423 ;
  assign n38109 = n38107 & ~n38108 ;
  assign n38110 = x26 & ~n38109 ;
  assign n38111 = x26 & ~n38110 ;
  assign n38112 = ~n38109 & ~n38110 ;
  assign n38113 = ~n38111 & ~n38112 ;
  assign n38114 = ~n37479 & ~n37701 ;
  assign n38115 = n38113 & n38114 ;
  assign n38116 = ~n38113 & ~n38114 ;
  assign n38117 = ~n38115 & ~n38116 ;
  assign n38118 = x116 & n5560 ;
  assign n38119 = x114 & n5943 ;
  assign n38120 = x115 & n5555 ;
  assign n38121 = ~n38119 & ~n38120 ;
  assign n38122 = ~n38118 & n38121 ;
  assign n38123 = n5563 & n18336 ;
  assign n38124 = n38122 & ~n38123 ;
  assign n38125 = x29 & ~n38124 ;
  assign n38126 = x29 & ~n38125 ;
  assign n38127 = ~n38124 & ~n38125 ;
  assign n38128 = ~n38126 & ~n38127 ;
  assign n38129 = ~n37694 & ~n37698 ;
  assign n38130 = ~n38128 & ~n38129 ;
  assign n38131 = ~n38128 & ~n38130 ;
  assign n38132 = ~n38129 & ~n38130 ;
  assign n38133 = ~n38131 & ~n38132 ;
  assign n38134 = x113 & n6725 ;
  assign n38135 = x111 & n7129 ;
  assign n38136 = x112 & n6720 ;
  assign n38137 = ~n38135 & ~n38136 ;
  assign n38138 = ~n38134 & n38137 ;
  assign n38139 = n6728 & n16361 ;
  assign n38140 = n38138 & ~n38139 ;
  assign n38141 = x32 & ~n38140 ;
  assign n38142 = x32 & ~n38141 ;
  assign n38143 = ~n38140 & ~n38141 ;
  assign n38144 = ~n38142 & ~n38143 ;
  assign n38145 = ~n37674 & ~n37680 ;
  assign n38146 = n38144 & n38145 ;
  assign n38147 = ~n38144 & ~n38145 ;
  assign n38148 = ~n38146 & ~n38147 ;
  assign n38149 = ~n37482 & ~n37642 ;
  assign n38150 = ~n37639 & ~n38149 ;
  assign n38151 = x104 & n10905 ;
  assign n38152 = x102 & n11466 ;
  assign n38153 = x103 & n10900 ;
  assign n38154 = ~n38152 & ~n38153 ;
  assign n38155 = ~n38151 & n38154 ;
  assign n38156 = n10908 & n11116 ;
  assign n38157 = n38155 & ~n38156 ;
  assign n38158 = x41 & ~n38157 ;
  assign n38159 = x41 & ~n38158 ;
  assign n38160 = ~n38157 & ~n38158 ;
  assign n38161 = ~n38159 & ~n38160 ;
  assign n38162 = ~n37622 & ~n37626 ;
  assign n38163 = x101 & n12506 ;
  assign n38164 = x99 & n13131 ;
  assign n38165 = x100 & n12501 ;
  assign n38166 = ~n38164 & ~n38165 ;
  assign n38167 = ~n38163 & n38166 ;
  assign n38168 = n9601 & n12509 ;
  assign n38169 = n38167 & ~n38168 ;
  assign n38170 = x44 & ~n38169 ;
  assign n38171 = x44 & ~n38170 ;
  assign n38172 = ~n38169 & ~n38170 ;
  assign n38173 = ~n38171 & ~n38172 ;
  assign n38174 = ~n37485 & ~n37607 ;
  assign n38175 = ~n37604 & ~n38174 ;
  assign n38176 = ~n37509 & ~n37515 ;
  assign n38177 = x79 & n27024 ;
  assign n38178 = x80 & ~n26217 ;
  assign n38179 = ~n38177 & ~n38178 ;
  assign n38180 = ~n37490 & ~n37494 ;
  assign n38181 = ~n38179 & n38180 ;
  assign n38182 = n38179 & ~n38180 ;
  assign n38183 = ~n38181 & ~n38182 ;
  assign n38184 = x83 & n24612 ;
  assign n38185 = x81 & n25390 ;
  assign n38186 = x82 & n24607 ;
  assign n38187 = ~n38185 & ~n38186 ;
  assign n38188 = ~n38184 & n38187 ;
  assign n38189 = ~n24615 & n38188 ;
  assign n38190 = ~n2843 & n38188 ;
  assign n38191 = ~n38189 & ~n38190 ;
  assign n38192 = x62 & ~n38191 ;
  assign n38193 = ~x62 & n38191 ;
  assign n38194 = ~n38192 & ~n38193 ;
  assign n38195 = n38183 & ~n38194 ;
  assign n38196 = ~n38183 & n38194 ;
  assign n38197 = ~n38195 & ~n38196 ;
  assign n38198 = ~n38176 & n38197 ;
  assign n38199 = n38176 & ~n38197 ;
  assign n38200 = ~n38198 & ~n38199 ;
  assign n38201 = x86 & n22325 ;
  assign n38202 = x84 & n23066 ;
  assign n38203 = x85 & n22320 ;
  assign n38204 = ~n38202 & ~n38203 ;
  assign n38205 = ~n38201 & n38204 ;
  assign n38206 = n3686 & n22328 ;
  assign n38207 = n38205 & ~n38206 ;
  assign n38208 = x59 & ~n38207 ;
  assign n38209 = x59 & ~n38208 ;
  assign n38210 = ~n38207 & ~n38208 ;
  assign n38211 = ~n38209 & ~n38210 ;
  assign n38212 = n38200 & ~n38211 ;
  assign n38213 = n38200 & ~n38212 ;
  assign n38214 = ~n38211 & ~n38212 ;
  assign n38215 = ~n38213 & ~n38214 ;
  assign n38216 = ~n37528 & ~n37534 ;
  assign n38217 = n38215 & n38216 ;
  assign n38218 = ~n38215 & ~n38216 ;
  assign n38219 = ~n38217 & ~n38218 ;
  assign n38220 = x89 & n20143 ;
  assign n38221 = x87 & n20854 ;
  assign n38222 = x88 & n20138 ;
  assign n38223 = ~n38221 & ~n38222 ;
  assign n38224 = ~n38220 & n38223 ;
  assign n38225 = n4488 & n20146 ;
  assign n38226 = n38224 & ~n38225 ;
  assign n38227 = x56 & ~n38226 ;
  assign n38228 = x56 & ~n38227 ;
  assign n38229 = ~n38226 & ~n38227 ;
  assign n38230 = ~n38228 & ~n38229 ;
  assign n38231 = n38219 & ~n38230 ;
  assign n38232 = n38219 & ~n38231 ;
  assign n38233 = ~n38230 & ~n38231 ;
  assign n38234 = ~n38232 & ~n38233 ;
  assign n38235 = ~n37552 & n38234 ;
  assign n38236 = n37552 & ~n38234 ;
  assign n38237 = ~n38235 & ~n38236 ;
  assign n38238 = x92 & n18025 ;
  assign n38239 = x90 & n18764 ;
  assign n38240 = x91 & n18020 ;
  assign n38241 = ~n38239 & ~n38240 ;
  assign n38242 = ~n38238 & n38241 ;
  assign n38243 = n5710 & n18028 ;
  assign n38244 = n38242 & ~n38243 ;
  assign n38245 = x53 & ~n38244 ;
  assign n38246 = x53 & ~n38245 ;
  assign n38247 = ~n38244 & ~n38245 ;
  assign n38248 = ~n38246 & ~n38247 ;
  assign n38249 = n38237 & n38248 ;
  assign n38250 = ~n38237 & ~n38248 ;
  assign n38251 = ~n38249 & ~n38250 ;
  assign n38252 = ~n37566 & ~n37572 ;
  assign n38253 = n38251 & ~n38252 ;
  assign n38254 = ~n38251 & n38252 ;
  assign n38255 = ~n38253 & ~n38254 ;
  assign n38256 = x95 & n16076 ;
  assign n38257 = x93 & n16756 ;
  assign n38258 = x94 & n16071 ;
  assign n38259 = ~n38257 & ~n38258 ;
  assign n38260 = ~n38256 & n38259 ;
  assign n38261 = n6894 & n16079 ;
  assign n38262 = n38260 & ~n38261 ;
  assign n38263 = x50 & ~n38262 ;
  assign n38264 = x50 & ~n38263 ;
  assign n38265 = ~n38262 & ~n38263 ;
  assign n38266 = ~n38264 & ~n38265 ;
  assign n38267 = n38255 & ~n38266 ;
  assign n38268 = n38255 & ~n38267 ;
  assign n38269 = ~n38266 & ~n38267 ;
  assign n38270 = ~n38268 & ~n38269 ;
  assign n38271 = ~n37585 & ~n37591 ;
  assign n38272 = n38270 & n38271 ;
  assign n38273 = ~n38270 & ~n38271 ;
  assign n38274 = ~n38272 & ~n38273 ;
  assign n38275 = x98 & n14233 ;
  assign n38276 = x96 & n14876 ;
  assign n38277 = x97 & n14228 ;
  assign n38278 = ~n38276 & ~n38277 ;
  assign n38279 = ~n38275 & n38278 ;
  assign n38280 = n8196 & n14236 ;
  assign n38281 = n38279 & ~n38280 ;
  assign n38282 = x47 & ~n38281 ;
  assign n38283 = x47 & ~n38282 ;
  assign n38284 = ~n38281 & ~n38282 ;
  assign n38285 = ~n38283 & ~n38284 ;
  assign n38286 = ~n38274 & n38285 ;
  assign n38287 = n38274 & ~n38285 ;
  assign n38288 = ~n38286 & ~n38287 ;
  assign n38289 = ~n38175 & n38288 ;
  assign n38290 = ~n38175 & ~n38289 ;
  assign n38291 = n38288 & ~n38289 ;
  assign n38292 = ~n38290 & ~n38291 ;
  assign n38293 = ~n38173 & ~n38292 ;
  assign n38294 = n38173 & ~n38291 ;
  assign n38295 = ~n38290 & n38294 ;
  assign n38296 = ~n38293 & ~n38295 ;
  assign n38297 = ~n38162 & n38296 ;
  assign n38298 = ~n38162 & ~n38297 ;
  assign n38299 = n38296 & ~n38297 ;
  assign n38300 = ~n38298 & ~n38299 ;
  assign n38301 = ~n38161 & ~n38300 ;
  assign n38302 = n38161 & ~n38299 ;
  assign n38303 = ~n38298 & n38302 ;
  assign n38304 = ~n38301 & ~n38303 ;
  assign n38305 = ~n38150 & n38304 ;
  assign n38306 = n38150 & ~n38304 ;
  assign n38307 = ~n38305 & ~n38306 ;
  assign n38308 = x107 & n9433 ;
  assign n38309 = x105 & n9915 ;
  assign n38310 = x106 & n9428 ;
  assign n38311 = ~n38309 & ~n38310 ;
  assign n38312 = ~n38308 & n38311 ;
  assign n38313 = n9436 & n12749 ;
  assign n38314 = n38312 & ~n38313 ;
  assign n38315 = x38 & ~n38314 ;
  assign n38316 = x38 & ~n38315 ;
  assign n38317 = ~n38314 & ~n38315 ;
  assign n38318 = ~n38316 & ~n38317 ;
  assign n38319 = n38307 & ~n38318 ;
  assign n38320 = n38307 & ~n38319 ;
  assign n38321 = ~n38318 & ~n38319 ;
  assign n38322 = ~n38320 & ~n38321 ;
  assign n38323 = ~n37657 & ~n37661 ;
  assign n38324 = n38322 & n38323 ;
  assign n38325 = ~n38322 & ~n38323 ;
  assign n38326 = ~n38324 & ~n38325 ;
  assign n38327 = x110 & n8006 ;
  assign n38328 = x108 & n8474 ;
  assign n38329 = x109 & n8001 ;
  assign n38330 = ~n38328 & ~n38329 ;
  assign n38331 = ~n38327 & n38330 ;
  assign n38332 = n8009 & n14497 ;
  assign n38333 = n38331 & ~n38332 ;
  assign n38334 = x35 & ~n38333 ;
  assign n38335 = x35 & ~n38334 ;
  assign n38336 = ~n38333 & ~n38334 ;
  assign n38337 = ~n38335 & ~n38336 ;
  assign n38338 = n38326 & ~n38337 ;
  assign n38339 = n38326 & ~n38338 ;
  assign n38340 = ~n38337 & ~n38338 ;
  assign n38341 = ~n38339 & ~n38340 ;
  assign n38342 = n38148 & ~n38341 ;
  assign n38343 = ~n38148 & n38341 ;
  assign n38344 = ~n38133 & ~n38343 ;
  assign n38345 = ~n38342 & n38344 ;
  assign n38346 = ~n38133 & ~n38345 ;
  assign n38347 = ~n38343 & ~n38345 ;
  assign n38348 = ~n38342 & n38347 ;
  assign n38349 = ~n38346 & ~n38348 ;
  assign n38350 = n38117 & ~n38349 ;
  assign n38351 = ~n38117 & n38349 ;
  assign n38352 = n38102 & ~n38351 ;
  assign n38353 = ~n38350 & n38352 ;
  assign n38354 = n38102 & ~n38353 ;
  assign n38355 = ~n38351 & ~n38353 ;
  assign n38356 = ~n38350 & n38355 ;
  assign n38357 = ~n38354 & ~n38356 ;
  assign n38358 = n38087 & ~n38357 ;
  assign n38359 = ~n38087 & n38357 ;
  assign n38360 = n38071 & ~n38359 ;
  assign n38361 = ~n38358 & n38360 ;
  assign n38362 = n38071 & ~n38361 ;
  assign n38363 = ~n38359 & ~n38361 ;
  assign n38364 = ~n38358 & n38363 ;
  assign n38365 = ~n38362 & ~n38364 ;
  assign n38366 = ~n37417 & ~n37717 ;
  assign n38367 = n38365 & n38366 ;
  assign n38368 = ~n38365 & ~n38366 ;
  assign n38369 = ~n38367 & ~n38368 ;
  assign n38370 = ~n37724 & ~n37727 ;
  assign n38371 = n38369 & ~n38370 ;
  assign n38372 = ~n38369 & n38370 ;
  assign n38373 = ~n38371 & ~n38372 ;
  assign n38690 = n38373 & x207 ;
  assign n38374 = ~n37759 & ~n38039 ;
  assign n38375 = ~x126 & n2275 ;
  assign n38376 = ~x127 & n2088 ;
  assign n38377 = ~n38375 & ~n38376 ;
  assign n38378 = ~n2096 & n38377 ;
  assign n38379 = n27368 & n38377 ;
  assign n38380 = ~n38378 & ~n38379 ;
  assign n38381 = ~x17 & ~n38380 ;
  assign n38382 = x17 & n38380 ;
  assign n38383 = ~n38381 & ~n38382 ;
  assign n38384 = ~n38374 & ~n38383 ;
  assign n38385 = n38374 & n38383 ;
  assign n38386 = ~n38384 & ~n38385 ;
  assign n38387 = ~x125 & n2751 ;
  assign n38388 = ~x123 & n3020 ;
  assign n38389 = ~x124 & n2746 ;
  assign n38390 = ~n38388 & ~n38389 ;
  assign n38391 = ~n38387 & n38390 ;
  assign n38392 = n2754 & n25330 ;
  assign n38393 = n38391 & ~n38392 ;
  assign n38394 = ~x20 & ~n38393 ;
  assign n38395 = ~x20 & ~n38394 ;
  assign n38396 = ~n38393 & ~n38394 ;
  assign n38397 = ~n38395 & ~n38396 ;
  assign n38398 = ~n37761 & ~n37772 ;
  assign n38399 = ~n38034 & ~n38398 ;
  assign n38400 = n38397 & n38399 ;
  assign n38401 = ~n38397 & ~n38399 ;
  assign n38402 = ~n38400 & ~n38401 ;
  assign n38403 = ~n37789 & ~n38031 ;
  assign n38404 = ~x122 & n3589 ;
  assign n38405 = ~x120 & n3878 ;
  assign n38406 = ~x121 & n3584 ;
  assign n38407 = ~n38405 & ~n38406 ;
  assign n38408 = ~n38404 & n38407 ;
  assign n38409 = ~n3592 & n38408 ;
  assign n38410 = ~n22998 & n38408 ;
  assign n38411 = ~n38409 & ~n38410 ;
  assign n38412 = ~x23 & ~n38411 ;
  assign n38413 = x23 & n38411 ;
  assign n38414 = ~n38412 & ~n38413 ;
  assign n38415 = ~n38403 & ~n38414 ;
  assign n38416 = n38403 & n38414 ;
  assign n38417 = ~n38415 & ~n38416 ;
  assign n38418 = ~x119 & n4531 ;
  assign n38419 = ~x117 & n4847 ;
  assign n38420 = ~x118 & n4526 ;
  assign n38421 = ~n38419 & ~n38420 ;
  assign n38422 = ~n38418 & n38421 ;
  assign n38423 = n4534 & n20778 ;
  assign n38424 = n38422 & ~n38423 ;
  assign n38425 = ~x26 & ~n38424 ;
  assign n38426 = ~x26 & ~n38425 ;
  assign n38427 = ~n38424 & ~n38425 ;
  assign n38428 = ~n38426 & ~n38427 ;
  assign n38429 = ~n37804 & ~n38026 ;
  assign n38430 = n38428 & n38429 ;
  assign n38431 = ~n38428 & ~n38429 ;
  assign n38432 = ~n38430 & ~n38431 ;
  assign n38433 = ~x116 & n5560 ;
  assign n38434 = ~x114 & n5943 ;
  assign n38435 = ~x115 & n5555 ;
  assign n38436 = ~n38434 & ~n38435 ;
  assign n38437 = ~n38433 & n38436 ;
  assign n38438 = n5563 & n18678 ;
  assign n38439 = n38437 & ~n38438 ;
  assign n38440 = ~x29 & ~n38439 ;
  assign n38441 = ~x29 & ~n38440 ;
  assign n38442 = ~n38439 & ~n38440 ;
  assign n38443 = ~n38441 & ~n38442 ;
  assign n38444 = ~n38019 & ~n38023 ;
  assign n38445 = ~n38443 & ~n38444 ;
  assign n38446 = ~n38443 & ~n38445 ;
  assign n38447 = ~n38444 & ~n38445 ;
  assign n38448 = ~n38446 & ~n38447 ;
  assign n38449 = ~x113 & n6725 ;
  assign n38450 = ~x111 & n7129 ;
  assign n38451 = ~x112 & n6720 ;
  assign n38452 = ~n38450 & ~n38451 ;
  assign n38453 = ~n38449 & n38452 ;
  assign n38454 = n6728 & n16684 ;
  assign n38455 = n38453 & ~n38454 ;
  assign n38456 = ~x32 & ~n38455 ;
  assign n38457 = ~x32 & ~n38456 ;
  assign n38458 = ~n38455 & ~n38456 ;
  assign n38459 = ~n38457 & ~n38458 ;
  assign n38460 = ~n37999 & ~n38005 ;
  assign n38461 = n38459 & n38460 ;
  assign n38462 = ~n38459 & ~n38460 ;
  assign n38463 = ~n38461 & ~n38462 ;
  assign n38464 = ~n37807 & ~n37967 ;
  assign n38465 = ~n37964 & ~n38464 ;
  assign n38466 = ~x104 & n10905 ;
  assign n38467 = ~x102 & n11466 ;
  assign n38468 = ~x103 & n10900 ;
  assign n38469 = ~n38467 & ~n38468 ;
  assign n38470 = ~n38466 & n38469 ;
  assign n38471 = n10908 & n11380 ;
  assign n38472 = n38470 & ~n38471 ;
  assign n38473 = ~x41 & ~n38472 ;
  assign n38474 = ~x41 & ~n38473 ;
  assign n38475 = ~n38472 & ~n38473 ;
  assign n38476 = ~n38474 & ~n38475 ;
  assign n38477 = ~n37947 & ~n37951 ;
  assign n38478 = ~x101 & n12506 ;
  assign n38479 = ~x99 & n13131 ;
  assign n38480 = ~x100 & n12501 ;
  assign n38481 = ~n38479 & ~n38480 ;
  assign n38482 = ~n38478 & n38481 ;
  assign n38483 = n9844 & n12509 ;
  assign n38484 = n38482 & ~n38483 ;
  assign n38485 = ~x44 & ~n38484 ;
  assign n38486 = ~x44 & ~n38485 ;
  assign n38487 = ~n38484 & ~n38485 ;
  assign n38488 = ~n38486 & ~n38487 ;
  assign n38489 = ~n37810 & ~n37932 ;
  assign n38490 = ~n37929 & ~n38489 ;
  assign n38491 = ~n37834 & ~n37840 ;
  assign n38492 = ~x79 & n27427 ;
  assign n38493 = ~x80 & ~n26217 ;
  assign n38494 = ~n38492 & ~n38493 ;
  assign n38495 = ~n37815 & ~n37819 ;
  assign n38496 = ~n38494 & n38495 ;
  assign n38497 = n38494 & ~n38495 ;
  assign n38498 = ~n38496 & ~n38497 ;
  assign n38499 = ~x83 & n24612 ;
  assign n38500 = ~x81 & n25390 ;
  assign n38501 = ~x82 & n24607 ;
  assign n38502 = ~n38500 & ~n38501 ;
  assign n38503 = ~n38499 & n38502 ;
  assign n38504 = ~n24615 & n38503 ;
  assign n38505 = ~n2972 & n38503 ;
  assign n38506 = ~n38504 & ~n38505 ;
  assign n38507 = ~x62 & ~n38506 ;
  assign n38508 = x62 & n38506 ;
  assign n38509 = ~n38507 & ~n38508 ;
  assign n38510 = n38498 & ~n38509 ;
  assign n38511 = ~n38498 & n38509 ;
  assign n38512 = ~n38510 & ~n38511 ;
  assign n38513 = ~n38491 & n38512 ;
  assign n38514 = n38491 & ~n38512 ;
  assign n38515 = ~n38513 & ~n38514 ;
  assign n38516 = ~x86 & n22325 ;
  assign n38517 = ~x84 & n23066 ;
  assign n38518 = ~x85 & n22320 ;
  assign n38519 = ~n38517 & ~n38518 ;
  assign n38520 = ~n38516 & n38519 ;
  assign n38521 = n3832 & n22328 ;
  assign n38522 = n38520 & ~n38521 ;
  assign n38523 = ~x59 & ~n38522 ;
  assign n38524 = ~x59 & ~n38523 ;
  assign n38525 = ~n38522 & ~n38523 ;
  assign n38526 = ~n38524 & ~n38525 ;
  assign n38527 = n38515 & ~n38526 ;
  assign n38528 = n38515 & ~n38527 ;
  assign n38529 = ~n38526 & ~n38527 ;
  assign n38530 = ~n38528 & ~n38529 ;
  assign n38531 = ~n37853 & ~n37859 ;
  assign n38532 = n38530 & n38531 ;
  assign n38533 = ~n38530 & ~n38531 ;
  assign n38534 = ~n38532 & ~n38533 ;
  assign n38535 = ~x89 & n20143 ;
  assign n38536 = ~x87 & n20854 ;
  assign n38537 = ~x88 & n20138 ;
  assign n38538 = ~n38536 & ~n38537 ;
  assign n38539 = ~n38535 & n38538 ;
  assign n38540 = n4664 & n20146 ;
  assign n38541 = n38539 & ~n38540 ;
  assign n38542 = ~x56 & ~n38541 ;
  assign n38543 = ~x56 & ~n38542 ;
  assign n38544 = ~n38541 & ~n38542 ;
  assign n38545 = ~n38543 & ~n38544 ;
  assign n38546 = n38534 & ~n38545 ;
  assign n38547 = n38534 & ~n38546 ;
  assign n38548 = ~n38545 & ~n38546 ;
  assign n38549 = ~n38547 & ~n38548 ;
  assign n38550 = ~n37877 & n38549 ;
  assign n38551 = n37877 & ~n38549 ;
  assign n38552 = ~n38550 & ~n38551 ;
  assign n38553 = ~x92 & n18025 ;
  assign n38554 = ~x90 & n18764 ;
  assign n38555 = ~x91 & n18020 ;
  assign n38556 = ~n38554 & ~n38555 ;
  assign n38557 = ~n38553 & n38556 ;
  assign n38558 = n5896 & n18028 ;
  assign n38559 = n38557 & ~n38558 ;
  assign n38560 = ~x53 & ~n38559 ;
  assign n38561 = ~x53 & ~n38560 ;
  assign n38562 = ~n38559 & ~n38560 ;
  assign n38563 = ~n38561 & ~n38562 ;
  assign n38564 = n38552 & n38563 ;
  assign n38565 = ~n38552 & ~n38563 ;
  assign n38566 = ~n38564 & ~n38565 ;
  assign n38567 = ~n37891 & ~n37897 ;
  assign n38568 = n38566 & ~n38567 ;
  assign n38569 = ~n38566 & n38567 ;
  assign n38570 = ~n38568 & ~n38569 ;
  assign n38571 = ~x95 & n16076 ;
  assign n38572 = ~x93 & n16756 ;
  assign n38573 = ~x94 & n16071 ;
  assign n38574 = ~n38572 & ~n38573 ;
  assign n38575 = ~n38571 & n38574 ;
  assign n38576 = n7100 & n16079 ;
  assign n38577 = n38575 & ~n38576 ;
  assign n38578 = ~x50 & ~n38577 ;
  assign n38579 = ~x50 & ~n38578 ;
  assign n38580 = ~n38577 & ~n38578 ;
  assign n38581 = ~n38579 & ~n38580 ;
  assign n38582 = n38570 & ~n38581 ;
  assign n38583 = n38570 & ~n38582 ;
  assign n38584 = ~n38581 & ~n38582 ;
  assign n38585 = ~n38583 & ~n38584 ;
  assign n38586 = ~n37910 & ~n37916 ;
  assign n38587 = n38585 & n38586 ;
  assign n38588 = ~n38585 & ~n38586 ;
  assign n38589 = ~n38587 & ~n38588 ;
  assign n38590 = ~x98 & n14233 ;
  assign n38591 = ~x96 & n14876 ;
  assign n38592 = ~x97 & n14228 ;
  assign n38593 = ~n38591 & ~n38592 ;
  assign n38594 = ~n38590 & n38593 ;
  assign n38595 = n8426 & n14236 ;
  assign n38596 = n38594 & ~n38595 ;
  assign n38597 = ~x47 & ~n38596 ;
  assign n38598 = ~x47 & ~n38597 ;
  assign n38599 = ~n38596 & ~n38597 ;
  assign n38600 = ~n38598 & ~n38599 ;
  assign n38601 = ~n38589 & n38600 ;
  assign n38602 = n38589 & ~n38600 ;
  assign n38603 = ~n38601 & ~n38602 ;
  assign n38604 = ~n38490 & n38603 ;
  assign n38605 = ~n38490 & ~n38604 ;
  assign n38606 = n38603 & ~n38604 ;
  assign n38607 = ~n38605 & ~n38606 ;
  assign n38608 = ~n38488 & ~n38607 ;
  assign n38609 = n38488 & ~n38606 ;
  assign n38610 = ~n38605 & n38609 ;
  assign n38611 = ~n38608 & ~n38610 ;
  assign n38612 = ~n38477 & n38611 ;
  assign n38613 = ~n38477 & ~n38612 ;
  assign n38614 = n38611 & ~n38612 ;
  assign n38615 = ~n38613 & ~n38614 ;
  assign n38616 = ~n38476 & ~n38615 ;
  assign n38617 = n38476 & ~n38614 ;
  assign n38618 = ~n38613 & n38617 ;
  assign n38619 = ~n38616 & ~n38618 ;
  assign n38620 = ~n38465 & n38619 ;
  assign n38621 = n38465 & ~n38619 ;
  assign n38622 = ~n38620 & ~n38621 ;
  assign n38623 = ~x107 & n9433 ;
  assign n38624 = ~x105 & n9915 ;
  assign n38625 = ~x106 & n9428 ;
  assign n38626 = ~n38624 & ~n38625 ;
  assign n38627 = ~n38623 & n38626 ;
  assign n38628 = n9436 & n13034 ;
  assign n38629 = n38627 & ~n38628 ;
  assign n38630 = ~x38 & ~n38629 ;
  assign n38631 = ~x38 & ~n38630 ;
  assign n38632 = ~n38629 & ~n38630 ;
  assign n38633 = ~n38631 & ~n38632 ;
  assign n38634 = n38622 & ~n38633 ;
  assign n38635 = n38622 & ~n38634 ;
  assign n38636 = ~n38633 & ~n38634 ;
  assign n38637 = ~n38635 & ~n38636 ;
  assign n38638 = ~n37982 & ~n37986 ;
  assign n38639 = n38637 & n38638 ;
  assign n38640 = ~n38637 & ~n38638 ;
  assign n38641 = ~n38639 & ~n38640 ;
  assign n38642 = ~x110 & n8006 ;
  assign n38643 = ~x108 & n8474 ;
  assign n38644 = ~x109 & n8001 ;
  assign n38645 = ~n38643 & ~n38644 ;
  assign n38646 = ~n38642 & n38645 ;
  assign n38647 = n8009 & n14802 ;
  assign n38648 = n38646 & ~n38647 ;
  assign n38649 = ~x35 & ~n38648 ;
  assign n38650 = ~x35 & ~n38649 ;
  assign n38651 = ~n38648 & ~n38649 ;
  assign n38652 = ~n38650 & ~n38651 ;
  assign n38653 = n38641 & ~n38652 ;
  assign n38654 = n38641 & ~n38653 ;
  assign n38655 = ~n38652 & ~n38653 ;
  assign n38656 = ~n38654 & ~n38655 ;
  assign n38657 = n38463 & ~n38656 ;
  assign n38658 = ~n38463 & n38656 ;
  assign n38659 = ~n38448 & ~n38658 ;
  assign n38660 = ~n38657 & n38659 ;
  assign n38661 = ~n38448 & ~n38660 ;
  assign n38662 = ~n38658 & ~n38660 ;
  assign n38663 = ~n38657 & n38662 ;
  assign n38664 = ~n38661 & ~n38663 ;
  assign n38665 = n38432 & ~n38664 ;
  assign n38666 = ~n38432 & n38664 ;
  assign n38667 = n38417 & ~n38666 ;
  assign n38668 = ~n38665 & n38667 ;
  assign n38669 = n38417 & ~n38668 ;
  assign n38670 = ~n38666 & ~n38668 ;
  assign n38671 = ~n38665 & n38670 ;
  assign n38672 = ~n38669 & ~n38671 ;
  assign n38673 = n38402 & ~n38672 ;
  assign n38674 = ~n38402 & n38672 ;
  assign n38675 = n38386 & ~n38674 ;
  assign n38676 = ~n38673 & n38675 ;
  assign n38677 = n38386 & ~n38676 ;
  assign n38678 = ~n38674 & ~n38676 ;
  assign n38679 = ~n38673 & n38678 ;
  assign n38680 = ~n38677 & ~n38679 ;
  assign n38681 = ~n37742 & ~n38042 ;
  assign n38682 = n38680 & n38681 ;
  assign n38683 = ~n38680 & ~n38681 ;
  assign n38684 = ~n38682 & ~n38683 ;
  assign n38685 = ~n38049 & ~n38052 ;
  assign n38686 = n38684 & ~n38685 ;
  assign n38687 = ~n38684 & n38685 ;
  assign n38688 = ~n38686 & ~n38687 ;
  assign n38691 = ~n38688 & ~x207 ;
  assign n38692 = ~n38690 & ~n38691 ;
  assign n38693 = ~n38368 & ~n38371 ;
  assign n38694 = ~n38069 & ~n38361 ;
  assign n38695 = ~n38086 & ~n38358 ;
  assign n38696 = x127 & n2275 ;
  assign n38697 = n2096 & n26962 ;
  assign n38698 = ~n38696 & ~n38697 ;
  assign n38699 = x17 & ~n38698 ;
  assign n38700 = x17 & ~n38699 ;
  assign n38701 = ~n38698 & ~n38699 ;
  assign n38702 = ~n38700 & ~n38701 ;
  assign n38703 = ~n38695 & ~n38702 ;
  assign n38704 = ~n38695 & ~n38703 ;
  assign n38705 = ~n38702 & ~n38703 ;
  assign n38706 = ~n38704 & ~n38705 ;
  assign n38707 = x126 & n2751 ;
  assign n38708 = x124 & n3020 ;
  assign n38709 = x125 & n2746 ;
  assign n38710 = ~n38708 & ~n38709 ;
  assign n38711 = ~n38707 & n38710 ;
  assign n38712 = n2754 & n25735 ;
  assign n38713 = n38711 & ~n38712 ;
  assign n38714 = x20 & ~n38713 ;
  assign n38715 = x20 & ~n38714 ;
  assign n38716 = ~n38713 & ~n38714 ;
  assign n38717 = ~n38715 & ~n38716 ;
  assign n38718 = ~n38100 & ~n38353 ;
  assign n38719 = n38717 & n38718 ;
  assign n38720 = ~n38717 & ~n38718 ;
  assign n38721 = ~n38719 & ~n38720 ;
  assign n38722 = x123 & n3589 ;
  assign n38723 = x121 & n3878 ;
  assign n38724 = x122 & n3584 ;
  assign n38725 = ~n38723 & ~n38724 ;
  assign n38726 = ~n38722 & n38725 ;
  assign n38727 = n3592 & n23382 ;
  assign n38728 = n38726 & ~n38727 ;
  assign n38729 = x23 & ~n38728 ;
  assign n38730 = x23 & ~n38729 ;
  assign n38731 = ~n38728 & ~n38729 ;
  assign n38732 = ~n38730 & ~n38731 ;
  assign n38733 = ~n38116 & ~n38350 ;
  assign n38734 = ~n38732 & ~n38733 ;
  assign n38735 = ~n38732 & ~n38734 ;
  assign n38736 = ~n38733 & ~n38734 ;
  assign n38737 = ~n38735 & ~n38736 ;
  assign n38738 = x120 & n4531 ;
  assign n38739 = x118 & n4847 ;
  assign n38740 = x119 & n4526 ;
  assign n38741 = ~n38739 & ~n38740 ;
  assign n38742 = ~n38738 & n38741 ;
  assign n38743 = n4534 & n21143 ;
  assign n38744 = n38742 & ~n38743 ;
  assign n38745 = x26 & ~n38744 ;
  assign n38746 = x26 & ~n38745 ;
  assign n38747 = ~n38744 & ~n38745 ;
  assign n38748 = ~n38746 & ~n38747 ;
  assign n38749 = ~n38130 & ~n38345 ;
  assign n38750 = n38748 & n38749 ;
  assign n38751 = ~n38748 & ~n38749 ;
  assign n38752 = ~n38750 & ~n38751 ;
  assign n38753 = x117 & n5560 ;
  assign n38754 = x115 & n5943 ;
  assign n38755 = x116 & n5555 ;
  assign n38756 = ~n38754 & ~n38755 ;
  assign n38757 = ~n38753 & n38756 ;
  assign n38758 = n5563 & n19026 ;
  assign n38759 = n38757 & ~n38758 ;
  assign n38760 = x29 & ~n38759 ;
  assign n38761 = x29 & ~n38760 ;
  assign n38762 = ~n38759 & ~n38760 ;
  assign n38763 = ~n38761 & ~n38762 ;
  assign n38764 = ~n38147 & ~n38342 ;
  assign n38765 = ~n38763 & ~n38764 ;
  assign n38766 = ~n38763 & ~n38765 ;
  assign n38767 = ~n38764 & ~n38765 ;
  assign n38768 = ~n38766 & ~n38767 ;
  assign n38769 = x114 & n6725 ;
  assign n38770 = x112 & n7129 ;
  assign n38771 = x113 & n6720 ;
  assign n38772 = ~n38770 & ~n38771 ;
  assign n38773 = ~n38769 & n38772 ;
  assign n38774 = n6728 & n17012 ;
  assign n38775 = n38773 & ~n38774 ;
  assign n38776 = x32 & ~n38775 ;
  assign n38777 = x32 & ~n38776 ;
  assign n38778 = ~n38775 & ~n38776 ;
  assign n38779 = ~n38777 & ~n38778 ;
  assign n38780 = ~n38325 & ~n38338 ;
  assign n38781 = n38779 & n38780 ;
  assign n38782 = ~n38779 & ~n38780 ;
  assign n38783 = ~n38781 & ~n38782 ;
  assign n38784 = ~n38305 & ~n38319 ;
  assign n38785 = x108 & n9433 ;
  assign n38786 = x106 & n9915 ;
  assign n38787 = x107 & n9428 ;
  assign n38788 = ~n38786 & ~n38787 ;
  assign n38789 = ~n38785 & n38788 ;
  assign n38790 = n9436 & n13323 ;
  assign n38791 = n38789 & ~n38790 ;
  assign n38792 = x38 & ~n38791 ;
  assign n38793 = x38 & ~n38792 ;
  assign n38794 = ~n38791 & ~n38792 ;
  assign n38795 = ~n38793 & ~n38794 ;
  assign n38796 = ~n38297 & ~n38301 ;
  assign n38797 = x105 & n10905 ;
  assign n38798 = x103 & n11466 ;
  assign n38799 = x104 & n10900 ;
  assign n38800 = ~n38798 & ~n38799 ;
  assign n38801 = ~n38797 & n38800 ;
  assign n38802 = n10908 & n11648 ;
  assign n38803 = n38801 & ~n38802 ;
  assign n38804 = x41 & ~n38803 ;
  assign n38805 = x41 & ~n38804 ;
  assign n38806 = ~n38803 & ~n38804 ;
  assign n38807 = ~n38805 & ~n38806 ;
  assign n38808 = ~n38289 & ~n38293 ;
  assign n38809 = ~n38218 & ~n38231 ;
  assign n38810 = x90 & n20143 ;
  assign n38811 = x88 & n20854 ;
  assign n38812 = x89 & n20138 ;
  assign n38813 = ~n38811 & ~n38812 ;
  assign n38814 = ~n38810 & n38813 ;
  assign n38815 = n4986 & n20146 ;
  assign n38816 = n38814 & ~n38815 ;
  assign n38817 = x56 & ~n38816 ;
  assign n38818 = x56 & ~n38817 ;
  assign n38819 = ~n38816 & ~n38817 ;
  assign n38820 = ~n38818 & ~n38819 ;
  assign n38821 = ~n38198 & ~n38212 ;
  assign n38822 = x84 & n24612 ;
  assign n38823 = x82 & n25390 ;
  assign n38824 = x83 & n24607 ;
  assign n38825 = ~n38823 & ~n38824 ;
  assign n38826 = ~n38822 & n38825 ;
  assign n38827 = n3114 & n24615 ;
  assign n38828 = n38826 & ~n38827 ;
  assign n38829 = x62 & ~n38828 ;
  assign n38830 = x62 & ~n38829 ;
  assign n38831 = ~n38828 & ~n38829 ;
  assign n38832 = ~n38830 & ~n38831 ;
  assign n38833 = x80 & n27024 ;
  assign n38834 = x81 & ~n26217 ;
  assign n38835 = ~n38833 & ~n38834 ;
  assign n38836 = n38179 & ~n38835 ;
  assign n38837 = ~n38179 & n38835 ;
  assign n38838 = ~n38832 & ~n38837 ;
  assign n38839 = ~n38836 & n38838 ;
  assign n38840 = ~n38832 & ~n38839 ;
  assign n38841 = ~n38837 & ~n38839 ;
  assign n38842 = ~n38836 & n38841 ;
  assign n38843 = ~n38840 & ~n38842 ;
  assign n38844 = ~n38182 & ~n38195 ;
  assign n38845 = n38843 & n38844 ;
  assign n38846 = ~n38843 & ~n38844 ;
  assign n38847 = ~n38845 & ~n38846 ;
  assign n38848 = x87 & n22325 ;
  assign n38849 = x85 & n23066 ;
  assign n38850 = x86 & n22320 ;
  assign n38851 = ~n38849 & ~n38850 ;
  assign n38852 = ~n38848 & n38851 ;
  assign n38853 = n3991 & n22328 ;
  assign n38854 = n38852 & ~n38853 ;
  assign n38855 = x59 & ~n38854 ;
  assign n38856 = x59 & ~n38855 ;
  assign n38857 = ~n38854 & ~n38855 ;
  assign n38858 = ~n38856 & ~n38857 ;
  assign n38859 = ~n38847 & n38858 ;
  assign n38860 = n38847 & ~n38858 ;
  assign n38861 = ~n38859 & ~n38860 ;
  assign n38862 = ~n38821 & n38861 ;
  assign n38863 = n38821 & ~n38861 ;
  assign n38864 = ~n38862 & ~n38863 ;
  assign n38865 = ~n38820 & n38864 ;
  assign n38866 = n38820 & ~n38864 ;
  assign n38867 = ~n38865 & ~n38866 ;
  assign n38868 = ~n38809 & n38867 ;
  assign n38869 = n38809 & ~n38867 ;
  assign n38870 = ~n38868 & ~n38869 ;
  assign n38871 = x93 & n18025 ;
  assign n38872 = x91 & n18764 ;
  assign n38873 = x92 & n18020 ;
  assign n38874 = ~n38872 & ~n38873 ;
  assign n38875 = ~n38871 & n38874 ;
  assign n38876 = n6094 & n18028 ;
  assign n38877 = n38875 & ~n38876 ;
  assign n38878 = x53 & ~n38877 ;
  assign n38879 = x53 & ~n38878 ;
  assign n38880 = ~n38877 & ~n38878 ;
  assign n38881 = ~n38879 & ~n38880 ;
  assign n38882 = n38870 & ~n38881 ;
  assign n38883 = n38870 & ~n38882 ;
  assign n38884 = ~n38881 & ~n38882 ;
  assign n38885 = ~n38883 & ~n38884 ;
  assign n38886 = ~n37552 & ~n38234 ;
  assign n38887 = ~n38250 & ~n38886 ;
  assign n38888 = ~n38885 & ~n38887 ;
  assign n38889 = ~n38885 & ~n38888 ;
  assign n38890 = ~n38887 & ~n38888 ;
  assign n38891 = ~n38889 & ~n38890 ;
  assign n38892 = x96 & n16076 ;
  assign n38893 = x94 & n16756 ;
  assign n38894 = x95 & n16071 ;
  assign n38895 = ~n38893 & ~n38894 ;
  assign n38896 = ~n38892 & n38895 ;
  assign n38897 = n7321 & n16079 ;
  assign n38898 = n38896 & ~n38897 ;
  assign n38899 = x50 & ~n38898 ;
  assign n38900 = x50 & ~n38899 ;
  assign n38901 = ~n38898 & ~n38899 ;
  assign n38902 = ~n38900 & ~n38901 ;
  assign n38903 = ~n38891 & n38902 ;
  assign n38904 = n38891 & ~n38902 ;
  assign n38905 = ~n38903 & ~n38904 ;
  assign n38906 = ~n38253 & ~n38267 ;
  assign n38907 = n38905 & n38906 ;
  assign n38908 = ~n38905 & ~n38906 ;
  assign n38909 = ~n38907 & ~n38908 ;
  assign n38910 = x99 & n14233 ;
  assign n38911 = x97 & n14876 ;
  assign n38912 = x98 & n14228 ;
  assign n38913 = ~n38911 & ~n38912 ;
  assign n38914 = ~n38910 & n38913 ;
  assign n38915 = n8660 & n14236 ;
  assign n38916 = n38914 & ~n38915 ;
  assign n38917 = x47 & ~n38916 ;
  assign n38918 = x47 & ~n38917 ;
  assign n38919 = ~n38916 & ~n38917 ;
  assign n38920 = ~n38918 & ~n38919 ;
  assign n38921 = n38909 & ~n38920 ;
  assign n38922 = n38909 & ~n38921 ;
  assign n38923 = ~n38920 & ~n38921 ;
  assign n38924 = ~n38922 & ~n38923 ;
  assign n38925 = ~n38273 & ~n38287 ;
  assign n38926 = ~n38924 & ~n38925 ;
  assign n38927 = ~n38924 & ~n38926 ;
  assign n38928 = ~n38925 & ~n38926 ;
  assign n38929 = ~n38927 & ~n38928 ;
  assign n38930 = x102 & n12506 ;
  assign n38931 = x100 & n13131 ;
  assign n38932 = x101 & n12501 ;
  assign n38933 = ~n38931 & ~n38932 ;
  assign n38934 = ~n38930 & n38933 ;
  assign n38935 = n10092 & n12509 ;
  assign n38936 = n38934 & ~n38935 ;
  assign n38937 = x44 & ~n38936 ;
  assign n38938 = x44 & ~n38937 ;
  assign n38939 = ~n38936 & ~n38937 ;
  assign n38940 = ~n38938 & ~n38939 ;
  assign n38941 = ~n38929 & n38940 ;
  assign n38942 = n38929 & ~n38940 ;
  assign n38943 = ~n38941 & ~n38942 ;
  assign n38944 = ~n38808 & ~n38943 ;
  assign n38945 = n38808 & n38943 ;
  assign n38946 = ~n38944 & ~n38945 ;
  assign n38947 = ~n38807 & n38946 ;
  assign n38948 = n38807 & ~n38946 ;
  assign n38949 = ~n38947 & ~n38948 ;
  assign n38950 = ~n38796 & n38949 ;
  assign n38951 = n38796 & ~n38949 ;
  assign n38952 = ~n38950 & ~n38951 ;
  assign n38953 = ~n38795 & n38952 ;
  assign n38954 = n38795 & ~n38952 ;
  assign n38955 = ~n38953 & ~n38954 ;
  assign n38956 = ~n38784 & n38955 ;
  assign n38957 = n38784 & ~n38955 ;
  assign n38958 = ~n38956 & ~n38957 ;
  assign n38959 = x111 & n8006 ;
  assign n38960 = x109 & n8474 ;
  assign n38961 = x110 & n8001 ;
  assign n38962 = ~n38960 & ~n38961 ;
  assign n38963 = ~n38959 & n38962 ;
  assign n38964 = n8009 & n15111 ;
  assign n38965 = n38963 & ~n38964 ;
  assign n38966 = x35 & ~n38965 ;
  assign n38967 = x35 & ~n38966 ;
  assign n38968 = ~n38965 & ~n38966 ;
  assign n38969 = ~n38967 & ~n38968 ;
  assign n38970 = n38958 & ~n38969 ;
  assign n38971 = n38958 & ~n38970 ;
  assign n38972 = ~n38969 & ~n38970 ;
  assign n38973 = ~n38971 & ~n38972 ;
  assign n38974 = n38783 & ~n38973 ;
  assign n38975 = ~n38783 & n38973 ;
  assign n38976 = ~n38768 & ~n38975 ;
  assign n38977 = ~n38974 & n38976 ;
  assign n38978 = ~n38768 & ~n38977 ;
  assign n38979 = ~n38975 & ~n38977 ;
  assign n38980 = ~n38974 & n38979 ;
  assign n38981 = ~n38978 & ~n38980 ;
  assign n38982 = n38752 & ~n38981 ;
  assign n38983 = ~n38752 & n38981 ;
  assign n38984 = ~n38737 & ~n38983 ;
  assign n38985 = ~n38982 & n38984 ;
  assign n38986 = ~n38737 & ~n38985 ;
  assign n38987 = ~n38983 & ~n38985 ;
  assign n38988 = ~n38982 & n38987 ;
  assign n38989 = ~n38986 & ~n38988 ;
  assign n38990 = ~n38721 & n38989 ;
  assign n38991 = n38721 & ~n38989 ;
  assign n38992 = ~n38990 & ~n38991 ;
  assign n38993 = ~n38706 & n38992 ;
  assign n38994 = n38706 & ~n38992 ;
  assign n38995 = ~n38993 & ~n38994 ;
  assign n38996 = ~n38694 & n38995 ;
  assign n38997 = ~n38694 & ~n38996 ;
  assign n38998 = n38995 & ~n38996 ;
  assign n38999 = ~n38997 & ~n38998 ;
  assign n39000 = ~n38693 & ~n38999 ;
  assign n39001 = n38693 & ~n38998 ;
  assign n39002 = ~n38997 & n39001 ;
  assign n39003 = ~n39000 & ~n39002 ;
  assign n39316 = n39003 & x208 ;
  assign n39004 = ~n38683 & ~n38686 ;
  assign n39005 = ~n38384 & ~n38676 ;
  assign n39006 = ~n38401 & ~n38673 ;
  assign n39007 = ~x127 & n2275 ;
  assign n39008 = n2096 & n27365 ;
  assign n39009 = ~n39007 & ~n39008 ;
  assign n39010 = ~x17 & ~n39009 ;
  assign n39011 = ~x17 & ~n39010 ;
  assign n39012 = ~n39009 & ~n39010 ;
  assign n39013 = ~n39011 & ~n39012 ;
  assign n39014 = ~n39006 & ~n39013 ;
  assign n39015 = ~n39006 & ~n39014 ;
  assign n39016 = ~n39013 & ~n39014 ;
  assign n39017 = ~n39015 & ~n39016 ;
  assign n39018 = ~x126 & n2751 ;
  assign n39019 = ~x124 & n3020 ;
  assign n39020 = ~x125 & n2746 ;
  assign n39021 = ~n39019 & ~n39020 ;
  assign n39022 = ~n39018 & n39021 ;
  assign n39023 = n2754 & n26128 ;
  assign n39024 = n39022 & ~n39023 ;
  assign n39025 = ~x20 & ~n39024 ;
  assign n39026 = ~x20 & ~n39025 ;
  assign n39027 = ~n39024 & ~n39025 ;
  assign n39028 = ~n39026 & ~n39027 ;
  assign n39029 = ~n38415 & ~n38668 ;
  assign n39030 = n39028 & n39029 ;
  assign n39031 = ~n39028 & ~n39029 ;
  assign n39032 = ~n39030 & ~n39031 ;
  assign n39033 = ~x123 & n3589 ;
  assign n39034 = ~x121 & n3878 ;
  assign n39035 = ~x122 & n3584 ;
  assign n39036 = ~n39034 & ~n39035 ;
  assign n39037 = ~n39033 & n39036 ;
  assign n39038 = n3592 & n23760 ;
  assign n39039 = n39037 & ~n39038 ;
  assign n39040 = ~x23 & ~n39039 ;
  assign n39041 = ~x23 & ~n39040 ;
  assign n39042 = ~n39039 & ~n39040 ;
  assign n39043 = ~n39041 & ~n39042 ;
  assign n39044 = ~n38431 & ~n38665 ;
  assign n39045 = ~n39043 & ~n39044 ;
  assign n39046 = ~n39043 & ~n39045 ;
  assign n39047 = ~n39044 & ~n39045 ;
  assign n39048 = ~n39046 & ~n39047 ;
  assign n39049 = ~x120 & n4531 ;
  assign n39050 = ~x118 & n4847 ;
  assign n39051 = ~x119 & n4526 ;
  assign n39052 = ~n39050 & ~n39051 ;
  assign n39053 = ~n39049 & n39052 ;
  assign n39054 = n4534 & n21501 ;
  assign n39055 = n39053 & ~n39054 ;
  assign n39056 = ~x26 & ~n39055 ;
  assign n39057 = ~x26 & ~n39056 ;
  assign n39058 = ~n39055 & ~n39056 ;
  assign n39059 = ~n39057 & ~n39058 ;
  assign n39060 = ~n38445 & ~n38660 ;
  assign n39061 = n39059 & n39060 ;
  assign n39062 = ~n39059 & ~n39060 ;
  assign n39063 = ~n39061 & ~n39062 ;
  assign n39064 = ~x117 & n5560 ;
  assign n39065 = ~x115 & n5943 ;
  assign n39066 = ~x116 & n5555 ;
  assign n39067 = ~n39065 & ~n39066 ;
  assign n39068 = ~n39064 & n39067 ;
  assign n39069 = n5563 & n19365 ;
  assign n39070 = n39068 & ~n39069 ;
  assign n39071 = ~x29 & ~n39070 ;
  assign n39072 = ~x29 & ~n39071 ;
  assign n39073 = ~n39070 & ~n39071 ;
  assign n39074 = ~n39072 & ~n39073 ;
  assign n39075 = ~n38462 & ~n38657 ;
  assign n39076 = ~n39074 & ~n39075 ;
  assign n39077 = ~n39074 & ~n39076 ;
  assign n39078 = ~n39075 & ~n39076 ;
  assign n39079 = ~n39077 & ~n39078 ;
  assign n39080 = ~x114 & n6725 ;
  assign n39081 = ~x112 & n7129 ;
  assign n39082 = ~x113 & n6720 ;
  assign n39083 = ~n39081 & ~n39082 ;
  assign n39084 = ~n39080 & n39083 ;
  assign n39085 = n6728 & n17333 ;
  assign n39086 = n39084 & ~n39085 ;
  assign n39087 = ~x32 & ~n39086 ;
  assign n39088 = ~x32 & ~n39087 ;
  assign n39089 = ~n39086 & ~n39087 ;
  assign n39090 = ~n39088 & ~n39089 ;
  assign n39091 = ~n38640 & ~n38653 ;
  assign n39092 = n39090 & n39091 ;
  assign n39093 = ~n39090 & ~n39091 ;
  assign n39094 = ~n39092 & ~n39093 ;
  assign n39095 = ~n38620 & ~n38634 ;
  assign n39096 = ~x108 & n9433 ;
  assign n39097 = ~x106 & n9915 ;
  assign n39098 = ~x107 & n9428 ;
  assign n39099 = ~n39097 & ~n39098 ;
  assign n39100 = ~n39096 & n39099 ;
  assign n39101 = n9436 & n13601 ;
  assign n39102 = n39100 & ~n39101 ;
  assign n39103 = ~x38 & ~n39102 ;
  assign n39104 = ~x38 & ~n39103 ;
  assign n39105 = ~n39102 & ~n39103 ;
  assign n39106 = ~n39104 & ~n39105 ;
  assign n39107 = ~n38612 & ~n38616 ;
  assign n39108 = ~x105 & n10905 ;
  assign n39109 = ~x103 & n11466 ;
  assign n39110 = ~x104 & n10900 ;
  assign n39111 = ~n39109 & ~n39110 ;
  assign n39112 = ~n39108 & n39111 ;
  assign n39113 = n10908 & n11907 ;
  assign n39114 = n39112 & ~n39113 ;
  assign n39115 = ~x41 & ~n39114 ;
  assign n39116 = ~x41 & ~n39115 ;
  assign n39117 = ~n39114 & ~n39115 ;
  assign n39118 = ~n39116 & ~n39117 ;
  assign n39119 = ~n38604 & ~n38608 ;
  assign n39120 = ~n38533 & ~n38546 ;
  assign n39121 = ~x90 & n20143 ;
  assign n39122 = ~x88 & n20854 ;
  assign n39123 = ~x89 & n20138 ;
  assign n39124 = ~n39122 & ~n39123 ;
  assign n39125 = ~n39121 & n39124 ;
  assign n39126 = n5155 & n20146 ;
  assign n39127 = n39125 & ~n39126 ;
  assign n39128 = ~x56 & ~n39127 ;
  assign n39129 = ~x56 & ~n39128 ;
  assign n39130 = ~n39127 & ~n39128 ;
  assign n39131 = ~n39129 & ~n39130 ;
  assign n39132 = ~n38513 & ~n38527 ;
  assign n39133 = ~x84 & n24612 ;
  assign n39134 = ~x82 & n25390 ;
  assign n39135 = ~x83 & n24607 ;
  assign n39136 = ~n39134 & ~n39135 ;
  assign n39137 = ~n39133 & n39136 ;
  assign n39138 = n3247 & n24615 ;
  assign n39139 = n39137 & ~n39138 ;
  assign n39140 = ~x62 & ~n39139 ;
  assign n39141 = ~x62 & ~n39140 ;
  assign n39142 = ~n39139 & ~n39140 ;
  assign n39143 = ~n39141 & ~n39142 ;
  assign n39144 = ~x80 & n27427 ;
  assign n39145 = ~x81 & ~n26217 ;
  assign n39146 = ~n39144 & ~n39145 ;
  assign n39147 = n38494 & ~n39146 ;
  assign n39148 = ~n38494 & n39146 ;
  assign n39149 = ~n39143 & ~n39148 ;
  assign n39150 = ~n39147 & n39149 ;
  assign n39151 = ~n39143 & ~n39150 ;
  assign n39152 = ~n39148 & ~n39150 ;
  assign n39153 = ~n39147 & n39152 ;
  assign n39154 = ~n39151 & ~n39153 ;
  assign n39155 = ~n38497 & ~n38510 ;
  assign n39156 = n39154 & n39155 ;
  assign n39157 = ~n39154 & ~n39155 ;
  assign n39158 = ~n39156 & ~n39157 ;
  assign n39159 = ~x87 & n22325 ;
  assign n39160 = ~x85 & n23066 ;
  assign n39161 = ~x86 & n22320 ;
  assign n39162 = ~n39160 & ~n39161 ;
  assign n39163 = ~n39159 & n39162 ;
  assign n39164 = n4143 & n22328 ;
  assign n39165 = n39163 & ~n39164 ;
  assign n39166 = ~x59 & ~n39165 ;
  assign n39167 = ~x59 & ~n39166 ;
  assign n39168 = ~n39165 & ~n39166 ;
  assign n39169 = ~n39167 & ~n39168 ;
  assign n39170 = ~n39158 & n39169 ;
  assign n39171 = n39158 & ~n39169 ;
  assign n39172 = ~n39170 & ~n39171 ;
  assign n39173 = ~n39132 & n39172 ;
  assign n39174 = n39132 & ~n39172 ;
  assign n39175 = ~n39173 & ~n39174 ;
  assign n39176 = ~n39131 & n39175 ;
  assign n39177 = n39131 & ~n39175 ;
  assign n39178 = ~n39176 & ~n39177 ;
  assign n39179 = ~n39120 & n39178 ;
  assign n39180 = n39120 & ~n39178 ;
  assign n39181 = ~n39179 & ~n39180 ;
  assign n39182 = ~x93 & n18025 ;
  assign n39183 = ~x91 & n18764 ;
  assign n39184 = ~x92 & n18020 ;
  assign n39185 = ~n39183 & ~n39184 ;
  assign n39186 = ~n39182 & n39185 ;
  assign n39187 = n6285 & n18028 ;
  assign n39188 = n39186 & ~n39187 ;
  assign n39189 = ~x53 & ~n39188 ;
  assign n39190 = ~x53 & ~n39189 ;
  assign n39191 = ~n39188 & ~n39189 ;
  assign n39192 = ~n39190 & ~n39191 ;
  assign n39193 = n39181 & ~n39192 ;
  assign n39194 = n39181 & ~n39193 ;
  assign n39195 = ~n39192 & ~n39193 ;
  assign n39196 = ~n39194 & ~n39195 ;
  assign n39197 = ~n37877 & ~n38549 ;
  assign n39198 = ~n38565 & ~n39197 ;
  assign n39199 = ~n39196 & ~n39198 ;
  assign n39200 = ~n39196 & ~n39199 ;
  assign n39201 = ~n39198 & ~n39199 ;
  assign n39202 = ~n39200 & ~n39201 ;
  assign n39203 = ~x96 & n16076 ;
  assign n39204 = ~x94 & n16756 ;
  assign n39205 = ~x95 & n16071 ;
  assign n39206 = ~n39204 & ~n39205 ;
  assign n39207 = ~n39203 & n39206 ;
  assign n39208 = n7531 & n16079 ;
  assign n39209 = n39207 & ~n39208 ;
  assign n39210 = ~x50 & ~n39209 ;
  assign n39211 = ~x50 & ~n39210 ;
  assign n39212 = ~n39209 & ~n39210 ;
  assign n39213 = ~n39211 & ~n39212 ;
  assign n39214 = ~n39202 & n39213 ;
  assign n39215 = n39202 & ~n39213 ;
  assign n39216 = ~n39214 & ~n39215 ;
  assign n39217 = ~n38568 & ~n38582 ;
  assign n39218 = n39216 & n39217 ;
  assign n39219 = ~n39216 & ~n39217 ;
  assign n39220 = ~n39218 & ~n39219 ;
  assign n39221 = ~x99 & n14233 ;
  assign n39222 = ~x97 & n14876 ;
  assign n39223 = ~x98 & n14228 ;
  assign n39224 = ~n39222 & ~n39223 ;
  assign n39225 = ~n39221 & n39224 ;
  assign n39226 = n8885 & n14236 ;
  assign n39227 = n39225 & ~n39226 ;
  assign n39228 = ~x47 & ~n39227 ;
  assign n39229 = ~x47 & ~n39228 ;
  assign n39230 = ~n39227 & ~n39228 ;
  assign n39231 = ~n39229 & ~n39230 ;
  assign n39232 = n39220 & ~n39231 ;
  assign n39233 = n39220 & ~n39232 ;
  assign n39234 = ~n39231 & ~n39232 ;
  assign n39235 = ~n39233 & ~n39234 ;
  assign n39236 = ~n38588 & ~n38602 ;
  assign n39237 = ~n39235 & ~n39236 ;
  assign n39238 = ~n39235 & ~n39237 ;
  assign n39239 = ~n39236 & ~n39237 ;
  assign n39240 = ~n39238 & ~n39239 ;
  assign n39241 = ~x102 & n12506 ;
  assign n39242 = ~x100 & n13131 ;
  assign n39243 = ~x101 & n12501 ;
  assign n39244 = ~n39242 & ~n39243 ;
  assign n39245 = ~n39241 & n39244 ;
  assign n39246 = n10333 & n12509 ;
  assign n39247 = n39245 & ~n39246 ;
  assign n39248 = ~x44 & ~n39247 ;
  assign n39249 = ~x44 & ~n39248 ;
  assign n39250 = ~n39247 & ~n39248 ;
  assign n39251 = ~n39249 & ~n39250 ;
  assign n39252 = ~n39240 & n39251 ;
  assign n39253 = n39240 & ~n39251 ;
  assign n39254 = ~n39252 & ~n39253 ;
  assign n39255 = ~n39119 & ~n39254 ;
  assign n39256 = n39119 & n39254 ;
  assign n39257 = ~n39255 & ~n39256 ;
  assign n39258 = ~n39118 & n39257 ;
  assign n39259 = n39118 & ~n39257 ;
  assign n39260 = ~n39258 & ~n39259 ;
  assign n39261 = ~n39107 & n39260 ;
  assign n39262 = n39107 & ~n39260 ;
  assign n39263 = ~n39261 & ~n39262 ;
  assign n39264 = ~n39106 & n39263 ;
  assign n39265 = n39106 & ~n39263 ;
  assign n39266 = ~n39264 & ~n39265 ;
  assign n39267 = ~n39095 & n39266 ;
  assign n39268 = n39095 & ~n39266 ;
  assign n39269 = ~n39267 & ~n39268 ;
  assign n39270 = ~x111 & n8006 ;
  assign n39271 = ~x109 & n8474 ;
  assign n39272 = ~x110 & n8001 ;
  assign n39273 = ~n39271 & ~n39272 ;
  assign n39274 = ~n39270 & n39273 ;
  assign n39275 = n8009 & n15411 ;
  assign n39276 = n39274 & ~n39275 ;
  assign n39277 = ~x35 & ~n39276 ;
  assign n39278 = ~x35 & ~n39277 ;
  assign n39279 = ~n39276 & ~n39277 ;
  assign n39280 = ~n39278 & ~n39279 ;
  assign n39281 = n39269 & ~n39280 ;
  assign n39282 = n39269 & ~n39281 ;
  assign n39283 = ~n39280 & ~n39281 ;
  assign n39284 = ~n39282 & ~n39283 ;
  assign n39285 = n39094 & ~n39284 ;
  assign n39286 = ~n39094 & n39284 ;
  assign n39287 = ~n39079 & ~n39286 ;
  assign n39288 = ~n39285 & n39287 ;
  assign n39289 = ~n39079 & ~n39288 ;
  assign n39290 = ~n39286 & ~n39288 ;
  assign n39291 = ~n39285 & n39290 ;
  assign n39292 = ~n39289 & ~n39291 ;
  assign n39293 = n39063 & ~n39292 ;
  assign n39294 = ~n39063 & n39292 ;
  assign n39295 = ~n39048 & ~n39294 ;
  assign n39296 = ~n39293 & n39295 ;
  assign n39297 = ~n39048 & ~n39296 ;
  assign n39298 = ~n39294 & ~n39296 ;
  assign n39299 = ~n39293 & n39298 ;
  assign n39300 = ~n39297 & ~n39299 ;
  assign n39301 = ~n39032 & n39300 ;
  assign n39302 = n39032 & ~n39300 ;
  assign n39303 = ~n39301 & ~n39302 ;
  assign n39304 = ~n39017 & n39303 ;
  assign n39305 = n39017 & ~n39303 ;
  assign n39306 = ~n39304 & ~n39305 ;
  assign n39307 = ~n39005 & n39306 ;
  assign n39308 = ~n39005 & ~n39307 ;
  assign n39309 = n39306 & ~n39307 ;
  assign n39310 = ~n39308 & ~n39309 ;
  assign n39311 = ~n39004 & ~n39310 ;
  assign n39312 = n39004 & ~n39309 ;
  assign n39313 = ~n39308 & n39312 ;
  assign n39314 = ~n39311 & ~n39313 ;
  assign n39317 = ~n39314 & ~x208 ;
  assign n39318 = ~n39316 & ~n39317 ;
  assign n39319 = ~n38996 & ~n39000 ;
  assign n39320 = ~n38703 & ~n38993 ;
  assign n39321 = ~n38720 & ~n38991 ;
  assign n39322 = x127 & n2751 ;
  assign n39323 = x125 & n3020 ;
  assign n39324 = x126 & n2746 ;
  assign n39325 = ~n39323 & ~n39324 ;
  assign n39326 = ~n39322 & n39325 ;
  assign n39327 = n2754 & n26533 ;
  assign n39328 = n39326 & ~n39327 ;
  assign n39329 = x20 & ~n39328 ;
  assign n39330 = x20 & ~n39329 ;
  assign n39331 = ~n39328 & ~n39329 ;
  assign n39332 = ~n39330 & ~n39331 ;
  assign n39333 = ~n39321 & ~n39332 ;
  assign n39334 = ~n39321 & ~n39333 ;
  assign n39335 = ~n39332 & ~n39333 ;
  assign n39336 = ~n39334 & ~n39335 ;
  assign n39337 = x124 & n3589 ;
  assign n39338 = x122 & n3878 ;
  assign n39339 = x123 & n3584 ;
  assign n39340 = ~n39338 & ~n39339 ;
  assign n39341 = ~n39337 & n39340 ;
  assign n39342 = n3592 & n23796 ;
  assign n39343 = n39341 & ~n39342 ;
  assign n39344 = x23 & ~n39343 ;
  assign n39345 = x23 & ~n39344 ;
  assign n39346 = ~n39343 & ~n39344 ;
  assign n39347 = ~n39345 & ~n39346 ;
  assign n39348 = ~n38734 & ~n38985 ;
  assign n39349 = n39347 & n39348 ;
  assign n39350 = ~n39347 & ~n39348 ;
  assign n39351 = ~n39349 & ~n39350 ;
  assign n39352 = x118 & n5560 ;
  assign n39353 = x116 & n5943 ;
  assign n39354 = x117 & n5555 ;
  assign n39355 = ~n39353 & ~n39354 ;
  assign n39356 = ~n39352 & n39355 ;
  assign n39357 = n5563 & n19395 ;
  assign n39358 = n39356 & ~n39357 ;
  assign n39359 = x29 & ~n39358 ;
  assign n39360 = x29 & ~n39359 ;
  assign n39361 = ~n39358 & ~n39359 ;
  assign n39362 = ~n39360 & ~n39361 ;
  assign n39363 = ~n38765 & ~n38977 ;
  assign n39364 = n39362 & n39363 ;
  assign n39365 = ~n39362 & ~n39363 ;
  assign n39366 = ~n39364 & ~n39365 ;
  assign n39367 = ~n38944 & ~n38947 ;
  assign n39368 = ~n38929 & ~n38940 ;
  assign n39369 = ~n38926 & ~n39368 ;
  assign n39370 = ~n38908 & ~n38921 ;
  assign n39371 = ~n38846 & ~n38860 ;
  assign n39372 = x85 & n24612 ;
  assign n39373 = x83 & n25390 ;
  assign n39374 = x84 & n24607 ;
  assign n39375 = ~n39373 & ~n39374 ;
  assign n39376 = ~n39372 & n39375 ;
  assign n39377 = n3389 & n24615 ;
  assign n39378 = n39376 & ~n39377 ;
  assign n39379 = x62 & ~n39378 ;
  assign n39380 = x62 & ~n39379 ;
  assign n39381 = ~n39378 & ~n39379 ;
  assign n39382 = ~n39380 & ~n39381 ;
  assign n39383 = x81 & n27024 ;
  assign n39384 = x82 & ~n26217 ;
  assign n39385 = ~n39383 & ~n39384 ;
  assign n39386 = ~x17 & ~n39385 ;
  assign n39387 = x17 & n39385 ;
  assign n39388 = ~n39386 & ~n39387 ;
  assign n39389 = ~n38835 & n39388 ;
  assign n39390 = n38835 & ~n39388 ;
  assign n39391 = ~n39389 & ~n39390 ;
  assign n39392 = ~n39382 & n39391 ;
  assign n39393 = ~n39382 & ~n39392 ;
  assign n39394 = n39391 & ~n39392 ;
  assign n39395 = ~n39393 & ~n39394 ;
  assign n39396 = ~n38841 & ~n39395 ;
  assign n39397 = ~n38841 & ~n39396 ;
  assign n39398 = ~n39395 & ~n39396 ;
  assign n39399 = ~n39397 & ~n39398 ;
  assign n39400 = x88 & n22325 ;
  assign n39401 = x86 & n23066 ;
  assign n39402 = x87 & n22320 ;
  assign n39403 = ~n39401 & ~n39402 ;
  assign n39404 = ~n39400 & n39403 ;
  assign n39405 = n4305 & n22328 ;
  assign n39406 = n39404 & ~n39405 ;
  assign n39407 = x59 & ~n39406 ;
  assign n39408 = x59 & ~n39407 ;
  assign n39409 = ~n39406 & ~n39407 ;
  assign n39410 = ~n39408 & ~n39409 ;
  assign n39411 = n39399 & n39410 ;
  assign n39412 = ~n39399 & ~n39410 ;
  assign n39413 = ~n39411 & ~n39412 ;
  assign n39414 = ~n39371 & n39413 ;
  assign n39415 = n39371 & ~n39413 ;
  assign n39416 = ~n39414 & ~n39415 ;
  assign n39417 = x91 & n20143 ;
  assign n39418 = x89 & n20854 ;
  assign n39419 = x90 & n20138 ;
  assign n39420 = ~n39418 & ~n39419 ;
  assign n39421 = ~n39417 & n39420 ;
  assign n39422 = n5336 & n20146 ;
  assign n39423 = n39421 & ~n39422 ;
  assign n39424 = x56 & ~n39423 ;
  assign n39425 = x56 & ~n39424 ;
  assign n39426 = ~n39423 & ~n39424 ;
  assign n39427 = ~n39425 & ~n39426 ;
  assign n39428 = n39416 & ~n39427 ;
  assign n39429 = n39416 & ~n39428 ;
  assign n39430 = ~n39427 & ~n39428 ;
  assign n39431 = ~n39429 & ~n39430 ;
  assign n39432 = ~n38862 & ~n38865 ;
  assign n39433 = n39431 & n39432 ;
  assign n39434 = ~n39431 & ~n39432 ;
  assign n39435 = ~n39433 & ~n39434 ;
  assign n39436 = x94 & n18025 ;
  assign n39437 = x92 & n18764 ;
  assign n39438 = x93 & n18020 ;
  assign n39439 = ~n39437 & ~n39438 ;
  assign n39440 = ~n39436 & n39439 ;
  assign n39441 = n6483 & n18028 ;
  assign n39442 = n39440 & ~n39441 ;
  assign n39443 = x53 & ~n39442 ;
  assign n39444 = x53 & ~n39443 ;
  assign n39445 = ~n39442 & ~n39443 ;
  assign n39446 = ~n39444 & ~n39445 ;
  assign n39447 = n39435 & ~n39446 ;
  assign n39448 = n39435 & ~n39447 ;
  assign n39449 = ~n39446 & ~n39447 ;
  assign n39450 = ~n39448 & ~n39449 ;
  assign n39451 = ~n38868 & ~n38882 ;
  assign n39452 = n39450 & n39451 ;
  assign n39453 = ~n39450 & ~n39451 ;
  assign n39454 = ~n39452 & ~n39453 ;
  assign n39455 = x97 & n16076 ;
  assign n39456 = x95 & n16756 ;
  assign n39457 = x96 & n16071 ;
  assign n39458 = ~n39456 & ~n39457 ;
  assign n39459 = ~n39455 & n39458 ;
  assign n39460 = n7745 & n16079 ;
  assign n39461 = n39459 & ~n39460 ;
  assign n39462 = x50 & ~n39461 ;
  assign n39463 = x50 & ~n39462 ;
  assign n39464 = ~n39461 & ~n39462 ;
  assign n39465 = ~n39463 & ~n39464 ;
  assign n39466 = ~n38891 & ~n38902 ;
  assign n39467 = ~n38888 & ~n39466 ;
  assign n39468 = ~n39465 & ~n39467 ;
  assign n39469 = n39465 & n39467 ;
  assign n39470 = ~n39468 & ~n39469 ;
  assign n39471 = ~n39454 & n39470 ;
  assign n39472 = n39454 & ~n39470 ;
  assign n39473 = ~n39471 & ~n39472 ;
  assign n39474 = x100 & n14233 ;
  assign n39475 = x98 & n14876 ;
  assign n39476 = x99 & n14228 ;
  assign n39477 = ~n39475 & ~n39476 ;
  assign n39478 = ~n39474 & n39477 ;
  assign n39479 = n9115 & n14236 ;
  assign n39480 = n39478 & ~n39479 ;
  assign n39481 = x47 & ~n39480 ;
  assign n39482 = x47 & ~n39481 ;
  assign n39483 = ~n39480 & ~n39481 ;
  assign n39484 = ~n39482 & ~n39483 ;
  assign n39485 = ~n39473 & ~n39484 ;
  assign n39486 = n39473 & n39484 ;
  assign n39487 = ~n39485 & ~n39486 ;
  assign n39488 = n39370 & ~n39487 ;
  assign n39489 = ~n39370 & n39487 ;
  assign n39490 = ~n39488 & ~n39489 ;
  assign n39491 = x103 & n12506 ;
  assign n39492 = x101 & n13131 ;
  assign n39493 = x102 & n12501 ;
  assign n39494 = ~n39492 & ~n39493 ;
  assign n39495 = ~n39491 & n39494 ;
  assign n39496 = n10588 & n12509 ;
  assign n39497 = n39495 & ~n39496 ;
  assign n39498 = x44 & ~n39497 ;
  assign n39499 = x44 & ~n39498 ;
  assign n39500 = ~n39497 & ~n39498 ;
  assign n39501 = ~n39499 & ~n39500 ;
  assign n39502 = n39490 & ~n39501 ;
  assign n39503 = n39490 & ~n39502 ;
  assign n39504 = ~n39501 & ~n39502 ;
  assign n39505 = ~n39503 & ~n39504 ;
  assign n39506 = ~n39369 & n39505 ;
  assign n39507 = n39369 & ~n39505 ;
  assign n39508 = ~n39506 & ~n39507 ;
  assign n39509 = x106 & n10905 ;
  assign n39510 = x104 & n11466 ;
  assign n39511 = x105 & n10900 ;
  assign n39512 = ~n39510 & ~n39511 ;
  assign n39513 = ~n39509 & n39512 ;
  assign n39514 = n10908 & n12181 ;
  assign n39515 = n39513 & ~n39514 ;
  assign n39516 = x41 & ~n39515 ;
  assign n39517 = x41 & ~n39516 ;
  assign n39518 = ~n39515 & ~n39516 ;
  assign n39519 = ~n39517 & ~n39518 ;
  assign n39520 = ~n39508 & ~n39519 ;
  assign n39521 = n39508 & n39519 ;
  assign n39522 = ~n39520 & ~n39521 ;
  assign n39523 = n39367 & ~n39522 ;
  assign n39524 = ~n39367 & n39522 ;
  assign n39525 = ~n39523 & ~n39524 ;
  assign n39526 = x109 & n9433 ;
  assign n39527 = x107 & n9915 ;
  assign n39528 = x108 & n9428 ;
  assign n39529 = ~n39527 & ~n39528 ;
  assign n39530 = ~n39526 & n39529 ;
  assign n39531 = n9436 & n13894 ;
  assign n39532 = n39530 & ~n39531 ;
  assign n39533 = x38 & ~n39532 ;
  assign n39534 = x38 & ~n39533 ;
  assign n39535 = ~n39532 & ~n39533 ;
  assign n39536 = ~n39534 & ~n39535 ;
  assign n39537 = n39525 & ~n39536 ;
  assign n39538 = n39525 & ~n39537 ;
  assign n39539 = ~n39536 & ~n39537 ;
  assign n39540 = ~n39538 & ~n39539 ;
  assign n39541 = ~n38950 & ~n38953 ;
  assign n39542 = n39540 & n39541 ;
  assign n39543 = ~n39540 & ~n39541 ;
  assign n39544 = ~n39542 & ~n39543 ;
  assign n39545 = x112 & n8006 ;
  assign n39546 = x110 & n8474 ;
  assign n39547 = x111 & n8001 ;
  assign n39548 = ~n39546 & ~n39547 ;
  assign n39549 = ~n39545 & n39548 ;
  assign n39550 = n8009 & n15442 ;
  assign n39551 = n39549 & ~n39550 ;
  assign n39552 = x35 & ~n39551 ;
  assign n39553 = x35 & ~n39552 ;
  assign n39554 = ~n39551 & ~n39552 ;
  assign n39555 = ~n39553 & ~n39554 ;
  assign n39556 = n39544 & ~n39555 ;
  assign n39557 = n39544 & ~n39556 ;
  assign n39558 = ~n39555 & ~n39556 ;
  assign n39559 = ~n39557 & ~n39558 ;
  assign n39560 = ~n38956 & ~n38970 ;
  assign n39561 = n39559 & n39560 ;
  assign n39562 = ~n39559 & ~n39560 ;
  assign n39563 = ~n39561 & ~n39562 ;
  assign n39564 = x115 & n6725 ;
  assign n39565 = x113 & n7129 ;
  assign n39566 = x114 & n6720 ;
  assign n39567 = ~n39565 & ~n39566 ;
  assign n39568 = ~n39564 & n39567 ;
  assign n39569 = n6728 & n17364 ;
  assign n39570 = n39568 & ~n39569 ;
  assign n39571 = x32 & ~n39570 ;
  assign n39572 = x32 & ~n39571 ;
  assign n39573 = ~n39570 & ~n39571 ;
  assign n39574 = ~n39572 & ~n39573 ;
  assign n39575 = ~n38782 & ~n38974 ;
  assign n39576 = ~n39574 & ~n39575 ;
  assign n39577 = n39574 & n39575 ;
  assign n39578 = ~n39576 & ~n39577 ;
  assign n39579 = n39563 & n39578 ;
  assign n39580 = n39563 & ~n39579 ;
  assign n39581 = n39578 & ~n39579 ;
  assign n39582 = ~n39580 & ~n39581 ;
  assign n39583 = n39366 & ~n39582 ;
  assign n39584 = n39366 & ~n39583 ;
  assign n39585 = ~n39582 & ~n39583 ;
  assign n39586 = ~n39584 & ~n39585 ;
  assign n39587 = x121 & n4531 ;
  assign n39588 = x119 & n4847 ;
  assign n39589 = x120 & n4526 ;
  assign n39590 = ~n39588 & ~n39589 ;
  assign n39591 = ~n39587 & n39590 ;
  assign n39592 = n4534 & n21870 ;
  assign n39593 = n39591 & ~n39592 ;
  assign n39594 = x26 & ~n39593 ;
  assign n39595 = x26 & ~n39594 ;
  assign n39596 = ~n39593 & ~n39594 ;
  assign n39597 = ~n39595 & ~n39596 ;
  assign n39598 = ~n38751 & ~n38982 ;
  assign n39599 = ~n39597 & ~n39598 ;
  assign n39600 = n39597 & n39598 ;
  assign n39601 = ~n39599 & ~n39600 ;
  assign n39602 = ~n39586 & n39601 ;
  assign n39603 = ~n39586 & ~n39602 ;
  assign n39604 = n39601 & ~n39602 ;
  assign n39605 = ~n39603 & ~n39604 ;
  assign n39606 = n39351 & ~n39605 ;
  assign n39607 = n39351 & ~n39606 ;
  assign n39608 = ~n39605 & ~n39606 ;
  assign n39609 = ~n39607 & ~n39608 ;
  assign n39610 = ~n39336 & n39609 ;
  assign n39611 = n39336 & ~n39609 ;
  assign n39612 = ~n39610 & ~n39611 ;
  assign n39613 = ~n39320 & ~n39612 ;
  assign n39614 = ~n39320 & ~n39613 ;
  assign n39615 = ~n39612 & ~n39613 ;
  assign n39616 = ~n39614 & ~n39615 ;
  assign n39617 = ~n39319 & ~n39616 ;
  assign n39618 = n39319 & ~n39615 ;
  assign n39619 = ~n39614 & n39618 ;
  assign n39620 = ~n39617 & ~n39619 ;
  assign n39924 = n39620 & x209 ;
  assign n39621 = ~n39307 & ~n39311 ;
  assign n39622 = ~n39014 & ~n39304 ;
  assign n39623 = ~n39031 & ~n39302 ;
  assign n39624 = ~x127 & n2751 ;
  assign n39625 = ~x125 & n3020 ;
  assign n39626 = ~x126 & n2746 ;
  assign n39627 = ~n39625 & ~n39626 ;
  assign n39628 = ~n39624 & n39627 ;
  assign n39629 = n2754 & n26932 ;
  assign n39630 = n39628 & ~n39629 ;
  assign n39631 = ~x20 & ~n39630 ;
  assign n39632 = ~x20 & ~n39631 ;
  assign n39633 = ~n39630 & ~n39631 ;
  assign n39634 = ~n39632 & ~n39633 ;
  assign n39635 = ~n39623 & ~n39634 ;
  assign n39636 = ~n39623 & ~n39635 ;
  assign n39637 = ~n39634 & ~n39635 ;
  assign n39638 = ~n39636 & ~n39637 ;
  assign n39639 = ~x124 & n3589 ;
  assign n39640 = ~x122 & n3878 ;
  assign n39641 = ~x123 & n3584 ;
  assign n39642 = ~n39640 & ~n39641 ;
  assign n39643 = ~n39639 & n39642 ;
  assign n39644 = n3592 & n24176 ;
  assign n39645 = n39643 & ~n39644 ;
  assign n39646 = ~x23 & ~n39645 ;
  assign n39647 = ~x23 & ~n39646 ;
  assign n39648 = ~n39645 & ~n39646 ;
  assign n39649 = ~n39647 & ~n39648 ;
  assign n39650 = ~n39045 & ~n39296 ;
  assign n39651 = n39649 & n39650 ;
  assign n39652 = ~n39649 & ~n39650 ;
  assign n39653 = ~n39651 & ~n39652 ;
  assign n39654 = ~x118 & n5560 ;
  assign n39655 = ~x116 & n5943 ;
  assign n39656 = ~x117 & n5555 ;
  assign n39657 = ~n39655 & ~n39656 ;
  assign n39658 = ~n39654 & n39657 ;
  assign n39659 = n5563 & n19736 ;
  assign n39660 = n39658 & ~n39659 ;
  assign n39661 = ~x29 & ~n39660 ;
  assign n39662 = ~x29 & ~n39661 ;
  assign n39663 = ~n39660 & ~n39661 ;
  assign n39664 = ~n39662 & ~n39663 ;
  assign n39665 = ~n39076 & ~n39288 ;
  assign n39666 = n39664 & n39665 ;
  assign n39667 = ~n39664 & ~n39665 ;
  assign n39668 = ~n39666 & ~n39667 ;
  assign n39669 = ~n39255 & ~n39258 ;
  assign n39670 = ~n39240 & ~n39251 ;
  assign n39671 = ~n39237 & ~n39670 ;
  assign n39672 = ~n39219 & ~n39232 ;
  assign n39673 = ~n39157 & ~n39171 ;
  assign n39674 = ~x85 & n24612 ;
  assign n39675 = ~x83 & n25390 ;
  assign n39676 = ~x84 & n24607 ;
  assign n39677 = ~n39675 & ~n39676 ;
  assign n39678 = ~n39674 & n39677 ;
  assign n39679 = n3521 & n24615 ;
  assign n39680 = n39678 & ~n39679 ;
  assign n39681 = ~x62 & ~n39680 ;
  assign n39682 = ~x62 & ~n39681 ;
  assign n39683 = ~n39680 & ~n39681 ;
  assign n39684 = ~n39682 & ~n39683 ;
  assign n39685 = ~x81 & n27427 ;
  assign n39686 = ~x82 & ~n26217 ;
  assign n39687 = ~n39685 & ~n39686 ;
  assign n39688 = x17 & ~n39687 ;
  assign n39689 = ~x17 & n39687 ;
  assign n39690 = ~n39688 & ~n39689 ;
  assign n39691 = ~n39146 & n39690 ;
  assign n39692 = n39146 & ~n39690 ;
  assign n39693 = ~n39691 & ~n39692 ;
  assign n39694 = ~n39684 & n39693 ;
  assign n39695 = ~n39684 & ~n39694 ;
  assign n39696 = n39693 & ~n39694 ;
  assign n39697 = ~n39695 & ~n39696 ;
  assign n39698 = ~n39152 & ~n39697 ;
  assign n39699 = ~n39152 & ~n39698 ;
  assign n39700 = ~n39697 & ~n39698 ;
  assign n39701 = ~n39699 & ~n39700 ;
  assign n39702 = ~x88 & n22325 ;
  assign n39703 = ~x86 & n23066 ;
  assign n39704 = ~x87 & n22320 ;
  assign n39705 = ~n39703 & ~n39704 ;
  assign n39706 = ~n39702 & n39705 ;
  assign n39707 = n4457 & n22328 ;
  assign n39708 = n39706 & ~n39707 ;
  assign n39709 = ~x59 & ~n39708 ;
  assign n39710 = ~x59 & ~n39709 ;
  assign n39711 = ~n39708 & ~n39709 ;
  assign n39712 = ~n39710 & ~n39711 ;
  assign n39713 = n39701 & n39712 ;
  assign n39714 = ~n39701 & ~n39712 ;
  assign n39715 = ~n39713 & ~n39714 ;
  assign n39716 = ~n39673 & n39715 ;
  assign n39717 = n39673 & ~n39715 ;
  assign n39718 = ~n39716 & ~n39717 ;
  assign n39719 = ~x91 & n20143 ;
  assign n39720 = ~x89 & n20854 ;
  assign n39721 = ~x90 & n20138 ;
  assign n39722 = ~n39720 & ~n39721 ;
  assign n39723 = ~n39719 & n39722 ;
  assign n39724 = n5507 & n20146 ;
  assign n39725 = n39723 & ~n39724 ;
  assign n39726 = ~x56 & ~n39725 ;
  assign n39727 = ~x56 & ~n39726 ;
  assign n39728 = ~n39725 & ~n39726 ;
  assign n39729 = ~n39727 & ~n39728 ;
  assign n39730 = n39718 & ~n39729 ;
  assign n39731 = n39718 & ~n39730 ;
  assign n39732 = ~n39729 & ~n39730 ;
  assign n39733 = ~n39731 & ~n39732 ;
  assign n39734 = ~n39173 & ~n39176 ;
  assign n39735 = n39733 & n39734 ;
  assign n39736 = ~n39733 & ~n39734 ;
  assign n39737 = ~n39735 & ~n39736 ;
  assign n39738 = ~x94 & n18025 ;
  assign n39739 = ~x92 & n18764 ;
  assign n39740 = ~x93 & n18020 ;
  assign n39741 = ~n39739 & ~n39740 ;
  assign n39742 = ~n39738 & n39741 ;
  assign n39743 = n6671 & n18028 ;
  assign n39744 = n39742 & ~n39743 ;
  assign n39745 = ~x53 & ~n39744 ;
  assign n39746 = ~x53 & ~n39745 ;
  assign n39747 = ~n39744 & ~n39745 ;
  assign n39748 = ~n39746 & ~n39747 ;
  assign n39749 = n39737 & ~n39748 ;
  assign n39750 = n39737 & ~n39749 ;
  assign n39751 = ~n39748 & ~n39749 ;
  assign n39752 = ~n39750 & ~n39751 ;
  assign n39753 = ~n39179 & ~n39193 ;
  assign n39754 = n39752 & n39753 ;
  assign n39755 = ~n39752 & ~n39753 ;
  assign n39756 = ~n39754 & ~n39755 ;
  assign n39757 = ~x97 & n16076 ;
  assign n39758 = ~x95 & n16756 ;
  assign n39759 = ~x96 & n16071 ;
  assign n39760 = ~n39758 & ~n39759 ;
  assign n39761 = ~n39757 & n39760 ;
  assign n39762 = n7949 & n16079 ;
  assign n39763 = n39761 & ~n39762 ;
  assign n39764 = ~x50 & ~n39763 ;
  assign n39765 = ~x50 & ~n39764 ;
  assign n39766 = ~n39763 & ~n39764 ;
  assign n39767 = ~n39765 & ~n39766 ;
  assign n39768 = ~n39202 & ~n39213 ;
  assign n39769 = ~n39199 & ~n39768 ;
  assign n39770 = ~n39767 & ~n39769 ;
  assign n39771 = n39767 & n39769 ;
  assign n39772 = ~n39770 & ~n39771 ;
  assign n39773 = ~n39756 & n39772 ;
  assign n39774 = n39756 & ~n39772 ;
  assign n39775 = ~n39773 & ~n39774 ;
  assign n39776 = ~x100 & n14233 ;
  assign n39777 = ~x98 & n14876 ;
  assign n39778 = ~x99 & n14228 ;
  assign n39779 = ~n39777 & ~n39778 ;
  assign n39780 = ~n39776 & n39779 ;
  assign n39781 = n9338 & n14236 ;
  assign n39782 = n39780 & ~n39781 ;
  assign n39783 = ~x47 & ~n39782 ;
  assign n39784 = ~x47 & ~n39783 ;
  assign n39785 = ~n39782 & ~n39783 ;
  assign n39786 = ~n39784 & ~n39785 ;
  assign n39787 = ~n39775 & ~n39786 ;
  assign n39788 = n39775 & n39786 ;
  assign n39789 = ~n39787 & ~n39788 ;
  assign n39790 = n39672 & ~n39789 ;
  assign n39791 = ~n39672 & n39789 ;
  assign n39792 = ~n39790 & ~n39791 ;
  assign n39793 = ~x103 & n12506 ;
  assign n39794 = ~x101 & n13131 ;
  assign n39795 = ~x102 & n12501 ;
  assign n39796 = ~n39794 & ~n39795 ;
  assign n39797 = ~n39793 & n39796 ;
  assign n39798 = n10833 & n12509 ;
  assign n39799 = n39797 & ~n39798 ;
  assign n39800 = ~x44 & ~n39799 ;
  assign n39801 = ~x44 & ~n39800 ;
  assign n39802 = ~n39799 & ~n39800 ;
  assign n39803 = ~n39801 & ~n39802 ;
  assign n39804 = n39792 & ~n39803 ;
  assign n39805 = n39792 & ~n39804 ;
  assign n39806 = ~n39803 & ~n39804 ;
  assign n39807 = ~n39805 & ~n39806 ;
  assign n39808 = ~n39671 & n39807 ;
  assign n39809 = n39671 & ~n39807 ;
  assign n39810 = ~n39808 & ~n39809 ;
  assign n39811 = ~x106 & n10905 ;
  assign n39812 = ~x104 & n11466 ;
  assign n39813 = ~x105 & n10900 ;
  assign n39814 = ~n39812 & ~n39813 ;
  assign n39815 = ~n39811 & n39814 ;
  assign n39816 = n10908 & n12447 ;
  assign n39817 = n39815 & ~n39816 ;
  assign n39818 = ~x41 & ~n39817 ;
  assign n39819 = ~x41 & ~n39818 ;
  assign n39820 = ~n39817 & ~n39818 ;
  assign n39821 = ~n39819 & ~n39820 ;
  assign n39822 = ~n39810 & ~n39821 ;
  assign n39823 = n39810 & n39821 ;
  assign n39824 = ~n39822 & ~n39823 ;
  assign n39825 = n39669 & ~n39824 ;
  assign n39826 = ~n39669 & n39824 ;
  assign n39827 = ~n39825 & ~n39826 ;
  assign n39828 = ~x109 & n9433 ;
  assign n39829 = ~x107 & n9915 ;
  assign n39830 = ~x108 & n9428 ;
  assign n39831 = ~n39829 & ~n39830 ;
  assign n39832 = ~n39828 & n39831 ;
  assign n39833 = n9436 & n14177 ;
  assign n39834 = n39832 & ~n39833 ;
  assign n39835 = ~x38 & ~n39834 ;
  assign n39836 = ~x38 & ~n39835 ;
  assign n39837 = ~n39834 & ~n39835 ;
  assign n39838 = ~n39836 & ~n39837 ;
  assign n39839 = n39827 & ~n39838 ;
  assign n39840 = n39827 & ~n39839 ;
  assign n39841 = ~n39838 & ~n39839 ;
  assign n39842 = ~n39840 & ~n39841 ;
  assign n39843 = ~n39261 & ~n39264 ;
  assign n39844 = n39842 & n39843 ;
  assign n39845 = ~n39842 & ~n39843 ;
  assign n39846 = ~n39844 & ~n39845 ;
  assign n39847 = ~x112 & n8006 ;
  assign n39848 = ~x110 & n8474 ;
  assign n39849 = ~x111 & n8001 ;
  assign n39850 = ~n39848 & ~n39849 ;
  assign n39851 = ~n39847 & n39850 ;
  assign n39852 = n8009 & n15744 ;
  assign n39853 = n39851 & ~n39852 ;
  assign n39854 = ~x35 & ~n39853 ;
  assign n39855 = ~x35 & ~n39854 ;
  assign n39856 = ~n39853 & ~n39854 ;
  assign n39857 = ~n39855 & ~n39856 ;
  assign n39858 = n39846 & ~n39857 ;
  assign n39859 = n39846 & ~n39858 ;
  assign n39860 = ~n39857 & ~n39858 ;
  assign n39861 = ~n39859 & ~n39860 ;
  assign n39862 = ~n39267 & ~n39281 ;
  assign n39863 = n39861 & n39862 ;
  assign n39864 = ~n39861 & ~n39862 ;
  assign n39865 = ~n39863 & ~n39864 ;
  assign n39866 = ~x115 & n6725 ;
  assign n39867 = ~x113 & n7129 ;
  assign n39868 = ~x114 & n6720 ;
  assign n39869 = ~n39867 & ~n39868 ;
  assign n39870 = ~n39866 & n39869 ;
  assign n39871 = n6728 & n17683 ;
  assign n39872 = n39870 & ~n39871 ;
  assign n39873 = ~x32 & ~n39872 ;
  assign n39874 = ~x32 & ~n39873 ;
  assign n39875 = ~n39872 & ~n39873 ;
  assign n39876 = ~n39874 & ~n39875 ;
  assign n39877 = ~n39093 & ~n39285 ;
  assign n39878 = ~n39876 & ~n39877 ;
  assign n39879 = n39876 & n39877 ;
  assign n39880 = ~n39878 & ~n39879 ;
  assign n39881 = n39865 & n39880 ;
  assign n39882 = n39865 & ~n39881 ;
  assign n39883 = n39880 & ~n39881 ;
  assign n39884 = ~n39882 & ~n39883 ;
  assign n39885 = n39668 & ~n39884 ;
  assign n39886 = n39668 & ~n39885 ;
  assign n39887 = ~n39884 & ~n39885 ;
  assign n39888 = ~n39886 & ~n39887 ;
  assign n39889 = ~x121 & n4531 ;
  assign n39890 = ~x119 & n4847 ;
  assign n39891 = ~x120 & n4526 ;
  assign n39892 = ~n39890 & ~n39891 ;
  assign n39893 = ~n39889 & n39892 ;
  assign n39894 = n4534 & n22229 ;
  assign n39895 = n39893 & ~n39894 ;
  assign n39896 = ~x26 & ~n39895 ;
  assign n39897 = ~x26 & ~n39896 ;
  assign n39898 = ~n39895 & ~n39896 ;
  assign n39899 = ~n39897 & ~n39898 ;
  assign n39900 = ~n39062 & ~n39293 ;
  assign n39901 = ~n39899 & ~n39900 ;
  assign n39902 = n39899 & n39900 ;
  assign n39903 = ~n39901 & ~n39902 ;
  assign n39904 = ~n39888 & n39903 ;
  assign n39905 = ~n39888 & ~n39904 ;
  assign n39906 = n39903 & ~n39904 ;
  assign n39907 = ~n39905 & ~n39906 ;
  assign n39908 = n39653 & ~n39907 ;
  assign n39909 = n39653 & ~n39908 ;
  assign n39910 = ~n39907 & ~n39908 ;
  assign n39911 = ~n39909 & ~n39910 ;
  assign n39912 = ~n39638 & n39911 ;
  assign n39913 = n39638 & ~n39911 ;
  assign n39914 = ~n39912 & ~n39913 ;
  assign n39915 = ~n39622 & ~n39914 ;
  assign n39916 = ~n39622 & ~n39915 ;
  assign n39917 = ~n39914 & ~n39915 ;
  assign n39918 = ~n39916 & ~n39917 ;
  assign n39919 = ~n39621 & ~n39918 ;
  assign n39920 = n39621 & ~n39917 ;
  assign n39921 = ~n39916 & n39920 ;
  assign n39922 = ~n39919 & ~n39921 ;
  assign n39925 = ~n39922 & ~x209 ;
  assign n39926 = ~n39924 & ~n39925 ;
  assign n39927 = ~n39613 & ~n39617 ;
  assign n39928 = ~n39336 & ~n39609 ;
  assign n39929 = ~n39333 & ~n39928 ;
  assign n39930 = x125 & n3589 ;
  assign n39931 = x123 & n3878 ;
  assign n39932 = x124 & n3584 ;
  assign n39933 = ~n39931 & ~n39932 ;
  assign n39934 = ~n39930 & n39933 ;
  assign n39935 = n3592 & n24935 ;
  assign n39936 = n39934 & ~n39935 ;
  assign n39937 = x23 & ~n39936 ;
  assign n39938 = x23 & ~n39937 ;
  assign n39939 = ~n39936 & ~n39937 ;
  assign n39940 = ~n39938 & ~n39939 ;
  assign n39941 = ~n39599 & ~n39602 ;
  assign n39942 = n39940 & n39941 ;
  assign n39943 = ~n39940 & ~n39941 ;
  assign n39944 = ~n39942 & ~n39943 ;
  assign n39945 = x122 & n4531 ;
  assign n39946 = x120 & n4847 ;
  assign n39947 = x121 & n4526 ;
  assign n39948 = ~n39946 & ~n39947 ;
  assign n39949 = ~n39945 & n39948 ;
  assign n39950 = n4534 & n22622 ;
  assign n39951 = n39949 & ~n39950 ;
  assign n39952 = x26 & ~n39951 ;
  assign n39953 = x26 & ~n39952 ;
  assign n39954 = ~n39951 & ~n39952 ;
  assign n39955 = ~n39953 & ~n39954 ;
  assign n39956 = ~n39365 & ~n39583 ;
  assign n39957 = n39955 & n39956 ;
  assign n39958 = ~n39955 & ~n39956 ;
  assign n39959 = ~n39957 & ~n39958 ;
  assign n39960 = x119 & n5560 ;
  assign n39961 = x117 & n5943 ;
  assign n39962 = x118 & n5555 ;
  assign n39963 = ~n39961 & ~n39962 ;
  assign n39964 = ~n39960 & n39963 ;
  assign n39965 = n5563 & n20423 ;
  assign n39966 = n39964 & ~n39965 ;
  assign n39967 = x29 & ~n39966 ;
  assign n39968 = x29 & ~n39967 ;
  assign n39969 = ~n39966 & ~n39967 ;
  assign n39970 = ~n39968 & ~n39969 ;
  assign n39971 = ~n39576 & ~n39579 ;
  assign n39972 = n39970 & n39971 ;
  assign n39973 = ~n39970 & ~n39971 ;
  assign n39974 = ~n39972 & ~n39973 ;
  assign n39975 = x116 & n6725 ;
  assign n39976 = x114 & n7129 ;
  assign n39977 = x115 & n6720 ;
  assign n39978 = ~n39976 & ~n39977 ;
  assign n39979 = ~n39975 & n39978 ;
  assign n39980 = n6728 & n18336 ;
  assign n39981 = n39979 & ~n39980 ;
  assign n39982 = x32 & ~n39981 ;
  assign n39983 = x32 & ~n39982 ;
  assign n39984 = ~n39981 & ~n39982 ;
  assign n39985 = ~n39983 & ~n39984 ;
  assign n39986 = ~n39556 & ~n39562 ;
  assign n39987 = n39985 & n39986 ;
  assign n39988 = ~n39985 & ~n39986 ;
  assign n39989 = ~n39987 & ~n39988 ;
  assign n39990 = ~n39369 & ~n39505 ;
  assign n39991 = ~n39502 & ~n39990 ;
  assign n39992 = x104 & n12506 ;
  assign n39993 = x102 & n13131 ;
  assign n39994 = x103 & n12501 ;
  assign n39995 = ~n39993 & ~n39994 ;
  assign n39996 = ~n39992 & n39995 ;
  assign n39997 = n11116 & n12509 ;
  assign n39998 = n39996 & ~n39997 ;
  assign n39999 = x44 & ~n39998 ;
  assign n40000 = x44 & ~n39999 ;
  assign n40001 = ~n39998 & ~n39999 ;
  assign n40002 = ~n40000 & ~n40001 ;
  assign n40003 = ~n39485 & ~n39489 ;
  assign n40004 = ~n39412 & ~n39414 ;
  assign n40005 = x82 & n27024 ;
  assign n40006 = x83 & ~n26217 ;
  assign n40007 = ~n40005 & ~n40006 ;
  assign n40008 = ~n39386 & ~n39389 ;
  assign n40009 = ~n40007 & n40008 ;
  assign n40010 = n40007 & ~n40008 ;
  assign n40011 = ~n40009 & ~n40010 ;
  assign n40012 = x86 & n24612 ;
  assign n40013 = x84 & n25390 ;
  assign n40014 = x85 & n24607 ;
  assign n40015 = ~n40013 & ~n40014 ;
  assign n40016 = ~n40012 & n40015 ;
  assign n40017 = n3686 & n24615 ;
  assign n40018 = n40016 & ~n40017 ;
  assign n40019 = x62 & ~n40018 ;
  assign n40020 = x62 & ~n40019 ;
  assign n40021 = ~n40018 & ~n40019 ;
  assign n40022 = ~n40020 & ~n40021 ;
  assign n40023 = ~n40011 & n40022 ;
  assign n40024 = n40011 & ~n40022 ;
  assign n40025 = ~n40023 & ~n40024 ;
  assign n40026 = ~n39392 & ~n39396 ;
  assign n40027 = n40025 & ~n40026 ;
  assign n40028 = ~n40025 & n40026 ;
  assign n40029 = ~n40027 & ~n40028 ;
  assign n40030 = x89 & n22325 ;
  assign n40031 = x87 & n23066 ;
  assign n40032 = x88 & n22320 ;
  assign n40033 = ~n40031 & ~n40032 ;
  assign n40034 = ~n40030 & n40033 ;
  assign n40035 = n4488 & n22328 ;
  assign n40036 = n40034 & ~n40035 ;
  assign n40037 = x59 & ~n40036 ;
  assign n40038 = x59 & ~n40037 ;
  assign n40039 = ~n40036 & ~n40037 ;
  assign n40040 = ~n40038 & ~n40039 ;
  assign n40041 = n40029 & ~n40040 ;
  assign n40042 = n40029 & ~n40041 ;
  assign n40043 = ~n40040 & ~n40041 ;
  assign n40044 = ~n40042 & ~n40043 ;
  assign n40045 = ~n40004 & n40044 ;
  assign n40046 = n40004 & ~n40044 ;
  assign n40047 = ~n40045 & ~n40046 ;
  assign n40048 = x92 & n20143 ;
  assign n40049 = x90 & n20854 ;
  assign n40050 = x91 & n20138 ;
  assign n40051 = ~n40049 & ~n40050 ;
  assign n40052 = ~n40048 & n40051 ;
  assign n40053 = n5710 & n20146 ;
  assign n40054 = n40052 & ~n40053 ;
  assign n40055 = x56 & ~n40054 ;
  assign n40056 = x56 & ~n40055 ;
  assign n40057 = ~n40054 & ~n40055 ;
  assign n40058 = ~n40056 & ~n40057 ;
  assign n40059 = n40047 & n40058 ;
  assign n40060 = ~n40047 & ~n40058 ;
  assign n40061 = ~n40059 & ~n40060 ;
  assign n40062 = ~n39428 & ~n39434 ;
  assign n40063 = n40061 & ~n40062 ;
  assign n40064 = ~n40061 & n40062 ;
  assign n40065 = ~n40063 & ~n40064 ;
  assign n40066 = x95 & n18025 ;
  assign n40067 = x93 & n18764 ;
  assign n40068 = x94 & n18020 ;
  assign n40069 = ~n40067 & ~n40068 ;
  assign n40070 = ~n40066 & n40069 ;
  assign n40071 = n6894 & n18028 ;
  assign n40072 = n40070 & ~n40071 ;
  assign n40073 = x53 & ~n40072 ;
  assign n40074 = x53 & ~n40073 ;
  assign n40075 = ~n40072 & ~n40073 ;
  assign n40076 = ~n40074 & ~n40075 ;
  assign n40077 = n40065 & ~n40076 ;
  assign n40078 = n40065 & ~n40077 ;
  assign n40079 = ~n40076 & ~n40077 ;
  assign n40080 = ~n40078 & ~n40079 ;
  assign n40081 = ~n39447 & ~n39453 ;
  assign n40082 = n40080 & n40081 ;
  assign n40083 = ~n40080 & ~n40081 ;
  assign n40084 = ~n40082 & ~n40083 ;
  assign n40085 = x98 & n16076 ;
  assign n40086 = x96 & n16756 ;
  assign n40087 = x97 & n16071 ;
  assign n40088 = ~n40086 & ~n40087 ;
  assign n40089 = ~n40085 & n40088 ;
  assign n40090 = n8196 & n16079 ;
  assign n40091 = n40089 & ~n40090 ;
  assign n40092 = x50 & ~n40091 ;
  assign n40093 = x50 & ~n40092 ;
  assign n40094 = ~n40091 & ~n40092 ;
  assign n40095 = ~n40093 & ~n40094 ;
  assign n40096 = n40084 & ~n40095 ;
  assign n40097 = n40084 & ~n40096 ;
  assign n40098 = ~n40095 & ~n40096 ;
  assign n40099 = ~n40097 & ~n40098 ;
  assign n40100 = n39454 & n39470 ;
  assign n40101 = ~n39468 & ~n40100 ;
  assign n40102 = n40099 & n40101 ;
  assign n40103 = ~n40099 & ~n40101 ;
  assign n40104 = ~n40102 & ~n40103 ;
  assign n40105 = x101 & n14233 ;
  assign n40106 = x99 & n14876 ;
  assign n40107 = x100 & n14228 ;
  assign n40108 = ~n40106 & ~n40107 ;
  assign n40109 = ~n40105 & n40108 ;
  assign n40110 = n9601 & n14236 ;
  assign n40111 = n40109 & ~n40110 ;
  assign n40112 = x47 & ~n40111 ;
  assign n40113 = x47 & ~n40112 ;
  assign n40114 = ~n40111 & ~n40112 ;
  assign n40115 = ~n40113 & ~n40114 ;
  assign n40116 = ~n40104 & n40115 ;
  assign n40117 = n40104 & ~n40115 ;
  assign n40118 = ~n40116 & ~n40117 ;
  assign n40119 = ~n40003 & n40118 ;
  assign n40120 = ~n40003 & ~n40119 ;
  assign n40121 = n40118 & ~n40119 ;
  assign n40122 = ~n40120 & ~n40121 ;
  assign n40123 = ~n40002 & ~n40122 ;
  assign n40124 = n40002 & ~n40121 ;
  assign n40125 = ~n40120 & n40124 ;
  assign n40126 = ~n40123 & ~n40125 ;
  assign n40127 = ~n39991 & n40126 ;
  assign n40128 = n39991 & ~n40126 ;
  assign n40129 = ~n40127 & ~n40128 ;
  assign n40130 = x107 & n10905 ;
  assign n40131 = x105 & n11466 ;
  assign n40132 = x106 & n10900 ;
  assign n40133 = ~n40131 & ~n40132 ;
  assign n40134 = ~n40130 & n40133 ;
  assign n40135 = n10908 & n12749 ;
  assign n40136 = n40134 & ~n40135 ;
  assign n40137 = x41 & ~n40136 ;
  assign n40138 = x41 & ~n40137 ;
  assign n40139 = ~n40136 & ~n40137 ;
  assign n40140 = ~n40138 & ~n40139 ;
  assign n40141 = n40129 & ~n40140 ;
  assign n40142 = n40129 & ~n40141 ;
  assign n40143 = ~n40140 & ~n40141 ;
  assign n40144 = ~n40142 & ~n40143 ;
  assign n40145 = ~n39520 & ~n39524 ;
  assign n40146 = n40144 & n40145 ;
  assign n40147 = ~n40144 & ~n40145 ;
  assign n40148 = ~n40146 & ~n40147 ;
  assign n40149 = x110 & n9433 ;
  assign n40150 = x108 & n9915 ;
  assign n40151 = x109 & n9428 ;
  assign n40152 = ~n40150 & ~n40151 ;
  assign n40153 = ~n40149 & n40152 ;
  assign n40154 = n9436 & n14497 ;
  assign n40155 = n40153 & ~n40154 ;
  assign n40156 = x38 & ~n40155 ;
  assign n40157 = x38 & ~n40156 ;
  assign n40158 = ~n40155 & ~n40156 ;
  assign n40159 = ~n40157 & ~n40158 ;
  assign n40160 = n40148 & ~n40159 ;
  assign n40161 = n40148 & ~n40160 ;
  assign n40162 = ~n40159 & ~n40160 ;
  assign n40163 = ~n40161 & ~n40162 ;
  assign n40164 = ~n39537 & ~n39543 ;
  assign n40165 = n40163 & n40164 ;
  assign n40166 = ~n40163 & ~n40164 ;
  assign n40167 = ~n40165 & ~n40166 ;
  assign n40168 = x113 & n8006 ;
  assign n40169 = x111 & n8474 ;
  assign n40170 = x112 & n8001 ;
  assign n40171 = ~n40169 & ~n40170 ;
  assign n40172 = ~n40168 & n40171 ;
  assign n40173 = n8009 & n16361 ;
  assign n40174 = n40172 & ~n40173 ;
  assign n40175 = x35 & ~n40174 ;
  assign n40176 = x35 & ~n40175 ;
  assign n40177 = ~n40174 & ~n40175 ;
  assign n40178 = ~n40176 & ~n40177 ;
  assign n40179 = n40167 & ~n40178 ;
  assign n40180 = n40167 & ~n40179 ;
  assign n40181 = ~n40178 & ~n40179 ;
  assign n40182 = ~n40180 & ~n40181 ;
  assign n40183 = n39989 & ~n40182 ;
  assign n40184 = ~n39989 & n40182 ;
  assign n40185 = n39974 & ~n40184 ;
  assign n40186 = ~n40183 & n40185 ;
  assign n40187 = n39974 & ~n40186 ;
  assign n40188 = ~n40184 & ~n40186 ;
  assign n40189 = ~n40183 & n40188 ;
  assign n40190 = ~n40187 & ~n40189 ;
  assign n40191 = n39959 & ~n40190 ;
  assign n40192 = ~n39959 & n40190 ;
  assign n40193 = n39944 & ~n40192 ;
  assign n40194 = ~n40191 & n40193 ;
  assign n40195 = n39944 & ~n40194 ;
  assign n40196 = ~n40192 & ~n40194 ;
  assign n40197 = ~n40191 & n40196 ;
  assign n40198 = ~n40195 & ~n40197 ;
  assign n40199 = ~n39350 & ~n39606 ;
  assign n40200 = x126 & n3020 ;
  assign n40201 = x127 & n2746 ;
  assign n40202 = ~n40200 & ~n40201 ;
  assign n40203 = ~n2754 & n40202 ;
  assign n40204 = n26965 & n40202 ;
  assign n40205 = ~n40203 & ~n40204 ;
  assign n40206 = x20 & ~n40205 ;
  assign n40207 = ~x20 & n40205 ;
  assign n40208 = ~n40206 & ~n40207 ;
  assign n40209 = ~n40199 & ~n40208 ;
  assign n40210 = ~n40199 & ~n40209 ;
  assign n40211 = ~n40208 & ~n40209 ;
  assign n40212 = ~n40210 & ~n40211 ;
  assign n40213 = ~n40198 & ~n40212 ;
  assign n40214 = n40198 & ~n40211 ;
  assign n40215 = ~n40210 & n40214 ;
  assign n40216 = ~n40213 & ~n40215 ;
  assign n40217 = ~n39929 & n40216 ;
  assign n40218 = ~n39929 & ~n40217 ;
  assign n40219 = n40216 & ~n40217 ;
  assign n40220 = ~n40218 & ~n40219 ;
  assign n40221 = ~n39927 & ~n40220 ;
  assign n40222 = n39927 & ~n40219 ;
  assign n40223 = ~n40218 & n40222 ;
  assign n40224 = ~n40221 & ~n40223 ;
  assign n40524 = n40224 & x210 ;
  assign n40225 = ~n39915 & ~n39919 ;
  assign n40226 = ~n39638 & ~n39911 ;
  assign n40227 = ~n39635 & ~n40226 ;
  assign n40228 = ~x125 & n3589 ;
  assign n40229 = ~x123 & n3878 ;
  assign n40230 = ~x124 & n3584 ;
  assign n40231 = ~n40229 & ~n40230 ;
  assign n40232 = ~n40228 & n40231 ;
  assign n40233 = n3592 & n25330 ;
  assign n40234 = n40232 & ~n40233 ;
  assign n40235 = ~x23 & ~n40234 ;
  assign n40236 = ~x23 & ~n40235 ;
  assign n40237 = ~n40234 & ~n40235 ;
  assign n40238 = ~n40236 & ~n40237 ;
  assign n40239 = ~n39901 & ~n39904 ;
  assign n40240 = n40238 & n40239 ;
  assign n40241 = ~n40238 & ~n40239 ;
  assign n40242 = ~n40240 & ~n40241 ;
  assign n40243 = ~x122 & n4531 ;
  assign n40244 = ~x120 & n4847 ;
  assign n40245 = ~x121 & n4526 ;
  assign n40246 = ~n40244 & ~n40245 ;
  assign n40247 = ~n40243 & n40246 ;
  assign n40248 = n4534 & n22998 ;
  assign n40249 = n40247 & ~n40248 ;
  assign n40250 = ~x26 & ~n40249 ;
  assign n40251 = ~x26 & ~n40250 ;
  assign n40252 = ~n40249 & ~n40250 ;
  assign n40253 = ~n40251 & ~n40252 ;
  assign n40254 = ~n39667 & ~n39885 ;
  assign n40255 = n40253 & n40254 ;
  assign n40256 = ~n40253 & ~n40254 ;
  assign n40257 = ~n40255 & ~n40256 ;
  assign n40258 = ~x119 & n5560 ;
  assign n40259 = ~x117 & n5943 ;
  assign n40260 = ~x118 & n5555 ;
  assign n40261 = ~n40259 & ~n40260 ;
  assign n40262 = ~n40258 & n40261 ;
  assign n40263 = n5563 & n20778 ;
  assign n40264 = n40262 & ~n40263 ;
  assign n40265 = ~x29 & ~n40264 ;
  assign n40266 = ~x29 & ~n40265 ;
  assign n40267 = ~n40264 & ~n40265 ;
  assign n40268 = ~n40266 & ~n40267 ;
  assign n40269 = ~n39878 & ~n39881 ;
  assign n40270 = n40268 & n40269 ;
  assign n40271 = ~n40268 & ~n40269 ;
  assign n40272 = ~n40270 & ~n40271 ;
  assign n40273 = ~x116 & n6725 ;
  assign n40274 = ~x114 & n7129 ;
  assign n40275 = ~x115 & n6720 ;
  assign n40276 = ~n40274 & ~n40275 ;
  assign n40277 = ~n40273 & n40276 ;
  assign n40278 = n6728 & n18678 ;
  assign n40279 = n40277 & ~n40278 ;
  assign n40280 = ~x32 & ~n40279 ;
  assign n40281 = ~x32 & ~n40280 ;
  assign n40282 = ~n40279 & ~n40280 ;
  assign n40283 = ~n40281 & ~n40282 ;
  assign n40284 = ~n39858 & ~n39864 ;
  assign n40285 = n40283 & n40284 ;
  assign n40286 = ~n40283 & ~n40284 ;
  assign n40287 = ~n40285 & ~n40286 ;
  assign n40288 = ~n39671 & ~n39807 ;
  assign n40289 = ~n39804 & ~n40288 ;
  assign n40290 = ~x104 & n12506 ;
  assign n40291 = ~x102 & n13131 ;
  assign n40292 = ~x103 & n12501 ;
  assign n40293 = ~n40291 & ~n40292 ;
  assign n40294 = ~n40290 & n40293 ;
  assign n40295 = n11380 & n12509 ;
  assign n40296 = n40294 & ~n40295 ;
  assign n40297 = ~x44 & ~n40296 ;
  assign n40298 = ~x44 & ~n40297 ;
  assign n40299 = ~n40296 & ~n40297 ;
  assign n40300 = ~n40298 & ~n40299 ;
  assign n40301 = ~n39787 & ~n39791 ;
  assign n40302 = ~n39714 & ~n39716 ;
  assign n40303 = ~x82 & n27427 ;
  assign n40304 = ~x83 & ~n26217 ;
  assign n40305 = ~n40303 & ~n40304 ;
  assign n40306 = ~n39688 & ~n39691 ;
  assign n40307 = ~n40305 & n40306 ;
  assign n40308 = n40305 & ~n40306 ;
  assign n40309 = ~n40307 & ~n40308 ;
  assign n40310 = ~x86 & n24612 ;
  assign n40311 = ~x84 & n25390 ;
  assign n40312 = ~x85 & n24607 ;
  assign n40313 = ~n40311 & ~n40312 ;
  assign n40314 = ~n40310 & n40313 ;
  assign n40315 = n3832 & n24615 ;
  assign n40316 = n40314 & ~n40315 ;
  assign n40317 = ~x62 & ~n40316 ;
  assign n40318 = ~x62 & ~n40317 ;
  assign n40319 = ~n40316 & ~n40317 ;
  assign n40320 = ~n40318 & ~n40319 ;
  assign n40321 = ~n40309 & n40320 ;
  assign n40322 = n40309 & ~n40320 ;
  assign n40323 = ~n40321 & ~n40322 ;
  assign n40324 = ~n39694 & ~n39698 ;
  assign n40325 = n40323 & ~n40324 ;
  assign n40326 = ~n40323 & n40324 ;
  assign n40327 = ~n40325 & ~n40326 ;
  assign n40328 = ~x89 & n22325 ;
  assign n40329 = ~x87 & n23066 ;
  assign n40330 = ~x88 & n22320 ;
  assign n40331 = ~n40329 & ~n40330 ;
  assign n40332 = ~n40328 & n40331 ;
  assign n40333 = n4664 & n22328 ;
  assign n40334 = n40332 & ~n40333 ;
  assign n40335 = ~x59 & ~n40334 ;
  assign n40336 = ~x59 & ~n40335 ;
  assign n40337 = ~n40334 & ~n40335 ;
  assign n40338 = ~n40336 & ~n40337 ;
  assign n40339 = n40327 & ~n40338 ;
  assign n40340 = n40327 & ~n40339 ;
  assign n40341 = ~n40338 & ~n40339 ;
  assign n40342 = ~n40340 & ~n40341 ;
  assign n40343 = ~n40302 & n40342 ;
  assign n40344 = n40302 & ~n40342 ;
  assign n40345 = ~n40343 & ~n40344 ;
  assign n40346 = ~x92 & n20143 ;
  assign n40347 = ~x90 & n20854 ;
  assign n40348 = ~x91 & n20138 ;
  assign n40349 = ~n40347 & ~n40348 ;
  assign n40350 = ~n40346 & n40349 ;
  assign n40351 = n5896 & n20146 ;
  assign n40352 = n40350 & ~n40351 ;
  assign n40353 = ~x56 & ~n40352 ;
  assign n40354 = ~x56 & ~n40353 ;
  assign n40355 = ~n40352 & ~n40353 ;
  assign n40356 = ~n40354 & ~n40355 ;
  assign n40357 = n40345 & n40356 ;
  assign n40358 = ~n40345 & ~n40356 ;
  assign n40359 = ~n40357 & ~n40358 ;
  assign n40360 = ~n39730 & ~n39736 ;
  assign n40361 = n40359 & ~n40360 ;
  assign n40362 = ~n40359 & n40360 ;
  assign n40363 = ~n40361 & ~n40362 ;
  assign n40364 = ~x95 & n18025 ;
  assign n40365 = ~x93 & n18764 ;
  assign n40366 = ~x94 & n18020 ;
  assign n40367 = ~n40365 & ~n40366 ;
  assign n40368 = ~n40364 & n40367 ;
  assign n40369 = n7100 & n18028 ;
  assign n40370 = n40368 & ~n40369 ;
  assign n40371 = ~x53 & ~n40370 ;
  assign n40372 = ~x53 & ~n40371 ;
  assign n40373 = ~n40370 & ~n40371 ;
  assign n40374 = ~n40372 & ~n40373 ;
  assign n40375 = n40363 & ~n40374 ;
  assign n40376 = n40363 & ~n40375 ;
  assign n40377 = ~n40374 & ~n40375 ;
  assign n40378 = ~n40376 & ~n40377 ;
  assign n40379 = ~n39749 & ~n39755 ;
  assign n40380 = n40378 & n40379 ;
  assign n40381 = ~n40378 & ~n40379 ;
  assign n40382 = ~n40380 & ~n40381 ;
  assign n40383 = ~x98 & n16076 ;
  assign n40384 = ~x96 & n16756 ;
  assign n40385 = ~x97 & n16071 ;
  assign n40386 = ~n40384 & ~n40385 ;
  assign n40387 = ~n40383 & n40386 ;
  assign n40388 = n8426 & n16079 ;
  assign n40389 = n40387 & ~n40388 ;
  assign n40390 = ~x50 & ~n40389 ;
  assign n40391 = ~x50 & ~n40390 ;
  assign n40392 = ~n40389 & ~n40390 ;
  assign n40393 = ~n40391 & ~n40392 ;
  assign n40394 = n40382 & ~n40393 ;
  assign n40395 = n40382 & ~n40394 ;
  assign n40396 = ~n40393 & ~n40394 ;
  assign n40397 = ~n40395 & ~n40396 ;
  assign n40398 = n39756 & n39772 ;
  assign n40399 = ~n39770 & ~n40398 ;
  assign n40400 = n40397 & n40399 ;
  assign n40401 = ~n40397 & ~n40399 ;
  assign n40402 = ~n40400 & ~n40401 ;
  assign n40403 = ~x101 & n14233 ;
  assign n40404 = ~x99 & n14876 ;
  assign n40405 = ~x100 & n14228 ;
  assign n40406 = ~n40404 & ~n40405 ;
  assign n40407 = ~n40403 & n40406 ;
  assign n40408 = n9844 & n14236 ;
  assign n40409 = n40407 & ~n40408 ;
  assign n40410 = ~x47 & ~n40409 ;
  assign n40411 = ~x47 & ~n40410 ;
  assign n40412 = ~n40409 & ~n40410 ;
  assign n40413 = ~n40411 & ~n40412 ;
  assign n40414 = ~n40402 & n40413 ;
  assign n40415 = n40402 & ~n40413 ;
  assign n40416 = ~n40414 & ~n40415 ;
  assign n40417 = ~n40301 & n40416 ;
  assign n40418 = ~n40301 & ~n40417 ;
  assign n40419 = n40416 & ~n40417 ;
  assign n40420 = ~n40418 & ~n40419 ;
  assign n40421 = ~n40300 & ~n40420 ;
  assign n40422 = n40300 & ~n40419 ;
  assign n40423 = ~n40418 & n40422 ;
  assign n40424 = ~n40421 & ~n40423 ;
  assign n40425 = ~n40289 & n40424 ;
  assign n40426 = n40289 & ~n40424 ;
  assign n40427 = ~n40425 & ~n40426 ;
  assign n40428 = ~x107 & n10905 ;
  assign n40429 = ~x105 & n11466 ;
  assign n40430 = ~x106 & n10900 ;
  assign n40431 = ~n40429 & ~n40430 ;
  assign n40432 = ~n40428 & n40431 ;
  assign n40433 = n10908 & n13034 ;
  assign n40434 = n40432 & ~n40433 ;
  assign n40435 = ~x41 & ~n40434 ;
  assign n40436 = ~x41 & ~n40435 ;
  assign n40437 = ~n40434 & ~n40435 ;
  assign n40438 = ~n40436 & ~n40437 ;
  assign n40439 = n40427 & ~n40438 ;
  assign n40440 = n40427 & ~n40439 ;
  assign n40441 = ~n40438 & ~n40439 ;
  assign n40442 = ~n40440 & ~n40441 ;
  assign n40443 = ~n39822 & ~n39826 ;
  assign n40444 = n40442 & n40443 ;
  assign n40445 = ~n40442 & ~n40443 ;
  assign n40446 = ~n40444 & ~n40445 ;
  assign n40447 = ~x110 & n9433 ;
  assign n40448 = ~x108 & n9915 ;
  assign n40449 = ~x109 & n9428 ;
  assign n40450 = ~n40448 & ~n40449 ;
  assign n40451 = ~n40447 & n40450 ;
  assign n40452 = n9436 & n14802 ;
  assign n40453 = n40451 & ~n40452 ;
  assign n40454 = ~x38 & ~n40453 ;
  assign n40455 = ~x38 & ~n40454 ;
  assign n40456 = ~n40453 & ~n40454 ;
  assign n40457 = ~n40455 & ~n40456 ;
  assign n40458 = n40446 & ~n40457 ;
  assign n40459 = n40446 & ~n40458 ;
  assign n40460 = ~n40457 & ~n40458 ;
  assign n40461 = ~n40459 & ~n40460 ;
  assign n40462 = ~n39839 & ~n39845 ;
  assign n40463 = n40461 & n40462 ;
  assign n40464 = ~n40461 & ~n40462 ;
  assign n40465 = ~n40463 & ~n40464 ;
  assign n40466 = ~x113 & n8006 ;
  assign n40467 = ~x111 & n8474 ;
  assign n40468 = ~x112 & n8001 ;
  assign n40469 = ~n40467 & ~n40468 ;
  assign n40470 = ~n40466 & n40469 ;
  assign n40471 = n8009 & n16684 ;
  assign n40472 = n40470 & ~n40471 ;
  assign n40473 = ~x35 & ~n40472 ;
  assign n40474 = ~x35 & ~n40473 ;
  assign n40475 = ~n40472 & ~n40473 ;
  assign n40476 = ~n40474 & ~n40475 ;
  assign n40477 = n40465 & ~n40476 ;
  assign n40478 = n40465 & ~n40477 ;
  assign n40479 = ~n40476 & ~n40477 ;
  assign n40480 = ~n40478 & ~n40479 ;
  assign n40481 = n40287 & ~n40480 ;
  assign n40482 = ~n40287 & n40480 ;
  assign n40483 = n40272 & ~n40482 ;
  assign n40484 = ~n40481 & n40483 ;
  assign n40485 = n40272 & ~n40484 ;
  assign n40486 = ~n40482 & ~n40484 ;
  assign n40487 = ~n40481 & n40486 ;
  assign n40488 = ~n40485 & ~n40487 ;
  assign n40489 = n40257 & ~n40488 ;
  assign n40490 = ~n40257 & n40488 ;
  assign n40491 = n40242 & ~n40490 ;
  assign n40492 = ~n40489 & n40491 ;
  assign n40493 = n40242 & ~n40492 ;
  assign n40494 = ~n40490 & ~n40492 ;
  assign n40495 = ~n40489 & n40494 ;
  assign n40496 = ~n40493 & ~n40495 ;
  assign n40497 = ~n39652 & ~n39908 ;
  assign n40498 = ~x126 & n3020 ;
  assign n40499 = ~x127 & n2746 ;
  assign n40500 = ~n40498 & ~n40499 ;
  assign n40501 = ~n2754 & n40500 ;
  assign n40502 = n27368 & n40500 ;
  assign n40503 = ~n40501 & ~n40502 ;
  assign n40504 = ~x20 & ~n40503 ;
  assign n40505 = x20 & n40503 ;
  assign n40506 = ~n40504 & ~n40505 ;
  assign n40507 = ~n40497 & ~n40506 ;
  assign n40508 = ~n40497 & ~n40507 ;
  assign n40509 = ~n40506 & ~n40507 ;
  assign n40510 = ~n40508 & ~n40509 ;
  assign n40511 = ~n40496 & ~n40510 ;
  assign n40512 = n40496 & ~n40509 ;
  assign n40513 = ~n40508 & n40512 ;
  assign n40514 = ~n40511 & ~n40513 ;
  assign n40515 = ~n40227 & n40514 ;
  assign n40516 = ~n40227 & ~n40515 ;
  assign n40517 = n40514 & ~n40515 ;
  assign n40518 = ~n40516 & ~n40517 ;
  assign n40519 = ~n40225 & ~n40518 ;
  assign n40520 = n40225 & ~n40517 ;
  assign n40521 = ~n40516 & n40520 ;
  assign n40522 = ~n40519 & ~n40521 ;
  assign n40525 = ~n40522 & ~x210 ;
  assign n40526 = ~n40524 & ~n40525 ;
  assign n40527 = ~n40217 & ~n40221 ;
  assign n40528 = ~n40209 & ~n40213 ;
  assign n40529 = ~n39943 & ~n40194 ;
  assign n40530 = x127 & n3020 ;
  assign n40531 = n2754 & n26962 ;
  assign n40532 = ~n40530 & ~n40531 ;
  assign n40533 = x20 & ~n40532 ;
  assign n40534 = x20 & ~n40533 ;
  assign n40535 = ~n40532 & ~n40533 ;
  assign n40536 = ~n40534 & ~n40535 ;
  assign n40537 = ~n40529 & ~n40536 ;
  assign n40538 = ~n40529 & ~n40537 ;
  assign n40539 = ~n40536 & ~n40537 ;
  assign n40540 = ~n40538 & ~n40539 ;
  assign n40541 = x126 & n3589 ;
  assign n40542 = x124 & n3878 ;
  assign n40543 = x125 & n3584 ;
  assign n40544 = ~n40542 & ~n40543 ;
  assign n40545 = ~n40541 & n40544 ;
  assign n40546 = n3592 & n25735 ;
  assign n40547 = n40545 & ~n40546 ;
  assign n40548 = x23 & ~n40547 ;
  assign n40549 = x23 & ~n40548 ;
  assign n40550 = ~n40547 & ~n40548 ;
  assign n40551 = ~n40549 & ~n40550 ;
  assign n40552 = ~n39958 & ~n40191 ;
  assign n40553 = ~n40551 & ~n40552 ;
  assign n40554 = ~n40551 & ~n40553 ;
  assign n40555 = ~n40552 & ~n40553 ;
  assign n40556 = ~n40554 & ~n40555 ;
  assign n40557 = x123 & n4531 ;
  assign n40558 = x121 & n4847 ;
  assign n40559 = x122 & n4526 ;
  assign n40560 = ~n40558 & ~n40559 ;
  assign n40561 = ~n40557 & n40560 ;
  assign n40562 = n4534 & n23382 ;
  assign n40563 = n40561 & ~n40562 ;
  assign n40564 = x26 & ~n40563 ;
  assign n40565 = x26 & ~n40564 ;
  assign n40566 = ~n40563 & ~n40564 ;
  assign n40567 = ~n40565 & ~n40566 ;
  assign n40568 = ~n39973 & ~n40186 ;
  assign n40569 = n40567 & n40568 ;
  assign n40570 = ~n40567 & ~n40568 ;
  assign n40571 = ~n40569 & ~n40570 ;
  assign n40572 = x120 & n5560 ;
  assign n40573 = x118 & n5943 ;
  assign n40574 = x119 & n5555 ;
  assign n40575 = ~n40573 & ~n40574 ;
  assign n40576 = ~n40572 & n40575 ;
  assign n40577 = n5563 & n21143 ;
  assign n40578 = n40576 & ~n40577 ;
  assign n40579 = x29 & ~n40578 ;
  assign n40580 = x29 & ~n40579 ;
  assign n40581 = ~n40578 & ~n40579 ;
  assign n40582 = ~n40580 & ~n40581 ;
  assign n40583 = ~n39988 & ~n40183 ;
  assign n40584 = ~n40582 & ~n40583 ;
  assign n40585 = ~n40582 & ~n40584 ;
  assign n40586 = ~n40583 & ~n40584 ;
  assign n40587 = ~n40585 & ~n40586 ;
  assign n40588 = x117 & n6725 ;
  assign n40589 = x115 & n7129 ;
  assign n40590 = x116 & n6720 ;
  assign n40591 = ~n40589 & ~n40590 ;
  assign n40592 = ~n40588 & n40591 ;
  assign n40593 = n6728 & n19026 ;
  assign n40594 = n40592 & ~n40593 ;
  assign n40595 = x32 & ~n40594 ;
  assign n40596 = x32 & ~n40595 ;
  assign n40597 = ~n40594 & ~n40595 ;
  assign n40598 = ~n40596 & ~n40597 ;
  assign n40599 = ~n40166 & ~n40179 ;
  assign n40600 = n40598 & n40599 ;
  assign n40601 = ~n40598 & ~n40599 ;
  assign n40602 = ~n40600 & ~n40601 ;
  assign n40603 = ~n40127 & ~n40141 ;
  assign n40604 = x108 & n10905 ;
  assign n40605 = x106 & n11466 ;
  assign n40606 = x107 & n10900 ;
  assign n40607 = ~n40605 & ~n40606 ;
  assign n40608 = ~n40604 & n40607 ;
  assign n40609 = n10908 & n13323 ;
  assign n40610 = n40608 & ~n40609 ;
  assign n40611 = x41 & ~n40610 ;
  assign n40612 = x41 & ~n40611 ;
  assign n40613 = ~n40610 & ~n40611 ;
  assign n40614 = ~n40612 & ~n40613 ;
  assign n40615 = ~n40119 & ~n40123 ;
  assign n40616 = x105 & n12506 ;
  assign n40617 = x103 & n13131 ;
  assign n40618 = x104 & n12501 ;
  assign n40619 = ~n40617 & ~n40618 ;
  assign n40620 = ~n40616 & n40619 ;
  assign n40621 = n11648 & n12509 ;
  assign n40622 = n40620 & ~n40621 ;
  assign n40623 = x44 & ~n40622 ;
  assign n40624 = x44 & ~n40623 ;
  assign n40625 = ~n40622 & ~n40623 ;
  assign n40626 = ~n40624 & ~n40625 ;
  assign n40627 = ~n40103 & ~n40117 ;
  assign n40628 = x102 & n14233 ;
  assign n40629 = x100 & n14876 ;
  assign n40630 = x101 & n14228 ;
  assign n40631 = ~n40629 & ~n40630 ;
  assign n40632 = ~n40628 & n40631 ;
  assign n40633 = n10092 & n14236 ;
  assign n40634 = n40632 & ~n40633 ;
  assign n40635 = x47 & ~n40634 ;
  assign n40636 = x47 & ~n40635 ;
  assign n40637 = ~n40634 & ~n40635 ;
  assign n40638 = ~n40636 & ~n40637 ;
  assign n40639 = ~n40083 & ~n40096 ;
  assign n40640 = x99 & n16076 ;
  assign n40641 = x97 & n16756 ;
  assign n40642 = x98 & n16071 ;
  assign n40643 = ~n40641 & ~n40642 ;
  assign n40644 = ~n40640 & n40643 ;
  assign n40645 = n8660 & n16079 ;
  assign n40646 = n40644 & ~n40645 ;
  assign n40647 = x50 & ~n40646 ;
  assign n40648 = x50 & ~n40647 ;
  assign n40649 = ~n40646 & ~n40647 ;
  assign n40650 = ~n40648 & ~n40649 ;
  assign n40651 = ~n40063 & ~n40077 ;
  assign n40652 = ~n40027 & ~n40041 ;
  assign n40653 = x90 & n22325 ;
  assign n40654 = x88 & n23066 ;
  assign n40655 = x89 & n22320 ;
  assign n40656 = ~n40654 & ~n40655 ;
  assign n40657 = ~n40653 & n40656 ;
  assign n40658 = n4986 & n22328 ;
  assign n40659 = n40657 & ~n40658 ;
  assign n40660 = x59 & ~n40659 ;
  assign n40661 = x59 & ~n40660 ;
  assign n40662 = ~n40659 & ~n40660 ;
  assign n40663 = ~n40661 & ~n40662 ;
  assign n40664 = ~n40010 & ~n40024 ;
  assign n40665 = x83 & n27024 ;
  assign n40666 = x84 & ~n26217 ;
  assign n40667 = ~n40665 & ~n40666 ;
  assign n40668 = ~n40007 & n40667 ;
  assign n40669 = n40007 & ~n40667 ;
  assign n40670 = ~n40668 & ~n40669 ;
  assign n40671 = x87 & n24612 ;
  assign n40672 = x85 & n25390 ;
  assign n40673 = x86 & n24607 ;
  assign n40674 = ~n40672 & ~n40673 ;
  assign n40675 = ~n40671 & n40674 ;
  assign n40676 = ~n24615 & n40675 ;
  assign n40677 = ~n3991 & n40675 ;
  assign n40678 = ~n40676 & ~n40677 ;
  assign n40679 = x62 & ~n40678 ;
  assign n40680 = ~x62 & n40678 ;
  assign n40681 = ~n40679 & ~n40680 ;
  assign n40682 = n40670 & ~n40681 ;
  assign n40683 = ~n40670 & n40681 ;
  assign n40684 = ~n40682 & ~n40683 ;
  assign n40685 = ~n40664 & n40684 ;
  assign n40686 = n40664 & ~n40684 ;
  assign n40687 = ~n40685 & ~n40686 ;
  assign n40688 = ~n40663 & n40687 ;
  assign n40689 = n40663 & ~n40687 ;
  assign n40690 = ~n40688 & ~n40689 ;
  assign n40691 = ~n40652 & n40690 ;
  assign n40692 = n40652 & ~n40690 ;
  assign n40693 = ~n40691 & ~n40692 ;
  assign n40694 = x93 & n20143 ;
  assign n40695 = x91 & n20854 ;
  assign n40696 = x92 & n20138 ;
  assign n40697 = ~n40695 & ~n40696 ;
  assign n40698 = ~n40694 & n40697 ;
  assign n40699 = n6094 & n20146 ;
  assign n40700 = n40698 & ~n40699 ;
  assign n40701 = x56 & ~n40700 ;
  assign n40702 = x56 & ~n40701 ;
  assign n40703 = ~n40700 & ~n40701 ;
  assign n40704 = ~n40702 & ~n40703 ;
  assign n40705 = n40693 & ~n40704 ;
  assign n40706 = n40693 & ~n40705 ;
  assign n40707 = ~n40704 & ~n40705 ;
  assign n40708 = ~n40706 & ~n40707 ;
  assign n40709 = ~n40004 & ~n40044 ;
  assign n40710 = ~n40060 & ~n40709 ;
  assign n40711 = ~n40708 & ~n40710 ;
  assign n40712 = ~n40708 & ~n40711 ;
  assign n40713 = ~n40710 & ~n40711 ;
  assign n40714 = ~n40712 & ~n40713 ;
  assign n40715 = x96 & n18025 ;
  assign n40716 = x94 & n18764 ;
  assign n40717 = x95 & n18020 ;
  assign n40718 = ~n40716 & ~n40717 ;
  assign n40719 = ~n40715 & n40718 ;
  assign n40720 = n7321 & n18028 ;
  assign n40721 = n40719 & ~n40720 ;
  assign n40722 = x53 & ~n40721 ;
  assign n40723 = x53 & ~n40722 ;
  assign n40724 = ~n40721 & ~n40722 ;
  assign n40725 = ~n40723 & ~n40724 ;
  assign n40726 = ~n40714 & n40725 ;
  assign n40727 = n40714 & ~n40725 ;
  assign n40728 = ~n40726 & ~n40727 ;
  assign n40729 = ~n40651 & ~n40728 ;
  assign n40730 = n40651 & n40728 ;
  assign n40731 = ~n40729 & ~n40730 ;
  assign n40732 = ~n40650 & n40731 ;
  assign n40733 = n40650 & ~n40731 ;
  assign n40734 = ~n40732 & ~n40733 ;
  assign n40735 = ~n40639 & n40734 ;
  assign n40736 = n40639 & ~n40734 ;
  assign n40737 = ~n40735 & ~n40736 ;
  assign n40738 = ~n40638 & n40737 ;
  assign n40739 = n40638 & ~n40737 ;
  assign n40740 = ~n40738 & ~n40739 ;
  assign n40741 = ~n40627 & n40740 ;
  assign n40742 = n40627 & ~n40740 ;
  assign n40743 = ~n40741 & ~n40742 ;
  assign n40744 = ~n40626 & n40743 ;
  assign n40745 = n40626 & ~n40743 ;
  assign n40746 = ~n40744 & ~n40745 ;
  assign n40747 = ~n40615 & n40746 ;
  assign n40748 = n40615 & ~n40746 ;
  assign n40749 = ~n40747 & ~n40748 ;
  assign n40750 = ~n40614 & n40749 ;
  assign n40751 = n40614 & ~n40749 ;
  assign n40752 = ~n40750 & ~n40751 ;
  assign n40753 = ~n40603 & n40752 ;
  assign n40754 = n40603 & ~n40752 ;
  assign n40755 = ~n40753 & ~n40754 ;
  assign n40756 = x111 & n9433 ;
  assign n40757 = x109 & n9915 ;
  assign n40758 = x110 & n9428 ;
  assign n40759 = ~n40757 & ~n40758 ;
  assign n40760 = ~n40756 & n40759 ;
  assign n40761 = n9436 & n15111 ;
  assign n40762 = n40760 & ~n40761 ;
  assign n40763 = x38 & ~n40762 ;
  assign n40764 = x38 & ~n40763 ;
  assign n40765 = ~n40762 & ~n40763 ;
  assign n40766 = ~n40764 & ~n40765 ;
  assign n40767 = n40755 & ~n40766 ;
  assign n40768 = n40755 & ~n40767 ;
  assign n40769 = ~n40766 & ~n40767 ;
  assign n40770 = ~n40768 & ~n40769 ;
  assign n40771 = ~n40147 & ~n40160 ;
  assign n40772 = n40770 & n40771 ;
  assign n40773 = ~n40770 & ~n40771 ;
  assign n40774 = ~n40772 & ~n40773 ;
  assign n40775 = x114 & n8006 ;
  assign n40776 = x112 & n8474 ;
  assign n40777 = x113 & n8001 ;
  assign n40778 = ~n40776 & ~n40777 ;
  assign n40779 = ~n40775 & n40778 ;
  assign n40780 = n8009 & n17012 ;
  assign n40781 = n40779 & ~n40780 ;
  assign n40782 = x35 & ~n40781 ;
  assign n40783 = x35 & ~n40782 ;
  assign n40784 = ~n40781 & ~n40782 ;
  assign n40785 = ~n40783 & ~n40784 ;
  assign n40786 = n40774 & ~n40785 ;
  assign n40787 = ~n40774 & n40785 ;
  assign n40788 = n40602 & ~n40787 ;
  assign n40789 = ~n40786 & n40788 ;
  assign n40790 = n40602 & ~n40789 ;
  assign n40791 = ~n40787 & ~n40789 ;
  assign n40792 = ~n40786 & n40791 ;
  assign n40793 = ~n40790 & ~n40792 ;
  assign n40794 = ~n40587 & n40793 ;
  assign n40795 = n40587 & ~n40793 ;
  assign n40796 = ~n40794 & ~n40795 ;
  assign n40797 = n40571 & ~n40796 ;
  assign n40798 = n40571 & ~n40797 ;
  assign n40799 = ~n40796 & ~n40797 ;
  assign n40800 = ~n40798 & ~n40799 ;
  assign n40801 = ~n40556 & n40800 ;
  assign n40802 = n40556 & ~n40800 ;
  assign n40803 = ~n40801 & ~n40802 ;
  assign n40804 = ~n40540 & ~n40803 ;
  assign n40805 = n40540 & n40803 ;
  assign n40806 = ~n40804 & ~n40805 ;
  assign n40807 = ~n40528 & n40806 ;
  assign n40808 = n40528 & ~n40806 ;
  assign n40809 = ~n40807 & ~n40808 ;
  assign n40810 = ~n40527 & n40809 ;
  assign n40811 = n40527 & ~n40809 ;
  assign n40812 = ~n40810 & ~n40811 ;
  assign n41100 = n40812 & x211 ;
  assign n40813 = ~n40515 & ~n40519 ;
  assign n40814 = ~n40507 & ~n40511 ;
  assign n40815 = ~n40241 & ~n40492 ;
  assign n40816 = ~x127 & n3020 ;
  assign n40817 = n2754 & n27365 ;
  assign n40818 = ~n40816 & ~n40817 ;
  assign n40819 = ~x20 & ~n40818 ;
  assign n40820 = ~x20 & ~n40819 ;
  assign n40821 = ~n40818 & ~n40819 ;
  assign n40822 = ~n40820 & ~n40821 ;
  assign n40823 = ~n40815 & ~n40822 ;
  assign n40824 = ~n40815 & ~n40823 ;
  assign n40825 = ~n40822 & ~n40823 ;
  assign n40826 = ~n40824 & ~n40825 ;
  assign n40827 = ~x126 & n3589 ;
  assign n40828 = ~x124 & n3878 ;
  assign n40829 = ~x125 & n3584 ;
  assign n40830 = ~n40828 & ~n40829 ;
  assign n40831 = ~n40827 & n40830 ;
  assign n40832 = n3592 & n26128 ;
  assign n40833 = n40831 & ~n40832 ;
  assign n40834 = ~x23 & ~n40833 ;
  assign n40835 = ~x23 & ~n40834 ;
  assign n40836 = ~n40833 & ~n40834 ;
  assign n40837 = ~n40835 & ~n40836 ;
  assign n40838 = ~n40256 & ~n40489 ;
  assign n40839 = ~n40837 & ~n40838 ;
  assign n40840 = ~n40837 & ~n40839 ;
  assign n40841 = ~n40838 & ~n40839 ;
  assign n40842 = ~n40840 & ~n40841 ;
  assign n40843 = ~x123 & n4531 ;
  assign n40844 = ~x121 & n4847 ;
  assign n40845 = ~x122 & n4526 ;
  assign n40846 = ~n40844 & ~n40845 ;
  assign n40847 = ~n40843 & n40846 ;
  assign n40848 = n4534 & n23760 ;
  assign n40849 = n40847 & ~n40848 ;
  assign n40850 = ~x26 & ~n40849 ;
  assign n40851 = ~x26 & ~n40850 ;
  assign n40852 = ~n40849 & ~n40850 ;
  assign n40853 = ~n40851 & ~n40852 ;
  assign n40854 = ~n40271 & ~n40484 ;
  assign n40855 = n40853 & n40854 ;
  assign n40856 = ~n40853 & ~n40854 ;
  assign n40857 = ~n40855 & ~n40856 ;
  assign n40858 = ~x120 & n5560 ;
  assign n40859 = ~x118 & n5943 ;
  assign n40860 = ~x119 & n5555 ;
  assign n40861 = ~n40859 & ~n40860 ;
  assign n40862 = ~n40858 & n40861 ;
  assign n40863 = n5563 & n21501 ;
  assign n40864 = n40862 & ~n40863 ;
  assign n40865 = ~x29 & ~n40864 ;
  assign n40866 = ~x29 & ~n40865 ;
  assign n40867 = ~n40864 & ~n40865 ;
  assign n40868 = ~n40866 & ~n40867 ;
  assign n40869 = ~n40286 & ~n40481 ;
  assign n40870 = ~n40868 & ~n40869 ;
  assign n40871 = ~n40868 & ~n40870 ;
  assign n40872 = ~n40869 & ~n40870 ;
  assign n40873 = ~n40871 & ~n40872 ;
  assign n40874 = ~x117 & n6725 ;
  assign n40875 = ~x115 & n7129 ;
  assign n40876 = ~x116 & n6720 ;
  assign n40877 = ~n40875 & ~n40876 ;
  assign n40878 = ~n40874 & n40877 ;
  assign n40879 = n6728 & n19365 ;
  assign n40880 = n40878 & ~n40879 ;
  assign n40881 = ~x32 & ~n40880 ;
  assign n40882 = ~x32 & ~n40881 ;
  assign n40883 = ~n40880 & ~n40881 ;
  assign n40884 = ~n40882 & ~n40883 ;
  assign n40885 = ~n40464 & ~n40477 ;
  assign n40886 = n40884 & n40885 ;
  assign n40887 = ~n40884 & ~n40885 ;
  assign n40888 = ~n40886 & ~n40887 ;
  assign n40889 = ~n40425 & ~n40439 ;
  assign n40890 = ~x108 & n10905 ;
  assign n40891 = ~x106 & n11466 ;
  assign n40892 = ~x107 & n10900 ;
  assign n40893 = ~n40891 & ~n40892 ;
  assign n40894 = ~n40890 & n40893 ;
  assign n40895 = n10908 & n13601 ;
  assign n40896 = n40894 & ~n40895 ;
  assign n40897 = ~x41 & ~n40896 ;
  assign n40898 = ~x41 & ~n40897 ;
  assign n40899 = ~n40896 & ~n40897 ;
  assign n40900 = ~n40898 & ~n40899 ;
  assign n40901 = ~n40417 & ~n40421 ;
  assign n40902 = ~x105 & n12506 ;
  assign n40903 = ~x103 & n13131 ;
  assign n40904 = ~x104 & n12501 ;
  assign n40905 = ~n40903 & ~n40904 ;
  assign n40906 = ~n40902 & n40905 ;
  assign n40907 = n11907 & n12509 ;
  assign n40908 = n40906 & ~n40907 ;
  assign n40909 = ~x44 & ~n40908 ;
  assign n40910 = ~x44 & ~n40909 ;
  assign n40911 = ~n40908 & ~n40909 ;
  assign n40912 = ~n40910 & ~n40911 ;
  assign n40913 = ~n40401 & ~n40415 ;
  assign n40914 = ~x102 & n14233 ;
  assign n40915 = ~x100 & n14876 ;
  assign n40916 = ~x101 & n14228 ;
  assign n40917 = ~n40915 & ~n40916 ;
  assign n40918 = ~n40914 & n40917 ;
  assign n40919 = n10333 & n14236 ;
  assign n40920 = n40918 & ~n40919 ;
  assign n40921 = ~x47 & ~n40920 ;
  assign n40922 = ~x47 & ~n40921 ;
  assign n40923 = ~n40920 & ~n40921 ;
  assign n40924 = ~n40922 & ~n40923 ;
  assign n40925 = ~n40381 & ~n40394 ;
  assign n40926 = ~x99 & n16076 ;
  assign n40927 = ~x97 & n16756 ;
  assign n40928 = ~x98 & n16071 ;
  assign n40929 = ~n40927 & ~n40928 ;
  assign n40930 = ~n40926 & n40929 ;
  assign n40931 = n8885 & n16079 ;
  assign n40932 = n40930 & ~n40931 ;
  assign n40933 = ~x50 & ~n40932 ;
  assign n40934 = ~x50 & ~n40933 ;
  assign n40935 = ~n40932 & ~n40933 ;
  assign n40936 = ~n40934 & ~n40935 ;
  assign n40937 = ~n40361 & ~n40375 ;
  assign n40938 = ~n40325 & ~n40339 ;
  assign n40939 = ~x90 & n22325 ;
  assign n40940 = ~x88 & n23066 ;
  assign n40941 = ~x89 & n22320 ;
  assign n40942 = ~n40940 & ~n40941 ;
  assign n40943 = ~n40939 & n40942 ;
  assign n40944 = n5155 & n22328 ;
  assign n40945 = n40943 & ~n40944 ;
  assign n40946 = ~x59 & ~n40945 ;
  assign n40947 = ~x59 & ~n40946 ;
  assign n40948 = ~n40945 & ~n40946 ;
  assign n40949 = ~n40947 & ~n40948 ;
  assign n40950 = ~n40308 & ~n40322 ;
  assign n40951 = ~x83 & n27427 ;
  assign n40952 = ~x84 & ~n26217 ;
  assign n40953 = ~n40951 & ~n40952 ;
  assign n40954 = ~n40305 & n40953 ;
  assign n40955 = n40305 & ~n40953 ;
  assign n40956 = ~n40954 & ~n40955 ;
  assign n40957 = ~x87 & n24612 ;
  assign n40958 = ~x85 & n25390 ;
  assign n40959 = ~x86 & n24607 ;
  assign n40960 = ~n40958 & ~n40959 ;
  assign n40961 = ~n40957 & n40960 ;
  assign n40962 = ~n24615 & n40961 ;
  assign n40963 = ~n4143 & n40961 ;
  assign n40964 = ~n40962 & ~n40963 ;
  assign n40965 = ~x62 & ~n40964 ;
  assign n40966 = x62 & n40964 ;
  assign n40967 = ~n40965 & ~n40966 ;
  assign n40968 = n40956 & ~n40967 ;
  assign n40969 = ~n40956 & n40967 ;
  assign n40970 = ~n40968 & ~n40969 ;
  assign n40971 = ~n40950 & n40970 ;
  assign n40972 = n40950 & ~n40970 ;
  assign n40973 = ~n40971 & ~n40972 ;
  assign n40974 = ~n40949 & n40973 ;
  assign n40975 = n40949 & ~n40973 ;
  assign n40976 = ~n40974 & ~n40975 ;
  assign n40977 = ~n40938 & n40976 ;
  assign n40978 = n40938 & ~n40976 ;
  assign n40979 = ~n40977 & ~n40978 ;
  assign n40980 = ~x93 & n20143 ;
  assign n40981 = ~x91 & n20854 ;
  assign n40982 = ~x92 & n20138 ;
  assign n40983 = ~n40981 & ~n40982 ;
  assign n40984 = ~n40980 & n40983 ;
  assign n40985 = n6285 & n20146 ;
  assign n40986 = n40984 & ~n40985 ;
  assign n40987 = ~x56 & ~n40986 ;
  assign n40988 = ~x56 & ~n40987 ;
  assign n40989 = ~n40986 & ~n40987 ;
  assign n40990 = ~n40988 & ~n40989 ;
  assign n40991 = n40979 & ~n40990 ;
  assign n40992 = n40979 & ~n40991 ;
  assign n40993 = ~n40990 & ~n40991 ;
  assign n40994 = ~n40992 & ~n40993 ;
  assign n40995 = ~n40302 & ~n40342 ;
  assign n40996 = ~n40358 & ~n40995 ;
  assign n40997 = ~n40994 & ~n40996 ;
  assign n40998 = ~n40994 & ~n40997 ;
  assign n40999 = ~n40996 & ~n40997 ;
  assign n41000 = ~n40998 & ~n40999 ;
  assign n41001 = ~x96 & n18025 ;
  assign n41002 = ~x94 & n18764 ;
  assign n41003 = ~x95 & n18020 ;
  assign n41004 = ~n41002 & ~n41003 ;
  assign n41005 = ~n41001 & n41004 ;
  assign n41006 = n7531 & n18028 ;
  assign n41007 = n41005 & ~n41006 ;
  assign n41008 = ~x53 & ~n41007 ;
  assign n41009 = ~x53 & ~n41008 ;
  assign n41010 = ~n41007 & ~n41008 ;
  assign n41011 = ~n41009 & ~n41010 ;
  assign n41012 = ~n41000 & n41011 ;
  assign n41013 = n41000 & ~n41011 ;
  assign n41014 = ~n41012 & ~n41013 ;
  assign n41015 = ~n40937 & ~n41014 ;
  assign n41016 = n40937 & n41014 ;
  assign n41017 = ~n41015 & ~n41016 ;
  assign n41018 = ~n40936 & n41017 ;
  assign n41019 = n40936 & ~n41017 ;
  assign n41020 = ~n41018 & ~n41019 ;
  assign n41021 = ~n40925 & n41020 ;
  assign n41022 = n40925 & ~n41020 ;
  assign n41023 = ~n41021 & ~n41022 ;
  assign n41024 = ~n40924 & n41023 ;
  assign n41025 = n40924 & ~n41023 ;
  assign n41026 = ~n41024 & ~n41025 ;
  assign n41027 = ~n40913 & n41026 ;
  assign n41028 = n40913 & ~n41026 ;
  assign n41029 = ~n41027 & ~n41028 ;
  assign n41030 = ~n40912 & n41029 ;
  assign n41031 = n40912 & ~n41029 ;
  assign n41032 = ~n41030 & ~n41031 ;
  assign n41033 = ~n40901 & n41032 ;
  assign n41034 = n40901 & ~n41032 ;
  assign n41035 = ~n41033 & ~n41034 ;
  assign n41036 = ~n40900 & n41035 ;
  assign n41037 = n40900 & ~n41035 ;
  assign n41038 = ~n41036 & ~n41037 ;
  assign n41039 = ~n40889 & n41038 ;
  assign n41040 = n40889 & ~n41038 ;
  assign n41041 = ~n41039 & ~n41040 ;
  assign n41042 = ~x111 & n9433 ;
  assign n41043 = ~x109 & n9915 ;
  assign n41044 = ~x110 & n9428 ;
  assign n41045 = ~n41043 & ~n41044 ;
  assign n41046 = ~n41042 & n41045 ;
  assign n41047 = n9436 & n15411 ;
  assign n41048 = n41046 & ~n41047 ;
  assign n41049 = ~x38 & ~n41048 ;
  assign n41050 = ~x38 & ~n41049 ;
  assign n41051 = ~n41048 & ~n41049 ;
  assign n41052 = ~n41050 & ~n41051 ;
  assign n41053 = n41041 & ~n41052 ;
  assign n41054 = n41041 & ~n41053 ;
  assign n41055 = ~n41052 & ~n41053 ;
  assign n41056 = ~n41054 & ~n41055 ;
  assign n41057 = ~n40445 & ~n40458 ;
  assign n41058 = n41056 & n41057 ;
  assign n41059 = ~n41056 & ~n41057 ;
  assign n41060 = ~n41058 & ~n41059 ;
  assign n41061 = ~x114 & n8006 ;
  assign n41062 = ~x112 & n8474 ;
  assign n41063 = ~x113 & n8001 ;
  assign n41064 = ~n41062 & ~n41063 ;
  assign n41065 = ~n41061 & n41064 ;
  assign n41066 = n8009 & n17333 ;
  assign n41067 = n41065 & ~n41066 ;
  assign n41068 = ~x35 & ~n41067 ;
  assign n41069 = ~x35 & ~n41068 ;
  assign n41070 = ~n41067 & ~n41068 ;
  assign n41071 = ~n41069 & ~n41070 ;
  assign n41072 = n41060 & ~n41071 ;
  assign n41073 = ~n41060 & n41071 ;
  assign n41074 = n40888 & ~n41073 ;
  assign n41075 = ~n41072 & n41074 ;
  assign n41076 = n40888 & ~n41075 ;
  assign n41077 = ~n41073 & ~n41075 ;
  assign n41078 = ~n41072 & n41077 ;
  assign n41079 = ~n41076 & ~n41078 ;
  assign n41080 = ~n40873 & n41079 ;
  assign n41081 = n40873 & ~n41079 ;
  assign n41082 = ~n41080 & ~n41081 ;
  assign n41083 = n40857 & ~n41082 ;
  assign n41084 = n40857 & ~n41083 ;
  assign n41085 = ~n41082 & ~n41083 ;
  assign n41086 = ~n41084 & ~n41085 ;
  assign n41087 = ~n40842 & n41086 ;
  assign n41088 = n40842 & ~n41086 ;
  assign n41089 = ~n41087 & ~n41088 ;
  assign n41090 = ~n40826 & ~n41089 ;
  assign n41091 = n40826 & n41089 ;
  assign n41092 = ~n41090 & ~n41091 ;
  assign n41093 = ~n40814 & n41092 ;
  assign n41094 = n40814 & ~n41092 ;
  assign n41095 = ~n41093 & ~n41094 ;
  assign n41096 = ~n40813 & n41095 ;
  assign n41097 = n40813 & ~n41095 ;
  assign n41098 = ~n41096 & ~n41097 ;
  assign n41101 = ~n41098 & ~x211 ;
  assign n41102 = ~n41100 & ~n41101 ;
  assign n41103 = ~n40556 & ~n40800 ;
  assign n41104 = ~n40553 & ~n41103 ;
  assign n41105 = x127 & n3589 ;
  assign n41106 = x125 & n3878 ;
  assign n41107 = x126 & n3584 ;
  assign n41108 = ~n41106 & ~n41107 ;
  assign n41109 = ~n41105 & n41108 ;
  assign n41110 = n3592 & n26533 ;
  assign n41111 = n41109 & ~n41110 ;
  assign n41112 = x23 & ~n41111 ;
  assign n41113 = x23 & ~n41112 ;
  assign n41114 = ~n41111 & ~n41112 ;
  assign n41115 = ~n41113 & ~n41114 ;
  assign n41116 = ~n41104 & ~n41115 ;
  assign n41117 = ~n41104 & ~n41116 ;
  assign n41118 = ~n41115 & ~n41116 ;
  assign n41119 = ~n41117 & ~n41118 ;
  assign n41120 = x124 & n4531 ;
  assign n41121 = x122 & n4847 ;
  assign n41122 = x123 & n4526 ;
  assign n41123 = ~n41121 & ~n41122 ;
  assign n41124 = ~n41120 & n41123 ;
  assign n41125 = n4534 & n23796 ;
  assign n41126 = n41124 & ~n41125 ;
  assign n41127 = x26 & ~n41126 ;
  assign n41128 = x26 & ~n41127 ;
  assign n41129 = ~n41126 & ~n41127 ;
  assign n41130 = ~n41128 & ~n41129 ;
  assign n41131 = ~n40570 & ~n40797 ;
  assign n41132 = n41130 & n41131 ;
  assign n41133 = ~n41130 & ~n41131 ;
  assign n41134 = ~n41132 & ~n41133 ;
  assign n41135 = ~n40587 & ~n40793 ;
  assign n41136 = ~n40584 & ~n41135 ;
  assign n41137 = x121 & n5560 ;
  assign n41138 = x119 & n5943 ;
  assign n41139 = x120 & n5555 ;
  assign n41140 = ~n41138 & ~n41139 ;
  assign n41141 = ~n41137 & n41140 ;
  assign n41142 = n5563 & n21870 ;
  assign n41143 = n41141 & ~n41142 ;
  assign n41144 = x29 & ~n41143 ;
  assign n41145 = x29 & ~n41144 ;
  assign n41146 = ~n41143 & ~n41144 ;
  assign n41147 = ~n41145 & ~n41146 ;
  assign n41148 = ~n41136 & n41147 ;
  assign n41149 = n41136 & ~n41147 ;
  assign n41150 = ~n41148 & ~n41149 ;
  assign n41151 = x118 & n6725 ;
  assign n41152 = x116 & n7129 ;
  assign n41153 = x117 & n6720 ;
  assign n41154 = ~n41152 & ~n41153 ;
  assign n41155 = ~n41151 & n41154 ;
  assign n41156 = n6728 & n19395 ;
  assign n41157 = n41155 & ~n41156 ;
  assign n41158 = x32 & ~n41157 ;
  assign n41159 = x32 & ~n41158 ;
  assign n41160 = ~n41157 & ~n41158 ;
  assign n41161 = ~n41159 & ~n41160 ;
  assign n41162 = ~n40601 & ~n40789 ;
  assign n41163 = n41161 & n41162 ;
  assign n41164 = ~n41161 & ~n41162 ;
  assign n41165 = ~n41163 & ~n41164 ;
  assign n41166 = ~n40773 & ~n40786 ;
  assign n41167 = ~n40729 & ~n40732 ;
  assign n41168 = x84 & n27024 ;
  assign n41169 = x85 & ~n26217 ;
  assign n41170 = ~n41168 & ~n41169 ;
  assign n41171 = ~x20 & ~n41170 ;
  assign n41172 = x20 & n41170 ;
  assign n41173 = ~n41171 & ~n41172 ;
  assign n41174 = ~n40667 & n41173 ;
  assign n41175 = n40667 & ~n41173 ;
  assign n41176 = ~n41174 & ~n41175 ;
  assign n41177 = x88 & n24612 ;
  assign n41178 = x86 & n25390 ;
  assign n41179 = x87 & n24607 ;
  assign n41180 = ~n41178 & ~n41179 ;
  assign n41181 = ~n41177 & n41180 ;
  assign n41182 = n4305 & n24615 ;
  assign n41183 = n41181 & ~n41182 ;
  assign n41184 = x62 & ~n41183 ;
  assign n41185 = x62 & ~n41184 ;
  assign n41186 = ~n41183 & ~n41184 ;
  assign n41187 = ~n41185 & ~n41186 ;
  assign n41188 = n41176 & ~n41187 ;
  assign n41189 = n41176 & ~n41188 ;
  assign n41190 = ~n41187 & ~n41188 ;
  assign n41191 = ~n41189 & ~n41190 ;
  assign n41192 = ~n40668 & ~n40682 ;
  assign n41193 = ~n41191 & ~n41192 ;
  assign n41194 = ~n41191 & ~n41193 ;
  assign n41195 = ~n41192 & ~n41193 ;
  assign n41196 = ~n41194 & ~n41195 ;
  assign n41197 = x91 & n22325 ;
  assign n41198 = x89 & n23066 ;
  assign n41199 = x90 & n22320 ;
  assign n41200 = ~n41198 & ~n41199 ;
  assign n41201 = ~n41197 & n41200 ;
  assign n41202 = n5336 & n22328 ;
  assign n41203 = n41201 & ~n41202 ;
  assign n41204 = x59 & ~n41203 ;
  assign n41205 = x59 & ~n41204 ;
  assign n41206 = ~n41203 & ~n41204 ;
  assign n41207 = ~n41205 & ~n41206 ;
  assign n41208 = ~n41196 & ~n41207 ;
  assign n41209 = ~n41196 & ~n41208 ;
  assign n41210 = ~n41207 & ~n41208 ;
  assign n41211 = ~n41209 & ~n41210 ;
  assign n41212 = ~n40685 & ~n40688 ;
  assign n41213 = n41211 & n41212 ;
  assign n41214 = ~n41211 & ~n41212 ;
  assign n41215 = ~n41213 & ~n41214 ;
  assign n41216 = x94 & n20143 ;
  assign n41217 = x92 & n20854 ;
  assign n41218 = x93 & n20138 ;
  assign n41219 = ~n41217 & ~n41218 ;
  assign n41220 = ~n41216 & n41219 ;
  assign n41221 = n6483 & n20146 ;
  assign n41222 = n41220 & ~n41221 ;
  assign n41223 = x56 & ~n41222 ;
  assign n41224 = x56 & ~n41223 ;
  assign n41225 = ~n41222 & ~n41223 ;
  assign n41226 = ~n41224 & ~n41225 ;
  assign n41227 = n41215 & ~n41226 ;
  assign n41228 = n41215 & ~n41227 ;
  assign n41229 = ~n41226 & ~n41227 ;
  assign n41230 = ~n41228 & ~n41229 ;
  assign n41231 = ~n40691 & ~n40705 ;
  assign n41232 = n41230 & n41231 ;
  assign n41233 = ~n41230 & ~n41231 ;
  assign n41234 = ~n41232 & ~n41233 ;
  assign n41235 = x97 & n18025 ;
  assign n41236 = x95 & n18764 ;
  assign n41237 = x96 & n18020 ;
  assign n41238 = ~n41236 & ~n41237 ;
  assign n41239 = ~n41235 & n41238 ;
  assign n41240 = n7745 & n18028 ;
  assign n41241 = n41239 & ~n41240 ;
  assign n41242 = x53 & ~n41241 ;
  assign n41243 = x53 & ~n41242 ;
  assign n41244 = ~n41241 & ~n41242 ;
  assign n41245 = ~n41243 & ~n41244 ;
  assign n41246 = ~n40714 & ~n40725 ;
  assign n41247 = ~n40711 & ~n41246 ;
  assign n41248 = ~n41245 & ~n41247 ;
  assign n41249 = n41245 & n41247 ;
  assign n41250 = ~n41248 & ~n41249 ;
  assign n41251 = ~n41234 & n41250 ;
  assign n41252 = n41234 & ~n41250 ;
  assign n41253 = ~n41251 & ~n41252 ;
  assign n41254 = x100 & n16076 ;
  assign n41255 = x98 & n16756 ;
  assign n41256 = x99 & n16071 ;
  assign n41257 = ~n41255 & ~n41256 ;
  assign n41258 = ~n41254 & n41257 ;
  assign n41259 = n9115 & n16079 ;
  assign n41260 = n41258 & ~n41259 ;
  assign n41261 = x50 & ~n41260 ;
  assign n41262 = x50 & ~n41261 ;
  assign n41263 = ~n41260 & ~n41261 ;
  assign n41264 = ~n41262 & ~n41263 ;
  assign n41265 = ~n41253 & ~n41264 ;
  assign n41266 = n41253 & n41264 ;
  assign n41267 = ~n41265 & ~n41266 ;
  assign n41268 = n41167 & ~n41267 ;
  assign n41269 = ~n41167 & n41267 ;
  assign n41270 = ~n41268 & ~n41269 ;
  assign n41271 = x103 & n14233 ;
  assign n41272 = x101 & n14876 ;
  assign n41273 = x102 & n14228 ;
  assign n41274 = ~n41272 & ~n41273 ;
  assign n41275 = ~n41271 & n41274 ;
  assign n41276 = n10588 & n14236 ;
  assign n41277 = n41275 & ~n41276 ;
  assign n41278 = x47 & ~n41277 ;
  assign n41279 = x47 & ~n41278 ;
  assign n41280 = ~n41277 & ~n41278 ;
  assign n41281 = ~n41279 & ~n41280 ;
  assign n41282 = n41270 & ~n41281 ;
  assign n41283 = n41270 & ~n41282 ;
  assign n41284 = ~n41281 & ~n41282 ;
  assign n41285 = ~n41283 & ~n41284 ;
  assign n41286 = ~n40735 & ~n40738 ;
  assign n41287 = n41285 & n41286 ;
  assign n41288 = ~n41285 & ~n41286 ;
  assign n41289 = ~n41287 & ~n41288 ;
  assign n41290 = x106 & n12506 ;
  assign n41291 = x104 & n13131 ;
  assign n41292 = x105 & n12501 ;
  assign n41293 = ~n41291 & ~n41292 ;
  assign n41294 = ~n41290 & n41293 ;
  assign n41295 = n12181 & n12509 ;
  assign n41296 = n41294 & ~n41295 ;
  assign n41297 = x44 & ~n41296 ;
  assign n41298 = x44 & ~n41297 ;
  assign n41299 = ~n41296 & ~n41297 ;
  assign n41300 = ~n41298 & ~n41299 ;
  assign n41301 = n41289 & ~n41300 ;
  assign n41302 = n41289 & ~n41301 ;
  assign n41303 = ~n41300 & ~n41301 ;
  assign n41304 = ~n41302 & ~n41303 ;
  assign n41305 = ~n40741 & ~n40744 ;
  assign n41306 = n41304 & n41305 ;
  assign n41307 = ~n41304 & ~n41305 ;
  assign n41308 = ~n41306 & ~n41307 ;
  assign n41309 = x109 & n10905 ;
  assign n41310 = x107 & n11466 ;
  assign n41311 = x108 & n10900 ;
  assign n41312 = ~n41310 & ~n41311 ;
  assign n41313 = ~n41309 & n41312 ;
  assign n41314 = n10908 & n13894 ;
  assign n41315 = n41313 & ~n41314 ;
  assign n41316 = x41 & ~n41315 ;
  assign n41317 = x41 & ~n41316 ;
  assign n41318 = ~n41315 & ~n41316 ;
  assign n41319 = ~n41317 & ~n41318 ;
  assign n41320 = n41308 & ~n41319 ;
  assign n41321 = n41308 & ~n41320 ;
  assign n41322 = ~n41319 & ~n41320 ;
  assign n41323 = ~n41321 & ~n41322 ;
  assign n41324 = ~n40747 & ~n40750 ;
  assign n41325 = n41323 & n41324 ;
  assign n41326 = ~n41323 & ~n41324 ;
  assign n41327 = ~n41325 & ~n41326 ;
  assign n41328 = x112 & n9433 ;
  assign n41329 = x110 & n9915 ;
  assign n41330 = x111 & n9428 ;
  assign n41331 = ~n41329 & ~n41330 ;
  assign n41332 = ~n41328 & n41331 ;
  assign n41333 = n9436 & n15442 ;
  assign n41334 = n41332 & ~n41333 ;
  assign n41335 = x38 & ~n41334 ;
  assign n41336 = x38 & ~n41335 ;
  assign n41337 = ~n41334 & ~n41335 ;
  assign n41338 = ~n41336 & ~n41337 ;
  assign n41339 = n41327 & ~n41338 ;
  assign n41340 = n41327 & ~n41339 ;
  assign n41341 = ~n41338 & ~n41339 ;
  assign n41342 = ~n41340 & ~n41341 ;
  assign n41343 = ~n40753 & ~n40767 ;
  assign n41344 = n41342 & n41343 ;
  assign n41345 = ~n41342 & ~n41343 ;
  assign n41346 = ~n41344 & ~n41345 ;
  assign n41347 = x115 & n8006 ;
  assign n41348 = x113 & n8474 ;
  assign n41349 = x114 & n8001 ;
  assign n41350 = ~n41348 & ~n41349 ;
  assign n41351 = ~n41347 & n41350 ;
  assign n41352 = n8009 & n17364 ;
  assign n41353 = n41351 & ~n41352 ;
  assign n41354 = x35 & ~n41353 ;
  assign n41355 = x35 & ~n41354 ;
  assign n41356 = ~n41353 & ~n41354 ;
  assign n41357 = ~n41355 & ~n41356 ;
  assign n41358 = n41346 & ~n41357 ;
  assign n41359 = ~n41346 & n41357 ;
  assign n41360 = ~n41166 & ~n41359 ;
  assign n41361 = ~n41358 & n41360 ;
  assign n41362 = ~n41166 & ~n41361 ;
  assign n41363 = ~n41358 & ~n41361 ;
  assign n41364 = ~n41359 & n41363 ;
  assign n41365 = ~n41362 & ~n41364 ;
  assign n41366 = n41165 & ~n41365 ;
  assign n41367 = ~n41165 & n41365 ;
  assign n41368 = ~n41150 & ~n41367 ;
  assign n41369 = ~n41366 & n41368 ;
  assign n41370 = ~n41150 & ~n41369 ;
  assign n41371 = ~n41367 & ~n41369 ;
  assign n41372 = ~n41366 & n41371 ;
  assign n41373 = ~n41370 & ~n41372 ;
  assign n41374 = n41134 & ~n41373 ;
  assign n41375 = ~n41134 & n41373 ;
  assign n41376 = ~n41119 & ~n41375 ;
  assign n41377 = ~n41374 & n41376 ;
  assign n41378 = ~n41119 & ~n41377 ;
  assign n41379 = ~n41375 & ~n41377 ;
  assign n41380 = ~n41374 & n41379 ;
  assign n41381 = ~n41378 & ~n41380 ;
  assign n41382 = ~n40537 & ~n40804 ;
  assign n41383 = n41381 & n41382 ;
  assign n41384 = ~n41381 & ~n41382 ;
  assign n41385 = ~n41383 & ~n41384 ;
  assign n41386 = ~n40807 & ~n40810 ;
  assign n41387 = n41385 & ~n41386 ;
  assign n41388 = ~n41385 & n41386 ;
  assign n41389 = ~n41387 & ~n41388 ;
  assign n41678 = n41389 & x212 ;
  assign n41390 = ~n40842 & ~n41086 ;
  assign n41391 = ~n40839 & ~n41390 ;
  assign n41392 = ~x127 & n3589 ;
  assign n41393 = ~x125 & n3878 ;
  assign n41394 = ~x126 & n3584 ;
  assign n41395 = ~n41393 & ~n41394 ;
  assign n41396 = ~n41392 & n41395 ;
  assign n41397 = n3592 & n26932 ;
  assign n41398 = n41396 & ~n41397 ;
  assign n41399 = ~x23 & ~n41398 ;
  assign n41400 = ~x23 & ~n41399 ;
  assign n41401 = ~n41398 & ~n41399 ;
  assign n41402 = ~n41400 & ~n41401 ;
  assign n41403 = ~n41391 & ~n41402 ;
  assign n41404 = ~n41391 & ~n41403 ;
  assign n41405 = ~n41402 & ~n41403 ;
  assign n41406 = ~n41404 & ~n41405 ;
  assign n41407 = ~x124 & n4531 ;
  assign n41408 = ~x122 & n4847 ;
  assign n41409 = ~x123 & n4526 ;
  assign n41410 = ~n41408 & ~n41409 ;
  assign n41411 = ~n41407 & n41410 ;
  assign n41412 = n4534 & n24176 ;
  assign n41413 = n41411 & ~n41412 ;
  assign n41414 = ~x26 & ~n41413 ;
  assign n41415 = ~x26 & ~n41414 ;
  assign n41416 = ~n41413 & ~n41414 ;
  assign n41417 = ~n41415 & ~n41416 ;
  assign n41418 = ~n40856 & ~n41083 ;
  assign n41419 = n41417 & n41418 ;
  assign n41420 = ~n41417 & ~n41418 ;
  assign n41421 = ~n41419 & ~n41420 ;
  assign n41422 = ~n40873 & ~n41079 ;
  assign n41423 = ~n40870 & ~n41422 ;
  assign n41424 = ~x121 & n5560 ;
  assign n41425 = ~x119 & n5943 ;
  assign n41426 = ~x120 & n5555 ;
  assign n41427 = ~n41425 & ~n41426 ;
  assign n41428 = ~n41424 & n41427 ;
  assign n41429 = n5563 & n22229 ;
  assign n41430 = n41428 & ~n41429 ;
  assign n41431 = ~x29 & ~n41430 ;
  assign n41432 = ~x29 & ~n41431 ;
  assign n41433 = ~n41430 & ~n41431 ;
  assign n41434 = ~n41432 & ~n41433 ;
  assign n41435 = ~n41423 & n41434 ;
  assign n41436 = n41423 & ~n41434 ;
  assign n41437 = ~n41435 & ~n41436 ;
  assign n41438 = ~x118 & n6725 ;
  assign n41439 = ~x116 & n7129 ;
  assign n41440 = ~x117 & n6720 ;
  assign n41441 = ~n41439 & ~n41440 ;
  assign n41442 = ~n41438 & n41441 ;
  assign n41443 = n6728 & n19736 ;
  assign n41444 = n41442 & ~n41443 ;
  assign n41445 = ~x32 & ~n41444 ;
  assign n41446 = ~x32 & ~n41445 ;
  assign n41447 = ~n41444 & ~n41445 ;
  assign n41448 = ~n41446 & ~n41447 ;
  assign n41449 = ~n40887 & ~n41075 ;
  assign n41450 = n41448 & n41449 ;
  assign n41451 = ~n41448 & ~n41449 ;
  assign n41452 = ~n41450 & ~n41451 ;
  assign n41453 = ~n41059 & ~n41072 ;
  assign n41454 = ~n41015 & ~n41018 ;
  assign n41455 = ~x84 & n27427 ;
  assign n41456 = ~x85 & ~n26217 ;
  assign n41457 = ~n41455 & ~n41456 ;
  assign n41458 = x20 & ~n41457 ;
  assign n41459 = ~x20 & n41457 ;
  assign n41460 = ~n41458 & ~n41459 ;
  assign n41461 = ~n40953 & n41460 ;
  assign n41462 = n40953 & ~n41460 ;
  assign n41463 = ~n41461 & ~n41462 ;
  assign n41464 = ~x88 & n24612 ;
  assign n41465 = ~x86 & n25390 ;
  assign n41466 = ~x87 & n24607 ;
  assign n41467 = ~n41465 & ~n41466 ;
  assign n41468 = ~n41464 & n41467 ;
  assign n41469 = n4457 & n24615 ;
  assign n41470 = n41468 & ~n41469 ;
  assign n41471 = ~x62 & ~n41470 ;
  assign n41472 = ~x62 & ~n41471 ;
  assign n41473 = ~n41470 & ~n41471 ;
  assign n41474 = ~n41472 & ~n41473 ;
  assign n41475 = n41463 & ~n41474 ;
  assign n41476 = n41463 & ~n41475 ;
  assign n41477 = ~n41474 & ~n41475 ;
  assign n41478 = ~n41476 & ~n41477 ;
  assign n41479 = ~n40954 & ~n40968 ;
  assign n41480 = ~n41478 & ~n41479 ;
  assign n41481 = ~n41478 & ~n41480 ;
  assign n41482 = ~n41479 & ~n41480 ;
  assign n41483 = ~n41481 & ~n41482 ;
  assign n41484 = ~x91 & n22325 ;
  assign n41485 = ~x89 & n23066 ;
  assign n41486 = ~x90 & n22320 ;
  assign n41487 = ~n41485 & ~n41486 ;
  assign n41488 = ~n41484 & n41487 ;
  assign n41489 = n5507 & n22328 ;
  assign n41490 = n41488 & ~n41489 ;
  assign n41491 = ~x59 & ~n41490 ;
  assign n41492 = ~x59 & ~n41491 ;
  assign n41493 = ~n41490 & ~n41491 ;
  assign n41494 = ~n41492 & ~n41493 ;
  assign n41495 = ~n41483 & ~n41494 ;
  assign n41496 = ~n41483 & ~n41495 ;
  assign n41497 = ~n41494 & ~n41495 ;
  assign n41498 = ~n41496 & ~n41497 ;
  assign n41499 = ~n40971 & ~n40974 ;
  assign n41500 = n41498 & n41499 ;
  assign n41501 = ~n41498 & ~n41499 ;
  assign n41502 = ~n41500 & ~n41501 ;
  assign n41503 = ~x94 & n20143 ;
  assign n41504 = ~x92 & n20854 ;
  assign n41505 = ~x93 & n20138 ;
  assign n41506 = ~n41504 & ~n41505 ;
  assign n41507 = ~n41503 & n41506 ;
  assign n41508 = n6671 & n20146 ;
  assign n41509 = n41507 & ~n41508 ;
  assign n41510 = ~x56 & ~n41509 ;
  assign n41511 = ~x56 & ~n41510 ;
  assign n41512 = ~n41509 & ~n41510 ;
  assign n41513 = ~n41511 & ~n41512 ;
  assign n41514 = n41502 & ~n41513 ;
  assign n41515 = n41502 & ~n41514 ;
  assign n41516 = ~n41513 & ~n41514 ;
  assign n41517 = ~n41515 & ~n41516 ;
  assign n41518 = ~n40977 & ~n40991 ;
  assign n41519 = n41517 & n41518 ;
  assign n41520 = ~n41517 & ~n41518 ;
  assign n41521 = ~n41519 & ~n41520 ;
  assign n41522 = ~x97 & n18025 ;
  assign n41523 = ~x95 & n18764 ;
  assign n41524 = ~x96 & n18020 ;
  assign n41525 = ~n41523 & ~n41524 ;
  assign n41526 = ~n41522 & n41525 ;
  assign n41527 = n7949 & n18028 ;
  assign n41528 = n41526 & ~n41527 ;
  assign n41529 = ~x53 & ~n41528 ;
  assign n41530 = ~x53 & ~n41529 ;
  assign n41531 = ~n41528 & ~n41529 ;
  assign n41532 = ~n41530 & ~n41531 ;
  assign n41533 = ~n41000 & ~n41011 ;
  assign n41534 = ~n40997 & ~n41533 ;
  assign n41535 = ~n41532 & ~n41534 ;
  assign n41536 = n41532 & n41534 ;
  assign n41537 = ~n41535 & ~n41536 ;
  assign n41538 = ~n41521 & n41537 ;
  assign n41539 = n41521 & ~n41537 ;
  assign n41540 = ~n41538 & ~n41539 ;
  assign n41541 = ~x100 & n16076 ;
  assign n41542 = ~x98 & n16756 ;
  assign n41543 = ~x99 & n16071 ;
  assign n41544 = ~n41542 & ~n41543 ;
  assign n41545 = ~n41541 & n41544 ;
  assign n41546 = n9338 & n16079 ;
  assign n41547 = n41545 & ~n41546 ;
  assign n41548 = ~x50 & ~n41547 ;
  assign n41549 = ~x50 & ~n41548 ;
  assign n41550 = ~n41547 & ~n41548 ;
  assign n41551 = ~n41549 & ~n41550 ;
  assign n41552 = ~n41540 & ~n41551 ;
  assign n41553 = n41540 & n41551 ;
  assign n41554 = ~n41552 & ~n41553 ;
  assign n41555 = n41454 & ~n41554 ;
  assign n41556 = ~n41454 & n41554 ;
  assign n41557 = ~n41555 & ~n41556 ;
  assign n41558 = ~x103 & n14233 ;
  assign n41559 = ~x101 & n14876 ;
  assign n41560 = ~x102 & n14228 ;
  assign n41561 = ~n41559 & ~n41560 ;
  assign n41562 = ~n41558 & n41561 ;
  assign n41563 = n10833 & n14236 ;
  assign n41564 = n41562 & ~n41563 ;
  assign n41565 = ~x47 & ~n41564 ;
  assign n41566 = ~x47 & ~n41565 ;
  assign n41567 = ~n41564 & ~n41565 ;
  assign n41568 = ~n41566 & ~n41567 ;
  assign n41569 = n41557 & ~n41568 ;
  assign n41570 = n41557 & ~n41569 ;
  assign n41571 = ~n41568 & ~n41569 ;
  assign n41572 = ~n41570 & ~n41571 ;
  assign n41573 = ~n41021 & ~n41024 ;
  assign n41574 = n41572 & n41573 ;
  assign n41575 = ~n41572 & ~n41573 ;
  assign n41576 = ~n41574 & ~n41575 ;
  assign n41577 = ~x106 & n12506 ;
  assign n41578 = ~x104 & n13131 ;
  assign n41579 = ~x105 & n12501 ;
  assign n41580 = ~n41578 & ~n41579 ;
  assign n41581 = ~n41577 & n41580 ;
  assign n41582 = n12447 & n12509 ;
  assign n41583 = n41581 & ~n41582 ;
  assign n41584 = ~x44 & ~n41583 ;
  assign n41585 = ~x44 & ~n41584 ;
  assign n41586 = ~n41583 & ~n41584 ;
  assign n41587 = ~n41585 & ~n41586 ;
  assign n41588 = n41576 & ~n41587 ;
  assign n41589 = n41576 & ~n41588 ;
  assign n41590 = ~n41587 & ~n41588 ;
  assign n41591 = ~n41589 & ~n41590 ;
  assign n41592 = ~n41027 & ~n41030 ;
  assign n41593 = n41591 & n41592 ;
  assign n41594 = ~n41591 & ~n41592 ;
  assign n41595 = ~n41593 & ~n41594 ;
  assign n41596 = ~x109 & n10905 ;
  assign n41597 = ~x107 & n11466 ;
  assign n41598 = ~x108 & n10900 ;
  assign n41599 = ~n41597 & ~n41598 ;
  assign n41600 = ~n41596 & n41599 ;
  assign n41601 = n10908 & n14177 ;
  assign n41602 = n41600 & ~n41601 ;
  assign n41603 = ~x41 & ~n41602 ;
  assign n41604 = ~x41 & ~n41603 ;
  assign n41605 = ~n41602 & ~n41603 ;
  assign n41606 = ~n41604 & ~n41605 ;
  assign n41607 = n41595 & ~n41606 ;
  assign n41608 = n41595 & ~n41607 ;
  assign n41609 = ~n41606 & ~n41607 ;
  assign n41610 = ~n41608 & ~n41609 ;
  assign n41611 = ~n41033 & ~n41036 ;
  assign n41612 = n41610 & n41611 ;
  assign n41613 = ~n41610 & ~n41611 ;
  assign n41614 = ~n41612 & ~n41613 ;
  assign n41615 = ~x112 & n9433 ;
  assign n41616 = ~x110 & n9915 ;
  assign n41617 = ~x111 & n9428 ;
  assign n41618 = ~n41616 & ~n41617 ;
  assign n41619 = ~n41615 & n41618 ;
  assign n41620 = n9436 & n15744 ;
  assign n41621 = n41619 & ~n41620 ;
  assign n41622 = ~x38 & ~n41621 ;
  assign n41623 = ~x38 & ~n41622 ;
  assign n41624 = ~n41621 & ~n41622 ;
  assign n41625 = ~n41623 & ~n41624 ;
  assign n41626 = n41614 & ~n41625 ;
  assign n41627 = n41614 & ~n41626 ;
  assign n41628 = ~n41625 & ~n41626 ;
  assign n41629 = ~n41627 & ~n41628 ;
  assign n41630 = ~n41039 & ~n41053 ;
  assign n41631 = n41629 & n41630 ;
  assign n41632 = ~n41629 & ~n41630 ;
  assign n41633 = ~n41631 & ~n41632 ;
  assign n41634 = ~x115 & n8006 ;
  assign n41635 = ~x113 & n8474 ;
  assign n41636 = ~x114 & n8001 ;
  assign n41637 = ~n41635 & ~n41636 ;
  assign n41638 = ~n41634 & n41637 ;
  assign n41639 = n8009 & n17683 ;
  assign n41640 = n41638 & ~n41639 ;
  assign n41641 = ~x35 & ~n41640 ;
  assign n41642 = ~x35 & ~n41641 ;
  assign n41643 = ~n41640 & ~n41641 ;
  assign n41644 = ~n41642 & ~n41643 ;
  assign n41645 = n41633 & ~n41644 ;
  assign n41646 = ~n41633 & n41644 ;
  assign n41647 = ~n41453 & ~n41646 ;
  assign n41648 = ~n41645 & n41647 ;
  assign n41649 = ~n41453 & ~n41648 ;
  assign n41650 = ~n41645 & ~n41648 ;
  assign n41651 = ~n41646 & n41650 ;
  assign n41652 = ~n41649 & ~n41651 ;
  assign n41653 = n41452 & ~n41652 ;
  assign n41654 = ~n41452 & n41652 ;
  assign n41655 = ~n41437 & ~n41654 ;
  assign n41656 = ~n41653 & n41655 ;
  assign n41657 = ~n41437 & ~n41656 ;
  assign n41658 = ~n41654 & ~n41656 ;
  assign n41659 = ~n41653 & n41658 ;
  assign n41660 = ~n41657 & ~n41659 ;
  assign n41661 = n41421 & ~n41660 ;
  assign n41662 = ~n41421 & n41660 ;
  assign n41663 = ~n41406 & ~n41662 ;
  assign n41664 = ~n41661 & n41663 ;
  assign n41665 = ~n41406 & ~n41664 ;
  assign n41666 = ~n41662 & ~n41664 ;
  assign n41667 = ~n41661 & n41666 ;
  assign n41668 = ~n41665 & ~n41667 ;
  assign n41669 = ~n40823 & ~n41090 ;
  assign n41670 = n41668 & n41669 ;
  assign n41671 = ~n41668 & ~n41669 ;
  assign n41672 = ~n41670 & ~n41671 ;
  assign n41673 = ~n41093 & ~n41096 ;
  assign n41674 = n41672 & ~n41673 ;
  assign n41675 = ~n41672 & n41673 ;
  assign n41676 = ~n41674 & ~n41675 ;
  assign n41679 = ~n41676 & ~x212 ;
  assign n41680 = ~n41678 & ~n41679 ;
  assign n41681 = ~n41133 & ~n41374 ;
  assign n41682 = x126 & n3878 ;
  assign n41683 = x127 & n3584 ;
  assign n41684 = ~n41682 & ~n41683 ;
  assign n41685 = ~n3592 & n41684 ;
  assign n41686 = n26965 & n41684 ;
  assign n41687 = ~n41685 & ~n41686 ;
  assign n41688 = x23 & ~n41687 ;
  assign n41689 = ~x23 & n41687 ;
  assign n41690 = ~n41688 & ~n41689 ;
  assign n41691 = ~n41681 & ~n41690 ;
  assign n41692 = n41681 & n41690 ;
  assign n41693 = ~n41691 & ~n41692 ;
  assign n41694 = x125 & n4531 ;
  assign n41695 = x123 & n4847 ;
  assign n41696 = x124 & n4526 ;
  assign n41697 = ~n41695 & ~n41696 ;
  assign n41698 = ~n41694 & n41697 ;
  assign n41699 = n4534 & n24935 ;
  assign n41700 = n41698 & ~n41699 ;
  assign n41701 = x26 & ~n41700 ;
  assign n41702 = x26 & ~n41701 ;
  assign n41703 = ~n41700 & ~n41701 ;
  assign n41704 = ~n41702 & ~n41703 ;
  assign n41705 = ~n41136 & ~n41147 ;
  assign n41706 = ~n41369 & ~n41705 ;
  assign n41707 = n41704 & n41706 ;
  assign n41708 = ~n41704 & ~n41706 ;
  assign n41709 = ~n41707 & ~n41708 ;
  assign n41710 = ~n41164 & ~n41366 ;
  assign n41711 = x122 & n5560 ;
  assign n41712 = x120 & n5943 ;
  assign n41713 = x121 & n5555 ;
  assign n41714 = ~n41712 & ~n41713 ;
  assign n41715 = ~n41711 & n41714 ;
  assign n41716 = ~n5563 & n41715 ;
  assign n41717 = ~n22622 & n41715 ;
  assign n41718 = ~n41716 & ~n41717 ;
  assign n41719 = x29 & ~n41718 ;
  assign n41720 = ~x29 & n41718 ;
  assign n41721 = ~n41719 & ~n41720 ;
  assign n41722 = ~n41710 & ~n41721 ;
  assign n41723 = n41710 & n41721 ;
  assign n41724 = ~n41722 & ~n41723 ;
  assign n41725 = x119 & n6725 ;
  assign n41726 = x117 & n7129 ;
  assign n41727 = x118 & n6720 ;
  assign n41728 = ~n41726 & ~n41727 ;
  assign n41729 = ~n41725 & n41728 ;
  assign n41730 = n6728 & n20423 ;
  assign n41731 = n41729 & ~n41730 ;
  assign n41732 = x32 & ~n41731 ;
  assign n41733 = x32 & ~n41732 ;
  assign n41734 = ~n41731 & ~n41732 ;
  assign n41735 = ~n41733 & ~n41734 ;
  assign n41736 = ~n41363 & n41735 ;
  assign n41737 = n41363 & ~n41735 ;
  assign n41738 = ~n41736 & ~n41737 ;
  assign n41739 = ~n41282 & ~n41288 ;
  assign n41740 = x104 & n14233 ;
  assign n41741 = x102 & n14876 ;
  assign n41742 = x103 & n14228 ;
  assign n41743 = ~n41741 & ~n41742 ;
  assign n41744 = ~n41740 & n41743 ;
  assign n41745 = n11116 & n14236 ;
  assign n41746 = n41744 & ~n41745 ;
  assign n41747 = x47 & ~n41746 ;
  assign n41748 = x47 & ~n41747 ;
  assign n41749 = ~n41746 & ~n41747 ;
  assign n41750 = ~n41748 & ~n41749 ;
  assign n41751 = ~n41265 & ~n41269 ;
  assign n41752 = ~n41208 & ~n41214 ;
  assign n41753 = x92 & n22325 ;
  assign n41754 = x90 & n23066 ;
  assign n41755 = x91 & n22320 ;
  assign n41756 = ~n41754 & ~n41755 ;
  assign n41757 = ~n41753 & n41756 ;
  assign n41758 = n5710 & n22328 ;
  assign n41759 = n41757 & ~n41758 ;
  assign n41760 = x59 & ~n41759 ;
  assign n41761 = x59 & ~n41760 ;
  assign n41762 = ~n41759 & ~n41760 ;
  assign n41763 = ~n41761 & ~n41762 ;
  assign n41764 = ~n41188 & ~n41193 ;
  assign n41765 = x85 & n27024 ;
  assign n41766 = x86 & ~n26217 ;
  assign n41767 = ~n41765 & ~n41766 ;
  assign n41768 = ~n41171 & ~n41174 ;
  assign n41769 = ~n41767 & n41768 ;
  assign n41770 = n41767 & ~n41768 ;
  assign n41771 = ~n41769 & ~n41770 ;
  assign n41772 = x89 & n24612 ;
  assign n41773 = x87 & n25390 ;
  assign n41774 = x88 & n24607 ;
  assign n41775 = ~n41773 & ~n41774 ;
  assign n41776 = ~n41772 & n41775 ;
  assign n41777 = ~n24615 & n41776 ;
  assign n41778 = ~n4488 & n41776 ;
  assign n41779 = ~n41777 & ~n41778 ;
  assign n41780 = x62 & ~n41779 ;
  assign n41781 = ~x62 & n41779 ;
  assign n41782 = ~n41780 & ~n41781 ;
  assign n41783 = n41771 & ~n41782 ;
  assign n41784 = ~n41771 & n41782 ;
  assign n41785 = ~n41783 & ~n41784 ;
  assign n41786 = ~n41764 & n41785 ;
  assign n41787 = n41764 & ~n41785 ;
  assign n41788 = ~n41786 & ~n41787 ;
  assign n41789 = ~n41763 & n41788 ;
  assign n41790 = n41763 & ~n41788 ;
  assign n41791 = ~n41789 & ~n41790 ;
  assign n41792 = ~n41752 & n41791 ;
  assign n41793 = n41752 & ~n41791 ;
  assign n41794 = ~n41792 & ~n41793 ;
  assign n41795 = x95 & n20143 ;
  assign n41796 = x93 & n20854 ;
  assign n41797 = x94 & n20138 ;
  assign n41798 = ~n41796 & ~n41797 ;
  assign n41799 = ~n41795 & n41798 ;
  assign n41800 = n6894 & n20146 ;
  assign n41801 = n41799 & ~n41800 ;
  assign n41802 = x56 & ~n41801 ;
  assign n41803 = x56 & ~n41802 ;
  assign n41804 = ~n41801 & ~n41802 ;
  assign n41805 = ~n41803 & ~n41804 ;
  assign n41806 = n41794 & ~n41805 ;
  assign n41807 = n41794 & ~n41806 ;
  assign n41808 = ~n41805 & ~n41806 ;
  assign n41809 = ~n41807 & ~n41808 ;
  assign n41810 = ~n41227 & ~n41233 ;
  assign n41811 = n41809 & n41810 ;
  assign n41812 = ~n41809 & ~n41810 ;
  assign n41813 = ~n41811 & ~n41812 ;
  assign n41814 = x98 & n18025 ;
  assign n41815 = x96 & n18764 ;
  assign n41816 = x97 & n18020 ;
  assign n41817 = ~n41815 & ~n41816 ;
  assign n41818 = ~n41814 & n41817 ;
  assign n41819 = n8196 & n18028 ;
  assign n41820 = n41818 & ~n41819 ;
  assign n41821 = x53 & ~n41820 ;
  assign n41822 = x53 & ~n41821 ;
  assign n41823 = ~n41820 & ~n41821 ;
  assign n41824 = ~n41822 & ~n41823 ;
  assign n41825 = n41813 & ~n41824 ;
  assign n41826 = n41813 & ~n41825 ;
  assign n41827 = ~n41824 & ~n41825 ;
  assign n41828 = ~n41826 & ~n41827 ;
  assign n41829 = n41234 & n41250 ;
  assign n41830 = ~n41248 & ~n41829 ;
  assign n41831 = n41828 & n41830 ;
  assign n41832 = ~n41828 & ~n41830 ;
  assign n41833 = ~n41831 & ~n41832 ;
  assign n41834 = x101 & n16076 ;
  assign n41835 = x99 & n16756 ;
  assign n41836 = x100 & n16071 ;
  assign n41837 = ~n41835 & ~n41836 ;
  assign n41838 = ~n41834 & n41837 ;
  assign n41839 = n9601 & n16079 ;
  assign n41840 = n41838 & ~n41839 ;
  assign n41841 = x50 & ~n41840 ;
  assign n41842 = x50 & ~n41841 ;
  assign n41843 = ~n41840 & ~n41841 ;
  assign n41844 = ~n41842 & ~n41843 ;
  assign n41845 = ~n41833 & n41844 ;
  assign n41846 = n41833 & ~n41844 ;
  assign n41847 = ~n41845 & ~n41846 ;
  assign n41848 = ~n41751 & n41847 ;
  assign n41849 = ~n41751 & ~n41848 ;
  assign n41850 = n41847 & ~n41848 ;
  assign n41851 = ~n41849 & ~n41850 ;
  assign n41852 = ~n41750 & ~n41851 ;
  assign n41853 = n41750 & ~n41850 ;
  assign n41854 = ~n41849 & n41853 ;
  assign n41855 = ~n41852 & ~n41854 ;
  assign n41856 = ~n41739 & n41855 ;
  assign n41857 = n41739 & ~n41855 ;
  assign n41858 = ~n41856 & ~n41857 ;
  assign n41859 = x107 & n12506 ;
  assign n41860 = x105 & n13131 ;
  assign n41861 = x106 & n12501 ;
  assign n41862 = ~n41860 & ~n41861 ;
  assign n41863 = ~n41859 & n41862 ;
  assign n41864 = n12509 & n12749 ;
  assign n41865 = n41863 & ~n41864 ;
  assign n41866 = x44 & ~n41865 ;
  assign n41867 = x44 & ~n41866 ;
  assign n41868 = ~n41865 & ~n41866 ;
  assign n41869 = ~n41867 & ~n41868 ;
  assign n41870 = n41858 & ~n41869 ;
  assign n41871 = n41858 & ~n41870 ;
  assign n41872 = ~n41869 & ~n41870 ;
  assign n41873 = ~n41871 & ~n41872 ;
  assign n41874 = ~n41301 & ~n41307 ;
  assign n41875 = n41873 & n41874 ;
  assign n41876 = ~n41873 & ~n41874 ;
  assign n41877 = ~n41875 & ~n41876 ;
  assign n41878 = x110 & n10905 ;
  assign n41879 = x108 & n11466 ;
  assign n41880 = x109 & n10900 ;
  assign n41881 = ~n41879 & ~n41880 ;
  assign n41882 = ~n41878 & n41881 ;
  assign n41883 = n10908 & n14497 ;
  assign n41884 = n41882 & ~n41883 ;
  assign n41885 = x41 & ~n41884 ;
  assign n41886 = x41 & ~n41885 ;
  assign n41887 = ~n41884 & ~n41885 ;
  assign n41888 = ~n41886 & ~n41887 ;
  assign n41889 = n41877 & ~n41888 ;
  assign n41890 = n41877 & ~n41889 ;
  assign n41891 = ~n41888 & ~n41889 ;
  assign n41892 = ~n41890 & ~n41891 ;
  assign n41893 = ~n41320 & ~n41326 ;
  assign n41894 = n41892 & n41893 ;
  assign n41895 = ~n41892 & ~n41893 ;
  assign n41896 = ~n41894 & ~n41895 ;
  assign n41897 = x113 & n9433 ;
  assign n41898 = x111 & n9915 ;
  assign n41899 = x112 & n9428 ;
  assign n41900 = ~n41898 & ~n41899 ;
  assign n41901 = ~n41897 & n41900 ;
  assign n41902 = n9436 & n16361 ;
  assign n41903 = n41901 & ~n41902 ;
  assign n41904 = x38 & ~n41903 ;
  assign n41905 = x38 & ~n41904 ;
  assign n41906 = ~n41903 & ~n41904 ;
  assign n41907 = ~n41905 & ~n41906 ;
  assign n41908 = n41896 & ~n41907 ;
  assign n41909 = n41896 & ~n41908 ;
  assign n41910 = ~n41907 & ~n41908 ;
  assign n41911 = ~n41909 & ~n41910 ;
  assign n41912 = ~n41339 & ~n41345 ;
  assign n41913 = n41911 & n41912 ;
  assign n41914 = ~n41911 & ~n41912 ;
  assign n41915 = ~n41913 & ~n41914 ;
  assign n41916 = x116 & n8006 ;
  assign n41917 = x114 & n8474 ;
  assign n41918 = x115 & n8001 ;
  assign n41919 = ~n41917 & ~n41918 ;
  assign n41920 = ~n41916 & n41919 ;
  assign n41921 = n8009 & n18336 ;
  assign n41922 = n41920 & ~n41921 ;
  assign n41923 = x35 & ~n41922 ;
  assign n41924 = x35 & ~n41923 ;
  assign n41925 = ~n41922 & ~n41923 ;
  assign n41926 = ~n41924 & ~n41925 ;
  assign n41927 = n41915 & ~n41926 ;
  assign n41928 = n41915 & ~n41927 ;
  assign n41929 = ~n41926 & ~n41927 ;
  assign n41930 = ~n41928 & ~n41929 ;
  assign n41931 = ~n41738 & ~n41930 ;
  assign n41932 = n41738 & n41930 ;
  assign n41933 = n41724 & ~n41932 ;
  assign n41934 = ~n41931 & n41933 ;
  assign n41935 = n41724 & ~n41934 ;
  assign n41936 = ~n41932 & ~n41934 ;
  assign n41937 = ~n41931 & n41936 ;
  assign n41938 = ~n41935 & ~n41937 ;
  assign n41939 = n41709 & ~n41938 ;
  assign n41940 = ~n41709 & n41938 ;
  assign n41941 = n41693 & ~n41940 ;
  assign n41942 = ~n41939 & n41941 ;
  assign n41943 = n41693 & ~n41942 ;
  assign n41944 = ~n41940 & ~n41942 ;
  assign n41945 = ~n41939 & n41944 ;
  assign n41946 = ~n41943 & ~n41945 ;
  assign n41947 = ~n41116 & ~n41377 ;
  assign n41948 = n41946 & n41947 ;
  assign n41949 = ~n41946 & ~n41947 ;
  assign n41950 = ~n41948 & ~n41949 ;
  assign n41951 = ~n41384 & ~n41387 ;
  assign n41952 = n41950 & ~n41951 ;
  assign n41953 = ~n41950 & n41951 ;
  assign n41954 = ~n41952 & ~n41953 ;
  assign n42230 = n41954 & x213 ;
  assign n41955 = ~n41420 & ~n41661 ;
  assign n41956 = ~x126 & n3878 ;
  assign n41957 = ~x127 & n3584 ;
  assign n41958 = ~n41956 & ~n41957 ;
  assign n41959 = ~n3592 & n41958 ;
  assign n41960 = n27368 & n41958 ;
  assign n41961 = ~n41959 & ~n41960 ;
  assign n41962 = ~x23 & ~n41961 ;
  assign n41963 = x23 & n41961 ;
  assign n41964 = ~n41962 & ~n41963 ;
  assign n41965 = ~n41955 & ~n41964 ;
  assign n41966 = n41955 & n41964 ;
  assign n41967 = ~n41965 & ~n41966 ;
  assign n41968 = ~x125 & n4531 ;
  assign n41969 = ~x123 & n4847 ;
  assign n41970 = ~x124 & n4526 ;
  assign n41971 = ~n41969 & ~n41970 ;
  assign n41972 = ~n41968 & n41971 ;
  assign n41973 = n4534 & n25330 ;
  assign n41974 = n41972 & ~n41973 ;
  assign n41975 = ~x26 & ~n41974 ;
  assign n41976 = ~x26 & ~n41975 ;
  assign n41977 = ~n41974 & ~n41975 ;
  assign n41978 = ~n41976 & ~n41977 ;
  assign n41979 = ~n41423 & ~n41434 ;
  assign n41980 = ~n41656 & ~n41979 ;
  assign n41981 = n41978 & n41980 ;
  assign n41982 = ~n41978 & ~n41980 ;
  assign n41983 = ~n41981 & ~n41982 ;
  assign n41984 = ~n41451 & ~n41653 ;
  assign n41985 = ~x122 & n5560 ;
  assign n41986 = ~x120 & n5943 ;
  assign n41987 = ~x121 & n5555 ;
  assign n41988 = ~n41986 & ~n41987 ;
  assign n41989 = ~n41985 & n41988 ;
  assign n41990 = ~n5563 & n41989 ;
  assign n41991 = ~n22998 & n41989 ;
  assign n41992 = ~n41990 & ~n41991 ;
  assign n41993 = ~x29 & ~n41992 ;
  assign n41994 = x29 & n41992 ;
  assign n41995 = ~n41993 & ~n41994 ;
  assign n41996 = ~n41984 & ~n41995 ;
  assign n41997 = n41984 & n41995 ;
  assign n41998 = ~n41996 & ~n41997 ;
  assign n41999 = ~x119 & n6725 ;
  assign n42000 = ~x117 & n7129 ;
  assign n42001 = ~x118 & n6720 ;
  assign n42002 = ~n42000 & ~n42001 ;
  assign n42003 = ~n41999 & n42002 ;
  assign n42004 = n6728 & n20778 ;
  assign n42005 = n42003 & ~n42004 ;
  assign n42006 = ~x32 & ~n42005 ;
  assign n42007 = ~x32 & ~n42006 ;
  assign n42008 = ~n42005 & ~n42006 ;
  assign n42009 = ~n42007 & ~n42008 ;
  assign n42010 = ~n41650 & n42009 ;
  assign n42011 = n41650 & ~n42009 ;
  assign n42012 = ~n42010 & ~n42011 ;
  assign n42013 = ~n41569 & ~n41575 ;
  assign n42014 = ~x104 & n14233 ;
  assign n42015 = ~x102 & n14876 ;
  assign n42016 = ~x103 & n14228 ;
  assign n42017 = ~n42015 & ~n42016 ;
  assign n42018 = ~n42014 & n42017 ;
  assign n42019 = n11380 & n14236 ;
  assign n42020 = n42018 & ~n42019 ;
  assign n42021 = ~x47 & ~n42020 ;
  assign n42022 = ~x47 & ~n42021 ;
  assign n42023 = ~n42020 & ~n42021 ;
  assign n42024 = ~n42022 & ~n42023 ;
  assign n42025 = ~n41552 & ~n41556 ;
  assign n42026 = ~n41495 & ~n41501 ;
  assign n42027 = ~x92 & n22325 ;
  assign n42028 = ~x90 & n23066 ;
  assign n42029 = ~x91 & n22320 ;
  assign n42030 = ~n42028 & ~n42029 ;
  assign n42031 = ~n42027 & n42030 ;
  assign n42032 = n5896 & n22328 ;
  assign n42033 = n42031 & ~n42032 ;
  assign n42034 = ~x59 & ~n42033 ;
  assign n42035 = ~x59 & ~n42034 ;
  assign n42036 = ~n42033 & ~n42034 ;
  assign n42037 = ~n42035 & ~n42036 ;
  assign n42038 = ~n41475 & ~n41480 ;
  assign n42039 = ~x85 & n27427 ;
  assign n42040 = ~x86 & ~n26217 ;
  assign n42041 = ~n42039 & ~n42040 ;
  assign n42042 = ~n41458 & ~n41461 ;
  assign n42043 = ~n42041 & n42042 ;
  assign n42044 = n42041 & ~n42042 ;
  assign n42045 = ~n42043 & ~n42044 ;
  assign n42046 = ~x89 & n24612 ;
  assign n42047 = ~x87 & n25390 ;
  assign n42048 = ~x88 & n24607 ;
  assign n42049 = ~n42047 & ~n42048 ;
  assign n42050 = ~n42046 & n42049 ;
  assign n42051 = ~n24615 & n42050 ;
  assign n42052 = ~n4664 & n42050 ;
  assign n42053 = ~n42051 & ~n42052 ;
  assign n42054 = ~x62 & ~n42053 ;
  assign n42055 = x62 & n42053 ;
  assign n42056 = ~n42054 & ~n42055 ;
  assign n42057 = n42045 & ~n42056 ;
  assign n42058 = ~n42045 & n42056 ;
  assign n42059 = ~n42057 & ~n42058 ;
  assign n42060 = ~n42038 & n42059 ;
  assign n42061 = n42038 & ~n42059 ;
  assign n42062 = ~n42060 & ~n42061 ;
  assign n42063 = ~n42037 & n42062 ;
  assign n42064 = n42037 & ~n42062 ;
  assign n42065 = ~n42063 & ~n42064 ;
  assign n42066 = ~n42026 & n42065 ;
  assign n42067 = n42026 & ~n42065 ;
  assign n42068 = ~n42066 & ~n42067 ;
  assign n42069 = ~x95 & n20143 ;
  assign n42070 = ~x93 & n20854 ;
  assign n42071 = ~x94 & n20138 ;
  assign n42072 = ~n42070 & ~n42071 ;
  assign n42073 = ~n42069 & n42072 ;
  assign n42074 = n7100 & n20146 ;
  assign n42075 = n42073 & ~n42074 ;
  assign n42076 = ~x56 & ~n42075 ;
  assign n42077 = ~x56 & ~n42076 ;
  assign n42078 = ~n42075 & ~n42076 ;
  assign n42079 = ~n42077 & ~n42078 ;
  assign n42080 = n42068 & ~n42079 ;
  assign n42081 = n42068 & ~n42080 ;
  assign n42082 = ~n42079 & ~n42080 ;
  assign n42083 = ~n42081 & ~n42082 ;
  assign n42084 = ~n41514 & ~n41520 ;
  assign n42085 = n42083 & n42084 ;
  assign n42086 = ~n42083 & ~n42084 ;
  assign n42087 = ~n42085 & ~n42086 ;
  assign n42088 = ~x98 & n18025 ;
  assign n42089 = ~x96 & n18764 ;
  assign n42090 = ~x97 & n18020 ;
  assign n42091 = ~n42089 & ~n42090 ;
  assign n42092 = ~n42088 & n42091 ;
  assign n42093 = n8426 & n18028 ;
  assign n42094 = n42092 & ~n42093 ;
  assign n42095 = ~x53 & ~n42094 ;
  assign n42096 = ~x53 & ~n42095 ;
  assign n42097 = ~n42094 & ~n42095 ;
  assign n42098 = ~n42096 & ~n42097 ;
  assign n42099 = n42087 & ~n42098 ;
  assign n42100 = n42087 & ~n42099 ;
  assign n42101 = ~n42098 & ~n42099 ;
  assign n42102 = ~n42100 & ~n42101 ;
  assign n42103 = n41521 & n41537 ;
  assign n42104 = ~n41535 & ~n42103 ;
  assign n42105 = n42102 & n42104 ;
  assign n42106 = ~n42102 & ~n42104 ;
  assign n42107 = ~n42105 & ~n42106 ;
  assign n42108 = ~x101 & n16076 ;
  assign n42109 = ~x99 & n16756 ;
  assign n42110 = ~x100 & n16071 ;
  assign n42111 = ~n42109 & ~n42110 ;
  assign n42112 = ~n42108 & n42111 ;
  assign n42113 = n9844 & n16079 ;
  assign n42114 = n42112 & ~n42113 ;
  assign n42115 = ~x50 & ~n42114 ;
  assign n42116 = ~x50 & ~n42115 ;
  assign n42117 = ~n42114 & ~n42115 ;
  assign n42118 = ~n42116 & ~n42117 ;
  assign n42119 = ~n42107 & n42118 ;
  assign n42120 = n42107 & ~n42118 ;
  assign n42121 = ~n42119 & ~n42120 ;
  assign n42122 = ~n42025 & n42121 ;
  assign n42123 = ~n42025 & ~n42122 ;
  assign n42124 = n42121 & ~n42122 ;
  assign n42125 = ~n42123 & ~n42124 ;
  assign n42126 = ~n42024 & ~n42125 ;
  assign n42127 = n42024 & ~n42124 ;
  assign n42128 = ~n42123 & n42127 ;
  assign n42129 = ~n42126 & ~n42128 ;
  assign n42130 = ~n42013 & n42129 ;
  assign n42131 = n42013 & ~n42129 ;
  assign n42132 = ~n42130 & ~n42131 ;
  assign n42133 = ~x107 & n12506 ;
  assign n42134 = ~x105 & n13131 ;
  assign n42135 = ~x106 & n12501 ;
  assign n42136 = ~n42134 & ~n42135 ;
  assign n42137 = ~n42133 & n42136 ;
  assign n42138 = n12509 & n13034 ;
  assign n42139 = n42137 & ~n42138 ;
  assign n42140 = ~x44 & ~n42139 ;
  assign n42141 = ~x44 & ~n42140 ;
  assign n42142 = ~n42139 & ~n42140 ;
  assign n42143 = ~n42141 & ~n42142 ;
  assign n42144 = n42132 & ~n42143 ;
  assign n42145 = n42132 & ~n42144 ;
  assign n42146 = ~n42143 & ~n42144 ;
  assign n42147 = ~n42145 & ~n42146 ;
  assign n42148 = ~n41588 & ~n41594 ;
  assign n42149 = n42147 & n42148 ;
  assign n42150 = ~n42147 & ~n42148 ;
  assign n42151 = ~n42149 & ~n42150 ;
  assign n42152 = ~x110 & n10905 ;
  assign n42153 = ~x108 & n11466 ;
  assign n42154 = ~x109 & n10900 ;
  assign n42155 = ~n42153 & ~n42154 ;
  assign n42156 = ~n42152 & n42155 ;
  assign n42157 = n10908 & n14802 ;
  assign n42158 = n42156 & ~n42157 ;
  assign n42159 = ~x41 & ~n42158 ;
  assign n42160 = ~x41 & ~n42159 ;
  assign n42161 = ~n42158 & ~n42159 ;
  assign n42162 = ~n42160 & ~n42161 ;
  assign n42163 = n42151 & ~n42162 ;
  assign n42164 = n42151 & ~n42163 ;
  assign n42165 = ~n42162 & ~n42163 ;
  assign n42166 = ~n42164 & ~n42165 ;
  assign n42167 = ~n41607 & ~n41613 ;
  assign n42168 = n42166 & n42167 ;
  assign n42169 = ~n42166 & ~n42167 ;
  assign n42170 = ~n42168 & ~n42169 ;
  assign n42171 = ~x113 & n9433 ;
  assign n42172 = ~x111 & n9915 ;
  assign n42173 = ~x112 & n9428 ;
  assign n42174 = ~n42172 & ~n42173 ;
  assign n42175 = ~n42171 & n42174 ;
  assign n42176 = n9436 & n16684 ;
  assign n42177 = n42175 & ~n42176 ;
  assign n42178 = ~x38 & ~n42177 ;
  assign n42179 = ~x38 & ~n42178 ;
  assign n42180 = ~n42177 & ~n42178 ;
  assign n42181 = ~n42179 & ~n42180 ;
  assign n42182 = n42170 & ~n42181 ;
  assign n42183 = n42170 & ~n42182 ;
  assign n42184 = ~n42181 & ~n42182 ;
  assign n42185 = ~n42183 & ~n42184 ;
  assign n42186 = ~n41626 & ~n41632 ;
  assign n42187 = n42185 & n42186 ;
  assign n42188 = ~n42185 & ~n42186 ;
  assign n42189 = ~n42187 & ~n42188 ;
  assign n42190 = ~x116 & n8006 ;
  assign n42191 = ~x114 & n8474 ;
  assign n42192 = ~x115 & n8001 ;
  assign n42193 = ~n42191 & ~n42192 ;
  assign n42194 = ~n42190 & n42193 ;
  assign n42195 = n8009 & n18678 ;
  assign n42196 = n42194 & ~n42195 ;
  assign n42197 = ~x35 & ~n42196 ;
  assign n42198 = ~x35 & ~n42197 ;
  assign n42199 = ~n42196 & ~n42197 ;
  assign n42200 = ~n42198 & ~n42199 ;
  assign n42201 = n42189 & ~n42200 ;
  assign n42202 = n42189 & ~n42201 ;
  assign n42203 = ~n42200 & ~n42201 ;
  assign n42204 = ~n42202 & ~n42203 ;
  assign n42205 = ~n42012 & ~n42204 ;
  assign n42206 = n42012 & n42204 ;
  assign n42207 = n41998 & ~n42206 ;
  assign n42208 = ~n42205 & n42207 ;
  assign n42209 = n41998 & ~n42208 ;
  assign n42210 = ~n42206 & ~n42208 ;
  assign n42211 = ~n42205 & n42210 ;
  assign n42212 = ~n42209 & ~n42211 ;
  assign n42213 = n41983 & ~n42212 ;
  assign n42214 = ~n41983 & n42212 ;
  assign n42215 = n41967 & ~n42214 ;
  assign n42216 = ~n42213 & n42215 ;
  assign n42217 = n41967 & ~n42216 ;
  assign n42218 = ~n42214 & ~n42216 ;
  assign n42219 = ~n42213 & n42218 ;
  assign n42220 = ~n42217 & ~n42219 ;
  assign n42221 = ~n41403 & ~n41664 ;
  assign n42222 = n42220 & n42221 ;
  assign n42223 = ~n42220 & ~n42221 ;
  assign n42224 = ~n42222 & ~n42223 ;
  assign n42225 = ~n41671 & ~n41674 ;
  assign n42226 = n42224 & ~n42225 ;
  assign n42227 = ~n42224 & n42225 ;
  assign n42228 = ~n42226 & ~n42227 ;
  assign n42231 = ~n42228 & ~x213 ;
  assign n42232 = ~n42230 & ~n42231 ;
  assign n42233 = ~n41949 & ~n41952 ;
  assign n42234 = ~n41691 & ~n41942 ;
  assign n42235 = ~n41708 & ~n41939 ;
  assign n42236 = x127 & n3878 ;
  assign n42237 = n3592 & n26962 ;
  assign n42238 = ~n42236 & ~n42237 ;
  assign n42239 = x23 & ~n42238 ;
  assign n42240 = x23 & ~n42239 ;
  assign n42241 = ~n42238 & ~n42239 ;
  assign n42242 = ~n42240 & ~n42241 ;
  assign n42243 = ~n42235 & ~n42242 ;
  assign n42244 = ~n42235 & ~n42243 ;
  assign n42245 = ~n42242 & ~n42243 ;
  assign n42246 = ~n42244 & ~n42245 ;
  assign n42247 = x126 & n4531 ;
  assign n42248 = x124 & n4847 ;
  assign n42249 = x125 & n4526 ;
  assign n42250 = ~n42248 & ~n42249 ;
  assign n42251 = ~n42247 & n42250 ;
  assign n42252 = n4534 & n25735 ;
  assign n42253 = n42251 & ~n42252 ;
  assign n42254 = x26 & ~n42253 ;
  assign n42255 = x26 & ~n42254 ;
  assign n42256 = ~n42253 & ~n42254 ;
  assign n42257 = ~n42255 & ~n42256 ;
  assign n42258 = ~n41722 & ~n41934 ;
  assign n42259 = n42257 & n42258 ;
  assign n42260 = ~n42257 & ~n42258 ;
  assign n42261 = ~n42259 & ~n42260 ;
  assign n42262 = x123 & n5560 ;
  assign n42263 = x121 & n5943 ;
  assign n42264 = x122 & n5555 ;
  assign n42265 = ~n42263 & ~n42264 ;
  assign n42266 = ~n42262 & n42265 ;
  assign n42267 = n5563 & n23382 ;
  assign n42268 = n42266 & ~n42267 ;
  assign n42269 = x29 & ~n42268 ;
  assign n42270 = x29 & ~n42269 ;
  assign n42271 = ~n42268 & ~n42269 ;
  assign n42272 = ~n42270 & ~n42271 ;
  assign n42273 = ~n41363 & ~n41735 ;
  assign n42274 = ~n41931 & ~n42273 ;
  assign n42275 = ~n42272 & ~n42274 ;
  assign n42276 = ~n42272 & ~n42275 ;
  assign n42277 = ~n42274 & ~n42275 ;
  assign n42278 = ~n42276 & ~n42277 ;
  assign n42279 = x120 & n6725 ;
  assign n42280 = x118 & n7129 ;
  assign n42281 = x119 & n6720 ;
  assign n42282 = ~n42280 & ~n42281 ;
  assign n42283 = ~n42279 & n42282 ;
  assign n42284 = n6728 & n21143 ;
  assign n42285 = n42283 & ~n42284 ;
  assign n42286 = x32 & ~n42285 ;
  assign n42287 = x32 & ~n42286 ;
  assign n42288 = ~n42285 & ~n42286 ;
  assign n42289 = ~n42287 & ~n42288 ;
  assign n42290 = ~n41914 & ~n41927 ;
  assign n42291 = n42289 & n42290 ;
  assign n42292 = ~n42289 & ~n42290 ;
  assign n42293 = ~n42291 & ~n42292 ;
  assign n42294 = x117 & n8006 ;
  assign n42295 = x115 & n8474 ;
  assign n42296 = x116 & n8001 ;
  assign n42297 = ~n42295 & ~n42296 ;
  assign n42298 = ~n42294 & n42297 ;
  assign n42299 = n8009 & n19026 ;
  assign n42300 = n42298 & ~n42299 ;
  assign n42301 = x35 & ~n42300 ;
  assign n42302 = x35 & ~n42301 ;
  assign n42303 = ~n42300 & ~n42301 ;
  assign n42304 = ~n42302 & ~n42303 ;
  assign n42305 = ~n41895 & ~n41908 ;
  assign n42306 = ~n41856 & ~n41870 ;
  assign n42307 = x108 & n12506 ;
  assign n42308 = x106 & n13131 ;
  assign n42309 = x107 & n12501 ;
  assign n42310 = ~n42308 & ~n42309 ;
  assign n42311 = ~n42307 & n42310 ;
  assign n42312 = n12509 & n13323 ;
  assign n42313 = n42311 & ~n42312 ;
  assign n42314 = x44 & ~n42313 ;
  assign n42315 = x44 & ~n42314 ;
  assign n42316 = ~n42313 & ~n42314 ;
  assign n42317 = ~n42315 & ~n42316 ;
  assign n42318 = ~n41848 & ~n41852 ;
  assign n42319 = ~n41812 & ~n41825 ;
  assign n42320 = x99 & n18025 ;
  assign n42321 = x97 & n18764 ;
  assign n42322 = x98 & n18020 ;
  assign n42323 = ~n42321 & ~n42322 ;
  assign n42324 = ~n42320 & n42323 ;
  assign n42325 = n8660 & n18028 ;
  assign n42326 = n42324 & ~n42325 ;
  assign n42327 = x53 & ~n42326 ;
  assign n42328 = x53 & ~n42327 ;
  assign n42329 = ~n42326 & ~n42327 ;
  assign n42330 = ~n42328 & ~n42329 ;
  assign n42331 = ~n41792 & ~n41806 ;
  assign n42332 = ~n41770 & ~n41783 ;
  assign n42333 = x86 & n27024 ;
  assign n42334 = x87 & ~n26217 ;
  assign n42335 = ~n42333 & ~n42334 ;
  assign n42336 = ~n41767 & n42335 ;
  assign n42337 = n41767 & ~n42335 ;
  assign n42338 = ~n42336 & ~n42337 ;
  assign n42339 = x90 & n24612 ;
  assign n42340 = x88 & n25390 ;
  assign n42341 = x89 & n24607 ;
  assign n42342 = ~n42340 & ~n42341 ;
  assign n42343 = ~n42339 & n42342 ;
  assign n42344 = ~n24615 & n42343 ;
  assign n42345 = ~n4986 & n42343 ;
  assign n42346 = ~n42344 & ~n42345 ;
  assign n42347 = x62 & ~n42346 ;
  assign n42348 = ~x62 & n42346 ;
  assign n42349 = ~n42347 & ~n42348 ;
  assign n42350 = n42338 & ~n42349 ;
  assign n42351 = ~n42338 & n42349 ;
  assign n42352 = ~n42350 & ~n42351 ;
  assign n42353 = ~n42332 & n42352 ;
  assign n42354 = n42332 & ~n42352 ;
  assign n42355 = ~n42353 & ~n42354 ;
  assign n42356 = x93 & n22325 ;
  assign n42357 = x91 & n23066 ;
  assign n42358 = x92 & n22320 ;
  assign n42359 = ~n42357 & ~n42358 ;
  assign n42360 = ~n42356 & n42359 ;
  assign n42361 = n6094 & n22328 ;
  assign n42362 = n42360 & ~n42361 ;
  assign n42363 = x59 & ~n42362 ;
  assign n42364 = x59 & ~n42363 ;
  assign n42365 = ~n42362 & ~n42363 ;
  assign n42366 = ~n42364 & ~n42365 ;
  assign n42367 = n42355 & ~n42366 ;
  assign n42368 = n42355 & ~n42367 ;
  assign n42369 = ~n42366 & ~n42367 ;
  assign n42370 = ~n42368 & ~n42369 ;
  assign n42371 = ~n41786 & ~n41789 ;
  assign n42372 = n42370 & n42371 ;
  assign n42373 = ~n42370 & ~n42371 ;
  assign n42374 = ~n42372 & ~n42373 ;
  assign n42375 = x96 & n20143 ;
  assign n42376 = x94 & n20854 ;
  assign n42377 = x95 & n20138 ;
  assign n42378 = ~n42376 & ~n42377 ;
  assign n42379 = ~n42375 & n42378 ;
  assign n42380 = n7321 & n20146 ;
  assign n42381 = n42379 & ~n42380 ;
  assign n42382 = x56 & ~n42381 ;
  assign n42383 = x56 & ~n42382 ;
  assign n42384 = ~n42381 & ~n42382 ;
  assign n42385 = ~n42383 & ~n42384 ;
  assign n42386 = ~n42374 & n42385 ;
  assign n42387 = n42374 & ~n42385 ;
  assign n42388 = ~n42386 & ~n42387 ;
  assign n42389 = ~n42331 & n42388 ;
  assign n42390 = n42331 & ~n42388 ;
  assign n42391 = ~n42389 & ~n42390 ;
  assign n42392 = ~n42330 & n42391 ;
  assign n42393 = n42330 & ~n42391 ;
  assign n42394 = ~n42392 & ~n42393 ;
  assign n42395 = ~n42319 & n42394 ;
  assign n42396 = n42319 & ~n42394 ;
  assign n42397 = ~n42395 & ~n42396 ;
  assign n42398 = x102 & n16076 ;
  assign n42399 = x100 & n16756 ;
  assign n42400 = x101 & n16071 ;
  assign n42401 = ~n42399 & ~n42400 ;
  assign n42402 = ~n42398 & n42401 ;
  assign n42403 = n10092 & n16079 ;
  assign n42404 = n42402 & ~n42403 ;
  assign n42405 = x50 & ~n42404 ;
  assign n42406 = x50 & ~n42405 ;
  assign n42407 = ~n42404 & ~n42405 ;
  assign n42408 = ~n42406 & ~n42407 ;
  assign n42409 = n42397 & ~n42408 ;
  assign n42410 = n42397 & ~n42409 ;
  assign n42411 = ~n42408 & ~n42409 ;
  assign n42412 = ~n42410 & ~n42411 ;
  assign n42413 = ~n41832 & ~n41846 ;
  assign n42414 = ~n42412 & ~n42413 ;
  assign n42415 = ~n42412 & ~n42414 ;
  assign n42416 = ~n42413 & ~n42414 ;
  assign n42417 = ~n42415 & ~n42416 ;
  assign n42418 = x105 & n14233 ;
  assign n42419 = x103 & n14876 ;
  assign n42420 = x104 & n14228 ;
  assign n42421 = ~n42419 & ~n42420 ;
  assign n42422 = ~n42418 & n42421 ;
  assign n42423 = n11648 & n14236 ;
  assign n42424 = n42422 & ~n42423 ;
  assign n42425 = x47 & ~n42424 ;
  assign n42426 = x47 & ~n42425 ;
  assign n42427 = ~n42424 & ~n42425 ;
  assign n42428 = ~n42426 & ~n42427 ;
  assign n42429 = ~n42417 & n42428 ;
  assign n42430 = n42417 & ~n42428 ;
  assign n42431 = ~n42429 & ~n42430 ;
  assign n42432 = ~n42318 & ~n42431 ;
  assign n42433 = n42318 & n42431 ;
  assign n42434 = ~n42432 & ~n42433 ;
  assign n42435 = ~n42317 & n42434 ;
  assign n42436 = n42317 & ~n42434 ;
  assign n42437 = ~n42435 & ~n42436 ;
  assign n42438 = ~n42306 & n42437 ;
  assign n42439 = n42306 & ~n42437 ;
  assign n42440 = ~n42438 & ~n42439 ;
  assign n42441 = x111 & n10905 ;
  assign n42442 = x109 & n11466 ;
  assign n42443 = x110 & n10900 ;
  assign n42444 = ~n42442 & ~n42443 ;
  assign n42445 = ~n42441 & n42444 ;
  assign n42446 = n10908 & n15111 ;
  assign n42447 = n42445 & ~n42446 ;
  assign n42448 = x41 & ~n42447 ;
  assign n42449 = x41 & ~n42448 ;
  assign n42450 = ~n42447 & ~n42448 ;
  assign n42451 = ~n42449 & ~n42450 ;
  assign n42452 = n42440 & ~n42451 ;
  assign n42453 = n42440 & ~n42452 ;
  assign n42454 = ~n42451 & ~n42452 ;
  assign n42455 = ~n42453 & ~n42454 ;
  assign n42456 = ~n41876 & ~n41889 ;
  assign n42457 = n42455 & n42456 ;
  assign n42458 = ~n42455 & ~n42456 ;
  assign n42459 = ~n42457 & ~n42458 ;
  assign n42460 = x114 & n9433 ;
  assign n42461 = x112 & n9915 ;
  assign n42462 = x113 & n9428 ;
  assign n42463 = ~n42461 & ~n42462 ;
  assign n42464 = ~n42460 & n42463 ;
  assign n42465 = n9436 & n17012 ;
  assign n42466 = n42464 & ~n42465 ;
  assign n42467 = x38 & ~n42466 ;
  assign n42468 = x38 & ~n42467 ;
  assign n42469 = ~n42466 & ~n42467 ;
  assign n42470 = ~n42468 & ~n42469 ;
  assign n42471 = ~n42459 & n42470 ;
  assign n42472 = n42459 & ~n42470 ;
  assign n42473 = ~n42471 & ~n42472 ;
  assign n42474 = ~n42305 & n42473 ;
  assign n42475 = ~n42305 & ~n42474 ;
  assign n42476 = n42473 & ~n42474 ;
  assign n42477 = ~n42475 & ~n42476 ;
  assign n42478 = ~n42304 & ~n42477 ;
  assign n42479 = ~n42304 & ~n42478 ;
  assign n42480 = ~n42477 & ~n42478 ;
  assign n42481 = ~n42479 & ~n42480 ;
  assign n42482 = n42293 & ~n42481 ;
  assign n42483 = n42293 & ~n42482 ;
  assign n42484 = ~n42481 & ~n42482 ;
  assign n42485 = ~n42483 & ~n42484 ;
  assign n42486 = ~n42278 & n42485 ;
  assign n42487 = n42278 & ~n42485 ;
  assign n42488 = ~n42486 & ~n42487 ;
  assign n42489 = n42261 & ~n42488 ;
  assign n42490 = n42261 & ~n42489 ;
  assign n42491 = ~n42488 & ~n42489 ;
  assign n42492 = ~n42490 & ~n42491 ;
  assign n42493 = ~n42246 & n42492 ;
  assign n42494 = n42246 & ~n42492 ;
  assign n42495 = ~n42493 & ~n42494 ;
  assign n42496 = ~n42234 & ~n42495 ;
  assign n42497 = ~n42234 & ~n42496 ;
  assign n42498 = ~n42495 & ~n42496 ;
  assign n42499 = ~n42497 & ~n42498 ;
  assign n42500 = ~n42233 & ~n42499 ;
  assign n42501 = n42233 & ~n42498 ;
  assign n42502 = ~n42497 & n42501 ;
  assign n42503 = ~n42500 & ~n42502 ;
  assign n42776 = n42503 & x214 ;
  assign n42504 = ~n42223 & ~n42226 ;
  assign n42505 = ~n41965 & ~n42216 ;
  assign n42506 = ~n41982 & ~n42213 ;
  assign n42507 = ~x127 & n3878 ;
  assign n42508 = n3592 & n27365 ;
  assign n42509 = ~n42507 & ~n42508 ;
  assign n42510 = ~x23 & ~n42509 ;
  assign n42511 = ~x23 & ~n42510 ;
  assign n42512 = ~n42509 & ~n42510 ;
  assign n42513 = ~n42511 & ~n42512 ;
  assign n42514 = ~n42506 & ~n42513 ;
  assign n42515 = ~n42506 & ~n42514 ;
  assign n42516 = ~n42513 & ~n42514 ;
  assign n42517 = ~n42515 & ~n42516 ;
  assign n42518 = ~x126 & n4531 ;
  assign n42519 = ~x124 & n4847 ;
  assign n42520 = ~x125 & n4526 ;
  assign n42521 = ~n42519 & ~n42520 ;
  assign n42522 = ~n42518 & n42521 ;
  assign n42523 = n4534 & n26128 ;
  assign n42524 = n42522 & ~n42523 ;
  assign n42525 = ~x26 & ~n42524 ;
  assign n42526 = ~x26 & ~n42525 ;
  assign n42527 = ~n42524 & ~n42525 ;
  assign n42528 = ~n42526 & ~n42527 ;
  assign n42529 = ~n41996 & ~n42208 ;
  assign n42530 = n42528 & n42529 ;
  assign n42531 = ~n42528 & ~n42529 ;
  assign n42532 = ~n42530 & ~n42531 ;
  assign n42533 = ~x123 & n5560 ;
  assign n42534 = ~x121 & n5943 ;
  assign n42535 = ~x122 & n5555 ;
  assign n42536 = ~n42534 & ~n42535 ;
  assign n42537 = ~n42533 & n42536 ;
  assign n42538 = n5563 & n23760 ;
  assign n42539 = n42537 & ~n42538 ;
  assign n42540 = ~x29 & ~n42539 ;
  assign n42541 = ~x29 & ~n42540 ;
  assign n42542 = ~n42539 & ~n42540 ;
  assign n42543 = ~n42541 & ~n42542 ;
  assign n42544 = ~n41650 & ~n42009 ;
  assign n42545 = ~n42205 & ~n42544 ;
  assign n42546 = ~n42543 & ~n42545 ;
  assign n42547 = ~n42543 & ~n42546 ;
  assign n42548 = ~n42545 & ~n42546 ;
  assign n42549 = ~n42547 & ~n42548 ;
  assign n42550 = ~x120 & n6725 ;
  assign n42551 = ~x118 & n7129 ;
  assign n42552 = ~x119 & n6720 ;
  assign n42553 = ~n42551 & ~n42552 ;
  assign n42554 = ~n42550 & n42553 ;
  assign n42555 = n6728 & n21501 ;
  assign n42556 = n42554 & ~n42555 ;
  assign n42557 = ~x32 & ~n42556 ;
  assign n42558 = ~x32 & ~n42557 ;
  assign n42559 = ~n42556 & ~n42557 ;
  assign n42560 = ~n42558 & ~n42559 ;
  assign n42561 = ~n42188 & ~n42201 ;
  assign n42562 = n42560 & n42561 ;
  assign n42563 = ~n42560 & ~n42561 ;
  assign n42564 = ~n42562 & ~n42563 ;
  assign n42565 = ~x117 & n8006 ;
  assign n42566 = ~x115 & n8474 ;
  assign n42567 = ~x116 & n8001 ;
  assign n42568 = ~n42566 & ~n42567 ;
  assign n42569 = ~n42565 & n42568 ;
  assign n42570 = n8009 & n19365 ;
  assign n42571 = n42569 & ~n42570 ;
  assign n42572 = ~x35 & ~n42571 ;
  assign n42573 = ~x35 & ~n42572 ;
  assign n42574 = ~n42571 & ~n42572 ;
  assign n42575 = ~n42573 & ~n42574 ;
  assign n42576 = ~n42169 & ~n42182 ;
  assign n42577 = ~n42130 & ~n42144 ;
  assign n42578 = ~x108 & n12506 ;
  assign n42579 = ~x106 & n13131 ;
  assign n42580 = ~x107 & n12501 ;
  assign n42581 = ~n42579 & ~n42580 ;
  assign n42582 = ~n42578 & n42581 ;
  assign n42583 = n12509 & n13601 ;
  assign n42584 = n42582 & ~n42583 ;
  assign n42585 = ~x44 & ~n42584 ;
  assign n42586 = ~x44 & ~n42585 ;
  assign n42587 = ~n42584 & ~n42585 ;
  assign n42588 = ~n42586 & ~n42587 ;
  assign n42589 = ~n42122 & ~n42126 ;
  assign n42590 = ~n42086 & ~n42099 ;
  assign n42591 = ~x99 & n18025 ;
  assign n42592 = ~x97 & n18764 ;
  assign n42593 = ~x98 & n18020 ;
  assign n42594 = ~n42592 & ~n42593 ;
  assign n42595 = ~n42591 & n42594 ;
  assign n42596 = n8885 & n18028 ;
  assign n42597 = n42595 & ~n42596 ;
  assign n42598 = ~x53 & ~n42597 ;
  assign n42599 = ~x53 & ~n42598 ;
  assign n42600 = ~n42597 & ~n42598 ;
  assign n42601 = ~n42599 & ~n42600 ;
  assign n42602 = ~n42066 & ~n42080 ;
  assign n42603 = ~n42044 & ~n42057 ;
  assign n42604 = ~x86 & n27427 ;
  assign n42605 = ~x87 & ~n26217 ;
  assign n42606 = ~n42604 & ~n42605 ;
  assign n42607 = ~n42041 & n42606 ;
  assign n42608 = n42041 & ~n42606 ;
  assign n42609 = ~n42607 & ~n42608 ;
  assign n42610 = ~x90 & n24612 ;
  assign n42611 = ~x88 & n25390 ;
  assign n42612 = ~x89 & n24607 ;
  assign n42613 = ~n42611 & ~n42612 ;
  assign n42614 = ~n42610 & n42613 ;
  assign n42615 = ~n24615 & n42614 ;
  assign n42616 = ~n5155 & n42614 ;
  assign n42617 = ~n42615 & ~n42616 ;
  assign n42618 = ~x62 & ~n42617 ;
  assign n42619 = x62 & n42617 ;
  assign n42620 = ~n42618 & ~n42619 ;
  assign n42621 = n42609 & ~n42620 ;
  assign n42622 = ~n42609 & n42620 ;
  assign n42623 = ~n42621 & ~n42622 ;
  assign n42624 = ~n42603 & n42623 ;
  assign n42625 = n42603 & ~n42623 ;
  assign n42626 = ~n42624 & ~n42625 ;
  assign n42627 = ~x93 & n22325 ;
  assign n42628 = ~x91 & n23066 ;
  assign n42629 = ~x92 & n22320 ;
  assign n42630 = ~n42628 & ~n42629 ;
  assign n42631 = ~n42627 & n42630 ;
  assign n42632 = n6285 & n22328 ;
  assign n42633 = n42631 & ~n42632 ;
  assign n42634 = ~x59 & ~n42633 ;
  assign n42635 = ~x59 & ~n42634 ;
  assign n42636 = ~n42633 & ~n42634 ;
  assign n42637 = ~n42635 & ~n42636 ;
  assign n42638 = n42626 & ~n42637 ;
  assign n42639 = n42626 & ~n42638 ;
  assign n42640 = ~n42637 & ~n42638 ;
  assign n42641 = ~n42639 & ~n42640 ;
  assign n42642 = ~n42060 & ~n42063 ;
  assign n42643 = n42641 & n42642 ;
  assign n42644 = ~n42641 & ~n42642 ;
  assign n42645 = ~n42643 & ~n42644 ;
  assign n42646 = ~x96 & n20143 ;
  assign n42647 = ~x94 & n20854 ;
  assign n42648 = ~x95 & n20138 ;
  assign n42649 = ~n42647 & ~n42648 ;
  assign n42650 = ~n42646 & n42649 ;
  assign n42651 = n7531 & n20146 ;
  assign n42652 = n42650 & ~n42651 ;
  assign n42653 = ~x56 & ~n42652 ;
  assign n42654 = ~x56 & ~n42653 ;
  assign n42655 = ~n42652 & ~n42653 ;
  assign n42656 = ~n42654 & ~n42655 ;
  assign n42657 = ~n42645 & n42656 ;
  assign n42658 = n42645 & ~n42656 ;
  assign n42659 = ~n42657 & ~n42658 ;
  assign n42660 = ~n42602 & n42659 ;
  assign n42661 = n42602 & ~n42659 ;
  assign n42662 = ~n42660 & ~n42661 ;
  assign n42663 = ~n42601 & n42662 ;
  assign n42664 = n42601 & ~n42662 ;
  assign n42665 = ~n42663 & ~n42664 ;
  assign n42666 = ~n42590 & n42665 ;
  assign n42667 = n42590 & ~n42665 ;
  assign n42668 = ~n42666 & ~n42667 ;
  assign n42669 = ~x102 & n16076 ;
  assign n42670 = ~x100 & n16756 ;
  assign n42671 = ~x101 & n16071 ;
  assign n42672 = ~n42670 & ~n42671 ;
  assign n42673 = ~n42669 & n42672 ;
  assign n42674 = n10333 & n16079 ;
  assign n42675 = n42673 & ~n42674 ;
  assign n42676 = ~x50 & ~n42675 ;
  assign n42677 = ~x50 & ~n42676 ;
  assign n42678 = ~n42675 & ~n42676 ;
  assign n42679 = ~n42677 & ~n42678 ;
  assign n42680 = n42668 & ~n42679 ;
  assign n42681 = n42668 & ~n42680 ;
  assign n42682 = ~n42679 & ~n42680 ;
  assign n42683 = ~n42681 & ~n42682 ;
  assign n42684 = ~n42106 & ~n42120 ;
  assign n42685 = ~n42683 & ~n42684 ;
  assign n42686 = ~n42683 & ~n42685 ;
  assign n42687 = ~n42684 & ~n42685 ;
  assign n42688 = ~n42686 & ~n42687 ;
  assign n42689 = ~x105 & n14233 ;
  assign n42690 = ~x103 & n14876 ;
  assign n42691 = ~x104 & n14228 ;
  assign n42692 = ~n42690 & ~n42691 ;
  assign n42693 = ~n42689 & n42692 ;
  assign n42694 = n11907 & n14236 ;
  assign n42695 = n42693 & ~n42694 ;
  assign n42696 = ~x47 & ~n42695 ;
  assign n42697 = ~x47 & ~n42696 ;
  assign n42698 = ~n42695 & ~n42696 ;
  assign n42699 = ~n42697 & ~n42698 ;
  assign n42700 = ~n42688 & n42699 ;
  assign n42701 = n42688 & ~n42699 ;
  assign n42702 = ~n42700 & ~n42701 ;
  assign n42703 = ~n42589 & ~n42702 ;
  assign n42704 = n42589 & n42702 ;
  assign n42705 = ~n42703 & ~n42704 ;
  assign n42706 = ~n42588 & n42705 ;
  assign n42707 = n42588 & ~n42705 ;
  assign n42708 = ~n42706 & ~n42707 ;
  assign n42709 = ~n42577 & n42708 ;
  assign n42710 = n42577 & ~n42708 ;
  assign n42711 = ~n42709 & ~n42710 ;
  assign n42712 = ~x111 & n10905 ;
  assign n42713 = ~x109 & n11466 ;
  assign n42714 = ~x110 & n10900 ;
  assign n42715 = ~n42713 & ~n42714 ;
  assign n42716 = ~n42712 & n42715 ;
  assign n42717 = n10908 & n15411 ;
  assign n42718 = n42716 & ~n42717 ;
  assign n42719 = ~x41 & ~n42718 ;
  assign n42720 = ~x41 & ~n42719 ;
  assign n42721 = ~n42718 & ~n42719 ;
  assign n42722 = ~n42720 & ~n42721 ;
  assign n42723 = n42711 & ~n42722 ;
  assign n42724 = n42711 & ~n42723 ;
  assign n42725 = ~n42722 & ~n42723 ;
  assign n42726 = ~n42724 & ~n42725 ;
  assign n42727 = ~n42150 & ~n42163 ;
  assign n42728 = n42726 & n42727 ;
  assign n42729 = ~n42726 & ~n42727 ;
  assign n42730 = ~n42728 & ~n42729 ;
  assign n42731 = ~x114 & n9433 ;
  assign n42732 = ~x112 & n9915 ;
  assign n42733 = ~x113 & n9428 ;
  assign n42734 = ~n42732 & ~n42733 ;
  assign n42735 = ~n42731 & n42734 ;
  assign n42736 = n9436 & n17333 ;
  assign n42737 = n42735 & ~n42736 ;
  assign n42738 = ~x38 & ~n42737 ;
  assign n42739 = ~x38 & ~n42738 ;
  assign n42740 = ~n42737 & ~n42738 ;
  assign n42741 = ~n42739 & ~n42740 ;
  assign n42742 = ~n42730 & n42741 ;
  assign n42743 = n42730 & ~n42741 ;
  assign n42744 = ~n42742 & ~n42743 ;
  assign n42745 = ~n42576 & n42744 ;
  assign n42746 = ~n42576 & ~n42745 ;
  assign n42747 = n42744 & ~n42745 ;
  assign n42748 = ~n42746 & ~n42747 ;
  assign n42749 = ~n42575 & ~n42748 ;
  assign n42750 = ~n42575 & ~n42749 ;
  assign n42751 = ~n42748 & ~n42749 ;
  assign n42752 = ~n42750 & ~n42751 ;
  assign n42753 = n42564 & ~n42752 ;
  assign n42754 = n42564 & ~n42753 ;
  assign n42755 = ~n42752 & ~n42753 ;
  assign n42756 = ~n42754 & ~n42755 ;
  assign n42757 = ~n42549 & n42756 ;
  assign n42758 = n42549 & ~n42756 ;
  assign n42759 = ~n42757 & ~n42758 ;
  assign n42760 = n42532 & ~n42759 ;
  assign n42761 = n42532 & ~n42760 ;
  assign n42762 = ~n42759 & ~n42760 ;
  assign n42763 = ~n42761 & ~n42762 ;
  assign n42764 = ~n42517 & n42763 ;
  assign n42765 = n42517 & ~n42763 ;
  assign n42766 = ~n42764 & ~n42765 ;
  assign n42767 = ~n42505 & ~n42766 ;
  assign n42768 = ~n42505 & ~n42767 ;
  assign n42769 = ~n42766 & ~n42767 ;
  assign n42770 = ~n42768 & ~n42769 ;
  assign n42771 = ~n42504 & ~n42770 ;
  assign n42772 = n42504 & ~n42769 ;
  assign n42773 = ~n42768 & n42772 ;
  assign n42774 = ~n42771 & ~n42773 ;
  assign n42777 = ~n42774 & ~x214 ;
  assign n42778 = ~n42776 & ~n42777 ;
  assign n42779 = ~n42496 & ~n42500 ;
  assign n42780 = ~n42246 & ~n42492 ;
  assign n42781 = ~n42243 & ~n42780 ;
  assign n42782 = ~n42260 & ~n42489 ;
  assign n42783 = x127 & n4531 ;
  assign n42784 = x125 & n4847 ;
  assign n42785 = x126 & n4526 ;
  assign n42786 = ~n42784 & ~n42785 ;
  assign n42787 = ~n42783 & n42786 ;
  assign n42788 = n4534 & n26533 ;
  assign n42789 = n42787 & ~n42788 ;
  assign n42790 = x26 & ~n42789 ;
  assign n42791 = x26 & ~n42790 ;
  assign n42792 = ~n42789 & ~n42790 ;
  assign n42793 = ~n42791 & ~n42792 ;
  assign n42794 = ~n42782 & ~n42793 ;
  assign n42795 = ~n42782 & ~n42794 ;
  assign n42796 = ~n42793 & ~n42794 ;
  assign n42797 = ~n42795 & ~n42796 ;
  assign n42798 = ~n42278 & ~n42485 ;
  assign n42799 = ~n42275 & ~n42798 ;
  assign n42800 = x124 & n5560 ;
  assign n42801 = x122 & n5943 ;
  assign n42802 = x123 & n5555 ;
  assign n42803 = ~n42801 & ~n42802 ;
  assign n42804 = ~n42800 & n42803 ;
  assign n42805 = n5563 & n23796 ;
  assign n42806 = n42804 & ~n42805 ;
  assign n42807 = x29 & ~n42806 ;
  assign n42808 = x29 & ~n42807 ;
  assign n42809 = ~n42806 & ~n42807 ;
  assign n42810 = ~n42808 & ~n42809 ;
  assign n42811 = ~n42799 & n42810 ;
  assign n42812 = n42799 & ~n42810 ;
  assign n42813 = ~n42811 & ~n42812 ;
  assign n42814 = x121 & n6725 ;
  assign n42815 = x119 & n7129 ;
  assign n42816 = x120 & n6720 ;
  assign n42817 = ~n42815 & ~n42816 ;
  assign n42818 = ~n42814 & n42817 ;
  assign n42819 = n6728 & n21870 ;
  assign n42820 = n42818 & ~n42819 ;
  assign n42821 = x32 & ~n42820 ;
  assign n42822 = x32 & ~n42821 ;
  assign n42823 = ~n42820 & ~n42821 ;
  assign n42824 = ~n42822 & ~n42823 ;
  assign n42825 = ~n42292 & ~n42482 ;
  assign n42826 = n42824 & n42825 ;
  assign n42827 = ~n42824 & ~n42825 ;
  assign n42828 = ~n42826 & ~n42827 ;
  assign n42829 = ~n42474 & ~n42478 ;
  assign n42830 = ~n42458 & ~n42472 ;
  assign n42831 = ~n42432 & ~n42435 ;
  assign n42832 = ~n42417 & ~n42428 ;
  assign n42833 = ~n42414 & ~n42832 ;
  assign n42834 = ~n42353 & ~n42367 ;
  assign n42835 = ~n42336 & ~n42350 ;
  assign n42836 = x87 & n27024 ;
  assign n42837 = x88 & ~n26217 ;
  assign n42838 = ~n42836 & ~n42837 ;
  assign n42839 = ~x23 & ~n42838 ;
  assign n42840 = x23 & n42838 ;
  assign n42841 = ~n42839 & ~n42840 ;
  assign n42842 = ~n42335 & n42841 ;
  assign n42843 = n42335 & ~n42841 ;
  assign n42844 = ~n42842 & ~n42843 ;
  assign n42845 = x91 & n24612 ;
  assign n42846 = x89 & n25390 ;
  assign n42847 = x90 & n24607 ;
  assign n42848 = ~n42846 & ~n42847 ;
  assign n42849 = ~n42845 & n42848 ;
  assign n42850 = n5336 & n24615 ;
  assign n42851 = n42849 & ~n42850 ;
  assign n42852 = x62 & ~n42851 ;
  assign n42853 = x62 & ~n42852 ;
  assign n42854 = ~n42851 & ~n42852 ;
  assign n42855 = ~n42853 & ~n42854 ;
  assign n42856 = n42844 & ~n42855 ;
  assign n42857 = n42844 & ~n42856 ;
  assign n42858 = ~n42855 & ~n42856 ;
  assign n42859 = ~n42857 & ~n42858 ;
  assign n42860 = ~n42835 & n42859 ;
  assign n42861 = n42835 & ~n42859 ;
  assign n42862 = ~n42860 & ~n42861 ;
  assign n42863 = x94 & n22325 ;
  assign n42864 = x92 & n23066 ;
  assign n42865 = x93 & n22320 ;
  assign n42866 = ~n42864 & ~n42865 ;
  assign n42867 = ~n42863 & n42866 ;
  assign n42868 = n6483 & n22328 ;
  assign n42869 = n42867 & ~n42868 ;
  assign n42870 = x59 & ~n42869 ;
  assign n42871 = x59 & ~n42870 ;
  assign n42872 = ~n42869 & ~n42870 ;
  assign n42873 = ~n42871 & ~n42872 ;
  assign n42874 = ~n42862 & ~n42873 ;
  assign n42875 = n42862 & n42873 ;
  assign n42876 = ~n42874 & ~n42875 ;
  assign n42877 = n42834 & ~n42876 ;
  assign n42878 = ~n42834 & n42876 ;
  assign n42879 = ~n42877 & ~n42878 ;
  assign n42880 = x97 & n20143 ;
  assign n42881 = x95 & n20854 ;
  assign n42882 = x96 & n20138 ;
  assign n42883 = ~n42881 & ~n42882 ;
  assign n42884 = ~n42880 & n42883 ;
  assign n42885 = n7745 & n20146 ;
  assign n42886 = n42884 & ~n42885 ;
  assign n42887 = x56 & ~n42886 ;
  assign n42888 = x56 & ~n42887 ;
  assign n42889 = ~n42886 & ~n42887 ;
  assign n42890 = ~n42888 & ~n42889 ;
  assign n42891 = ~n42373 & ~n42387 ;
  assign n42892 = ~n42890 & ~n42891 ;
  assign n42893 = n42890 & n42891 ;
  assign n42894 = ~n42892 & ~n42893 ;
  assign n42895 = n42879 & n42894 ;
  assign n42896 = ~n42879 & ~n42894 ;
  assign n42897 = ~n42895 & ~n42896 ;
  assign n42898 = x100 & n18025 ;
  assign n42899 = x98 & n18764 ;
  assign n42900 = x99 & n18020 ;
  assign n42901 = ~n42899 & ~n42900 ;
  assign n42902 = ~n42898 & n42901 ;
  assign n42903 = n9115 & n18028 ;
  assign n42904 = n42902 & ~n42903 ;
  assign n42905 = x53 & ~n42904 ;
  assign n42906 = x53 & ~n42905 ;
  assign n42907 = ~n42904 & ~n42905 ;
  assign n42908 = ~n42906 & ~n42907 ;
  assign n42909 = n42897 & ~n42908 ;
  assign n42910 = n42897 & ~n42909 ;
  assign n42911 = ~n42908 & ~n42909 ;
  assign n42912 = ~n42910 & ~n42911 ;
  assign n42913 = ~n42389 & ~n42392 ;
  assign n42914 = n42912 & n42913 ;
  assign n42915 = ~n42912 & ~n42913 ;
  assign n42916 = ~n42914 & ~n42915 ;
  assign n42917 = x103 & n16076 ;
  assign n42918 = x101 & n16756 ;
  assign n42919 = x102 & n16071 ;
  assign n42920 = ~n42918 & ~n42919 ;
  assign n42921 = ~n42917 & n42920 ;
  assign n42922 = n10588 & n16079 ;
  assign n42923 = n42921 & ~n42922 ;
  assign n42924 = x50 & ~n42923 ;
  assign n42925 = x50 & ~n42924 ;
  assign n42926 = ~n42923 & ~n42924 ;
  assign n42927 = ~n42925 & ~n42926 ;
  assign n42928 = n42916 & ~n42927 ;
  assign n42929 = n42916 & ~n42928 ;
  assign n42930 = ~n42927 & ~n42928 ;
  assign n42931 = ~n42929 & ~n42930 ;
  assign n42932 = ~n42395 & ~n42409 ;
  assign n42933 = n42931 & n42932 ;
  assign n42934 = ~n42931 & ~n42932 ;
  assign n42935 = ~n42933 & ~n42934 ;
  assign n42936 = x106 & n14233 ;
  assign n42937 = x104 & n14876 ;
  assign n42938 = x105 & n14228 ;
  assign n42939 = ~n42937 & ~n42938 ;
  assign n42940 = ~n42936 & n42939 ;
  assign n42941 = n12181 & n14236 ;
  assign n42942 = n42940 & ~n42941 ;
  assign n42943 = x47 & ~n42942 ;
  assign n42944 = x47 & ~n42943 ;
  assign n42945 = ~n42942 & ~n42943 ;
  assign n42946 = ~n42944 & ~n42945 ;
  assign n42947 = n42935 & ~n42946 ;
  assign n42948 = n42935 & ~n42947 ;
  assign n42949 = ~n42946 & ~n42947 ;
  assign n42950 = ~n42948 & ~n42949 ;
  assign n42951 = ~n42833 & n42950 ;
  assign n42952 = n42833 & ~n42950 ;
  assign n42953 = ~n42951 & ~n42952 ;
  assign n42954 = x109 & n12506 ;
  assign n42955 = x107 & n13131 ;
  assign n42956 = x108 & n12501 ;
  assign n42957 = ~n42955 & ~n42956 ;
  assign n42958 = ~n42954 & n42957 ;
  assign n42959 = n12509 & n13894 ;
  assign n42960 = n42958 & ~n42959 ;
  assign n42961 = x44 & ~n42960 ;
  assign n42962 = x44 & ~n42961 ;
  assign n42963 = ~n42960 & ~n42961 ;
  assign n42964 = ~n42962 & ~n42963 ;
  assign n42965 = ~n42953 & ~n42964 ;
  assign n42966 = n42953 & n42964 ;
  assign n42967 = ~n42965 & ~n42966 ;
  assign n42968 = n42831 & ~n42967 ;
  assign n42969 = ~n42831 & n42967 ;
  assign n42970 = ~n42968 & ~n42969 ;
  assign n42971 = x112 & n10905 ;
  assign n42972 = x110 & n11466 ;
  assign n42973 = x111 & n10900 ;
  assign n42974 = ~n42972 & ~n42973 ;
  assign n42975 = ~n42971 & n42974 ;
  assign n42976 = n10908 & n15442 ;
  assign n42977 = n42975 & ~n42976 ;
  assign n42978 = x41 & ~n42977 ;
  assign n42979 = x41 & ~n42978 ;
  assign n42980 = ~n42977 & ~n42978 ;
  assign n42981 = ~n42979 & ~n42980 ;
  assign n42982 = n42970 & ~n42981 ;
  assign n42983 = n42970 & ~n42982 ;
  assign n42984 = ~n42981 & ~n42982 ;
  assign n42985 = ~n42983 & ~n42984 ;
  assign n42986 = ~n42438 & ~n42452 ;
  assign n42987 = n42985 & n42986 ;
  assign n42988 = ~n42985 & ~n42986 ;
  assign n42989 = ~n42987 & ~n42988 ;
  assign n42990 = x115 & n9433 ;
  assign n42991 = x113 & n9915 ;
  assign n42992 = x114 & n9428 ;
  assign n42993 = ~n42991 & ~n42992 ;
  assign n42994 = ~n42990 & n42993 ;
  assign n42995 = n9436 & n17364 ;
  assign n42996 = n42994 & ~n42995 ;
  assign n42997 = x38 & ~n42996 ;
  assign n42998 = x38 & ~n42997 ;
  assign n42999 = ~n42996 & ~n42997 ;
  assign n43000 = ~n42998 & ~n42999 ;
  assign n43001 = n42989 & ~n43000 ;
  assign n43002 = ~n42989 & n43000 ;
  assign n43003 = ~n42830 & ~n43002 ;
  assign n43004 = ~n43001 & n43003 ;
  assign n43005 = ~n42830 & ~n43004 ;
  assign n43006 = ~n43001 & ~n43004 ;
  assign n43007 = ~n43002 & n43006 ;
  assign n43008 = ~n43005 & ~n43007 ;
  assign n43009 = x118 & n8006 ;
  assign n43010 = x116 & n8474 ;
  assign n43011 = x117 & n8001 ;
  assign n43012 = ~n43010 & ~n43011 ;
  assign n43013 = ~n43009 & n43012 ;
  assign n43014 = n8009 & n19395 ;
  assign n43015 = n43013 & ~n43014 ;
  assign n43016 = x35 & ~n43015 ;
  assign n43017 = x35 & ~n43016 ;
  assign n43018 = ~n43015 & ~n43016 ;
  assign n43019 = ~n43017 & ~n43018 ;
  assign n43020 = n43008 & n43019 ;
  assign n43021 = ~n43008 & ~n43019 ;
  assign n43022 = ~n43020 & ~n43021 ;
  assign n43023 = ~n42829 & n43022 ;
  assign n43024 = n42829 & ~n43022 ;
  assign n43025 = ~n43023 & ~n43024 ;
  assign n43026 = n42828 & n43025 ;
  assign n43027 = ~n42828 & ~n43025 ;
  assign n43028 = ~n42813 & ~n43027 ;
  assign n43029 = ~n43026 & n43028 ;
  assign n43030 = ~n42813 & ~n43029 ;
  assign n43031 = ~n43027 & ~n43029 ;
  assign n43032 = ~n43026 & n43031 ;
  assign n43033 = ~n43030 & ~n43032 ;
  assign n43034 = ~n42797 & n43033 ;
  assign n43035 = n42797 & ~n43033 ;
  assign n43036 = ~n43034 & ~n43035 ;
  assign n43037 = ~n42781 & ~n43036 ;
  assign n43038 = ~n42781 & ~n43037 ;
  assign n43039 = ~n43036 & ~n43037 ;
  assign n43040 = ~n43038 & ~n43039 ;
  assign n43041 = ~n42779 & ~n43040 ;
  assign n43042 = n42779 & ~n43039 ;
  assign n43043 = ~n43038 & n43042 ;
  assign n43044 = ~n43041 & ~n43043 ;
  assign n43312 = n43044 & x215 ;
  assign n43045 = ~n42767 & ~n42771 ;
  assign n43046 = ~n42517 & ~n42763 ;
  assign n43047 = ~n42514 & ~n43046 ;
  assign n43048 = ~n42531 & ~n42760 ;
  assign n43049 = ~x127 & n4531 ;
  assign n43050 = ~x125 & n4847 ;
  assign n43051 = ~x126 & n4526 ;
  assign n43052 = ~n43050 & ~n43051 ;
  assign n43053 = ~n43049 & n43052 ;
  assign n43054 = n4534 & n26932 ;
  assign n43055 = n43053 & ~n43054 ;
  assign n43056 = ~x26 & ~n43055 ;
  assign n43057 = ~x26 & ~n43056 ;
  assign n43058 = ~n43055 & ~n43056 ;
  assign n43059 = ~n43057 & ~n43058 ;
  assign n43060 = ~n43048 & ~n43059 ;
  assign n43061 = ~n43048 & ~n43060 ;
  assign n43062 = ~n43059 & ~n43060 ;
  assign n43063 = ~n43061 & ~n43062 ;
  assign n43064 = ~n42549 & ~n42756 ;
  assign n43065 = ~n42546 & ~n43064 ;
  assign n43066 = ~x124 & n5560 ;
  assign n43067 = ~x122 & n5943 ;
  assign n43068 = ~x123 & n5555 ;
  assign n43069 = ~n43067 & ~n43068 ;
  assign n43070 = ~n43066 & n43069 ;
  assign n43071 = n5563 & n24176 ;
  assign n43072 = n43070 & ~n43071 ;
  assign n43073 = ~x29 & ~n43072 ;
  assign n43074 = ~x29 & ~n43073 ;
  assign n43075 = ~n43072 & ~n43073 ;
  assign n43076 = ~n43074 & ~n43075 ;
  assign n43077 = ~n43065 & n43076 ;
  assign n43078 = n43065 & ~n43076 ;
  assign n43079 = ~n43077 & ~n43078 ;
  assign n43080 = ~x121 & n6725 ;
  assign n43081 = ~x119 & n7129 ;
  assign n43082 = ~x120 & n6720 ;
  assign n43083 = ~n43081 & ~n43082 ;
  assign n43084 = ~n43080 & n43083 ;
  assign n43085 = n6728 & n22229 ;
  assign n43086 = n43084 & ~n43085 ;
  assign n43087 = ~x32 & ~n43086 ;
  assign n43088 = ~x32 & ~n43087 ;
  assign n43089 = ~n43086 & ~n43087 ;
  assign n43090 = ~n43088 & ~n43089 ;
  assign n43091 = ~n42563 & ~n42753 ;
  assign n43092 = n43090 & n43091 ;
  assign n43093 = ~n43090 & ~n43091 ;
  assign n43094 = ~n43092 & ~n43093 ;
  assign n43095 = ~n42745 & ~n42749 ;
  assign n43096 = ~n42729 & ~n42743 ;
  assign n43097 = ~n42703 & ~n42706 ;
  assign n43098 = ~n42688 & ~n42699 ;
  assign n43099 = ~n42685 & ~n43098 ;
  assign n43100 = ~n42624 & ~n42638 ;
  assign n43101 = ~n42607 & ~n42621 ;
  assign n43102 = ~x87 & n27427 ;
  assign n43103 = ~x88 & ~n26217 ;
  assign n43104 = ~n43102 & ~n43103 ;
  assign n43105 = x23 & ~n43104 ;
  assign n43106 = ~x23 & n43104 ;
  assign n43107 = ~n43105 & ~n43106 ;
  assign n43108 = ~n42606 & n43107 ;
  assign n43109 = n42606 & ~n43107 ;
  assign n43110 = ~n43108 & ~n43109 ;
  assign n43111 = ~x91 & n24612 ;
  assign n43112 = ~x89 & n25390 ;
  assign n43113 = ~x90 & n24607 ;
  assign n43114 = ~n43112 & ~n43113 ;
  assign n43115 = ~n43111 & n43114 ;
  assign n43116 = n5507 & n24615 ;
  assign n43117 = n43115 & ~n43116 ;
  assign n43118 = ~x62 & ~n43117 ;
  assign n43119 = ~x62 & ~n43118 ;
  assign n43120 = ~n43117 & ~n43118 ;
  assign n43121 = ~n43119 & ~n43120 ;
  assign n43122 = n43110 & ~n43121 ;
  assign n43123 = n43110 & ~n43122 ;
  assign n43124 = ~n43121 & ~n43122 ;
  assign n43125 = ~n43123 & ~n43124 ;
  assign n43126 = ~n43101 & n43125 ;
  assign n43127 = n43101 & ~n43125 ;
  assign n43128 = ~n43126 & ~n43127 ;
  assign n43129 = ~x94 & n22325 ;
  assign n43130 = ~x92 & n23066 ;
  assign n43131 = ~x93 & n22320 ;
  assign n43132 = ~n43130 & ~n43131 ;
  assign n43133 = ~n43129 & n43132 ;
  assign n43134 = n6671 & n22328 ;
  assign n43135 = n43133 & ~n43134 ;
  assign n43136 = ~x59 & ~n43135 ;
  assign n43137 = ~x59 & ~n43136 ;
  assign n43138 = ~n43135 & ~n43136 ;
  assign n43139 = ~n43137 & ~n43138 ;
  assign n43140 = ~n43128 & ~n43139 ;
  assign n43141 = n43128 & n43139 ;
  assign n43142 = ~n43140 & ~n43141 ;
  assign n43143 = n43100 & ~n43142 ;
  assign n43144 = ~n43100 & n43142 ;
  assign n43145 = ~n43143 & ~n43144 ;
  assign n43146 = ~x97 & n20143 ;
  assign n43147 = ~x95 & n20854 ;
  assign n43148 = ~x96 & n20138 ;
  assign n43149 = ~n43147 & ~n43148 ;
  assign n43150 = ~n43146 & n43149 ;
  assign n43151 = n7949 & n20146 ;
  assign n43152 = n43150 & ~n43151 ;
  assign n43153 = ~x56 & ~n43152 ;
  assign n43154 = ~x56 & ~n43153 ;
  assign n43155 = ~n43152 & ~n43153 ;
  assign n43156 = ~n43154 & ~n43155 ;
  assign n43157 = ~n42644 & ~n42658 ;
  assign n43158 = ~n43156 & ~n43157 ;
  assign n43159 = n43156 & n43157 ;
  assign n43160 = ~n43158 & ~n43159 ;
  assign n43161 = n43145 & n43160 ;
  assign n43162 = ~n43145 & ~n43160 ;
  assign n43163 = ~n43161 & ~n43162 ;
  assign n43164 = ~x100 & n18025 ;
  assign n43165 = ~x98 & n18764 ;
  assign n43166 = ~x99 & n18020 ;
  assign n43167 = ~n43165 & ~n43166 ;
  assign n43168 = ~n43164 & n43167 ;
  assign n43169 = n9338 & n18028 ;
  assign n43170 = n43168 & ~n43169 ;
  assign n43171 = ~x53 & ~n43170 ;
  assign n43172 = ~x53 & ~n43171 ;
  assign n43173 = ~n43170 & ~n43171 ;
  assign n43174 = ~n43172 & ~n43173 ;
  assign n43175 = n43163 & ~n43174 ;
  assign n43176 = n43163 & ~n43175 ;
  assign n43177 = ~n43174 & ~n43175 ;
  assign n43178 = ~n43176 & ~n43177 ;
  assign n43179 = ~n42660 & ~n42663 ;
  assign n43180 = n43178 & n43179 ;
  assign n43181 = ~n43178 & ~n43179 ;
  assign n43182 = ~n43180 & ~n43181 ;
  assign n43183 = ~x103 & n16076 ;
  assign n43184 = ~x101 & n16756 ;
  assign n43185 = ~x102 & n16071 ;
  assign n43186 = ~n43184 & ~n43185 ;
  assign n43187 = ~n43183 & n43186 ;
  assign n43188 = n10833 & n16079 ;
  assign n43189 = n43187 & ~n43188 ;
  assign n43190 = ~x50 & ~n43189 ;
  assign n43191 = ~x50 & ~n43190 ;
  assign n43192 = ~n43189 & ~n43190 ;
  assign n43193 = ~n43191 & ~n43192 ;
  assign n43194 = n43182 & ~n43193 ;
  assign n43195 = n43182 & ~n43194 ;
  assign n43196 = ~n43193 & ~n43194 ;
  assign n43197 = ~n43195 & ~n43196 ;
  assign n43198 = ~n42666 & ~n42680 ;
  assign n43199 = n43197 & n43198 ;
  assign n43200 = ~n43197 & ~n43198 ;
  assign n43201 = ~n43199 & ~n43200 ;
  assign n43202 = ~x106 & n14233 ;
  assign n43203 = ~x104 & n14876 ;
  assign n43204 = ~x105 & n14228 ;
  assign n43205 = ~n43203 & ~n43204 ;
  assign n43206 = ~n43202 & n43205 ;
  assign n43207 = n12447 & n14236 ;
  assign n43208 = n43206 & ~n43207 ;
  assign n43209 = ~x47 & ~n43208 ;
  assign n43210 = ~x47 & ~n43209 ;
  assign n43211 = ~n43208 & ~n43209 ;
  assign n43212 = ~n43210 & ~n43211 ;
  assign n43213 = n43201 & ~n43212 ;
  assign n43214 = n43201 & ~n43213 ;
  assign n43215 = ~n43212 & ~n43213 ;
  assign n43216 = ~n43214 & ~n43215 ;
  assign n43217 = ~n43099 & n43216 ;
  assign n43218 = n43099 & ~n43216 ;
  assign n43219 = ~n43217 & ~n43218 ;
  assign n43220 = ~x109 & n12506 ;
  assign n43221 = ~x107 & n13131 ;
  assign n43222 = ~x108 & n12501 ;
  assign n43223 = ~n43221 & ~n43222 ;
  assign n43224 = ~n43220 & n43223 ;
  assign n43225 = n12509 & n14177 ;
  assign n43226 = n43224 & ~n43225 ;
  assign n43227 = ~x44 & ~n43226 ;
  assign n43228 = ~x44 & ~n43227 ;
  assign n43229 = ~n43226 & ~n43227 ;
  assign n43230 = ~n43228 & ~n43229 ;
  assign n43231 = ~n43219 & ~n43230 ;
  assign n43232 = n43219 & n43230 ;
  assign n43233 = ~n43231 & ~n43232 ;
  assign n43234 = n43097 & ~n43233 ;
  assign n43235 = ~n43097 & n43233 ;
  assign n43236 = ~n43234 & ~n43235 ;
  assign n43237 = ~x112 & n10905 ;
  assign n43238 = ~x110 & n11466 ;
  assign n43239 = ~x111 & n10900 ;
  assign n43240 = ~n43238 & ~n43239 ;
  assign n43241 = ~n43237 & n43240 ;
  assign n43242 = n10908 & n15744 ;
  assign n43243 = n43241 & ~n43242 ;
  assign n43244 = ~x41 & ~n43243 ;
  assign n43245 = ~x41 & ~n43244 ;
  assign n43246 = ~n43243 & ~n43244 ;
  assign n43247 = ~n43245 & ~n43246 ;
  assign n43248 = n43236 & ~n43247 ;
  assign n43249 = n43236 & ~n43248 ;
  assign n43250 = ~n43247 & ~n43248 ;
  assign n43251 = ~n43249 & ~n43250 ;
  assign n43252 = ~n42709 & ~n42723 ;
  assign n43253 = n43251 & n43252 ;
  assign n43254 = ~n43251 & ~n43252 ;
  assign n43255 = ~n43253 & ~n43254 ;
  assign n43256 = ~x115 & n9433 ;
  assign n43257 = ~x113 & n9915 ;
  assign n43258 = ~x114 & n9428 ;
  assign n43259 = ~n43257 & ~n43258 ;
  assign n43260 = ~n43256 & n43259 ;
  assign n43261 = n9436 & n17683 ;
  assign n43262 = n43260 & ~n43261 ;
  assign n43263 = ~x38 & ~n43262 ;
  assign n43264 = ~x38 & ~n43263 ;
  assign n43265 = ~n43262 & ~n43263 ;
  assign n43266 = ~n43264 & ~n43265 ;
  assign n43267 = n43255 & ~n43266 ;
  assign n43268 = ~n43255 & n43266 ;
  assign n43269 = ~n43096 & ~n43268 ;
  assign n43270 = ~n43267 & n43269 ;
  assign n43271 = ~n43096 & ~n43270 ;
  assign n43272 = ~n43267 & ~n43270 ;
  assign n43273 = ~n43268 & n43272 ;
  assign n43274 = ~n43271 & ~n43273 ;
  assign n43275 = ~x118 & n8006 ;
  assign n43276 = ~x116 & n8474 ;
  assign n43277 = ~x117 & n8001 ;
  assign n43278 = ~n43276 & ~n43277 ;
  assign n43279 = ~n43275 & n43278 ;
  assign n43280 = n8009 & n19736 ;
  assign n43281 = n43279 & ~n43280 ;
  assign n43282 = ~x35 & ~n43281 ;
  assign n43283 = ~x35 & ~n43282 ;
  assign n43284 = ~n43281 & ~n43282 ;
  assign n43285 = ~n43283 & ~n43284 ;
  assign n43286 = n43274 & n43285 ;
  assign n43287 = ~n43274 & ~n43285 ;
  assign n43288 = ~n43286 & ~n43287 ;
  assign n43289 = ~n43095 & n43288 ;
  assign n43290 = n43095 & ~n43288 ;
  assign n43291 = ~n43289 & ~n43290 ;
  assign n43292 = n43094 & n43291 ;
  assign n43293 = ~n43094 & ~n43291 ;
  assign n43294 = ~n43079 & ~n43293 ;
  assign n43295 = ~n43292 & n43294 ;
  assign n43296 = ~n43079 & ~n43295 ;
  assign n43297 = ~n43293 & ~n43295 ;
  assign n43298 = ~n43292 & n43297 ;
  assign n43299 = ~n43296 & ~n43298 ;
  assign n43300 = ~n43063 & n43299 ;
  assign n43301 = n43063 & ~n43299 ;
  assign n43302 = ~n43300 & ~n43301 ;
  assign n43303 = ~n43047 & ~n43302 ;
  assign n43304 = ~n43047 & ~n43303 ;
  assign n43305 = ~n43302 & ~n43303 ;
  assign n43306 = ~n43304 & ~n43305 ;
  assign n43307 = ~n43045 & ~n43306 ;
  assign n43308 = n43045 & ~n43305 ;
  assign n43309 = ~n43304 & n43308 ;
  assign n43310 = ~n43307 & ~n43309 ;
  assign n43313 = ~n43310 & ~x215 ;
  assign n43314 = ~n43312 & ~n43313 ;
  assign n43315 = ~n43037 & ~n43041 ;
  assign n43316 = ~n42797 & ~n43033 ;
  assign n43317 = ~n42794 & ~n43316 ;
  assign n43318 = x125 & n5560 ;
  assign n43319 = x123 & n5943 ;
  assign n43320 = x124 & n5555 ;
  assign n43321 = ~n43319 & ~n43320 ;
  assign n43322 = ~n43318 & n43321 ;
  assign n43323 = n5563 & n24935 ;
  assign n43324 = n43322 & ~n43323 ;
  assign n43325 = x29 & ~n43324 ;
  assign n43326 = x29 & ~n43325 ;
  assign n43327 = ~n43324 & ~n43325 ;
  assign n43328 = ~n43326 & ~n43327 ;
  assign n43329 = ~n42827 & ~n43026 ;
  assign n43330 = ~n43328 & ~n43329 ;
  assign n43331 = ~n43328 & ~n43330 ;
  assign n43332 = ~n43329 & ~n43330 ;
  assign n43333 = ~n43331 & ~n43332 ;
  assign n43334 = ~n43021 & ~n43023 ;
  assign n43335 = x122 & n6725 ;
  assign n43336 = x120 & n7129 ;
  assign n43337 = x121 & n6720 ;
  assign n43338 = ~n43336 & ~n43337 ;
  assign n43339 = ~n43335 & n43338 ;
  assign n43340 = ~n6728 & n43339 ;
  assign n43341 = ~n22622 & n43339 ;
  assign n43342 = ~n43340 & ~n43341 ;
  assign n43343 = x32 & ~n43342 ;
  assign n43344 = ~x32 & n43342 ;
  assign n43345 = ~n43343 & ~n43344 ;
  assign n43346 = ~n43334 & ~n43345 ;
  assign n43347 = n43334 & n43345 ;
  assign n43348 = ~n43346 & ~n43347 ;
  assign n43349 = ~n42928 & ~n42934 ;
  assign n43350 = x104 & n16076 ;
  assign n43351 = x102 & n16756 ;
  assign n43352 = x103 & n16071 ;
  assign n43353 = ~n43351 & ~n43352 ;
  assign n43354 = ~n43350 & n43353 ;
  assign n43355 = n11116 & n16079 ;
  assign n43356 = n43354 & ~n43355 ;
  assign n43357 = x50 & ~n43356 ;
  assign n43358 = x50 & ~n43357 ;
  assign n43359 = ~n43356 & ~n43357 ;
  assign n43360 = ~n43358 & ~n43359 ;
  assign n43361 = ~n42909 & ~n42915 ;
  assign n43362 = ~n42835 & ~n42859 ;
  assign n43363 = ~n42856 & ~n43362 ;
  assign n43364 = x88 & n27024 ;
  assign n43365 = x89 & ~n26217 ;
  assign n43366 = ~n43364 & ~n43365 ;
  assign n43367 = ~n42839 & ~n42842 ;
  assign n43368 = ~n43366 & n43367 ;
  assign n43369 = n43366 & ~n43367 ;
  assign n43370 = ~n43368 & ~n43369 ;
  assign n43371 = x92 & n24612 ;
  assign n43372 = x90 & n25390 ;
  assign n43373 = x91 & n24607 ;
  assign n43374 = ~n43372 & ~n43373 ;
  assign n43375 = ~n43371 & n43374 ;
  assign n43376 = ~n24615 & n43375 ;
  assign n43377 = ~n5710 & n43375 ;
  assign n43378 = ~n43376 & ~n43377 ;
  assign n43379 = x62 & ~n43378 ;
  assign n43380 = ~x62 & n43378 ;
  assign n43381 = ~n43379 & ~n43380 ;
  assign n43382 = n43370 & ~n43381 ;
  assign n43383 = ~n43370 & n43381 ;
  assign n43384 = ~n43382 & ~n43383 ;
  assign n43385 = ~n43363 & n43384 ;
  assign n43386 = n43363 & ~n43384 ;
  assign n43387 = ~n43385 & ~n43386 ;
  assign n43388 = x95 & n22325 ;
  assign n43389 = x93 & n23066 ;
  assign n43390 = x94 & n22320 ;
  assign n43391 = ~n43389 & ~n43390 ;
  assign n43392 = ~n43388 & n43391 ;
  assign n43393 = n6894 & n22328 ;
  assign n43394 = n43392 & ~n43393 ;
  assign n43395 = x59 & ~n43394 ;
  assign n43396 = x59 & ~n43395 ;
  assign n43397 = ~n43394 & ~n43395 ;
  assign n43398 = ~n43396 & ~n43397 ;
  assign n43399 = n43387 & ~n43398 ;
  assign n43400 = n43387 & ~n43399 ;
  assign n43401 = ~n43398 & ~n43399 ;
  assign n43402 = ~n43400 & ~n43401 ;
  assign n43403 = ~n42874 & ~n42878 ;
  assign n43404 = n43402 & n43403 ;
  assign n43405 = ~n43402 & ~n43403 ;
  assign n43406 = ~n43404 & ~n43405 ;
  assign n43407 = x98 & n20143 ;
  assign n43408 = x96 & n20854 ;
  assign n43409 = x97 & n20138 ;
  assign n43410 = ~n43408 & ~n43409 ;
  assign n43411 = ~n43407 & n43410 ;
  assign n43412 = n8196 & n20146 ;
  assign n43413 = n43411 & ~n43412 ;
  assign n43414 = x56 & ~n43413 ;
  assign n43415 = x56 & ~n43414 ;
  assign n43416 = ~n43413 & ~n43414 ;
  assign n43417 = ~n43415 & ~n43416 ;
  assign n43418 = n43406 & ~n43417 ;
  assign n43419 = n43406 & ~n43418 ;
  assign n43420 = ~n43417 & ~n43418 ;
  assign n43421 = ~n43419 & ~n43420 ;
  assign n43422 = ~n42892 & ~n42895 ;
  assign n43423 = n43421 & n43422 ;
  assign n43424 = ~n43421 & ~n43422 ;
  assign n43425 = ~n43423 & ~n43424 ;
  assign n43426 = x101 & n18025 ;
  assign n43427 = x99 & n18764 ;
  assign n43428 = x100 & n18020 ;
  assign n43429 = ~n43427 & ~n43428 ;
  assign n43430 = ~n43426 & n43429 ;
  assign n43431 = n9601 & n18028 ;
  assign n43432 = n43430 & ~n43431 ;
  assign n43433 = x53 & ~n43432 ;
  assign n43434 = x53 & ~n43433 ;
  assign n43435 = ~n43432 & ~n43433 ;
  assign n43436 = ~n43434 & ~n43435 ;
  assign n43437 = ~n43425 & n43436 ;
  assign n43438 = n43425 & ~n43436 ;
  assign n43439 = ~n43437 & ~n43438 ;
  assign n43440 = ~n43361 & n43439 ;
  assign n43441 = ~n43361 & ~n43440 ;
  assign n43442 = n43439 & ~n43440 ;
  assign n43443 = ~n43441 & ~n43442 ;
  assign n43444 = ~n43360 & ~n43443 ;
  assign n43445 = n43360 & ~n43442 ;
  assign n43446 = ~n43441 & n43445 ;
  assign n43447 = ~n43444 & ~n43446 ;
  assign n43448 = ~n43349 & n43447 ;
  assign n43449 = n43349 & ~n43447 ;
  assign n43450 = ~n43448 & ~n43449 ;
  assign n43451 = x107 & n14233 ;
  assign n43452 = x105 & n14876 ;
  assign n43453 = x106 & n14228 ;
  assign n43454 = ~n43452 & ~n43453 ;
  assign n43455 = ~n43451 & n43454 ;
  assign n43456 = n12749 & n14236 ;
  assign n43457 = n43455 & ~n43456 ;
  assign n43458 = x47 & ~n43457 ;
  assign n43459 = x47 & ~n43458 ;
  assign n43460 = ~n43457 & ~n43458 ;
  assign n43461 = ~n43459 & ~n43460 ;
  assign n43462 = n43450 & ~n43461 ;
  assign n43463 = n43450 & ~n43462 ;
  assign n43464 = ~n43461 & ~n43462 ;
  assign n43465 = ~n43463 & ~n43464 ;
  assign n43466 = ~n42833 & ~n42950 ;
  assign n43467 = ~n42947 & ~n43466 ;
  assign n43468 = n43465 & n43467 ;
  assign n43469 = ~n43465 & ~n43467 ;
  assign n43470 = ~n43468 & ~n43469 ;
  assign n43471 = x110 & n12506 ;
  assign n43472 = x108 & n13131 ;
  assign n43473 = x109 & n12501 ;
  assign n43474 = ~n43472 & ~n43473 ;
  assign n43475 = ~n43471 & n43474 ;
  assign n43476 = n12509 & n14497 ;
  assign n43477 = n43475 & ~n43476 ;
  assign n43478 = x44 & ~n43477 ;
  assign n43479 = x44 & ~n43478 ;
  assign n43480 = ~n43477 & ~n43478 ;
  assign n43481 = ~n43479 & ~n43480 ;
  assign n43482 = n43470 & ~n43481 ;
  assign n43483 = n43470 & ~n43482 ;
  assign n43484 = ~n43481 & ~n43482 ;
  assign n43485 = ~n43483 & ~n43484 ;
  assign n43486 = ~n42965 & ~n42969 ;
  assign n43487 = n43485 & n43486 ;
  assign n43488 = ~n43485 & ~n43486 ;
  assign n43489 = ~n43487 & ~n43488 ;
  assign n43490 = x113 & n10905 ;
  assign n43491 = x111 & n11466 ;
  assign n43492 = x112 & n10900 ;
  assign n43493 = ~n43491 & ~n43492 ;
  assign n43494 = ~n43490 & n43493 ;
  assign n43495 = n10908 & n16361 ;
  assign n43496 = n43494 & ~n43495 ;
  assign n43497 = x41 & ~n43496 ;
  assign n43498 = x41 & ~n43497 ;
  assign n43499 = ~n43496 & ~n43497 ;
  assign n43500 = ~n43498 & ~n43499 ;
  assign n43501 = n43489 & ~n43500 ;
  assign n43502 = n43489 & ~n43501 ;
  assign n43503 = ~n43500 & ~n43501 ;
  assign n43504 = ~n43502 & ~n43503 ;
  assign n43505 = ~n42982 & ~n42988 ;
  assign n43506 = n43504 & n43505 ;
  assign n43507 = ~n43504 & ~n43505 ;
  assign n43508 = ~n43506 & ~n43507 ;
  assign n43509 = x116 & n9433 ;
  assign n43510 = x114 & n9915 ;
  assign n43511 = x115 & n9428 ;
  assign n43512 = ~n43510 & ~n43511 ;
  assign n43513 = ~n43509 & n43512 ;
  assign n43514 = n9436 & n18336 ;
  assign n43515 = n43513 & ~n43514 ;
  assign n43516 = x38 & ~n43515 ;
  assign n43517 = x38 & ~n43516 ;
  assign n43518 = ~n43515 & ~n43516 ;
  assign n43519 = ~n43517 & ~n43518 ;
  assign n43520 = n43508 & ~n43519 ;
  assign n43521 = n43508 & ~n43520 ;
  assign n43522 = ~n43519 & ~n43520 ;
  assign n43523 = ~n43521 & ~n43522 ;
  assign n43524 = ~n43006 & n43523 ;
  assign n43525 = n43006 & ~n43523 ;
  assign n43526 = ~n43524 & ~n43525 ;
  assign n43527 = x119 & n8006 ;
  assign n43528 = x117 & n8474 ;
  assign n43529 = x118 & n8001 ;
  assign n43530 = ~n43528 & ~n43529 ;
  assign n43531 = ~n43527 & n43530 ;
  assign n43532 = n8009 & n20423 ;
  assign n43533 = n43531 & ~n43532 ;
  assign n43534 = x35 & ~n43533 ;
  assign n43535 = x35 & ~n43534 ;
  assign n43536 = ~n43533 & ~n43534 ;
  assign n43537 = ~n43535 & ~n43536 ;
  assign n43538 = ~n43526 & ~n43537 ;
  assign n43539 = n43526 & n43537 ;
  assign n43540 = ~n43538 & ~n43539 ;
  assign n43541 = n43348 & n43540 ;
  assign n43542 = ~n43348 & ~n43540 ;
  assign n43543 = ~n43541 & ~n43542 ;
  assign n43544 = ~n43333 & n43543 ;
  assign n43545 = ~n43333 & ~n43544 ;
  assign n43546 = n43543 & ~n43544 ;
  assign n43547 = ~n43545 & ~n43546 ;
  assign n43548 = ~n42799 & ~n42810 ;
  assign n43549 = ~n43029 & ~n43548 ;
  assign n43550 = x126 & n4847 ;
  assign n43551 = x127 & n4526 ;
  assign n43552 = ~n43550 & ~n43551 ;
  assign n43553 = ~n4534 & n43552 ;
  assign n43554 = n26965 & n43552 ;
  assign n43555 = ~n43553 & ~n43554 ;
  assign n43556 = x26 & ~n43555 ;
  assign n43557 = ~x26 & n43555 ;
  assign n43558 = ~n43556 & ~n43557 ;
  assign n43559 = ~n43549 & ~n43558 ;
  assign n43560 = ~n43549 & ~n43559 ;
  assign n43561 = ~n43558 & ~n43559 ;
  assign n43562 = ~n43560 & ~n43561 ;
  assign n43563 = ~n43547 & ~n43562 ;
  assign n43564 = n43547 & ~n43561 ;
  assign n43565 = ~n43560 & n43564 ;
  assign n43566 = ~n43563 & ~n43565 ;
  assign n43567 = ~n43317 & n43566 ;
  assign n43568 = ~n43317 & ~n43567 ;
  assign n43569 = n43566 & ~n43567 ;
  assign n43570 = ~n43568 & ~n43569 ;
  assign n43571 = ~n43315 & ~n43570 ;
  assign n43572 = n43315 & ~n43569 ;
  assign n43573 = ~n43568 & n43572 ;
  assign n43574 = ~n43571 & ~n43573 ;
  assign n43836 = n43574 & x216 ;
  assign n43575 = ~n43303 & ~n43307 ;
  assign n43576 = ~n43063 & ~n43299 ;
  assign n43577 = ~n43060 & ~n43576 ;
  assign n43578 = ~x125 & n5560 ;
  assign n43579 = ~x123 & n5943 ;
  assign n43580 = ~x124 & n5555 ;
  assign n43581 = ~n43579 & ~n43580 ;
  assign n43582 = ~n43578 & n43581 ;
  assign n43583 = n5563 & n25330 ;
  assign n43584 = n43582 & ~n43583 ;
  assign n43585 = ~x29 & ~n43584 ;
  assign n43586 = ~x29 & ~n43585 ;
  assign n43587 = ~n43584 & ~n43585 ;
  assign n43588 = ~n43586 & ~n43587 ;
  assign n43589 = ~n43093 & ~n43292 ;
  assign n43590 = ~n43588 & ~n43589 ;
  assign n43591 = ~n43588 & ~n43590 ;
  assign n43592 = ~n43589 & ~n43590 ;
  assign n43593 = ~n43591 & ~n43592 ;
  assign n43594 = ~n43287 & ~n43289 ;
  assign n43595 = ~x122 & n6725 ;
  assign n43596 = ~x120 & n7129 ;
  assign n43597 = ~x121 & n6720 ;
  assign n43598 = ~n43596 & ~n43597 ;
  assign n43599 = ~n43595 & n43598 ;
  assign n43600 = ~n6728 & n43599 ;
  assign n43601 = ~n22998 & n43599 ;
  assign n43602 = ~n43600 & ~n43601 ;
  assign n43603 = ~x32 & ~n43602 ;
  assign n43604 = x32 & n43602 ;
  assign n43605 = ~n43603 & ~n43604 ;
  assign n43606 = ~n43594 & ~n43605 ;
  assign n43607 = n43594 & n43605 ;
  assign n43608 = ~n43606 & ~n43607 ;
  assign n43609 = ~n43194 & ~n43200 ;
  assign n43610 = ~x104 & n16076 ;
  assign n43611 = ~x102 & n16756 ;
  assign n43612 = ~x103 & n16071 ;
  assign n43613 = ~n43611 & ~n43612 ;
  assign n43614 = ~n43610 & n43613 ;
  assign n43615 = n11380 & n16079 ;
  assign n43616 = n43614 & ~n43615 ;
  assign n43617 = ~x50 & ~n43616 ;
  assign n43618 = ~x50 & ~n43617 ;
  assign n43619 = ~n43616 & ~n43617 ;
  assign n43620 = ~n43618 & ~n43619 ;
  assign n43621 = ~n43175 & ~n43181 ;
  assign n43622 = ~n43101 & ~n43125 ;
  assign n43623 = ~n43122 & ~n43622 ;
  assign n43624 = ~x88 & n27427 ;
  assign n43625 = ~x89 & ~n26217 ;
  assign n43626 = ~n43624 & ~n43625 ;
  assign n43627 = ~n43105 & ~n43108 ;
  assign n43628 = ~n43626 & n43627 ;
  assign n43629 = n43626 & ~n43627 ;
  assign n43630 = ~n43628 & ~n43629 ;
  assign n43631 = ~x92 & n24612 ;
  assign n43632 = ~x90 & n25390 ;
  assign n43633 = ~x91 & n24607 ;
  assign n43634 = ~n43632 & ~n43633 ;
  assign n43635 = ~n43631 & n43634 ;
  assign n43636 = ~n24615 & n43635 ;
  assign n43637 = ~n5896 & n43635 ;
  assign n43638 = ~n43636 & ~n43637 ;
  assign n43639 = ~x62 & ~n43638 ;
  assign n43640 = x62 & n43638 ;
  assign n43641 = ~n43639 & ~n43640 ;
  assign n43642 = n43630 & ~n43641 ;
  assign n43643 = ~n43630 & n43641 ;
  assign n43644 = ~n43642 & ~n43643 ;
  assign n43645 = ~n43623 & n43644 ;
  assign n43646 = n43623 & ~n43644 ;
  assign n43647 = ~n43645 & ~n43646 ;
  assign n43648 = ~x95 & n22325 ;
  assign n43649 = ~x93 & n23066 ;
  assign n43650 = ~x94 & n22320 ;
  assign n43651 = ~n43649 & ~n43650 ;
  assign n43652 = ~n43648 & n43651 ;
  assign n43653 = n7100 & n22328 ;
  assign n43654 = n43652 & ~n43653 ;
  assign n43655 = ~x59 & ~n43654 ;
  assign n43656 = ~x59 & ~n43655 ;
  assign n43657 = ~n43654 & ~n43655 ;
  assign n43658 = ~n43656 & ~n43657 ;
  assign n43659 = n43647 & ~n43658 ;
  assign n43660 = n43647 & ~n43659 ;
  assign n43661 = ~n43658 & ~n43659 ;
  assign n43662 = ~n43660 & ~n43661 ;
  assign n43663 = ~n43140 & ~n43144 ;
  assign n43664 = n43662 & n43663 ;
  assign n43665 = ~n43662 & ~n43663 ;
  assign n43666 = ~n43664 & ~n43665 ;
  assign n43667 = ~x98 & n20143 ;
  assign n43668 = ~x96 & n20854 ;
  assign n43669 = ~x97 & n20138 ;
  assign n43670 = ~n43668 & ~n43669 ;
  assign n43671 = ~n43667 & n43670 ;
  assign n43672 = n8426 & n20146 ;
  assign n43673 = n43671 & ~n43672 ;
  assign n43674 = ~x56 & ~n43673 ;
  assign n43675 = ~x56 & ~n43674 ;
  assign n43676 = ~n43673 & ~n43674 ;
  assign n43677 = ~n43675 & ~n43676 ;
  assign n43678 = n43666 & ~n43677 ;
  assign n43679 = n43666 & ~n43678 ;
  assign n43680 = ~n43677 & ~n43678 ;
  assign n43681 = ~n43679 & ~n43680 ;
  assign n43682 = ~n43158 & ~n43161 ;
  assign n43683 = n43681 & n43682 ;
  assign n43684 = ~n43681 & ~n43682 ;
  assign n43685 = ~n43683 & ~n43684 ;
  assign n43686 = ~x101 & n18025 ;
  assign n43687 = ~x99 & n18764 ;
  assign n43688 = ~x100 & n18020 ;
  assign n43689 = ~n43687 & ~n43688 ;
  assign n43690 = ~n43686 & n43689 ;
  assign n43691 = n9844 & n18028 ;
  assign n43692 = n43690 & ~n43691 ;
  assign n43693 = ~x53 & ~n43692 ;
  assign n43694 = ~x53 & ~n43693 ;
  assign n43695 = ~n43692 & ~n43693 ;
  assign n43696 = ~n43694 & ~n43695 ;
  assign n43697 = ~n43685 & n43696 ;
  assign n43698 = n43685 & ~n43696 ;
  assign n43699 = ~n43697 & ~n43698 ;
  assign n43700 = ~n43621 & n43699 ;
  assign n43701 = ~n43621 & ~n43700 ;
  assign n43702 = n43699 & ~n43700 ;
  assign n43703 = ~n43701 & ~n43702 ;
  assign n43704 = ~n43620 & ~n43703 ;
  assign n43705 = n43620 & ~n43702 ;
  assign n43706 = ~n43701 & n43705 ;
  assign n43707 = ~n43704 & ~n43706 ;
  assign n43708 = ~n43609 & n43707 ;
  assign n43709 = n43609 & ~n43707 ;
  assign n43710 = ~n43708 & ~n43709 ;
  assign n43711 = ~x107 & n14233 ;
  assign n43712 = ~x105 & n14876 ;
  assign n43713 = ~x106 & n14228 ;
  assign n43714 = ~n43712 & ~n43713 ;
  assign n43715 = ~n43711 & n43714 ;
  assign n43716 = n13034 & n14236 ;
  assign n43717 = n43715 & ~n43716 ;
  assign n43718 = ~x47 & ~n43717 ;
  assign n43719 = ~x47 & ~n43718 ;
  assign n43720 = ~n43717 & ~n43718 ;
  assign n43721 = ~n43719 & ~n43720 ;
  assign n43722 = n43710 & ~n43721 ;
  assign n43723 = n43710 & ~n43722 ;
  assign n43724 = ~n43721 & ~n43722 ;
  assign n43725 = ~n43723 & ~n43724 ;
  assign n43726 = ~n43099 & ~n43216 ;
  assign n43727 = ~n43213 & ~n43726 ;
  assign n43728 = n43725 & n43727 ;
  assign n43729 = ~n43725 & ~n43727 ;
  assign n43730 = ~n43728 & ~n43729 ;
  assign n43731 = ~x110 & n12506 ;
  assign n43732 = ~x108 & n13131 ;
  assign n43733 = ~x109 & n12501 ;
  assign n43734 = ~n43732 & ~n43733 ;
  assign n43735 = ~n43731 & n43734 ;
  assign n43736 = n12509 & n14802 ;
  assign n43737 = n43735 & ~n43736 ;
  assign n43738 = ~x44 & ~n43737 ;
  assign n43739 = ~x44 & ~n43738 ;
  assign n43740 = ~n43737 & ~n43738 ;
  assign n43741 = ~n43739 & ~n43740 ;
  assign n43742 = n43730 & ~n43741 ;
  assign n43743 = n43730 & ~n43742 ;
  assign n43744 = ~n43741 & ~n43742 ;
  assign n43745 = ~n43743 & ~n43744 ;
  assign n43746 = ~n43231 & ~n43235 ;
  assign n43747 = n43745 & n43746 ;
  assign n43748 = ~n43745 & ~n43746 ;
  assign n43749 = ~n43747 & ~n43748 ;
  assign n43750 = ~x113 & n10905 ;
  assign n43751 = ~x111 & n11466 ;
  assign n43752 = ~x112 & n10900 ;
  assign n43753 = ~n43751 & ~n43752 ;
  assign n43754 = ~n43750 & n43753 ;
  assign n43755 = n10908 & n16684 ;
  assign n43756 = n43754 & ~n43755 ;
  assign n43757 = ~x41 & ~n43756 ;
  assign n43758 = ~x41 & ~n43757 ;
  assign n43759 = ~n43756 & ~n43757 ;
  assign n43760 = ~n43758 & ~n43759 ;
  assign n43761 = n43749 & ~n43760 ;
  assign n43762 = n43749 & ~n43761 ;
  assign n43763 = ~n43760 & ~n43761 ;
  assign n43764 = ~n43762 & ~n43763 ;
  assign n43765 = ~n43248 & ~n43254 ;
  assign n43766 = n43764 & n43765 ;
  assign n43767 = ~n43764 & ~n43765 ;
  assign n43768 = ~n43766 & ~n43767 ;
  assign n43769 = ~x116 & n9433 ;
  assign n43770 = ~x114 & n9915 ;
  assign n43771 = ~x115 & n9428 ;
  assign n43772 = ~n43770 & ~n43771 ;
  assign n43773 = ~n43769 & n43772 ;
  assign n43774 = n9436 & n18678 ;
  assign n43775 = n43773 & ~n43774 ;
  assign n43776 = ~x38 & ~n43775 ;
  assign n43777 = ~x38 & ~n43776 ;
  assign n43778 = ~n43775 & ~n43776 ;
  assign n43779 = ~n43777 & ~n43778 ;
  assign n43780 = n43768 & ~n43779 ;
  assign n43781 = n43768 & ~n43780 ;
  assign n43782 = ~n43779 & ~n43780 ;
  assign n43783 = ~n43781 & ~n43782 ;
  assign n43784 = ~n43272 & n43783 ;
  assign n43785 = n43272 & ~n43783 ;
  assign n43786 = ~n43784 & ~n43785 ;
  assign n43787 = ~x119 & n8006 ;
  assign n43788 = ~x117 & n8474 ;
  assign n43789 = ~x118 & n8001 ;
  assign n43790 = ~n43788 & ~n43789 ;
  assign n43791 = ~n43787 & n43790 ;
  assign n43792 = n8009 & n20778 ;
  assign n43793 = n43791 & ~n43792 ;
  assign n43794 = ~x35 & ~n43793 ;
  assign n43795 = ~x35 & ~n43794 ;
  assign n43796 = ~n43793 & ~n43794 ;
  assign n43797 = ~n43795 & ~n43796 ;
  assign n43798 = ~n43786 & ~n43797 ;
  assign n43799 = n43786 & n43797 ;
  assign n43800 = ~n43798 & ~n43799 ;
  assign n43801 = n43608 & n43800 ;
  assign n43802 = ~n43608 & ~n43800 ;
  assign n43803 = ~n43801 & ~n43802 ;
  assign n43804 = ~n43593 & n43803 ;
  assign n43805 = ~n43593 & ~n43804 ;
  assign n43806 = n43803 & ~n43804 ;
  assign n43807 = ~n43805 & ~n43806 ;
  assign n43808 = ~n43065 & ~n43076 ;
  assign n43809 = ~n43295 & ~n43808 ;
  assign n43810 = ~x126 & n4847 ;
  assign n43811 = ~x127 & n4526 ;
  assign n43812 = ~n43810 & ~n43811 ;
  assign n43813 = ~n4534 & n43812 ;
  assign n43814 = n27368 & n43812 ;
  assign n43815 = ~n43813 & ~n43814 ;
  assign n43816 = ~x26 & ~n43815 ;
  assign n43817 = x26 & n43815 ;
  assign n43818 = ~n43816 & ~n43817 ;
  assign n43819 = ~n43809 & ~n43818 ;
  assign n43820 = ~n43809 & ~n43819 ;
  assign n43821 = ~n43818 & ~n43819 ;
  assign n43822 = ~n43820 & ~n43821 ;
  assign n43823 = ~n43807 & ~n43822 ;
  assign n43824 = n43807 & ~n43821 ;
  assign n43825 = ~n43820 & n43824 ;
  assign n43826 = ~n43823 & ~n43825 ;
  assign n43827 = ~n43577 & n43826 ;
  assign n43828 = ~n43577 & ~n43827 ;
  assign n43829 = n43826 & ~n43827 ;
  assign n43830 = ~n43828 & ~n43829 ;
  assign n43831 = ~n43575 & ~n43830 ;
  assign n43832 = n43575 & ~n43829 ;
  assign n43833 = ~n43828 & n43832 ;
  assign n43834 = ~n43831 & ~n43833 ;
  assign n43837 = ~n43834 & ~x216 ;
  assign n43838 = ~n43836 & ~n43837 ;
  assign n43839 = ~n43567 & ~n43571 ;
  assign n43840 = ~n43559 & ~n43563 ;
  assign n43841 = ~n43330 & ~n43544 ;
  assign n43842 = x127 & n4847 ;
  assign n43843 = n4534 & n26962 ;
  assign n43844 = ~n43842 & ~n43843 ;
  assign n43845 = x26 & ~n43844 ;
  assign n43846 = x26 & ~n43845 ;
  assign n43847 = ~n43844 & ~n43845 ;
  assign n43848 = ~n43846 & ~n43847 ;
  assign n43849 = ~n43841 & ~n43848 ;
  assign n43850 = ~n43841 & ~n43849 ;
  assign n43851 = ~n43848 & ~n43849 ;
  assign n43852 = ~n43850 & ~n43851 ;
  assign n43853 = x126 & n5560 ;
  assign n43854 = x124 & n5943 ;
  assign n43855 = x125 & n5555 ;
  assign n43856 = ~n43854 & ~n43855 ;
  assign n43857 = ~n43853 & n43856 ;
  assign n43858 = n5563 & n25735 ;
  assign n43859 = n43857 & ~n43858 ;
  assign n43860 = x29 & ~n43859 ;
  assign n43861 = x29 & ~n43860 ;
  assign n43862 = ~n43859 & ~n43860 ;
  assign n43863 = ~n43861 & ~n43862 ;
  assign n43864 = ~n43346 & ~n43541 ;
  assign n43865 = n43863 & n43864 ;
  assign n43866 = ~n43863 & ~n43864 ;
  assign n43867 = ~n43865 & ~n43866 ;
  assign n43868 = x123 & n6725 ;
  assign n43869 = x121 & n7129 ;
  assign n43870 = x122 & n6720 ;
  assign n43871 = ~n43869 & ~n43870 ;
  assign n43872 = ~n43868 & n43871 ;
  assign n43873 = n6728 & n23382 ;
  assign n43874 = n43872 & ~n43873 ;
  assign n43875 = x32 & ~n43874 ;
  assign n43876 = x32 & ~n43875 ;
  assign n43877 = ~n43874 & ~n43875 ;
  assign n43878 = ~n43876 & ~n43877 ;
  assign n43879 = ~n43006 & ~n43523 ;
  assign n43880 = ~n43538 & ~n43879 ;
  assign n43881 = n43878 & n43880 ;
  assign n43882 = ~n43878 & ~n43880 ;
  assign n43883 = ~n43881 & ~n43882 ;
  assign n43884 = x120 & n8006 ;
  assign n43885 = x118 & n8474 ;
  assign n43886 = x119 & n8001 ;
  assign n43887 = ~n43885 & ~n43886 ;
  assign n43888 = ~n43884 & n43887 ;
  assign n43889 = n8009 & n21143 ;
  assign n43890 = n43888 & ~n43889 ;
  assign n43891 = x35 & ~n43890 ;
  assign n43892 = x35 & ~n43891 ;
  assign n43893 = ~n43890 & ~n43891 ;
  assign n43894 = ~n43892 & ~n43893 ;
  assign n43895 = ~n43507 & ~n43520 ;
  assign n43896 = x117 & n9433 ;
  assign n43897 = x115 & n9915 ;
  assign n43898 = x116 & n9428 ;
  assign n43899 = ~n43897 & ~n43898 ;
  assign n43900 = ~n43896 & n43899 ;
  assign n43901 = n9436 & n19026 ;
  assign n43902 = n43900 & ~n43901 ;
  assign n43903 = x38 & ~n43902 ;
  assign n43904 = x38 & ~n43903 ;
  assign n43905 = ~n43902 & ~n43903 ;
  assign n43906 = ~n43904 & ~n43905 ;
  assign n43907 = ~n43488 & ~n43501 ;
  assign n43908 = ~n43448 & ~n43462 ;
  assign n43909 = x108 & n14233 ;
  assign n43910 = x106 & n14876 ;
  assign n43911 = x107 & n14228 ;
  assign n43912 = ~n43910 & ~n43911 ;
  assign n43913 = ~n43909 & n43912 ;
  assign n43914 = n13323 & n14236 ;
  assign n43915 = n43913 & ~n43914 ;
  assign n43916 = x47 & ~n43915 ;
  assign n43917 = x47 & ~n43916 ;
  assign n43918 = ~n43915 & ~n43916 ;
  assign n43919 = ~n43917 & ~n43918 ;
  assign n43920 = ~n43440 & ~n43444 ;
  assign n43921 = ~n43405 & ~n43418 ;
  assign n43922 = x99 & n20143 ;
  assign n43923 = x97 & n20854 ;
  assign n43924 = x98 & n20138 ;
  assign n43925 = ~n43923 & ~n43924 ;
  assign n43926 = ~n43922 & n43925 ;
  assign n43927 = n8660 & n20146 ;
  assign n43928 = n43926 & ~n43927 ;
  assign n43929 = x56 & ~n43928 ;
  assign n43930 = x56 & ~n43929 ;
  assign n43931 = ~n43928 & ~n43929 ;
  assign n43932 = ~n43930 & ~n43931 ;
  assign n43933 = ~n43385 & ~n43399 ;
  assign n43934 = x96 & n22325 ;
  assign n43935 = x94 & n23066 ;
  assign n43936 = x95 & n22320 ;
  assign n43937 = ~n43935 & ~n43936 ;
  assign n43938 = ~n43934 & n43937 ;
  assign n43939 = n7321 & n22328 ;
  assign n43940 = n43938 & ~n43939 ;
  assign n43941 = x59 & ~n43940 ;
  assign n43942 = x59 & ~n43941 ;
  assign n43943 = ~n43940 & ~n43941 ;
  assign n43944 = ~n43942 & ~n43943 ;
  assign n43945 = ~n43369 & ~n43382 ;
  assign n43946 = x89 & n27024 ;
  assign n43947 = x90 & ~n26217 ;
  assign n43948 = ~n43946 & ~n43947 ;
  assign n43949 = ~n43366 & n43948 ;
  assign n43950 = n43366 & ~n43948 ;
  assign n43951 = ~n43949 & ~n43950 ;
  assign n43952 = x93 & n24612 ;
  assign n43953 = x91 & n25390 ;
  assign n43954 = x92 & n24607 ;
  assign n43955 = ~n43953 & ~n43954 ;
  assign n43956 = ~n43952 & n43955 ;
  assign n43957 = ~n24615 & n43956 ;
  assign n43958 = ~n6094 & n43956 ;
  assign n43959 = ~n43957 & ~n43958 ;
  assign n43960 = x62 & ~n43959 ;
  assign n43961 = ~x62 & n43959 ;
  assign n43962 = ~n43960 & ~n43961 ;
  assign n43963 = n43951 & ~n43962 ;
  assign n43964 = ~n43951 & n43962 ;
  assign n43965 = ~n43963 & ~n43964 ;
  assign n43966 = ~n43945 & n43965 ;
  assign n43967 = n43945 & ~n43965 ;
  assign n43968 = ~n43966 & ~n43967 ;
  assign n43969 = ~n43944 & n43968 ;
  assign n43970 = n43944 & ~n43968 ;
  assign n43971 = ~n43969 & ~n43970 ;
  assign n43972 = ~n43933 & n43971 ;
  assign n43973 = n43933 & ~n43971 ;
  assign n43974 = ~n43972 & ~n43973 ;
  assign n43975 = ~n43932 & n43974 ;
  assign n43976 = n43932 & ~n43974 ;
  assign n43977 = ~n43975 & ~n43976 ;
  assign n43978 = ~n43921 & n43977 ;
  assign n43979 = n43921 & ~n43977 ;
  assign n43980 = ~n43978 & ~n43979 ;
  assign n43981 = x102 & n18025 ;
  assign n43982 = x100 & n18764 ;
  assign n43983 = x101 & n18020 ;
  assign n43984 = ~n43982 & ~n43983 ;
  assign n43985 = ~n43981 & n43984 ;
  assign n43986 = n10092 & n18028 ;
  assign n43987 = n43985 & ~n43986 ;
  assign n43988 = x53 & ~n43987 ;
  assign n43989 = x53 & ~n43988 ;
  assign n43990 = ~n43987 & ~n43988 ;
  assign n43991 = ~n43989 & ~n43990 ;
  assign n43992 = n43980 & ~n43991 ;
  assign n43993 = n43980 & ~n43992 ;
  assign n43994 = ~n43991 & ~n43992 ;
  assign n43995 = ~n43993 & ~n43994 ;
  assign n43996 = ~n43424 & ~n43438 ;
  assign n43997 = ~n43995 & ~n43996 ;
  assign n43998 = ~n43995 & ~n43997 ;
  assign n43999 = ~n43996 & ~n43997 ;
  assign n44000 = ~n43998 & ~n43999 ;
  assign n44001 = x105 & n16076 ;
  assign n44002 = x103 & n16756 ;
  assign n44003 = x104 & n16071 ;
  assign n44004 = ~n44002 & ~n44003 ;
  assign n44005 = ~n44001 & n44004 ;
  assign n44006 = n11648 & n16079 ;
  assign n44007 = n44005 & ~n44006 ;
  assign n44008 = x50 & ~n44007 ;
  assign n44009 = x50 & ~n44008 ;
  assign n44010 = ~n44007 & ~n44008 ;
  assign n44011 = ~n44009 & ~n44010 ;
  assign n44012 = ~n44000 & n44011 ;
  assign n44013 = n44000 & ~n44011 ;
  assign n44014 = ~n44012 & ~n44013 ;
  assign n44015 = ~n43920 & ~n44014 ;
  assign n44016 = n43920 & n44014 ;
  assign n44017 = ~n44015 & ~n44016 ;
  assign n44018 = ~n43919 & n44017 ;
  assign n44019 = n43919 & ~n44017 ;
  assign n44020 = ~n44018 & ~n44019 ;
  assign n44021 = ~n43908 & n44020 ;
  assign n44022 = n43908 & ~n44020 ;
  assign n44023 = ~n44021 & ~n44022 ;
  assign n44024 = x111 & n12506 ;
  assign n44025 = x109 & n13131 ;
  assign n44026 = x110 & n12501 ;
  assign n44027 = ~n44025 & ~n44026 ;
  assign n44028 = ~n44024 & n44027 ;
  assign n44029 = n12509 & n15111 ;
  assign n44030 = n44028 & ~n44029 ;
  assign n44031 = x44 & ~n44030 ;
  assign n44032 = x44 & ~n44031 ;
  assign n44033 = ~n44030 & ~n44031 ;
  assign n44034 = ~n44032 & ~n44033 ;
  assign n44035 = n44023 & ~n44034 ;
  assign n44036 = n44023 & ~n44035 ;
  assign n44037 = ~n44034 & ~n44035 ;
  assign n44038 = ~n44036 & ~n44037 ;
  assign n44039 = ~n43469 & ~n43482 ;
  assign n44040 = n44038 & n44039 ;
  assign n44041 = ~n44038 & ~n44039 ;
  assign n44042 = ~n44040 & ~n44041 ;
  assign n44043 = x114 & n10905 ;
  assign n44044 = x112 & n11466 ;
  assign n44045 = x113 & n10900 ;
  assign n44046 = ~n44044 & ~n44045 ;
  assign n44047 = ~n44043 & n44046 ;
  assign n44048 = n10908 & n17012 ;
  assign n44049 = n44047 & ~n44048 ;
  assign n44050 = x41 & ~n44049 ;
  assign n44051 = x41 & ~n44050 ;
  assign n44052 = ~n44049 & ~n44050 ;
  assign n44053 = ~n44051 & ~n44052 ;
  assign n44054 = ~n44042 & n44053 ;
  assign n44055 = n44042 & ~n44053 ;
  assign n44056 = ~n44054 & ~n44055 ;
  assign n44057 = ~n43907 & n44056 ;
  assign n44058 = ~n43907 & ~n44057 ;
  assign n44059 = n44056 & ~n44057 ;
  assign n44060 = ~n44058 & ~n44059 ;
  assign n44061 = ~n43906 & ~n44060 ;
  assign n44062 = n43906 & ~n44059 ;
  assign n44063 = ~n44058 & n44062 ;
  assign n44064 = ~n44061 & ~n44063 ;
  assign n44065 = ~n43895 & n44064 ;
  assign n44066 = n43895 & ~n44064 ;
  assign n44067 = ~n44065 & ~n44066 ;
  assign n44068 = ~n43894 & n44067 ;
  assign n44069 = ~n43894 & ~n44068 ;
  assign n44070 = n44067 & ~n44068 ;
  assign n44071 = ~n44069 & ~n44070 ;
  assign n44072 = n43883 & ~n44071 ;
  assign n44073 = n43883 & ~n44072 ;
  assign n44074 = ~n44071 & ~n44072 ;
  assign n44075 = ~n44073 & ~n44074 ;
  assign n44076 = ~n43867 & n44075 ;
  assign n44077 = n43867 & ~n44075 ;
  assign n44078 = ~n44076 & ~n44077 ;
  assign n44079 = ~n43852 & n44078 ;
  assign n44080 = n43852 & ~n44078 ;
  assign n44081 = ~n44079 & ~n44080 ;
  assign n44082 = ~n43840 & n44081 ;
  assign n44083 = n43840 & ~n44081 ;
  assign n44084 = ~n44082 & ~n44083 ;
  assign n44085 = ~n43839 & n44084 ;
  assign n44086 = n43839 & ~n44084 ;
  assign n44087 = ~n44085 & ~n44086 ;
  assign n44338 = n44087 & x217 ;
  assign n44088 = ~n43827 & ~n43831 ;
  assign n44089 = ~n43819 & ~n43823 ;
  assign n44090 = ~n43590 & ~n43804 ;
  assign n44091 = ~x127 & n4847 ;
  assign n44092 = n4534 & n27365 ;
  assign n44093 = ~n44091 & ~n44092 ;
  assign n44094 = ~x26 & ~n44093 ;
  assign n44095 = ~x26 & ~n44094 ;
  assign n44096 = ~n44093 & ~n44094 ;
  assign n44097 = ~n44095 & ~n44096 ;
  assign n44098 = ~n44090 & ~n44097 ;
  assign n44099 = ~n44090 & ~n44098 ;
  assign n44100 = ~n44097 & ~n44098 ;
  assign n44101 = ~n44099 & ~n44100 ;
  assign n44102 = ~x126 & n5560 ;
  assign n44103 = ~x124 & n5943 ;
  assign n44104 = ~x125 & n5555 ;
  assign n44105 = ~n44103 & ~n44104 ;
  assign n44106 = ~n44102 & n44105 ;
  assign n44107 = n5563 & n26128 ;
  assign n44108 = n44106 & ~n44107 ;
  assign n44109 = ~x29 & ~n44108 ;
  assign n44110 = ~x29 & ~n44109 ;
  assign n44111 = ~n44108 & ~n44109 ;
  assign n44112 = ~n44110 & ~n44111 ;
  assign n44113 = ~n43606 & ~n43801 ;
  assign n44114 = n44112 & n44113 ;
  assign n44115 = ~n44112 & ~n44113 ;
  assign n44116 = ~n44114 & ~n44115 ;
  assign n44117 = ~x123 & n6725 ;
  assign n44118 = ~x121 & n7129 ;
  assign n44119 = ~x122 & n6720 ;
  assign n44120 = ~n44118 & ~n44119 ;
  assign n44121 = ~n44117 & n44120 ;
  assign n44122 = n6728 & n23760 ;
  assign n44123 = n44121 & ~n44122 ;
  assign n44124 = ~x32 & ~n44123 ;
  assign n44125 = ~x32 & ~n44124 ;
  assign n44126 = ~n44123 & ~n44124 ;
  assign n44127 = ~n44125 & ~n44126 ;
  assign n44128 = ~n43272 & ~n43783 ;
  assign n44129 = ~n43798 & ~n44128 ;
  assign n44130 = n44127 & n44129 ;
  assign n44131 = ~n44127 & ~n44129 ;
  assign n44132 = ~n44130 & ~n44131 ;
  assign n44133 = ~x120 & n8006 ;
  assign n44134 = ~x118 & n8474 ;
  assign n44135 = ~x119 & n8001 ;
  assign n44136 = ~n44134 & ~n44135 ;
  assign n44137 = ~n44133 & n44136 ;
  assign n44138 = n8009 & n21501 ;
  assign n44139 = n44137 & ~n44138 ;
  assign n44140 = ~x35 & ~n44139 ;
  assign n44141 = ~x35 & ~n44140 ;
  assign n44142 = ~n44139 & ~n44140 ;
  assign n44143 = ~n44141 & ~n44142 ;
  assign n44144 = ~n43767 & ~n43780 ;
  assign n44145 = ~x117 & n9433 ;
  assign n44146 = ~x115 & n9915 ;
  assign n44147 = ~x116 & n9428 ;
  assign n44148 = ~n44146 & ~n44147 ;
  assign n44149 = ~n44145 & n44148 ;
  assign n44150 = n9436 & n19365 ;
  assign n44151 = n44149 & ~n44150 ;
  assign n44152 = ~x38 & ~n44151 ;
  assign n44153 = ~x38 & ~n44152 ;
  assign n44154 = ~n44151 & ~n44152 ;
  assign n44155 = ~n44153 & ~n44154 ;
  assign n44156 = ~n43748 & ~n43761 ;
  assign n44157 = ~n43708 & ~n43722 ;
  assign n44158 = ~x108 & n14233 ;
  assign n44159 = ~x106 & n14876 ;
  assign n44160 = ~x107 & n14228 ;
  assign n44161 = ~n44159 & ~n44160 ;
  assign n44162 = ~n44158 & n44161 ;
  assign n44163 = n13601 & n14236 ;
  assign n44164 = n44162 & ~n44163 ;
  assign n44165 = ~x47 & ~n44164 ;
  assign n44166 = ~x47 & ~n44165 ;
  assign n44167 = ~n44164 & ~n44165 ;
  assign n44168 = ~n44166 & ~n44167 ;
  assign n44169 = ~n43700 & ~n43704 ;
  assign n44170 = ~n43665 & ~n43678 ;
  assign n44171 = ~x99 & n20143 ;
  assign n44172 = ~x97 & n20854 ;
  assign n44173 = ~x98 & n20138 ;
  assign n44174 = ~n44172 & ~n44173 ;
  assign n44175 = ~n44171 & n44174 ;
  assign n44176 = n8885 & n20146 ;
  assign n44177 = n44175 & ~n44176 ;
  assign n44178 = ~x56 & ~n44177 ;
  assign n44179 = ~x56 & ~n44178 ;
  assign n44180 = ~n44177 & ~n44178 ;
  assign n44181 = ~n44179 & ~n44180 ;
  assign n44182 = ~n43645 & ~n43659 ;
  assign n44183 = ~x96 & n22325 ;
  assign n44184 = ~x94 & n23066 ;
  assign n44185 = ~x95 & n22320 ;
  assign n44186 = ~n44184 & ~n44185 ;
  assign n44187 = ~n44183 & n44186 ;
  assign n44188 = n7531 & n22328 ;
  assign n44189 = n44187 & ~n44188 ;
  assign n44190 = ~x59 & ~n44189 ;
  assign n44191 = ~x59 & ~n44190 ;
  assign n44192 = ~n44189 & ~n44190 ;
  assign n44193 = ~n44191 & ~n44192 ;
  assign n44194 = ~n43629 & ~n43642 ;
  assign n44195 = ~x89 & n27427 ;
  assign n44196 = ~x90 & ~n26217 ;
  assign n44197 = ~n44195 & ~n44196 ;
  assign n44198 = ~n43626 & n44197 ;
  assign n44199 = n43626 & ~n44197 ;
  assign n44200 = ~n44198 & ~n44199 ;
  assign n44201 = ~x93 & n24612 ;
  assign n44202 = ~x91 & n25390 ;
  assign n44203 = ~x92 & n24607 ;
  assign n44204 = ~n44202 & ~n44203 ;
  assign n44205 = ~n44201 & n44204 ;
  assign n44206 = ~n24615 & n44205 ;
  assign n44207 = ~n6285 & n44205 ;
  assign n44208 = ~n44206 & ~n44207 ;
  assign n44209 = ~x62 & ~n44208 ;
  assign n44210 = x62 & n44208 ;
  assign n44211 = ~n44209 & ~n44210 ;
  assign n44212 = n44200 & ~n44211 ;
  assign n44213 = ~n44200 & n44211 ;
  assign n44214 = ~n44212 & ~n44213 ;
  assign n44215 = ~n44194 & n44214 ;
  assign n44216 = n44194 & ~n44214 ;
  assign n44217 = ~n44215 & ~n44216 ;
  assign n44218 = ~n44193 & n44217 ;
  assign n44219 = n44193 & ~n44217 ;
  assign n44220 = ~n44218 & ~n44219 ;
  assign n44221 = ~n44182 & n44220 ;
  assign n44222 = n44182 & ~n44220 ;
  assign n44223 = ~n44221 & ~n44222 ;
  assign n44224 = ~n44181 & n44223 ;
  assign n44225 = n44181 & ~n44223 ;
  assign n44226 = ~n44224 & ~n44225 ;
  assign n44227 = ~n44170 & n44226 ;
  assign n44228 = n44170 & ~n44226 ;
  assign n44229 = ~n44227 & ~n44228 ;
  assign n44230 = ~x102 & n18025 ;
  assign n44231 = ~x100 & n18764 ;
  assign n44232 = ~x101 & n18020 ;
  assign n44233 = ~n44231 & ~n44232 ;
  assign n44234 = ~n44230 & n44233 ;
  assign n44235 = n10333 & n18028 ;
  assign n44236 = n44234 & ~n44235 ;
  assign n44237 = ~x53 & ~n44236 ;
  assign n44238 = ~x53 & ~n44237 ;
  assign n44239 = ~n44236 & ~n44237 ;
  assign n44240 = ~n44238 & ~n44239 ;
  assign n44241 = n44229 & ~n44240 ;
  assign n44242 = n44229 & ~n44241 ;
  assign n44243 = ~n44240 & ~n44241 ;
  assign n44244 = ~n44242 & ~n44243 ;
  assign n44245 = ~n43684 & ~n43698 ;
  assign n44246 = ~n44244 & ~n44245 ;
  assign n44247 = ~n44244 & ~n44246 ;
  assign n44248 = ~n44245 & ~n44246 ;
  assign n44249 = ~n44247 & ~n44248 ;
  assign n44250 = ~x105 & n16076 ;
  assign n44251 = ~x103 & n16756 ;
  assign n44252 = ~x104 & n16071 ;
  assign n44253 = ~n44251 & ~n44252 ;
  assign n44254 = ~n44250 & n44253 ;
  assign n44255 = n11907 & n16079 ;
  assign n44256 = n44254 & ~n44255 ;
  assign n44257 = ~x50 & ~n44256 ;
  assign n44258 = ~x50 & ~n44257 ;
  assign n44259 = ~n44256 & ~n44257 ;
  assign n44260 = ~n44258 & ~n44259 ;
  assign n44261 = ~n44249 & n44260 ;
  assign n44262 = n44249 & ~n44260 ;
  assign n44263 = ~n44261 & ~n44262 ;
  assign n44264 = ~n44169 & ~n44263 ;
  assign n44265 = n44169 & n44263 ;
  assign n44266 = ~n44264 & ~n44265 ;
  assign n44267 = ~n44168 & n44266 ;
  assign n44268 = n44168 & ~n44266 ;
  assign n44269 = ~n44267 & ~n44268 ;
  assign n44270 = ~n44157 & n44269 ;
  assign n44271 = n44157 & ~n44269 ;
  assign n44272 = ~n44270 & ~n44271 ;
  assign n44273 = ~x111 & n12506 ;
  assign n44274 = ~x109 & n13131 ;
  assign n44275 = ~x110 & n12501 ;
  assign n44276 = ~n44274 & ~n44275 ;
  assign n44277 = ~n44273 & n44276 ;
  assign n44278 = n12509 & n15411 ;
  assign n44279 = n44277 & ~n44278 ;
  assign n44280 = ~x44 & ~n44279 ;
  assign n44281 = ~x44 & ~n44280 ;
  assign n44282 = ~n44279 & ~n44280 ;
  assign n44283 = ~n44281 & ~n44282 ;
  assign n44284 = n44272 & ~n44283 ;
  assign n44285 = n44272 & ~n44284 ;
  assign n44286 = ~n44283 & ~n44284 ;
  assign n44287 = ~n44285 & ~n44286 ;
  assign n44288 = ~n43729 & ~n43742 ;
  assign n44289 = n44287 & n44288 ;
  assign n44290 = ~n44287 & ~n44288 ;
  assign n44291 = ~n44289 & ~n44290 ;
  assign n44292 = ~x114 & n10905 ;
  assign n44293 = ~x112 & n11466 ;
  assign n44294 = ~x113 & n10900 ;
  assign n44295 = ~n44293 & ~n44294 ;
  assign n44296 = ~n44292 & n44295 ;
  assign n44297 = n10908 & n17333 ;
  assign n44298 = n44296 & ~n44297 ;
  assign n44299 = ~x41 & ~n44298 ;
  assign n44300 = ~x41 & ~n44299 ;
  assign n44301 = ~n44298 & ~n44299 ;
  assign n44302 = ~n44300 & ~n44301 ;
  assign n44303 = ~n44291 & n44302 ;
  assign n44304 = n44291 & ~n44302 ;
  assign n44305 = ~n44303 & ~n44304 ;
  assign n44306 = ~n44156 & n44305 ;
  assign n44307 = ~n44156 & ~n44306 ;
  assign n44308 = n44305 & ~n44306 ;
  assign n44309 = ~n44307 & ~n44308 ;
  assign n44310 = ~n44155 & ~n44309 ;
  assign n44311 = n44155 & ~n44308 ;
  assign n44312 = ~n44307 & n44311 ;
  assign n44313 = ~n44310 & ~n44312 ;
  assign n44314 = ~n44144 & n44313 ;
  assign n44315 = n44144 & ~n44313 ;
  assign n44316 = ~n44314 & ~n44315 ;
  assign n44317 = ~n44143 & n44316 ;
  assign n44318 = ~n44143 & ~n44317 ;
  assign n44319 = n44316 & ~n44317 ;
  assign n44320 = ~n44318 & ~n44319 ;
  assign n44321 = n44132 & ~n44320 ;
  assign n44322 = n44132 & ~n44321 ;
  assign n44323 = ~n44320 & ~n44321 ;
  assign n44324 = ~n44322 & ~n44323 ;
  assign n44325 = ~n44116 & n44324 ;
  assign n44326 = n44116 & ~n44324 ;
  assign n44327 = ~n44325 & ~n44326 ;
  assign n44328 = ~n44101 & n44327 ;
  assign n44329 = n44101 & ~n44327 ;
  assign n44330 = ~n44328 & ~n44329 ;
  assign n44331 = ~n44089 & n44330 ;
  assign n44332 = n44089 & ~n44330 ;
  assign n44333 = ~n44331 & ~n44332 ;
  assign n44334 = ~n44088 & n44333 ;
  assign n44335 = n44088 & ~n44333 ;
  assign n44336 = ~n44334 & ~n44335 ;
  assign n44339 = ~n44336 & ~x217 ;
  assign n44340 = ~n44338 & ~n44339 ;
  assign n44341 = ~n43849 & ~n44079 ;
  assign n44342 = ~n43866 & ~n44077 ;
  assign n44343 = x127 & n5560 ;
  assign n44344 = x125 & n5943 ;
  assign n44345 = x126 & n5555 ;
  assign n44346 = ~n44344 & ~n44345 ;
  assign n44347 = ~n44343 & n44346 ;
  assign n44348 = n5563 & n26533 ;
  assign n44349 = n44347 & ~n44348 ;
  assign n44350 = x29 & ~n44349 ;
  assign n44351 = x29 & ~n44350 ;
  assign n44352 = ~n44349 & ~n44350 ;
  assign n44353 = ~n44351 & ~n44352 ;
  assign n44354 = ~n44342 & ~n44353 ;
  assign n44355 = ~n44342 & ~n44354 ;
  assign n44356 = ~n44353 & ~n44354 ;
  assign n44357 = ~n44355 & ~n44356 ;
  assign n44358 = ~n44057 & ~n44061 ;
  assign n44359 = ~n44041 & ~n44055 ;
  assign n44360 = ~n44015 & ~n44018 ;
  assign n44361 = ~n44000 & ~n44011 ;
  assign n44362 = ~n43997 & ~n44361 ;
  assign n44363 = x97 & n22325 ;
  assign n44364 = x95 & n23066 ;
  assign n44365 = x96 & n22320 ;
  assign n44366 = ~n44364 & ~n44365 ;
  assign n44367 = ~n44363 & n44366 ;
  assign n44368 = n7745 & n22328 ;
  assign n44369 = n44367 & ~n44368 ;
  assign n44370 = x59 & ~n44369 ;
  assign n44371 = x59 & ~n44370 ;
  assign n44372 = ~n44369 & ~n44370 ;
  assign n44373 = ~n44371 & ~n44372 ;
  assign n44374 = ~n43966 & ~n43969 ;
  assign n44375 = n44373 & n44374 ;
  assign n44376 = ~n44373 & ~n44374 ;
  assign n44377 = ~n44375 & ~n44376 ;
  assign n44378 = ~n43949 & ~n43963 ;
  assign n44379 = x90 & n27024 ;
  assign n44380 = x91 & ~n26217 ;
  assign n44381 = ~n44379 & ~n44380 ;
  assign n44382 = ~x26 & ~n44381 ;
  assign n44383 = x26 & n44381 ;
  assign n44384 = ~n44382 & ~n44383 ;
  assign n44385 = ~n43948 & n44384 ;
  assign n44386 = n43948 & ~n44384 ;
  assign n44387 = ~n44385 & ~n44386 ;
  assign n44388 = ~n44378 & n44387 ;
  assign n44389 = n44378 & ~n44387 ;
  assign n44390 = ~n44388 & ~n44389 ;
  assign n44391 = x94 & n24612 ;
  assign n44392 = x92 & n25390 ;
  assign n44393 = x93 & n24607 ;
  assign n44394 = ~n44392 & ~n44393 ;
  assign n44395 = ~n44391 & n44394 ;
  assign n44396 = n6483 & n24615 ;
  assign n44397 = n44395 & ~n44396 ;
  assign n44398 = x62 & ~n44397 ;
  assign n44399 = x62 & ~n44398 ;
  assign n44400 = ~n44397 & ~n44398 ;
  assign n44401 = ~n44399 & ~n44400 ;
  assign n44402 = n44390 & ~n44401 ;
  assign n44403 = n44390 & ~n44402 ;
  assign n44404 = ~n44401 & ~n44402 ;
  assign n44405 = ~n44403 & ~n44404 ;
  assign n44406 = ~n44377 & n44405 ;
  assign n44407 = n44377 & ~n44405 ;
  assign n44408 = ~n44406 & ~n44407 ;
  assign n44409 = x100 & n20143 ;
  assign n44410 = x98 & n20854 ;
  assign n44411 = x99 & n20138 ;
  assign n44412 = ~n44410 & ~n44411 ;
  assign n44413 = ~n44409 & n44412 ;
  assign n44414 = n9115 & n20146 ;
  assign n44415 = n44413 & ~n44414 ;
  assign n44416 = x56 & ~n44415 ;
  assign n44417 = x56 & ~n44416 ;
  assign n44418 = ~n44415 & ~n44416 ;
  assign n44419 = ~n44417 & ~n44418 ;
  assign n44420 = n44408 & ~n44419 ;
  assign n44421 = n44408 & ~n44420 ;
  assign n44422 = ~n44419 & ~n44420 ;
  assign n44423 = ~n44421 & ~n44422 ;
  assign n44424 = ~n43972 & ~n43975 ;
  assign n44425 = n44423 & n44424 ;
  assign n44426 = ~n44423 & ~n44424 ;
  assign n44427 = ~n44425 & ~n44426 ;
  assign n44428 = x103 & n18025 ;
  assign n44429 = x101 & n18764 ;
  assign n44430 = x102 & n18020 ;
  assign n44431 = ~n44429 & ~n44430 ;
  assign n44432 = ~n44428 & n44431 ;
  assign n44433 = n10588 & n18028 ;
  assign n44434 = n44432 & ~n44433 ;
  assign n44435 = x53 & ~n44434 ;
  assign n44436 = x53 & ~n44435 ;
  assign n44437 = ~n44434 & ~n44435 ;
  assign n44438 = ~n44436 & ~n44437 ;
  assign n44439 = n44427 & ~n44438 ;
  assign n44440 = n44427 & ~n44439 ;
  assign n44441 = ~n44438 & ~n44439 ;
  assign n44442 = ~n44440 & ~n44441 ;
  assign n44443 = ~n43978 & ~n43992 ;
  assign n44444 = n44442 & n44443 ;
  assign n44445 = ~n44442 & ~n44443 ;
  assign n44446 = ~n44444 & ~n44445 ;
  assign n44447 = x106 & n16076 ;
  assign n44448 = x104 & n16756 ;
  assign n44449 = x105 & n16071 ;
  assign n44450 = ~n44448 & ~n44449 ;
  assign n44451 = ~n44447 & n44450 ;
  assign n44452 = n12181 & n16079 ;
  assign n44453 = n44451 & ~n44452 ;
  assign n44454 = x50 & ~n44453 ;
  assign n44455 = x50 & ~n44454 ;
  assign n44456 = ~n44453 & ~n44454 ;
  assign n44457 = ~n44455 & ~n44456 ;
  assign n44458 = n44446 & ~n44457 ;
  assign n44459 = n44446 & ~n44458 ;
  assign n44460 = ~n44457 & ~n44458 ;
  assign n44461 = ~n44459 & ~n44460 ;
  assign n44462 = ~n44362 & n44461 ;
  assign n44463 = n44362 & ~n44461 ;
  assign n44464 = ~n44462 & ~n44463 ;
  assign n44465 = x109 & n14233 ;
  assign n44466 = x107 & n14876 ;
  assign n44467 = x108 & n14228 ;
  assign n44468 = ~n44466 & ~n44467 ;
  assign n44469 = ~n44465 & n44468 ;
  assign n44470 = n13894 & n14236 ;
  assign n44471 = n44469 & ~n44470 ;
  assign n44472 = x47 & ~n44471 ;
  assign n44473 = x47 & ~n44472 ;
  assign n44474 = ~n44471 & ~n44472 ;
  assign n44475 = ~n44473 & ~n44474 ;
  assign n44476 = ~n44464 & ~n44475 ;
  assign n44477 = n44464 & n44475 ;
  assign n44478 = ~n44476 & ~n44477 ;
  assign n44479 = n44360 & ~n44478 ;
  assign n44480 = ~n44360 & n44478 ;
  assign n44481 = ~n44479 & ~n44480 ;
  assign n44482 = x112 & n12506 ;
  assign n44483 = x110 & n13131 ;
  assign n44484 = x111 & n12501 ;
  assign n44485 = ~n44483 & ~n44484 ;
  assign n44486 = ~n44482 & n44485 ;
  assign n44487 = n12509 & n15442 ;
  assign n44488 = n44486 & ~n44487 ;
  assign n44489 = x44 & ~n44488 ;
  assign n44490 = x44 & ~n44489 ;
  assign n44491 = ~n44488 & ~n44489 ;
  assign n44492 = ~n44490 & ~n44491 ;
  assign n44493 = n44481 & ~n44492 ;
  assign n44494 = n44481 & ~n44493 ;
  assign n44495 = ~n44492 & ~n44493 ;
  assign n44496 = ~n44494 & ~n44495 ;
  assign n44497 = ~n44021 & ~n44035 ;
  assign n44498 = n44496 & n44497 ;
  assign n44499 = ~n44496 & ~n44497 ;
  assign n44500 = ~n44498 & ~n44499 ;
  assign n44501 = x115 & n10905 ;
  assign n44502 = x113 & n11466 ;
  assign n44503 = x114 & n10900 ;
  assign n44504 = ~n44502 & ~n44503 ;
  assign n44505 = ~n44501 & n44504 ;
  assign n44506 = n10908 & n17364 ;
  assign n44507 = n44505 & ~n44506 ;
  assign n44508 = x41 & ~n44507 ;
  assign n44509 = x41 & ~n44508 ;
  assign n44510 = ~n44507 & ~n44508 ;
  assign n44511 = ~n44509 & ~n44510 ;
  assign n44512 = n44500 & ~n44511 ;
  assign n44513 = ~n44500 & n44511 ;
  assign n44514 = ~n44359 & ~n44513 ;
  assign n44515 = ~n44512 & n44514 ;
  assign n44516 = ~n44359 & ~n44515 ;
  assign n44517 = ~n44512 & ~n44515 ;
  assign n44518 = ~n44513 & n44517 ;
  assign n44519 = ~n44516 & ~n44518 ;
  assign n44520 = x118 & n9433 ;
  assign n44521 = x116 & n9915 ;
  assign n44522 = x117 & n9428 ;
  assign n44523 = ~n44521 & ~n44522 ;
  assign n44524 = ~n44520 & n44523 ;
  assign n44525 = n9436 & n19395 ;
  assign n44526 = n44524 & ~n44525 ;
  assign n44527 = x38 & ~n44526 ;
  assign n44528 = x38 & ~n44527 ;
  assign n44529 = ~n44526 & ~n44527 ;
  assign n44530 = ~n44528 & ~n44529 ;
  assign n44531 = n44519 & n44530 ;
  assign n44532 = ~n44519 & ~n44530 ;
  assign n44533 = ~n44531 & ~n44532 ;
  assign n44534 = ~n44358 & n44533 ;
  assign n44535 = n44358 & ~n44533 ;
  assign n44536 = ~n44534 & ~n44535 ;
  assign n44537 = x121 & n8006 ;
  assign n44538 = x119 & n8474 ;
  assign n44539 = x120 & n8001 ;
  assign n44540 = ~n44538 & ~n44539 ;
  assign n44541 = ~n44537 & n44540 ;
  assign n44542 = n8009 & n21870 ;
  assign n44543 = n44541 & ~n44542 ;
  assign n44544 = x35 & ~n44543 ;
  assign n44545 = x35 & ~n44544 ;
  assign n44546 = ~n44543 & ~n44544 ;
  assign n44547 = ~n44545 & ~n44546 ;
  assign n44548 = n44536 & ~n44547 ;
  assign n44549 = n44536 & ~n44548 ;
  assign n44550 = ~n44547 & ~n44548 ;
  assign n44551 = ~n44549 & ~n44550 ;
  assign n44552 = ~n44065 & ~n44068 ;
  assign n44553 = n44551 & n44552 ;
  assign n44554 = ~n44551 & ~n44552 ;
  assign n44555 = ~n44553 & ~n44554 ;
  assign n44556 = x124 & n6725 ;
  assign n44557 = x122 & n7129 ;
  assign n44558 = x123 & n6720 ;
  assign n44559 = ~n44557 & ~n44558 ;
  assign n44560 = ~n44556 & n44559 ;
  assign n44561 = n6728 & n23796 ;
  assign n44562 = n44560 & ~n44561 ;
  assign n44563 = x32 & ~n44562 ;
  assign n44564 = x32 & ~n44563 ;
  assign n44565 = ~n44562 & ~n44563 ;
  assign n44566 = ~n44564 & ~n44565 ;
  assign n44567 = ~n43882 & ~n44072 ;
  assign n44568 = n44566 & n44567 ;
  assign n44569 = ~n44566 & ~n44567 ;
  assign n44570 = ~n44568 & ~n44569 ;
  assign n44571 = n44555 & ~n44570 ;
  assign n44572 = ~n44555 & n44570 ;
  assign n44573 = ~n44571 & ~n44572 ;
  assign n44574 = ~n44357 & ~n44573 ;
  assign n44575 = n44357 & n44573 ;
  assign n44576 = ~n44574 & ~n44575 ;
  assign n44577 = n44341 & ~n44576 ;
  assign n44578 = ~n44341 & n44576 ;
  assign n44579 = ~n44577 & ~n44578 ;
  assign n44580 = ~n44082 & ~n44085 ;
  assign n44581 = n44579 & ~n44580 ;
  assign n44582 = ~n44579 & n44580 ;
  assign n44583 = ~n44581 & ~n44582 ;
  assign n44828 = n44583 & x218 ;
  assign n44584 = ~n44098 & ~n44328 ;
  assign n44585 = ~n44115 & ~n44326 ;
  assign n44586 = ~x127 & n5560 ;
  assign n44587 = ~x125 & n5943 ;
  assign n44588 = ~x126 & n5555 ;
  assign n44589 = ~n44587 & ~n44588 ;
  assign n44590 = ~n44586 & n44589 ;
  assign n44591 = n5563 & n26932 ;
  assign n44592 = n44590 & ~n44591 ;
  assign n44593 = ~x29 & ~n44592 ;
  assign n44594 = ~x29 & ~n44593 ;
  assign n44595 = ~n44592 & ~n44593 ;
  assign n44596 = ~n44594 & ~n44595 ;
  assign n44597 = ~n44585 & ~n44596 ;
  assign n44598 = ~n44585 & ~n44597 ;
  assign n44599 = ~n44596 & ~n44597 ;
  assign n44600 = ~n44598 & ~n44599 ;
  assign n44601 = ~n44306 & ~n44310 ;
  assign n44602 = ~n44290 & ~n44304 ;
  assign n44603 = ~n44264 & ~n44267 ;
  assign n44604 = ~n44249 & ~n44260 ;
  assign n44605 = ~n44246 & ~n44604 ;
  assign n44606 = ~x97 & n22325 ;
  assign n44607 = ~x95 & n23066 ;
  assign n44608 = ~x96 & n22320 ;
  assign n44609 = ~n44607 & ~n44608 ;
  assign n44610 = ~n44606 & n44609 ;
  assign n44611 = n7949 & n22328 ;
  assign n44612 = n44610 & ~n44611 ;
  assign n44613 = ~x59 & ~n44612 ;
  assign n44614 = ~x59 & ~n44613 ;
  assign n44615 = ~n44612 & ~n44613 ;
  assign n44616 = ~n44614 & ~n44615 ;
  assign n44617 = ~n44215 & ~n44218 ;
  assign n44618 = n44616 & n44617 ;
  assign n44619 = ~n44616 & ~n44617 ;
  assign n44620 = ~n44618 & ~n44619 ;
  assign n44621 = ~n44198 & ~n44212 ;
  assign n44622 = ~x90 & n27427 ;
  assign n44623 = ~x91 & ~n26217 ;
  assign n44624 = ~n44622 & ~n44623 ;
  assign n44625 = x26 & ~n44624 ;
  assign n44626 = ~x26 & n44624 ;
  assign n44627 = ~n44625 & ~n44626 ;
  assign n44628 = ~n44197 & n44627 ;
  assign n44629 = n44197 & ~n44627 ;
  assign n44630 = ~n44628 & ~n44629 ;
  assign n44631 = ~n44621 & n44630 ;
  assign n44632 = n44621 & ~n44630 ;
  assign n44633 = ~n44631 & ~n44632 ;
  assign n44634 = ~x94 & n24612 ;
  assign n44635 = ~x92 & n25390 ;
  assign n44636 = ~x93 & n24607 ;
  assign n44637 = ~n44635 & ~n44636 ;
  assign n44638 = ~n44634 & n44637 ;
  assign n44639 = n6671 & n24615 ;
  assign n44640 = n44638 & ~n44639 ;
  assign n44641 = ~x62 & ~n44640 ;
  assign n44642 = ~x62 & ~n44641 ;
  assign n44643 = ~n44640 & ~n44641 ;
  assign n44644 = ~n44642 & ~n44643 ;
  assign n44645 = n44633 & ~n44644 ;
  assign n44646 = n44633 & ~n44645 ;
  assign n44647 = ~n44644 & ~n44645 ;
  assign n44648 = ~n44646 & ~n44647 ;
  assign n44649 = ~n44620 & n44648 ;
  assign n44650 = n44620 & ~n44648 ;
  assign n44651 = ~n44649 & ~n44650 ;
  assign n44652 = ~x100 & n20143 ;
  assign n44653 = ~x98 & n20854 ;
  assign n44654 = ~x99 & n20138 ;
  assign n44655 = ~n44653 & ~n44654 ;
  assign n44656 = ~n44652 & n44655 ;
  assign n44657 = n9338 & n20146 ;
  assign n44658 = n44656 & ~n44657 ;
  assign n44659 = ~x56 & ~n44658 ;
  assign n44660 = ~x56 & ~n44659 ;
  assign n44661 = ~n44658 & ~n44659 ;
  assign n44662 = ~n44660 & ~n44661 ;
  assign n44663 = n44651 & ~n44662 ;
  assign n44664 = n44651 & ~n44663 ;
  assign n44665 = ~n44662 & ~n44663 ;
  assign n44666 = ~n44664 & ~n44665 ;
  assign n44667 = ~n44221 & ~n44224 ;
  assign n44668 = n44666 & n44667 ;
  assign n44669 = ~n44666 & ~n44667 ;
  assign n44670 = ~n44668 & ~n44669 ;
  assign n44671 = ~x103 & n18025 ;
  assign n44672 = ~x101 & n18764 ;
  assign n44673 = ~x102 & n18020 ;
  assign n44674 = ~n44672 & ~n44673 ;
  assign n44675 = ~n44671 & n44674 ;
  assign n44676 = n10833 & n18028 ;
  assign n44677 = n44675 & ~n44676 ;
  assign n44678 = ~x53 & ~n44677 ;
  assign n44679 = ~x53 & ~n44678 ;
  assign n44680 = ~n44677 & ~n44678 ;
  assign n44681 = ~n44679 & ~n44680 ;
  assign n44682 = n44670 & ~n44681 ;
  assign n44683 = n44670 & ~n44682 ;
  assign n44684 = ~n44681 & ~n44682 ;
  assign n44685 = ~n44683 & ~n44684 ;
  assign n44686 = ~n44227 & ~n44241 ;
  assign n44687 = n44685 & n44686 ;
  assign n44688 = ~n44685 & ~n44686 ;
  assign n44689 = ~n44687 & ~n44688 ;
  assign n44690 = ~x106 & n16076 ;
  assign n44691 = ~x104 & n16756 ;
  assign n44692 = ~x105 & n16071 ;
  assign n44693 = ~n44691 & ~n44692 ;
  assign n44694 = ~n44690 & n44693 ;
  assign n44695 = n12447 & n16079 ;
  assign n44696 = n44694 & ~n44695 ;
  assign n44697 = ~x50 & ~n44696 ;
  assign n44698 = ~x50 & ~n44697 ;
  assign n44699 = ~n44696 & ~n44697 ;
  assign n44700 = ~n44698 & ~n44699 ;
  assign n44701 = n44689 & ~n44700 ;
  assign n44702 = n44689 & ~n44701 ;
  assign n44703 = ~n44700 & ~n44701 ;
  assign n44704 = ~n44702 & ~n44703 ;
  assign n44705 = ~n44605 & n44704 ;
  assign n44706 = n44605 & ~n44704 ;
  assign n44707 = ~n44705 & ~n44706 ;
  assign n44708 = ~x109 & n14233 ;
  assign n44709 = ~x107 & n14876 ;
  assign n44710 = ~x108 & n14228 ;
  assign n44711 = ~n44709 & ~n44710 ;
  assign n44712 = ~n44708 & n44711 ;
  assign n44713 = n14177 & n14236 ;
  assign n44714 = n44712 & ~n44713 ;
  assign n44715 = ~x47 & ~n44714 ;
  assign n44716 = ~x47 & ~n44715 ;
  assign n44717 = ~n44714 & ~n44715 ;
  assign n44718 = ~n44716 & ~n44717 ;
  assign n44719 = ~n44707 & ~n44718 ;
  assign n44720 = n44707 & n44718 ;
  assign n44721 = ~n44719 & ~n44720 ;
  assign n44722 = n44603 & ~n44721 ;
  assign n44723 = ~n44603 & n44721 ;
  assign n44724 = ~n44722 & ~n44723 ;
  assign n44725 = ~x112 & n12506 ;
  assign n44726 = ~x110 & n13131 ;
  assign n44727 = ~x111 & n12501 ;
  assign n44728 = ~n44726 & ~n44727 ;
  assign n44729 = ~n44725 & n44728 ;
  assign n44730 = n12509 & n15744 ;
  assign n44731 = n44729 & ~n44730 ;
  assign n44732 = ~x44 & ~n44731 ;
  assign n44733 = ~x44 & ~n44732 ;
  assign n44734 = ~n44731 & ~n44732 ;
  assign n44735 = ~n44733 & ~n44734 ;
  assign n44736 = n44724 & ~n44735 ;
  assign n44737 = n44724 & ~n44736 ;
  assign n44738 = ~n44735 & ~n44736 ;
  assign n44739 = ~n44737 & ~n44738 ;
  assign n44740 = ~n44270 & ~n44284 ;
  assign n44741 = n44739 & n44740 ;
  assign n44742 = ~n44739 & ~n44740 ;
  assign n44743 = ~n44741 & ~n44742 ;
  assign n44744 = ~x115 & n10905 ;
  assign n44745 = ~x113 & n11466 ;
  assign n44746 = ~x114 & n10900 ;
  assign n44747 = ~n44745 & ~n44746 ;
  assign n44748 = ~n44744 & n44747 ;
  assign n44749 = n10908 & n17683 ;
  assign n44750 = n44748 & ~n44749 ;
  assign n44751 = ~x41 & ~n44750 ;
  assign n44752 = ~x41 & ~n44751 ;
  assign n44753 = ~n44750 & ~n44751 ;
  assign n44754 = ~n44752 & ~n44753 ;
  assign n44755 = n44743 & ~n44754 ;
  assign n44756 = ~n44743 & n44754 ;
  assign n44757 = ~n44602 & ~n44756 ;
  assign n44758 = ~n44755 & n44757 ;
  assign n44759 = ~n44602 & ~n44758 ;
  assign n44760 = ~n44755 & ~n44758 ;
  assign n44761 = ~n44756 & n44760 ;
  assign n44762 = ~n44759 & ~n44761 ;
  assign n44763 = ~x118 & n9433 ;
  assign n44764 = ~x116 & n9915 ;
  assign n44765 = ~x117 & n9428 ;
  assign n44766 = ~n44764 & ~n44765 ;
  assign n44767 = ~n44763 & n44766 ;
  assign n44768 = n9436 & n19736 ;
  assign n44769 = n44767 & ~n44768 ;
  assign n44770 = ~x38 & ~n44769 ;
  assign n44771 = ~x38 & ~n44770 ;
  assign n44772 = ~n44769 & ~n44770 ;
  assign n44773 = ~n44771 & ~n44772 ;
  assign n44774 = n44762 & n44773 ;
  assign n44775 = ~n44762 & ~n44773 ;
  assign n44776 = ~n44774 & ~n44775 ;
  assign n44777 = ~n44601 & n44776 ;
  assign n44778 = n44601 & ~n44776 ;
  assign n44779 = ~n44777 & ~n44778 ;
  assign n44780 = ~x121 & n8006 ;
  assign n44781 = ~x119 & n8474 ;
  assign n44782 = ~x120 & n8001 ;
  assign n44783 = ~n44781 & ~n44782 ;
  assign n44784 = ~n44780 & n44783 ;
  assign n44785 = n8009 & n22229 ;
  assign n44786 = n44784 & ~n44785 ;
  assign n44787 = ~x35 & ~n44786 ;
  assign n44788 = ~x35 & ~n44787 ;
  assign n44789 = ~n44786 & ~n44787 ;
  assign n44790 = ~n44788 & ~n44789 ;
  assign n44791 = n44779 & ~n44790 ;
  assign n44792 = n44779 & ~n44791 ;
  assign n44793 = ~n44790 & ~n44791 ;
  assign n44794 = ~n44792 & ~n44793 ;
  assign n44795 = ~n44314 & ~n44317 ;
  assign n44796 = n44794 & n44795 ;
  assign n44797 = ~n44794 & ~n44795 ;
  assign n44798 = ~n44796 & ~n44797 ;
  assign n44799 = ~x124 & n6725 ;
  assign n44800 = ~x122 & n7129 ;
  assign n44801 = ~x123 & n6720 ;
  assign n44802 = ~n44800 & ~n44801 ;
  assign n44803 = ~n44799 & n44802 ;
  assign n44804 = n6728 & n24176 ;
  assign n44805 = n44803 & ~n44804 ;
  assign n44806 = ~x32 & ~n44805 ;
  assign n44807 = ~x32 & ~n44806 ;
  assign n44808 = ~n44805 & ~n44806 ;
  assign n44809 = ~n44807 & ~n44808 ;
  assign n44810 = ~n44131 & ~n44321 ;
  assign n44811 = n44809 & n44810 ;
  assign n44812 = ~n44809 & ~n44810 ;
  assign n44813 = ~n44811 & ~n44812 ;
  assign n44814 = n44798 & ~n44813 ;
  assign n44815 = ~n44798 & n44813 ;
  assign n44816 = ~n44814 & ~n44815 ;
  assign n44817 = ~n44600 & ~n44816 ;
  assign n44818 = n44600 & n44816 ;
  assign n44819 = ~n44817 & ~n44818 ;
  assign n44820 = n44584 & ~n44819 ;
  assign n44821 = ~n44584 & n44819 ;
  assign n44822 = ~n44820 & ~n44821 ;
  assign n44823 = ~n44331 & ~n44334 ;
  assign n44824 = n44822 & ~n44823 ;
  assign n44825 = ~n44822 & n44823 ;
  assign n44826 = ~n44824 & ~n44825 ;
  assign n44829 = ~n44826 & ~x218 ;
  assign n44830 = ~n44828 & ~n44829 ;
  assign n44831 = n44555 & n44570 ;
  assign n44832 = ~n44569 & ~n44831 ;
  assign n44833 = x126 & n5943 ;
  assign n44834 = x127 & n5555 ;
  assign n44835 = ~n44833 & ~n44834 ;
  assign n44836 = ~n5563 & n44835 ;
  assign n44837 = n26965 & n44835 ;
  assign n44838 = ~n44836 & ~n44837 ;
  assign n44839 = x29 & ~n44838 ;
  assign n44840 = ~x29 & n44838 ;
  assign n44841 = ~n44839 & ~n44840 ;
  assign n44842 = ~n44832 & ~n44841 ;
  assign n44843 = n44832 & n44841 ;
  assign n44844 = ~n44842 & ~n44843 ;
  assign n44845 = x125 & n6725 ;
  assign n44846 = x123 & n7129 ;
  assign n44847 = x124 & n6720 ;
  assign n44848 = ~n44846 & ~n44847 ;
  assign n44849 = ~n44845 & n44848 ;
  assign n44850 = n6728 & n24935 ;
  assign n44851 = n44849 & ~n44850 ;
  assign n44852 = x32 & ~n44851 ;
  assign n44853 = x32 & ~n44852 ;
  assign n44854 = ~n44851 & ~n44852 ;
  assign n44855 = ~n44853 & ~n44854 ;
  assign n44856 = ~n44548 & ~n44554 ;
  assign n44857 = n44855 & n44856 ;
  assign n44858 = ~n44855 & ~n44856 ;
  assign n44859 = ~n44857 & ~n44858 ;
  assign n44860 = ~n44532 & ~n44534 ;
  assign n44861 = ~n44439 & ~n44445 ;
  assign n44862 = x104 & n18025 ;
  assign n44863 = x102 & n18764 ;
  assign n44864 = x103 & n18020 ;
  assign n44865 = ~n44863 & ~n44864 ;
  assign n44866 = ~n44862 & n44865 ;
  assign n44867 = n11116 & n18028 ;
  assign n44868 = n44866 & ~n44867 ;
  assign n44869 = x53 & ~n44868 ;
  assign n44870 = x53 & ~n44869 ;
  assign n44871 = ~n44868 & ~n44869 ;
  assign n44872 = ~n44870 & ~n44871 ;
  assign n44873 = ~n44420 & ~n44426 ;
  assign n44874 = x91 & n27024 ;
  assign n44875 = x92 & ~n26217 ;
  assign n44876 = ~n44874 & ~n44875 ;
  assign n44877 = ~n44382 & ~n44385 ;
  assign n44878 = ~n44876 & n44877 ;
  assign n44879 = n44876 & ~n44877 ;
  assign n44880 = ~n44878 & ~n44879 ;
  assign n44881 = x95 & n24612 ;
  assign n44882 = x93 & n25390 ;
  assign n44883 = x94 & n24607 ;
  assign n44884 = ~n44882 & ~n44883 ;
  assign n44885 = ~n44881 & n44884 ;
  assign n44886 = n6894 & n24615 ;
  assign n44887 = n44885 & ~n44886 ;
  assign n44888 = x62 & ~n44887 ;
  assign n44889 = x62 & ~n44888 ;
  assign n44890 = ~n44887 & ~n44888 ;
  assign n44891 = ~n44889 & ~n44890 ;
  assign n44892 = ~n44880 & n44891 ;
  assign n44893 = n44880 & ~n44891 ;
  assign n44894 = ~n44892 & ~n44893 ;
  assign n44895 = ~n44388 & ~n44402 ;
  assign n44896 = n44894 & ~n44895 ;
  assign n44897 = ~n44894 & n44895 ;
  assign n44898 = ~n44896 & ~n44897 ;
  assign n44899 = x98 & n22325 ;
  assign n44900 = x96 & n23066 ;
  assign n44901 = x97 & n22320 ;
  assign n44902 = ~n44900 & ~n44901 ;
  assign n44903 = ~n44899 & n44902 ;
  assign n44904 = n8196 & n22328 ;
  assign n44905 = n44903 & ~n44904 ;
  assign n44906 = x59 & ~n44905 ;
  assign n44907 = x59 & ~n44906 ;
  assign n44908 = ~n44905 & ~n44906 ;
  assign n44909 = ~n44907 & ~n44908 ;
  assign n44910 = n44898 & ~n44909 ;
  assign n44911 = n44898 & ~n44910 ;
  assign n44912 = ~n44909 & ~n44910 ;
  assign n44913 = ~n44911 & ~n44912 ;
  assign n44914 = ~n44376 & ~n44407 ;
  assign n44915 = ~n44913 & ~n44914 ;
  assign n44916 = ~n44913 & ~n44915 ;
  assign n44917 = ~n44914 & ~n44915 ;
  assign n44918 = ~n44916 & ~n44917 ;
  assign n44919 = x101 & n20143 ;
  assign n44920 = x99 & n20854 ;
  assign n44921 = x100 & n20138 ;
  assign n44922 = ~n44920 & ~n44921 ;
  assign n44923 = ~n44919 & n44922 ;
  assign n44924 = n9601 & n20146 ;
  assign n44925 = n44923 & ~n44924 ;
  assign n44926 = x56 & ~n44925 ;
  assign n44927 = x56 & ~n44926 ;
  assign n44928 = ~n44925 & ~n44926 ;
  assign n44929 = ~n44927 & ~n44928 ;
  assign n44930 = ~n44918 & n44929 ;
  assign n44931 = n44918 & ~n44929 ;
  assign n44932 = ~n44930 & ~n44931 ;
  assign n44933 = ~n44873 & ~n44932 ;
  assign n44934 = ~n44873 & ~n44933 ;
  assign n44935 = ~n44932 & ~n44933 ;
  assign n44936 = ~n44934 & ~n44935 ;
  assign n44937 = ~n44872 & ~n44936 ;
  assign n44938 = n44872 & ~n44935 ;
  assign n44939 = ~n44934 & n44938 ;
  assign n44940 = ~n44937 & ~n44939 ;
  assign n44941 = ~n44861 & n44940 ;
  assign n44942 = n44861 & ~n44940 ;
  assign n44943 = ~n44941 & ~n44942 ;
  assign n44944 = x107 & n16076 ;
  assign n44945 = x105 & n16756 ;
  assign n44946 = x106 & n16071 ;
  assign n44947 = ~n44945 & ~n44946 ;
  assign n44948 = ~n44944 & n44947 ;
  assign n44949 = n12749 & n16079 ;
  assign n44950 = n44948 & ~n44949 ;
  assign n44951 = x50 & ~n44950 ;
  assign n44952 = x50 & ~n44951 ;
  assign n44953 = ~n44950 & ~n44951 ;
  assign n44954 = ~n44952 & ~n44953 ;
  assign n44955 = n44943 & ~n44954 ;
  assign n44956 = n44943 & ~n44955 ;
  assign n44957 = ~n44954 & ~n44955 ;
  assign n44958 = ~n44956 & ~n44957 ;
  assign n44959 = ~n44362 & ~n44461 ;
  assign n44960 = ~n44458 & ~n44959 ;
  assign n44961 = n44958 & n44960 ;
  assign n44962 = ~n44958 & ~n44960 ;
  assign n44963 = ~n44961 & ~n44962 ;
  assign n44964 = x110 & n14233 ;
  assign n44965 = x108 & n14876 ;
  assign n44966 = x109 & n14228 ;
  assign n44967 = ~n44965 & ~n44966 ;
  assign n44968 = ~n44964 & n44967 ;
  assign n44969 = n14236 & n14497 ;
  assign n44970 = n44968 & ~n44969 ;
  assign n44971 = x47 & ~n44970 ;
  assign n44972 = x47 & ~n44971 ;
  assign n44973 = ~n44970 & ~n44971 ;
  assign n44974 = ~n44972 & ~n44973 ;
  assign n44975 = n44963 & ~n44974 ;
  assign n44976 = n44963 & ~n44975 ;
  assign n44977 = ~n44974 & ~n44975 ;
  assign n44978 = ~n44976 & ~n44977 ;
  assign n44979 = ~n44476 & ~n44480 ;
  assign n44980 = n44978 & n44979 ;
  assign n44981 = ~n44978 & ~n44979 ;
  assign n44982 = ~n44980 & ~n44981 ;
  assign n44983 = x113 & n12506 ;
  assign n44984 = x111 & n13131 ;
  assign n44985 = x112 & n12501 ;
  assign n44986 = ~n44984 & ~n44985 ;
  assign n44987 = ~n44983 & n44986 ;
  assign n44988 = n12509 & n16361 ;
  assign n44989 = n44987 & ~n44988 ;
  assign n44990 = x44 & ~n44989 ;
  assign n44991 = x44 & ~n44990 ;
  assign n44992 = ~n44989 & ~n44990 ;
  assign n44993 = ~n44991 & ~n44992 ;
  assign n44994 = n44982 & ~n44993 ;
  assign n44995 = n44982 & ~n44994 ;
  assign n44996 = ~n44993 & ~n44994 ;
  assign n44997 = ~n44995 & ~n44996 ;
  assign n44998 = ~n44493 & ~n44499 ;
  assign n44999 = n44997 & n44998 ;
  assign n45000 = ~n44997 & ~n44998 ;
  assign n45001 = ~n44999 & ~n45000 ;
  assign n45002 = x116 & n10905 ;
  assign n45003 = x114 & n11466 ;
  assign n45004 = x115 & n10900 ;
  assign n45005 = ~n45003 & ~n45004 ;
  assign n45006 = ~n45002 & n45005 ;
  assign n45007 = n10908 & n18336 ;
  assign n45008 = n45006 & ~n45007 ;
  assign n45009 = x41 & ~n45008 ;
  assign n45010 = x41 & ~n45009 ;
  assign n45011 = ~n45008 & ~n45009 ;
  assign n45012 = ~n45010 & ~n45011 ;
  assign n45013 = n45001 & ~n45012 ;
  assign n45014 = n45001 & ~n45013 ;
  assign n45015 = ~n45012 & ~n45013 ;
  assign n45016 = ~n45014 & ~n45015 ;
  assign n45017 = ~n44517 & n45016 ;
  assign n45018 = n44517 & ~n45016 ;
  assign n45019 = ~n45017 & ~n45018 ;
  assign n45020 = x119 & n9433 ;
  assign n45021 = x117 & n9915 ;
  assign n45022 = x118 & n9428 ;
  assign n45023 = ~n45021 & ~n45022 ;
  assign n45024 = ~n45020 & n45023 ;
  assign n45025 = n9436 & n20423 ;
  assign n45026 = n45024 & ~n45025 ;
  assign n45027 = x38 & ~n45026 ;
  assign n45028 = x38 & ~n45027 ;
  assign n45029 = ~n45026 & ~n45027 ;
  assign n45030 = ~n45028 & ~n45029 ;
  assign n45031 = ~n45019 & ~n45030 ;
  assign n45032 = n45019 & n45030 ;
  assign n45033 = ~n45031 & ~n45032 ;
  assign n45034 = ~n44860 & n45033 ;
  assign n45035 = n44860 & ~n45033 ;
  assign n45036 = ~n45034 & ~n45035 ;
  assign n45037 = x122 & n8006 ;
  assign n45038 = x120 & n8474 ;
  assign n45039 = x121 & n8001 ;
  assign n45040 = ~n45038 & ~n45039 ;
  assign n45041 = ~n45037 & n45040 ;
  assign n45042 = n8009 & n22622 ;
  assign n45043 = n45041 & ~n45042 ;
  assign n45044 = x35 & ~n45043 ;
  assign n45045 = x35 & ~n45044 ;
  assign n45046 = ~n45043 & ~n45044 ;
  assign n45047 = ~n45045 & ~n45046 ;
  assign n45048 = n45036 & ~n45047 ;
  assign n45049 = n45036 & ~n45048 ;
  assign n45050 = ~n45047 & ~n45048 ;
  assign n45051 = ~n45049 & ~n45050 ;
  assign n45052 = n44859 & ~n45051 ;
  assign n45053 = ~n44859 & n45051 ;
  assign n45054 = n44844 & ~n45053 ;
  assign n45055 = ~n45052 & n45054 ;
  assign n45056 = n44844 & ~n45055 ;
  assign n45057 = ~n45053 & ~n45055 ;
  assign n45058 = ~n45052 & n45057 ;
  assign n45059 = ~n45056 & ~n45058 ;
  assign n45060 = ~n44354 & ~n44574 ;
  assign n45061 = n45059 & n45060 ;
  assign n45062 = ~n45059 & ~n45060 ;
  assign n45063 = ~n45061 & ~n45062 ;
  assign n45064 = ~n44578 & ~n44581 ;
  assign n45065 = n45063 & ~n45064 ;
  assign n45066 = ~n45063 & n45064 ;
  assign n45067 = ~n45065 & ~n45066 ;
  assign n45306 = n45067 & x219 ;
  assign n45068 = n44798 & n44813 ;
  assign n45069 = ~n44812 & ~n45068 ;
  assign n45070 = ~x126 & n5943 ;
  assign n45071 = ~x127 & n5555 ;
  assign n45072 = ~n45070 & ~n45071 ;
  assign n45073 = ~n5563 & n45072 ;
  assign n45074 = n27368 & n45072 ;
  assign n45075 = ~n45073 & ~n45074 ;
  assign n45076 = ~x29 & ~n45075 ;
  assign n45077 = x29 & n45075 ;
  assign n45078 = ~n45076 & ~n45077 ;
  assign n45079 = ~n45069 & ~n45078 ;
  assign n45080 = n45069 & n45078 ;
  assign n45081 = ~n45079 & ~n45080 ;
  assign n45082 = ~x125 & n6725 ;
  assign n45083 = ~x123 & n7129 ;
  assign n45084 = ~x124 & n6720 ;
  assign n45085 = ~n45083 & ~n45084 ;
  assign n45086 = ~n45082 & n45085 ;
  assign n45087 = n6728 & n25330 ;
  assign n45088 = n45086 & ~n45087 ;
  assign n45089 = ~x32 & ~n45088 ;
  assign n45090 = ~x32 & ~n45089 ;
  assign n45091 = ~n45088 & ~n45089 ;
  assign n45092 = ~n45090 & ~n45091 ;
  assign n45093 = ~n44791 & ~n44797 ;
  assign n45094 = n45092 & n45093 ;
  assign n45095 = ~n45092 & ~n45093 ;
  assign n45096 = ~n45094 & ~n45095 ;
  assign n45097 = ~n44775 & ~n44777 ;
  assign n45098 = ~n44682 & ~n44688 ;
  assign n45099 = ~x104 & n18025 ;
  assign n45100 = ~x102 & n18764 ;
  assign n45101 = ~x103 & n18020 ;
  assign n45102 = ~n45100 & ~n45101 ;
  assign n45103 = ~n45099 & n45102 ;
  assign n45104 = n11380 & n18028 ;
  assign n45105 = n45103 & ~n45104 ;
  assign n45106 = ~x53 & ~n45105 ;
  assign n45107 = ~x53 & ~n45106 ;
  assign n45108 = ~n45105 & ~n45106 ;
  assign n45109 = ~n45107 & ~n45108 ;
  assign n45110 = ~n44663 & ~n44669 ;
  assign n45111 = ~x91 & n27427 ;
  assign n45112 = ~x92 & ~n26217 ;
  assign n45113 = ~n45111 & ~n45112 ;
  assign n45114 = ~n44625 & ~n44628 ;
  assign n45115 = ~n45113 & n45114 ;
  assign n45116 = n45113 & ~n45114 ;
  assign n45117 = ~n45115 & ~n45116 ;
  assign n45118 = ~x95 & n24612 ;
  assign n45119 = ~x93 & n25390 ;
  assign n45120 = ~x94 & n24607 ;
  assign n45121 = ~n45119 & ~n45120 ;
  assign n45122 = ~n45118 & n45121 ;
  assign n45123 = n7100 & n24615 ;
  assign n45124 = n45122 & ~n45123 ;
  assign n45125 = ~x62 & ~n45124 ;
  assign n45126 = ~x62 & ~n45125 ;
  assign n45127 = ~n45124 & ~n45125 ;
  assign n45128 = ~n45126 & ~n45127 ;
  assign n45129 = ~n45117 & n45128 ;
  assign n45130 = n45117 & ~n45128 ;
  assign n45131 = ~n45129 & ~n45130 ;
  assign n45132 = ~n44631 & ~n44645 ;
  assign n45133 = n45131 & ~n45132 ;
  assign n45134 = ~n45131 & n45132 ;
  assign n45135 = ~n45133 & ~n45134 ;
  assign n45136 = ~x98 & n22325 ;
  assign n45137 = ~x96 & n23066 ;
  assign n45138 = ~x97 & n22320 ;
  assign n45139 = ~n45137 & ~n45138 ;
  assign n45140 = ~n45136 & n45139 ;
  assign n45141 = n8426 & n22328 ;
  assign n45142 = n45140 & ~n45141 ;
  assign n45143 = ~x59 & ~n45142 ;
  assign n45144 = ~x59 & ~n45143 ;
  assign n45145 = ~n45142 & ~n45143 ;
  assign n45146 = ~n45144 & ~n45145 ;
  assign n45147 = n45135 & ~n45146 ;
  assign n45148 = n45135 & ~n45147 ;
  assign n45149 = ~n45146 & ~n45147 ;
  assign n45150 = ~n45148 & ~n45149 ;
  assign n45151 = ~n44619 & ~n44650 ;
  assign n45152 = ~n45150 & ~n45151 ;
  assign n45153 = ~n45150 & ~n45152 ;
  assign n45154 = ~n45151 & ~n45152 ;
  assign n45155 = ~n45153 & ~n45154 ;
  assign n45156 = ~x101 & n20143 ;
  assign n45157 = ~x99 & n20854 ;
  assign n45158 = ~x100 & n20138 ;
  assign n45159 = ~n45157 & ~n45158 ;
  assign n45160 = ~n45156 & n45159 ;
  assign n45161 = n9844 & n20146 ;
  assign n45162 = n45160 & ~n45161 ;
  assign n45163 = ~x56 & ~n45162 ;
  assign n45164 = ~x56 & ~n45163 ;
  assign n45165 = ~n45162 & ~n45163 ;
  assign n45166 = ~n45164 & ~n45165 ;
  assign n45167 = ~n45155 & n45166 ;
  assign n45168 = n45155 & ~n45166 ;
  assign n45169 = ~n45167 & ~n45168 ;
  assign n45170 = ~n45110 & ~n45169 ;
  assign n45171 = ~n45110 & ~n45170 ;
  assign n45172 = ~n45169 & ~n45170 ;
  assign n45173 = ~n45171 & ~n45172 ;
  assign n45174 = ~n45109 & ~n45173 ;
  assign n45175 = n45109 & ~n45172 ;
  assign n45176 = ~n45171 & n45175 ;
  assign n45177 = ~n45174 & ~n45176 ;
  assign n45178 = ~n45098 & n45177 ;
  assign n45179 = n45098 & ~n45177 ;
  assign n45180 = ~n45178 & ~n45179 ;
  assign n45181 = ~x107 & n16076 ;
  assign n45182 = ~x105 & n16756 ;
  assign n45183 = ~x106 & n16071 ;
  assign n45184 = ~n45182 & ~n45183 ;
  assign n45185 = ~n45181 & n45184 ;
  assign n45186 = n13034 & n16079 ;
  assign n45187 = n45185 & ~n45186 ;
  assign n45188 = ~x50 & ~n45187 ;
  assign n45189 = ~x50 & ~n45188 ;
  assign n45190 = ~n45187 & ~n45188 ;
  assign n45191 = ~n45189 & ~n45190 ;
  assign n45192 = n45180 & ~n45191 ;
  assign n45193 = n45180 & ~n45192 ;
  assign n45194 = ~n45191 & ~n45192 ;
  assign n45195 = ~n45193 & ~n45194 ;
  assign n45196 = ~n44605 & ~n44704 ;
  assign n45197 = ~n44701 & ~n45196 ;
  assign n45198 = n45195 & n45197 ;
  assign n45199 = ~n45195 & ~n45197 ;
  assign n45200 = ~n45198 & ~n45199 ;
  assign n45201 = ~x110 & n14233 ;
  assign n45202 = ~x108 & n14876 ;
  assign n45203 = ~x109 & n14228 ;
  assign n45204 = ~n45202 & ~n45203 ;
  assign n45205 = ~n45201 & n45204 ;
  assign n45206 = n14236 & n14802 ;
  assign n45207 = n45205 & ~n45206 ;
  assign n45208 = ~x47 & ~n45207 ;
  assign n45209 = ~x47 & ~n45208 ;
  assign n45210 = ~n45207 & ~n45208 ;
  assign n45211 = ~n45209 & ~n45210 ;
  assign n45212 = n45200 & ~n45211 ;
  assign n45213 = n45200 & ~n45212 ;
  assign n45214 = ~n45211 & ~n45212 ;
  assign n45215 = ~n45213 & ~n45214 ;
  assign n45216 = ~n44719 & ~n44723 ;
  assign n45217 = n45215 & n45216 ;
  assign n45218 = ~n45215 & ~n45216 ;
  assign n45219 = ~n45217 & ~n45218 ;
  assign n45220 = ~x113 & n12506 ;
  assign n45221 = ~x111 & n13131 ;
  assign n45222 = ~x112 & n12501 ;
  assign n45223 = ~n45221 & ~n45222 ;
  assign n45224 = ~n45220 & n45223 ;
  assign n45225 = n12509 & n16684 ;
  assign n45226 = n45224 & ~n45225 ;
  assign n45227 = ~x44 & ~n45226 ;
  assign n45228 = ~x44 & ~n45227 ;
  assign n45229 = ~n45226 & ~n45227 ;
  assign n45230 = ~n45228 & ~n45229 ;
  assign n45231 = n45219 & ~n45230 ;
  assign n45232 = n45219 & ~n45231 ;
  assign n45233 = ~n45230 & ~n45231 ;
  assign n45234 = ~n45232 & ~n45233 ;
  assign n45235 = ~n44736 & ~n44742 ;
  assign n45236 = n45234 & n45235 ;
  assign n45237 = ~n45234 & ~n45235 ;
  assign n45238 = ~n45236 & ~n45237 ;
  assign n45239 = ~x116 & n10905 ;
  assign n45240 = ~x114 & n11466 ;
  assign n45241 = ~x115 & n10900 ;
  assign n45242 = ~n45240 & ~n45241 ;
  assign n45243 = ~n45239 & n45242 ;
  assign n45244 = n10908 & n18678 ;
  assign n45245 = n45243 & ~n45244 ;
  assign n45246 = ~x41 & ~n45245 ;
  assign n45247 = ~x41 & ~n45246 ;
  assign n45248 = ~n45245 & ~n45246 ;
  assign n45249 = ~n45247 & ~n45248 ;
  assign n45250 = n45238 & ~n45249 ;
  assign n45251 = n45238 & ~n45250 ;
  assign n45252 = ~n45249 & ~n45250 ;
  assign n45253 = ~n45251 & ~n45252 ;
  assign n45254 = ~n44760 & n45253 ;
  assign n45255 = n44760 & ~n45253 ;
  assign n45256 = ~n45254 & ~n45255 ;
  assign n45257 = ~x119 & n9433 ;
  assign n45258 = ~x117 & n9915 ;
  assign n45259 = ~x118 & n9428 ;
  assign n45260 = ~n45258 & ~n45259 ;
  assign n45261 = ~n45257 & n45260 ;
  assign n45262 = n9436 & n20778 ;
  assign n45263 = n45261 & ~n45262 ;
  assign n45264 = ~x38 & ~n45263 ;
  assign n45265 = ~x38 & ~n45264 ;
  assign n45266 = ~n45263 & ~n45264 ;
  assign n45267 = ~n45265 & ~n45266 ;
  assign n45268 = ~n45256 & ~n45267 ;
  assign n45269 = n45256 & n45267 ;
  assign n45270 = ~n45268 & ~n45269 ;
  assign n45271 = ~n45097 & n45270 ;
  assign n45272 = n45097 & ~n45270 ;
  assign n45273 = ~n45271 & ~n45272 ;
  assign n45274 = ~x122 & n8006 ;
  assign n45275 = ~x120 & n8474 ;
  assign n45276 = ~x121 & n8001 ;
  assign n45277 = ~n45275 & ~n45276 ;
  assign n45278 = ~n45274 & n45277 ;
  assign n45279 = n8009 & n22998 ;
  assign n45280 = n45278 & ~n45279 ;
  assign n45281 = ~x35 & ~n45280 ;
  assign n45282 = ~x35 & ~n45281 ;
  assign n45283 = ~n45280 & ~n45281 ;
  assign n45284 = ~n45282 & ~n45283 ;
  assign n45285 = n45273 & ~n45284 ;
  assign n45286 = n45273 & ~n45285 ;
  assign n45287 = ~n45284 & ~n45285 ;
  assign n45288 = ~n45286 & ~n45287 ;
  assign n45289 = n45096 & ~n45288 ;
  assign n45290 = ~n45096 & n45288 ;
  assign n45291 = n45081 & ~n45290 ;
  assign n45292 = ~n45289 & n45291 ;
  assign n45293 = n45081 & ~n45292 ;
  assign n45294 = ~n45290 & ~n45292 ;
  assign n45295 = ~n45289 & n45294 ;
  assign n45296 = ~n45293 & ~n45295 ;
  assign n45297 = ~n44597 & ~n44817 ;
  assign n45298 = n45296 & n45297 ;
  assign n45299 = ~n45296 & ~n45297 ;
  assign n45300 = ~n45298 & ~n45299 ;
  assign n45301 = ~n44821 & ~n44824 ;
  assign n45302 = n45300 & ~n45301 ;
  assign n45303 = ~n45300 & n45301 ;
  assign n45304 = ~n45302 & ~n45303 ;
  assign n45307 = ~n45304 & ~x219 ;
  assign n45308 = ~n45306 & ~n45307 ;
  assign n45309 = ~n45062 & ~n45065 ;
  assign n45310 = ~n44842 & ~n45055 ;
  assign n45311 = ~n44858 & ~n45052 ;
  assign n45312 = x127 & n5943 ;
  assign n45313 = n5563 & n26962 ;
  assign n45314 = ~n45312 & ~n45313 ;
  assign n45315 = x29 & ~n45314 ;
  assign n45316 = x29 & ~n45315 ;
  assign n45317 = ~n45314 & ~n45315 ;
  assign n45318 = ~n45316 & ~n45317 ;
  assign n45319 = ~n45311 & ~n45318 ;
  assign n45320 = ~n45311 & ~n45319 ;
  assign n45321 = ~n45318 & ~n45319 ;
  assign n45322 = ~n45320 & ~n45321 ;
  assign n45323 = x126 & n6725 ;
  assign n45324 = x124 & n7129 ;
  assign n45325 = x125 & n6720 ;
  assign n45326 = ~n45324 & ~n45325 ;
  assign n45327 = ~n45323 & n45326 ;
  assign n45328 = n6728 & n25735 ;
  assign n45329 = n45327 & ~n45328 ;
  assign n45330 = x32 & ~n45329 ;
  assign n45331 = x32 & ~n45330 ;
  assign n45332 = ~n45329 & ~n45330 ;
  assign n45333 = ~n45331 & ~n45332 ;
  assign n45334 = ~n45034 & ~n45048 ;
  assign n45335 = n45333 & n45334 ;
  assign n45336 = ~n45333 & ~n45334 ;
  assign n45337 = ~n45335 & ~n45336 ;
  assign n45338 = ~n44517 & ~n45016 ;
  assign n45339 = ~n45031 & ~n45338 ;
  assign n45340 = x120 & n9433 ;
  assign n45341 = x118 & n9915 ;
  assign n45342 = x119 & n9428 ;
  assign n45343 = ~n45341 & ~n45342 ;
  assign n45344 = ~n45340 & n45343 ;
  assign n45345 = n9436 & n21143 ;
  assign n45346 = n45344 & ~n45345 ;
  assign n45347 = x38 & ~n45346 ;
  assign n45348 = x38 & ~n45347 ;
  assign n45349 = ~n45346 & ~n45347 ;
  assign n45350 = ~n45348 & ~n45349 ;
  assign n45351 = ~n45000 & ~n45013 ;
  assign n45352 = x117 & n10905 ;
  assign n45353 = x115 & n11466 ;
  assign n45354 = x116 & n10900 ;
  assign n45355 = ~n45353 & ~n45354 ;
  assign n45356 = ~n45352 & n45355 ;
  assign n45357 = n10908 & n19026 ;
  assign n45358 = n45356 & ~n45357 ;
  assign n45359 = x41 & ~n45358 ;
  assign n45360 = x41 & ~n45359 ;
  assign n45361 = ~n45358 & ~n45359 ;
  assign n45362 = ~n45360 & ~n45361 ;
  assign n45363 = ~n44981 & ~n44994 ;
  assign n45364 = ~n44941 & ~n44955 ;
  assign n45365 = x108 & n16076 ;
  assign n45366 = x106 & n16756 ;
  assign n45367 = x107 & n16071 ;
  assign n45368 = ~n45366 & ~n45367 ;
  assign n45369 = ~n45365 & n45368 ;
  assign n45370 = n13323 & n16079 ;
  assign n45371 = n45369 & ~n45370 ;
  assign n45372 = x50 & ~n45371 ;
  assign n45373 = x50 & ~n45372 ;
  assign n45374 = ~n45371 & ~n45372 ;
  assign n45375 = ~n45373 & ~n45374 ;
  assign n45376 = ~n44933 & ~n44937 ;
  assign n45377 = ~n44896 & ~n44910 ;
  assign n45378 = x99 & n22325 ;
  assign n45379 = x97 & n23066 ;
  assign n45380 = x98 & n22320 ;
  assign n45381 = ~n45379 & ~n45380 ;
  assign n45382 = ~n45378 & n45381 ;
  assign n45383 = n8660 & n22328 ;
  assign n45384 = n45382 & ~n45383 ;
  assign n45385 = x59 & ~n45384 ;
  assign n45386 = x59 & ~n45385 ;
  assign n45387 = ~n45384 & ~n45385 ;
  assign n45388 = ~n45386 & ~n45387 ;
  assign n45389 = ~n44879 & ~n44893 ;
  assign n45390 = x92 & n27024 ;
  assign n45391 = x93 & ~n26217 ;
  assign n45392 = ~n45390 & ~n45391 ;
  assign n45393 = n44876 & ~n45392 ;
  assign n45394 = ~n44876 & n45392 ;
  assign n45395 = ~n45389 & ~n45394 ;
  assign n45396 = ~n45393 & n45395 ;
  assign n45397 = ~n45389 & ~n45396 ;
  assign n45398 = ~n45394 & ~n45396 ;
  assign n45399 = ~n45393 & n45398 ;
  assign n45400 = ~n45397 & ~n45399 ;
  assign n45401 = x96 & n24612 ;
  assign n45402 = x94 & n25390 ;
  assign n45403 = x95 & n24607 ;
  assign n45404 = ~n45402 & ~n45403 ;
  assign n45405 = ~n45401 & n45404 ;
  assign n45406 = n7321 & n24615 ;
  assign n45407 = n45405 & ~n45406 ;
  assign n45408 = x62 & ~n45407 ;
  assign n45409 = x62 & ~n45408 ;
  assign n45410 = ~n45407 & ~n45408 ;
  assign n45411 = ~n45409 & ~n45410 ;
  assign n45412 = ~n45400 & n45411 ;
  assign n45413 = n45400 & ~n45411 ;
  assign n45414 = ~n45412 & ~n45413 ;
  assign n45415 = ~n45388 & ~n45414 ;
  assign n45416 = n45388 & n45414 ;
  assign n45417 = ~n45415 & ~n45416 ;
  assign n45418 = ~n45377 & n45417 ;
  assign n45419 = n45377 & ~n45417 ;
  assign n45420 = ~n45418 & ~n45419 ;
  assign n45421 = x102 & n20143 ;
  assign n45422 = x100 & n20854 ;
  assign n45423 = x101 & n20138 ;
  assign n45424 = ~n45422 & ~n45423 ;
  assign n45425 = ~n45421 & n45424 ;
  assign n45426 = n10092 & n20146 ;
  assign n45427 = n45425 & ~n45426 ;
  assign n45428 = x56 & ~n45427 ;
  assign n45429 = x56 & ~n45428 ;
  assign n45430 = ~n45427 & ~n45428 ;
  assign n45431 = ~n45429 & ~n45430 ;
  assign n45432 = n45420 & ~n45431 ;
  assign n45433 = n45420 & ~n45432 ;
  assign n45434 = ~n45431 & ~n45432 ;
  assign n45435 = ~n45433 & ~n45434 ;
  assign n45436 = ~n44918 & ~n44929 ;
  assign n45437 = ~n44915 & ~n45436 ;
  assign n45438 = ~n45435 & ~n45437 ;
  assign n45439 = ~n45435 & ~n45438 ;
  assign n45440 = ~n45437 & ~n45438 ;
  assign n45441 = ~n45439 & ~n45440 ;
  assign n45442 = x105 & n18025 ;
  assign n45443 = x103 & n18764 ;
  assign n45444 = x104 & n18020 ;
  assign n45445 = ~n45443 & ~n45444 ;
  assign n45446 = ~n45442 & n45445 ;
  assign n45447 = n11648 & n18028 ;
  assign n45448 = n45446 & ~n45447 ;
  assign n45449 = x53 & ~n45448 ;
  assign n45450 = x53 & ~n45449 ;
  assign n45451 = ~n45448 & ~n45449 ;
  assign n45452 = ~n45450 & ~n45451 ;
  assign n45453 = ~n45441 & n45452 ;
  assign n45454 = n45441 & ~n45452 ;
  assign n45455 = ~n45453 & ~n45454 ;
  assign n45456 = ~n45376 & ~n45455 ;
  assign n45457 = n45376 & n45455 ;
  assign n45458 = ~n45456 & ~n45457 ;
  assign n45459 = ~n45375 & n45458 ;
  assign n45460 = n45375 & ~n45458 ;
  assign n45461 = ~n45459 & ~n45460 ;
  assign n45462 = ~n45364 & n45461 ;
  assign n45463 = n45364 & ~n45461 ;
  assign n45464 = ~n45462 & ~n45463 ;
  assign n45465 = x111 & n14233 ;
  assign n45466 = x109 & n14876 ;
  assign n45467 = x110 & n14228 ;
  assign n45468 = ~n45466 & ~n45467 ;
  assign n45469 = ~n45465 & n45468 ;
  assign n45470 = n14236 & n15111 ;
  assign n45471 = n45469 & ~n45470 ;
  assign n45472 = x47 & ~n45471 ;
  assign n45473 = x47 & ~n45472 ;
  assign n45474 = ~n45471 & ~n45472 ;
  assign n45475 = ~n45473 & ~n45474 ;
  assign n45476 = n45464 & ~n45475 ;
  assign n45477 = n45464 & ~n45476 ;
  assign n45478 = ~n45475 & ~n45476 ;
  assign n45479 = ~n45477 & ~n45478 ;
  assign n45480 = ~n44962 & ~n44975 ;
  assign n45481 = n45479 & n45480 ;
  assign n45482 = ~n45479 & ~n45480 ;
  assign n45483 = ~n45481 & ~n45482 ;
  assign n45484 = x114 & n12506 ;
  assign n45485 = x112 & n13131 ;
  assign n45486 = x113 & n12501 ;
  assign n45487 = ~n45485 & ~n45486 ;
  assign n45488 = ~n45484 & n45487 ;
  assign n45489 = n12509 & n17012 ;
  assign n45490 = n45488 & ~n45489 ;
  assign n45491 = x44 & ~n45490 ;
  assign n45492 = x44 & ~n45491 ;
  assign n45493 = ~n45490 & ~n45491 ;
  assign n45494 = ~n45492 & ~n45493 ;
  assign n45495 = ~n45483 & n45494 ;
  assign n45496 = n45483 & ~n45494 ;
  assign n45497 = ~n45495 & ~n45496 ;
  assign n45498 = ~n45363 & n45497 ;
  assign n45499 = ~n45363 & ~n45498 ;
  assign n45500 = n45497 & ~n45498 ;
  assign n45501 = ~n45499 & ~n45500 ;
  assign n45502 = ~n45362 & ~n45501 ;
  assign n45503 = n45362 & ~n45500 ;
  assign n45504 = ~n45499 & n45503 ;
  assign n45505 = ~n45502 & ~n45504 ;
  assign n45506 = ~n45351 & n45505 ;
  assign n45507 = n45351 & ~n45505 ;
  assign n45508 = ~n45506 & ~n45507 ;
  assign n45509 = ~n45350 & n45508 ;
  assign n45510 = n45350 & ~n45508 ;
  assign n45511 = ~n45509 & ~n45510 ;
  assign n45512 = ~n45339 & n45511 ;
  assign n45513 = n45339 & ~n45511 ;
  assign n45514 = ~n45512 & ~n45513 ;
  assign n45515 = x123 & n8006 ;
  assign n45516 = x121 & n8474 ;
  assign n45517 = x122 & n8001 ;
  assign n45518 = ~n45516 & ~n45517 ;
  assign n45519 = ~n45515 & n45518 ;
  assign n45520 = n8009 & n23382 ;
  assign n45521 = n45519 & ~n45520 ;
  assign n45522 = x35 & ~n45521 ;
  assign n45523 = x35 & ~n45522 ;
  assign n45524 = ~n45521 & ~n45522 ;
  assign n45525 = ~n45523 & ~n45524 ;
  assign n45526 = n45514 & ~n45525 ;
  assign n45527 = n45514 & ~n45526 ;
  assign n45528 = ~n45525 & ~n45526 ;
  assign n45529 = ~n45527 & ~n45528 ;
  assign n45530 = ~n45337 & n45529 ;
  assign n45531 = n45337 & ~n45529 ;
  assign n45532 = ~n45530 & ~n45531 ;
  assign n45533 = ~n45322 & n45532 ;
  assign n45534 = n45322 & ~n45532 ;
  assign n45535 = ~n45533 & ~n45534 ;
  assign n45536 = ~n45310 & n45535 ;
  assign n45537 = ~n45310 & ~n45536 ;
  assign n45538 = n45535 & ~n45536 ;
  assign n45539 = ~n45537 & ~n45538 ;
  assign n45540 = ~n45309 & ~n45539 ;
  assign n45541 = n45309 & ~n45538 ;
  assign n45542 = ~n45537 & n45541 ;
  assign n45543 = ~n45540 & ~n45542 ;
  assign n45780 = n45543 & x220 ;
  assign n45544 = ~n45299 & ~n45302 ;
  assign n45545 = ~n45079 & ~n45292 ;
  assign n45546 = ~n45095 & ~n45289 ;
  assign n45547 = ~x127 & n5943 ;
  assign n45548 = n5563 & n27365 ;
  assign n45549 = ~n45547 & ~n45548 ;
  assign n45550 = ~x29 & ~n45549 ;
  assign n45551 = ~x29 & ~n45550 ;
  assign n45552 = ~n45549 & ~n45550 ;
  assign n45553 = ~n45551 & ~n45552 ;
  assign n45554 = ~n45546 & ~n45553 ;
  assign n45555 = ~n45546 & ~n45554 ;
  assign n45556 = ~n45553 & ~n45554 ;
  assign n45557 = ~n45555 & ~n45556 ;
  assign n45558 = ~x126 & n6725 ;
  assign n45559 = ~x124 & n7129 ;
  assign n45560 = ~x125 & n6720 ;
  assign n45561 = ~n45559 & ~n45560 ;
  assign n45562 = ~n45558 & n45561 ;
  assign n45563 = n6728 & n26128 ;
  assign n45564 = n45562 & ~n45563 ;
  assign n45565 = ~x32 & ~n45564 ;
  assign n45566 = ~x32 & ~n45565 ;
  assign n45567 = ~n45564 & ~n45565 ;
  assign n45568 = ~n45566 & ~n45567 ;
  assign n45569 = ~n45271 & ~n45285 ;
  assign n45570 = n45568 & n45569 ;
  assign n45571 = ~n45568 & ~n45569 ;
  assign n45572 = ~n45570 & ~n45571 ;
  assign n45573 = ~n44760 & ~n45253 ;
  assign n45574 = ~n45268 & ~n45573 ;
  assign n45575 = ~x120 & n9433 ;
  assign n45576 = ~x118 & n9915 ;
  assign n45577 = ~x119 & n9428 ;
  assign n45578 = ~n45576 & ~n45577 ;
  assign n45579 = ~n45575 & n45578 ;
  assign n45580 = n9436 & n21501 ;
  assign n45581 = n45579 & ~n45580 ;
  assign n45582 = ~x38 & ~n45581 ;
  assign n45583 = ~x38 & ~n45582 ;
  assign n45584 = ~n45581 & ~n45582 ;
  assign n45585 = ~n45583 & ~n45584 ;
  assign n45586 = ~n45237 & ~n45250 ;
  assign n45587 = ~x117 & n10905 ;
  assign n45588 = ~x115 & n11466 ;
  assign n45589 = ~x116 & n10900 ;
  assign n45590 = ~n45588 & ~n45589 ;
  assign n45591 = ~n45587 & n45590 ;
  assign n45592 = n10908 & n19365 ;
  assign n45593 = n45591 & ~n45592 ;
  assign n45594 = ~x41 & ~n45593 ;
  assign n45595 = ~x41 & ~n45594 ;
  assign n45596 = ~n45593 & ~n45594 ;
  assign n45597 = ~n45595 & ~n45596 ;
  assign n45598 = ~n45218 & ~n45231 ;
  assign n45599 = ~n45178 & ~n45192 ;
  assign n45600 = ~x108 & n16076 ;
  assign n45601 = ~x106 & n16756 ;
  assign n45602 = ~x107 & n16071 ;
  assign n45603 = ~n45601 & ~n45602 ;
  assign n45604 = ~n45600 & n45603 ;
  assign n45605 = n13601 & n16079 ;
  assign n45606 = n45604 & ~n45605 ;
  assign n45607 = ~x50 & ~n45606 ;
  assign n45608 = ~x50 & ~n45607 ;
  assign n45609 = ~n45606 & ~n45607 ;
  assign n45610 = ~n45608 & ~n45609 ;
  assign n45611 = ~n45170 & ~n45174 ;
  assign n45612 = ~n45133 & ~n45147 ;
  assign n45613 = ~x99 & n22325 ;
  assign n45614 = ~x97 & n23066 ;
  assign n45615 = ~x98 & n22320 ;
  assign n45616 = ~n45614 & ~n45615 ;
  assign n45617 = ~n45613 & n45616 ;
  assign n45618 = n8885 & n22328 ;
  assign n45619 = n45617 & ~n45618 ;
  assign n45620 = ~x59 & ~n45619 ;
  assign n45621 = ~x59 & ~n45620 ;
  assign n45622 = ~n45619 & ~n45620 ;
  assign n45623 = ~n45621 & ~n45622 ;
  assign n45624 = ~n45116 & ~n45130 ;
  assign n45625 = ~x92 & n27427 ;
  assign n45626 = ~x93 & ~n26217 ;
  assign n45627 = ~n45625 & ~n45626 ;
  assign n45628 = n45113 & ~n45627 ;
  assign n45629 = ~n45113 & n45627 ;
  assign n45630 = ~n45624 & ~n45629 ;
  assign n45631 = ~n45628 & n45630 ;
  assign n45632 = ~n45624 & ~n45631 ;
  assign n45633 = ~n45629 & ~n45631 ;
  assign n45634 = ~n45628 & n45633 ;
  assign n45635 = ~n45632 & ~n45634 ;
  assign n45636 = ~x96 & n24612 ;
  assign n45637 = ~x94 & n25390 ;
  assign n45638 = ~x95 & n24607 ;
  assign n45639 = ~n45637 & ~n45638 ;
  assign n45640 = ~n45636 & n45639 ;
  assign n45641 = n7531 & n24615 ;
  assign n45642 = n45640 & ~n45641 ;
  assign n45643 = ~x62 & ~n45642 ;
  assign n45644 = ~x62 & ~n45643 ;
  assign n45645 = ~n45642 & ~n45643 ;
  assign n45646 = ~n45644 & ~n45645 ;
  assign n45647 = ~n45635 & n45646 ;
  assign n45648 = n45635 & ~n45646 ;
  assign n45649 = ~n45647 & ~n45648 ;
  assign n45650 = ~n45623 & ~n45649 ;
  assign n45651 = n45623 & n45649 ;
  assign n45652 = ~n45650 & ~n45651 ;
  assign n45653 = ~n45612 & n45652 ;
  assign n45654 = n45612 & ~n45652 ;
  assign n45655 = ~n45653 & ~n45654 ;
  assign n45656 = ~x102 & n20143 ;
  assign n45657 = ~x100 & n20854 ;
  assign n45658 = ~x101 & n20138 ;
  assign n45659 = ~n45657 & ~n45658 ;
  assign n45660 = ~n45656 & n45659 ;
  assign n45661 = n10333 & n20146 ;
  assign n45662 = n45660 & ~n45661 ;
  assign n45663 = ~x56 & ~n45662 ;
  assign n45664 = ~x56 & ~n45663 ;
  assign n45665 = ~n45662 & ~n45663 ;
  assign n45666 = ~n45664 & ~n45665 ;
  assign n45667 = n45655 & ~n45666 ;
  assign n45668 = n45655 & ~n45667 ;
  assign n45669 = ~n45666 & ~n45667 ;
  assign n45670 = ~n45668 & ~n45669 ;
  assign n45671 = ~n45155 & ~n45166 ;
  assign n45672 = ~n45152 & ~n45671 ;
  assign n45673 = ~n45670 & ~n45672 ;
  assign n45674 = ~n45670 & ~n45673 ;
  assign n45675 = ~n45672 & ~n45673 ;
  assign n45676 = ~n45674 & ~n45675 ;
  assign n45677 = ~x105 & n18025 ;
  assign n45678 = ~x103 & n18764 ;
  assign n45679 = ~x104 & n18020 ;
  assign n45680 = ~n45678 & ~n45679 ;
  assign n45681 = ~n45677 & n45680 ;
  assign n45682 = n11907 & n18028 ;
  assign n45683 = n45681 & ~n45682 ;
  assign n45684 = ~x53 & ~n45683 ;
  assign n45685 = ~x53 & ~n45684 ;
  assign n45686 = ~n45683 & ~n45684 ;
  assign n45687 = ~n45685 & ~n45686 ;
  assign n45688 = ~n45676 & n45687 ;
  assign n45689 = n45676 & ~n45687 ;
  assign n45690 = ~n45688 & ~n45689 ;
  assign n45691 = ~n45611 & ~n45690 ;
  assign n45692 = n45611 & n45690 ;
  assign n45693 = ~n45691 & ~n45692 ;
  assign n45694 = ~n45610 & n45693 ;
  assign n45695 = n45610 & ~n45693 ;
  assign n45696 = ~n45694 & ~n45695 ;
  assign n45697 = ~n45599 & n45696 ;
  assign n45698 = n45599 & ~n45696 ;
  assign n45699 = ~n45697 & ~n45698 ;
  assign n45700 = ~x111 & n14233 ;
  assign n45701 = ~x109 & n14876 ;
  assign n45702 = ~x110 & n14228 ;
  assign n45703 = ~n45701 & ~n45702 ;
  assign n45704 = ~n45700 & n45703 ;
  assign n45705 = n14236 & n15411 ;
  assign n45706 = n45704 & ~n45705 ;
  assign n45707 = ~x47 & ~n45706 ;
  assign n45708 = ~x47 & ~n45707 ;
  assign n45709 = ~n45706 & ~n45707 ;
  assign n45710 = ~n45708 & ~n45709 ;
  assign n45711 = n45699 & ~n45710 ;
  assign n45712 = n45699 & ~n45711 ;
  assign n45713 = ~n45710 & ~n45711 ;
  assign n45714 = ~n45712 & ~n45713 ;
  assign n45715 = ~n45199 & ~n45212 ;
  assign n45716 = n45714 & n45715 ;
  assign n45717 = ~n45714 & ~n45715 ;
  assign n45718 = ~n45716 & ~n45717 ;
  assign n45719 = ~x114 & n12506 ;
  assign n45720 = ~x112 & n13131 ;
  assign n45721 = ~x113 & n12501 ;
  assign n45722 = ~n45720 & ~n45721 ;
  assign n45723 = ~n45719 & n45722 ;
  assign n45724 = n12509 & n17333 ;
  assign n45725 = n45723 & ~n45724 ;
  assign n45726 = ~x44 & ~n45725 ;
  assign n45727 = ~x44 & ~n45726 ;
  assign n45728 = ~n45725 & ~n45726 ;
  assign n45729 = ~n45727 & ~n45728 ;
  assign n45730 = ~n45718 & n45729 ;
  assign n45731 = n45718 & ~n45729 ;
  assign n45732 = ~n45730 & ~n45731 ;
  assign n45733 = ~n45598 & n45732 ;
  assign n45734 = ~n45598 & ~n45733 ;
  assign n45735 = n45732 & ~n45733 ;
  assign n45736 = ~n45734 & ~n45735 ;
  assign n45737 = ~n45597 & ~n45736 ;
  assign n45738 = n45597 & ~n45735 ;
  assign n45739 = ~n45734 & n45738 ;
  assign n45740 = ~n45737 & ~n45739 ;
  assign n45741 = ~n45586 & n45740 ;
  assign n45742 = n45586 & ~n45740 ;
  assign n45743 = ~n45741 & ~n45742 ;
  assign n45744 = ~n45585 & n45743 ;
  assign n45745 = n45585 & ~n45743 ;
  assign n45746 = ~n45744 & ~n45745 ;
  assign n45747 = ~n45574 & n45746 ;
  assign n45748 = n45574 & ~n45746 ;
  assign n45749 = ~n45747 & ~n45748 ;
  assign n45750 = ~x123 & n8006 ;
  assign n45751 = ~x121 & n8474 ;
  assign n45752 = ~x122 & n8001 ;
  assign n45753 = ~n45751 & ~n45752 ;
  assign n45754 = ~n45750 & n45753 ;
  assign n45755 = n8009 & n23760 ;
  assign n45756 = n45754 & ~n45755 ;
  assign n45757 = ~x35 & ~n45756 ;
  assign n45758 = ~x35 & ~n45757 ;
  assign n45759 = ~n45756 & ~n45757 ;
  assign n45760 = ~n45758 & ~n45759 ;
  assign n45761 = n45749 & ~n45760 ;
  assign n45762 = n45749 & ~n45761 ;
  assign n45763 = ~n45760 & ~n45761 ;
  assign n45764 = ~n45762 & ~n45763 ;
  assign n45765 = ~n45572 & n45764 ;
  assign n45766 = n45572 & ~n45764 ;
  assign n45767 = ~n45765 & ~n45766 ;
  assign n45768 = ~n45557 & n45767 ;
  assign n45769 = n45557 & ~n45767 ;
  assign n45770 = ~n45768 & ~n45769 ;
  assign n45771 = ~n45545 & n45770 ;
  assign n45772 = ~n45545 & ~n45771 ;
  assign n45773 = n45770 & ~n45771 ;
  assign n45774 = ~n45772 & ~n45773 ;
  assign n45775 = ~n45544 & ~n45774 ;
  assign n45776 = n45544 & ~n45773 ;
  assign n45777 = ~n45772 & n45776 ;
  assign n45778 = ~n45775 & ~n45777 ;
  assign n45781 = ~n45778 & ~x220 ;
  assign n45782 = ~n45780 & ~n45781 ;
  assign n45783 = ~n45536 & ~n45540 ;
  assign n45784 = ~n45319 & ~n45533 ;
  assign n45785 = ~n45498 & ~n45502 ;
  assign n45786 = ~n45482 & ~n45496 ;
  assign n45787 = ~n45456 & ~n45459 ;
  assign n45788 = ~n45441 & ~n45452 ;
  assign n45789 = ~n45438 & ~n45788 ;
  assign n45790 = ~n45400 & ~n45411 ;
  assign n45791 = ~n45415 & ~n45790 ;
  assign n45792 = x93 & n27024 ;
  assign n45793 = x94 & ~n26217 ;
  assign n45794 = ~n45792 & ~n45793 ;
  assign n45795 = ~x29 & ~n45794 ;
  assign n45796 = x29 & n45794 ;
  assign n45797 = ~n45795 & ~n45796 ;
  assign n45798 = ~n45392 & n45797 ;
  assign n45799 = ~n45392 & ~n45798 ;
  assign n45800 = n45797 & ~n45798 ;
  assign n45801 = ~n45799 & ~n45800 ;
  assign n45802 = ~n45398 & ~n45801 ;
  assign n45803 = ~n45398 & ~n45802 ;
  assign n45804 = ~n45801 & ~n45802 ;
  assign n45805 = ~n45803 & ~n45804 ;
  assign n45806 = x97 & n24612 ;
  assign n45807 = x95 & n25390 ;
  assign n45808 = x96 & n24607 ;
  assign n45809 = ~n45807 & ~n45808 ;
  assign n45810 = ~n45806 & n45809 ;
  assign n45811 = n7745 & n24615 ;
  assign n45812 = n45810 & ~n45811 ;
  assign n45813 = x62 & ~n45812 ;
  assign n45814 = x62 & ~n45813 ;
  assign n45815 = ~n45812 & ~n45813 ;
  assign n45816 = ~n45814 & ~n45815 ;
  assign n45817 = ~n45805 & n45816 ;
  assign n45818 = n45805 & ~n45816 ;
  assign n45819 = ~n45817 & ~n45818 ;
  assign n45820 = x100 & n22325 ;
  assign n45821 = x98 & n23066 ;
  assign n45822 = x99 & n22320 ;
  assign n45823 = ~n45821 & ~n45822 ;
  assign n45824 = ~n45820 & n45823 ;
  assign n45825 = n9115 & n22328 ;
  assign n45826 = n45824 & ~n45825 ;
  assign n45827 = x59 & ~n45826 ;
  assign n45828 = x59 & ~n45827 ;
  assign n45829 = ~n45826 & ~n45827 ;
  assign n45830 = ~n45828 & ~n45829 ;
  assign n45831 = ~n45819 & ~n45830 ;
  assign n45832 = n45819 & n45830 ;
  assign n45833 = ~n45831 & ~n45832 ;
  assign n45834 = ~n45791 & n45833 ;
  assign n45835 = n45791 & ~n45833 ;
  assign n45836 = ~n45834 & ~n45835 ;
  assign n45837 = x103 & n20143 ;
  assign n45838 = x101 & n20854 ;
  assign n45839 = x102 & n20138 ;
  assign n45840 = ~n45838 & ~n45839 ;
  assign n45841 = ~n45837 & n45840 ;
  assign n45842 = n10588 & n20146 ;
  assign n45843 = n45841 & ~n45842 ;
  assign n45844 = x56 & ~n45843 ;
  assign n45845 = x56 & ~n45844 ;
  assign n45846 = ~n45843 & ~n45844 ;
  assign n45847 = ~n45845 & ~n45846 ;
  assign n45848 = n45836 & ~n45847 ;
  assign n45849 = n45836 & ~n45848 ;
  assign n45850 = ~n45847 & ~n45848 ;
  assign n45851 = ~n45849 & ~n45850 ;
  assign n45852 = ~n45418 & ~n45432 ;
  assign n45853 = n45851 & n45852 ;
  assign n45854 = ~n45851 & ~n45852 ;
  assign n45855 = ~n45853 & ~n45854 ;
  assign n45856 = x106 & n18025 ;
  assign n45857 = x104 & n18764 ;
  assign n45858 = x105 & n18020 ;
  assign n45859 = ~n45857 & ~n45858 ;
  assign n45860 = ~n45856 & n45859 ;
  assign n45861 = n12181 & n18028 ;
  assign n45862 = n45860 & ~n45861 ;
  assign n45863 = x53 & ~n45862 ;
  assign n45864 = x53 & ~n45863 ;
  assign n45865 = ~n45862 & ~n45863 ;
  assign n45866 = ~n45864 & ~n45865 ;
  assign n45867 = n45855 & ~n45866 ;
  assign n45868 = n45855 & ~n45867 ;
  assign n45869 = ~n45866 & ~n45867 ;
  assign n45870 = ~n45868 & ~n45869 ;
  assign n45871 = ~n45789 & n45870 ;
  assign n45872 = n45789 & ~n45870 ;
  assign n45873 = ~n45871 & ~n45872 ;
  assign n45874 = x109 & n16076 ;
  assign n45875 = x107 & n16756 ;
  assign n45876 = x108 & n16071 ;
  assign n45877 = ~n45875 & ~n45876 ;
  assign n45878 = ~n45874 & n45877 ;
  assign n45879 = n13894 & n16079 ;
  assign n45880 = n45878 & ~n45879 ;
  assign n45881 = x50 & ~n45880 ;
  assign n45882 = x50 & ~n45881 ;
  assign n45883 = ~n45880 & ~n45881 ;
  assign n45884 = ~n45882 & ~n45883 ;
  assign n45885 = ~n45873 & ~n45884 ;
  assign n45886 = n45873 & n45884 ;
  assign n45887 = ~n45885 & ~n45886 ;
  assign n45888 = n45787 & ~n45887 ;
  assign n45889 = ~n45787 & n45887 ;
  assign n45890 = ~n45888 & ~n45889 ;
  assign n45891 = x112 & n14233 ;
  assign n45892 = x110 & n14876 ;
  assign n45893 = x111 & n14228 ;
  assign n45894 = ~n45892 & ~n45893 ;
  assign n45895 = ~n45891 & n45894 ;
  assign n45896 = n14236 & n15442 ;
  assign n45897 = n45895 & ~n45896 ;
  assign n45898 = x47 & ~n45897 ;
  assign n45899 = x47 & ~n45898 ;
  assign n45900 = ~n45897 & ~n45898 ;
  assign n45901 = ~n45899 & ~n45900 ;
  assign n45902 = n45890 & ~n45901 ;
  assign n45903 = n45890 & ~n45902 ;
  assign n45904 = ~n45901 & ~n45902 ;
  assign n45905 = ~n45903 & ~n45904 ;
  assign n45906 = ~n45462 & ~n45476 ;
  assign n45907 = n45905 & n45906 ;
  assign n45908 = ~n45905 & ~n45906 ;
  assign n45909 = ~n45907 & ~n45908 ;
  assign n45910 = x115 & n12506 ;
  assign n45911 = x113 & n13131 ;
  assign n45912 = x114 & n12501 ;
  assign n45913 = ~n45911 & ~n45912 ;
  assign n45914 = ~n45910 & n45913 ;
  assign n45915 = n12509 & n17364 ;
  assign n45916 = n45914 & ~n45915 ;
  assign n45917 = x44 & ~n45916 ;
  assign n45918 = x44 & ~n45917 ;
  assign n45919 = ~n45916 & ~n45917 ;
  assign n45920 = ~n45918 & ~n45919 ;
  assign n45921 = n45909 & ~n45920 ;
  assign n45922 = ~n45909 & n45920 ;
  assign n45923 = ~n45786 & ~n45922 ;
  assign n45924 = ~n45921 & n45923 ;
  assign n45925 = ~n45786 & ~n45924 ;
  assign n45926 = ~n45921 & ~n45924 ;
  assign n45927 = ~n45922 & n45926 ;
  assign n45928 = ~n45925 & ~n45927 ;
  assign n45929 = x118 & n10905 ;
  assign n45930 = x116 & n11466 ;
  assign n45931 = x117 & n10900 ;
  assign n45932 = ~n45930 & ~n45931 ;
  assign n45933 = ~n45929 & n45932 ;
  assign n45934 = n10908 & n19395 ;
  assign n45935 = n45933 & ~n45934 ;
  assign n45936 = x41 & ~n45935 ;
  assign n45937 = x41 & ~n45936 ;
  assign n45938 = ~n45935 & ~n45936 ;
  assign n45939 = ~n45937 & ~n45938 ;
  assign n45940 = n45928 & n45939 ;
  assign n45941 = ~n45928 & ~n45939 ;
  assign n45942 = ~n45940 & ~n45941 ;
  assign n45943 = ~n45785 & n45942 ;
  assign n45944 = n45785 & ~n45942 ;
  assign n45945 = ~n45943 & ~n45944 ;
  assign n45946 = x121 & n9433 ;
  assign n45947 = x119 & n9915 ;
  assign n45948 = x120 & n9428 ;
  assign n45949 = ~n45947 & ~n45948 ;
  assign n45950 = ~n45946 & n45949 ;
  assign n45951 = n9436 & n21870 ;
  assign n45952 = n45950 & ~n45951 ;
  assign n45953 = x38 & ~n45952 ;
  assign n45954 = x38 & ~n45953 ;
  assign n45955 = ~n45952 & ~n45953 ;
  assign n45956 = ~n45954 & ~n45955 ;
  assign n45957 = n45945 & ~n45956 ;
  assign n45958 = n45945 & ~n45957 ;
  assign n45959 = ~n45956 & ~n45957 ;
  assign n45960 = ~n45958 & ~n45959 ;
  assign n45961 = ~n45506 & ~n45509 ;
  assign n45962 = n45960 & n45961 ;
  assign n45963 = ~n45960 & ~n45961 ;
  assign n45964 = ~n45962 & ~n45963 ;
  assign n45965 = x124 & n8006 ;
  assign n45966 = x122 & n8474 ;
  assign n45967 = x123 & n8001 ;
  assign n45968 = ~n45966 & ~n45967 ;
  assign n45969 = ~n45965 & n45968 ;
  assign n45970 = n8009 & n23796 ;
  assign n45971 = n45969 & ~n45970 ;
  assign n45972 = x35 & ~n45971 ;
  assign n45973 = x35 & ~n45972 ;
  assign n45974 = ~n45971 & ~n45972 ;
  assign n45975 = ~n45973 & ~n45974 ;
  assign n45976 = n45964 & ~n45975 ;
  assign n45977 = n45964 & ~n45976 ;
  assign n45978 = ~n45975 & ~n45976 ;
  assign n45979 = ~n45977 & ~n45978 ;
  assign n45980 = ~n45512 & ~n45526 ;
  assign n45981 = n45979 & n45980 ;
  assign n45982 = ~n45979 & ~n45980 ;
  assign n45983 = ~n45981 & ~n45982 ;
  assign n45984 = ~n45336 & ~n45531 ;
  assign n45985 = x127 & n6725 ;
  assign n45986 = x125 & n7129 ;
  assign n45987 = x126 & n6720 ;
  assign n45988 = ~n45986 & ~n45987 ;
  assign n45989 = ~n45985 & n45988 ;
  assign n45990 = n6728 & n26533 ;
  assign n45991 = n45989 & ~n45990 ;
  assign n45992 = x32 & ~n45991 ;
  assign n45993 = x32 & ~n45992 ;
  assign n45994 = ~n45991 & ~n45992 ;
  assign n45995 = ~n45993 & ~n45994 ;
  assign n45996 = ~n45984 & ~n45995 ;
  assign n45997 = ~n45984 & ~n45996 ;
  assign n45998 = ~n45995 & ~n45996 ;
  assign n45999 = ~n45997 & ~n45998 ;
  assign n46000 = ~n45983 & n45999 ;
  assign n46001 = n45983 & ~n45999 ;
  assign n46002 = ~n46000 & ~n46001 ;
  assign n46003 = ~n45784 & n46002 ;
  assign n46004 = n45784 & ~n46002 ;
  assign n46005 = ~n46003 & ~n46004 ;
  assign n46006 = ~n45783 & n46005 ;
  assign n46007 = n45783 & ~n46005 ;
  assign n46008 = ~n46006 & ~n46007 ;
  assign n46236 = n46008 & x221 ;
  assign n46009 = ~n45771 & ~n45775 ;
  assign n46010 = ~n45554 & ~n45768 ;
  assign n46011 = ~n45733 & ~n45737 ;
  assign n46012 = ~n45717 & ~n45731 ;
  assign n46013 = ~n45691 & ~n45694 ;
  assign n46014 = ~n45676 & ~n45687 ;
  assign n46015 = ~n45673 & ~n46014 ;
  assign n46016 = ~n45635 & ~n45646 ;
  assign n46017 = ~n45650 & ~n46016 ;
  assign n46018 = ~x93 & n27427 ;
  assign n46019 = ~x94 & ~n26217 ;
  assign n46020 = ~n46018 & ~n46019 ;
  assign n46021 = x29 & ~n46020 ;
  assign n46022 = ~x29 & n46020 ;
  assign n46023 = ~n46021 & ~n46022 ;
  assign n46024 = ~n45627 & n46023 ;
  assign n46025 = ~n45627 & ~n46024 ;
  assign n46026 = n46023 & ~n46024 ;
  assign n46027 = ~n46025 & ~n46026 ;
  assign n46028 = ~n45633 & ~n46027 ;
  assign n46029 = ~n45633 & ~n46028 ;
  assign n46030 = ~n46027 & ~n46028 ;
  assign n46031 = ~n46029 & ~n46030 ;
  assign n46032 = ~x97 & n24612 ;
  assign n46033 = ~x95 & n25390 ;
  assign n46034 = ~x96 & n24607 ;
  assign n46035 = ~n46033 & ~n46034 ;
  assign n46036 = ~n46032 & n46035 ;
  assign n46037 = n7949 & n24615 ;
  assign n46038 = n46036 & ~n46037 ;
  assign n46039 = ~x62 & ~n46038 ;
  assign n46040 = ~x62 & ~n46039 ;
  assign n46041 = ~n46038 & ~n46039 ;
  assign n46042 = ~n46040 & ~n46041 ;
  assign n46043 = ~n46031 & n46042 ;
  assign n46044 = n46031 & ~n46042 ;
  assign n46045 = ~n46043 & ~n46044 ;
  assign n46046 = ~x100 & n22325 ;
  assign n46047 = ~x98 & n23066 ;
  assign n46048 = ~x99 & n22320 ;
  assign n46049 = ~n46047 & ~n46048 ;
  assign n46050 = ~n46046 & n46049 ;
  assign n46051 = n9338 & n22328 ;
  assign n46052 = n46050 & ~n46051 ;
  assign n46053 = ~x59 & ~n46052 ;
  assign n46054 = ~x59 & ~n46053 ;
  assign n46055 = ~n46052 & ~n46053 ;
  assign n46056 = ~n46054 & ~n46055 ;
  assign n46057 = ~n46045 & ~n46056 ;
  assign n46058 = n46045 & n46056 ;
  assign n46059 = ~n46057 & ~n46058 ;
  assign n46060 = ~n46017 & n46059 ;
  assign n46061 = n46017 & ~n46059 ;
  assign n46062 = ~n46060 & ~n46061 ;
  assign n46063 = ~x103 & n20143 ;
  assign n46064 = ~x101 & n20854 ;
  assign n46065 = ~x102 & n20138 ;
  assign n46066 = ~n46064 & ~n46065 ;
  assign n46067 = ~n46063 & n46066 ;
  assign n46068 = n10833 & n20146 ;
  assign n46069 = n46067 & ~n46068 ;
  assign n46070 = ~x56 & ~n46069 ;
  assign n46071 = ~x56 & ~n46070 ;
  assign n46072 = ~n46069 & ~n46070 ;
  assign n46073 = ~n46071 & ~n46072 ;
  assign n46074 = n46062 & ~n46073 ;
  assign n46075 = n46062 & ~n46074 ;
  assign n46076 = ~n46073 & ~n46074 ;
  assign n46077 = ~n46075 & ~n46076 ;
  assign n46078 = ~n45653 & ~n45667 ;
  assign n46079 = n46077 & n46078 ;
  assign n46080 = ~n46077 & ~n46078 ;
  assign n46081 = ~n46079 & ~n46080 ;
  assign n46082 = ~x106 & n18025 ;
  assign n46083 = ~x104 & n18764 ;
  assign n46084 = ~x105 & n18020 ;
  assign n46085 = ~n46083 & ~n46084 ;
  assign n46086 = ~n46082 & n46085 ;
  assign n46087 = n12447 & n18028 ;
  assign n46088 = n46086 & ~n46087 ;
  assign n46089 = ~x53 & ~n46088 ;
  assign n46090 = ~x53 & ~n46089 ;
  assign n46091 = ~n46088 & ~n46089 ;
  assign n46092 = ~n46090 & ~n46091 ;
  assign n46093 = n46081 & ~n46092 ;
  assign n46094 = n46081 & ~n46093 ;
  assign n46095 = ~n46092 & ~n46093 ;
  assign n46096 = ~n46094 & ~n46095 ;
  assign n46097 = ~n46015 & n46096 ;
  assign n46098 = n46015 & ~n46096 ;
  assign n46099 = ~n46097 & ~n46098 ;
  assign n46100 = ~x109 & n16076 ;
  assign n46101 = ~x107 & n16756 ;
  assign n46102 = ~x108 & n16071 ;
  assign n46103 = ~n46101 & ~n46102 ;
  assign n46104 = ~n46100 & n46103 ;
  assign n46105 = n14177 & n16079 ;
  assign n46106 = n46104 & ~n46105 ;
  assign n46107 = ~x50 & ~n46106 ;
  assign n46108 = ~x50 & ~n46107 ;
  assign n46109 = ~n46106 & ~n46107 ;
  assign n46110 = ~n46108 & ~n46109 ;
  assign n46111 = ~n46099 & ~n46110 ;
  assign n46112 = n46099 & n46110 ;
  assign n46113 = ~n46111 & ~n46112 ;
  assign n46114 = n46013 & ~n46113 ;
  assign n46115 = ~n46013 & n46113 ;
  assign n46116 = ~n46114 & ~n46115 ;
  assign n46117 = ~x112 & n14233 ;
  assign n46118 = ~x110 & n14876 ;
  assign n46119 = ~x111 & n14228 ;
  assign n46120 = ~n46118 & ~n46119 ;
  assign n46121 = ~n46117 & n46120 ;
  assign n46122 = n14236 & n15744 ;
  assign n46123 = n46121 & ~n46122 ;
  assign n46124 = ~x47 & ~n46123 ;
  assign n46125 = ~x47 & ~n46124 ;
  assign n46126 = ~n46123 & ~n46124 ;
  assign n46127 = ~n46125 & ~n46126 ;
  assign n46128 = n46116 & ~n46127 ;
  assign n46129 = n46116 & ~n46128 ;
  assign n46130 = ~n46127 & ~n46128 ;
  assign n46131 = ~n46129 & ~n46130 ;
  assign n46132 = ~n45697 & ~n45711 ;
  assign n46133 = n46131 & n46132 ;
  assign n46134 = ~n46131 & ~n46132 ;
  assign n46135 = ~n46133 & ~n46134 ;
  assign n46136 = ~x115 & n12506 ;
  assign n46137 = ~x113 & n13131 ;
  assign n46138 = ~x114 & n12501 ;
  assign n46139 = ~n46137 & ~n46138 ;
  assign n46140 = ~n46136 & n46139 ;
  assign n46141 = n12509 & n17683 ;
  assign n46142 = n46140 & ~n46141 ;
  assign n46143 = ~x44 & ~n46142 ;
  assign n46144 = ~x44 & ~n46143 ;
  assign n46145 = ~n46142 & ~n46143 ;
  assign n46146 = ~n46144 & ~n46145 ;
  assign n46147 = n46135 & ~n46146 ;
  assign n46148 = ~n46135 & n46146 ;
  assign n46149 = ~n46012 & ~n46148 ;
  assign n46150 = ~n46147 & n46149 ;
  assign n46151 = ~n46012 & ~n46150 ;
  assign n46152 = ~n46147 & ~n46150 ;
  assign n46153 = ~n46148 & n46152 ;
  assign n46154 = ~n46151 & ~n46153 ;
  assign n46155 = ~x118 & n10905 ;
  assign n46156 = ~x116 & n11466 ;
  assign n46157 = ~x117 & n10900 ;
  assign n46158 = ~n46156 & ~n46157 ;
  assign n46159 = ~n46155 & n46158 ;
  assign n46160 = n10908 & n19736 ;
  assign n46161 = n46159 & ~n46160 ;
  assign n46162 = ~x41 & ~n46161 ;
  assign n46163 = ~x41 & ~n46162 ;
  assign n46164 = ~n46161 & ~n46162 ;
  assign n46165 = ~n46163 & ~n46164 ;
  assign n46166 = n46154 & n46165 ;
  assign n46167 = ~n46154 & ~n46165 ;
  assign n46168 = ~n46166 & ~n46167 ;
  assign n46169 = ~n46011 & n46168 ;
  assign n46170 = n46011 & ~n46168 ;
  assign n46171 = ~n46169 & ~n46170 ;
  assign n46172 = ~x121 & n9433 ;
  assign n46173 = ~x119 & n9915 ;
  assign n46174 = ~x120 & n9428 ;
  assign n46175 = ~n46173 & ~n46174 ;
  assign n46176 = ~n46172 & n46175 ;
  assign n46177 = n9436 & n22229 ;
  assign n46178 = n46176 & ~n46177 ;
  assign n46179 = ~x38 & ~n46178 ;
  assign n46180 = ~x38 & ~n46179 ;
  assign n46181 = ~n46178 & ~n46179 ;
  assign n46182 = ~n46180 & ~n46181 ;
  assign n46183 = n46171 & ~n46182 ;
  assign n46184 = n46171 & ~n46183 ;
  assign n46185 = ~n46182 & ~n46183 ;
  assign n46186 = ~n46184 & ~n46185 ;
  assign n46187 = ~n45741 & ~n45744 ;
  assign n46188 = n46186 & n46187 ;
  assign n46189 = ~n46186 & ~n46187 ;
  assign n46190 = ~n46188 & ~n46189 ;
  assign n46191 = ~x124 & n8006 ;
  assign n46192 = ~x122 & n8474 ;
  assign n46193 = ~x123 & n8001 ;
  assign n46194 = ~n46192 & ~n46193 ;
  assign n46195 = ~n46191 & n46194 ;
  assign n46196 = n8009 & n24176 ;
  assign n46197 = n46195 & ~n46196 ;
  assign n46198 = ~x35 & ~n46197 ;
  assign n46199 = ~x35 & ~n46198 ;
  assign n46200 = ~n46197 & ~n46198 ;
  assign n46201 = ~n46199 & ~n46200 ;
  assign n46202 = n46190 & ~n46201 ;
  assign n46203 = n46190 & ~n46202 ;
  assign n46204 = ~n46201 & ~n46202 ;
  assign n46205 = ~n46203 & ~n46204 ;
  assign n46206 = ~n45747 & ~n45761 ;
  assign n46207 = n46205 & n46206 ;
  assign n46208 = ~n46205 & ~n46206 ;
  assign n46209 = ~n46207 & ~n46208 ;
  assign n46210 = ~n45571 & ~n45766 ;
  assign n46211 = ~x127 & n6725 ;
  assign n46212 = ~x125 & n7129 ;
  assign n46213 = ~x126 & n6720 ;
  assign n46214 = ~n46212 & ~n46213 ;
  assign n46215 = ~n46211 & n46214 ;
  assign n46216 = n6728 & n26932 ;
  assign n46217 = n46215 & ~n46216 ;
  assign n46218 = ~x32 & ~n46217 ;
  assign n46219 = ~x32 & ~n46218 ;
  assign n46220 = ~n46217 & ~n46218 ;
  assign n46221 = ~n46219 & ~n46220 ;
  assign n46222 = ~n46210 & ~n46221 ;
  assign n46223 = ~n46210 & ~n46222 ;
  assign n46224 = ~n46221 & ~n46222 ;
  assign n46225 = ~n46223 & ~n46224 ;
  assign n46226 = ~n46209 & n46225 ;
  assign n46227 = n46209 & ~n46225 ;
  assign n46228 = ~n46226 & ~n46227 ;
  assign n46229 = ~n46010 & n46228 ;
  assign n46230 = n46010 & ~n46228 ;
  assign n46231 = ~n46229 & ~n46230 ;
  assign n46232 = ~n46009 & n46231 ;
  assign n46233 = n46009 & ~n46231 ;
  assign n46234 = ~n46232 & ~n46233 ;
  assign n46237 = ~n46234 & ~x221 ;
  assign n46238 = ~n46236 & ~n46237 ;
  assign n46239 = ~n45976 & ~n45982 ;
  assign n46240 = x126 & n7129 ;
  assign n46241 = x127 & n6720 ;
  assign n46242 = ~n46240 & ~n46241 ;
  assign n46243 = ~n6728 & n46242 ;
  assign n46244 = n26965 & n46242 ;
  assign n46245 = ~n46243 & ~n46244 ;
  assign n46246 = x32 & ~n46245 ;
  assign n46247 = ~x32 & n46245 ;
  assign n46248 = ~n46246 & ~n46247 ;
  assign n46249 = ~n46239 & ~n46248 ;
  assign n46250 = n46239 & n46248 ;
  assign n46251 = ~n46249 & ~n46250 ;
  assign n46252 = ~n45941 & ~n45943 ;
  assign n46253 = ~n45848 & ~n45854 ;
  assign n46254 = x104 & n20143 ;
  assign n46255 = x102 & n20854 ;
  assign n46256 = x103 & n20138 ;
  assign n46257 = ~n46255 & ~n46256 ;
  assign n46258 = ~n46254 & n46257 ;
  assign n46259 = n11116 & n20146 ;
  assign n46260 = n46258 & ~n46259 ;
  assign n46261 = x56 & ~n46260 ;
  assign n46262 = x56 & ~n46261 ;
  assign n46263 = ~n46260 & ~n46261 ;
  assign n46264 = ~n46262 & ~n46263 ;
  assign n46265 = ~n45831 & ~n45834 ;
  assign n46266 = x101 & n22325 ;
  assign n46267 = x99 & n23066 ;
  assign n46268 = x100 & n22320 ;
  assign n46269 = ~n46267 & ~n46268 ;
  assign n46270 = ~n46266 & n46269 ;
  assign n46271 = n9601 & n22328 ;
  assign n46272 = n46270 & ~n46271 ;
  assign n46273 = x59 & ~n46272 ;
  assign n46274 = x59 & ~n46273 ;
  assign n46275 = ~n46272 & ~n46273 ;
  assign n46276 = ~n46274 & ~n46275 ;
  assign n46277 = ~n45805 & ~n45816 ;
  assign n46278 = ~n45802 & ~n46277 ;
  assign n46279 = x94 & n27024 ;
  assign n46280 = x95 & ~n26217 ;
  assign n46281 = ~n46279 & ~n46280 ;
  assign n46282 = ~n45795 & ~n45798 ;
  assign n46283 = ~n46281 & n46282 ;
  assign n46284 = n46281 & ~n46282 ;
  assign n46285 = ~n46283 & ~n46284 ;
  assign n46286 = x98 & n24612 ;
  assign n46287 = x96 & n25390 ;
  assign n46288 = x97 & n24607 ;
  assign n46289 = ~n46287 & ~n46288 ;
  assign n46290 = ~n46286 & n46289 ;
  assign n46291 = n8196 & n24615 ;
  assign n46292 = n46290 & ~n46291 ;
  assign n46293 = x62 & ~n46292 ;
  assign n46294 = x62 & ~n46293 ;
  assign n46295 = ~n46292 & ~n46293 ;
  assign n46296 = ~n46294 & ~n46295 ;
  assign n46297 = ~n46285 & n46296 ;
  assign n46298 = n46285 & ~n46296 ;
  assign n46299 = ~n46297 & ~n46298 ;
  assign n46300 = ~n46278 & n46299 ;
  assign n46301 = ~n46278 & ~n46300 ;
  assign n46302 = n46299 & ~n46300 ;
  assign n46303 = ~n46301 & ~n46302 ;
  assign n46304 = ~n46276 & ~n46303 ;
  assign n46305 = n46276 & ~n46302 ;
  assign n46306 = ~n46301 & n46305 ;
  assign n46307 = ~n46304 & ~n46306 ;
  assign n46308 = ~n46265 & n46307 ;
  assign n46309 = ~n46265 & ~n46308 ;
  assign n46310 = n46307 & ~n46308 ;
  assign n46311 = ~n46309 & ~n46310 ;
  assign n46312 = ~n46264 & ~n46311 ;
  assign n46313 = n46264 & ~n46310 ;
  assign n46314 = ~n46309 & n46313 ;
  assign n46315 = ~n46312 & ~n46314 ;
  assign n46316 = ~n46253 & n46315 ;
  assign n46317 = n46253 & ~n46315 ;
  assign n46318 = ~n46316 & ~n46317 ;
  assign n46319 = x107 & n18025 ;
  assign n46320 = x105 & n18764 ;
  assign n46321 = x106 & n18020 ;
  assign n46322 = ~n46320 & ~n46321 ;
  assign n46323 = ~n46319 & n46322 ;
  assign n46324 = n12749 & n18028 ;
  assign n46325 = n46323 & ~n46324 ;
  assign n46326 = x53 & ~n46325 ;
  assign n46327 = x53 & ~n46326 ;
  assign n46328 = ~n46325 & ~n46326 ;
  assign n46329 = ~n46327 & ~n46328 ;
  assign n46330 = n46318 & ~n46329 ;
  assign n46331 = n46318 & ~n46330 ;
  assign n46332 = ~n46329 & ~n46330 ;
  assign n46333 = ~n46331 & ~n46332 ;
  assign n46334 = ~n45789 & ~n45870 ;
  assign n46335 = ~n45867 & ~n46334 ;
  assign n46336 = n46333 & n46335 ;
  assign n46337 = ~n46333 & ~n46335 ;
  assign n46338 = ~n46336 & ~n46337 ;
  assign n46339 = x110 & n16076 ;
  assign n46340 = x108 & n16756 ;
  assign n46341 = x109 & n16071 ;
  assign n46342 = ~n46340 & ~n46341 ;
  assign n46343 = ~n46339 & n46342 ;
  assign n46344 = n14497 & n16079 ;
  assign n46345 = n46343 & ~n46344 ;
  assign n46346 = x50 & ~n46345 ;
  assign n46347 = x50 & ~n46346 ;
  assign n46348 = ~n46345 & ~n46346 ;
  assign n46349 = ~n46347 & ~n46348 ;
  assign n46350 = n46338 & ~n46349 ;
  assign n46351 = n46338 & ~n46350 ;
  assign n46352 = ~n46349 & ~n46350 ;
  assign n46353 = ~n46351 & ~n46352 ;
  assign n46354 = ~n45885 & ~n45889 ;
  assign n46355 = n46353 & n46354 ;
  assign n46356 = ~n46353 & ~n46354 ;
  assign n46357 = ~n46355 & ~n46356 ;
  assign n46358 = x113 & n14233 ;
  assign n46359 = x111 & n14876 ;
  assign n46360 = x112 & n14228 ;
  assign n46361 = ~n46359 & ~n46360 ;
  assign n46362 = ~n46358 & n46361 ;
  assign n46363 = n14236 & n16361 ;
  assign n46364 = n46362 & ~n46363 ;
  assign n46365 = x47 & ~n46364 ;
  assign n46366 = x47 & ~n46365 ;
  assign n46367 = ~n46364 & ~n46365 ;
  assign n46368 = ~n46366 & ~n46367 ;
  assign n46369 = n46357 & ~n46368 ;
  assign n46370 = n46357 & ~n46369 ;
  assign n46371 = ~n46368 & ~n46369 ;
  assign n46372 = ~n46370 & ~n46371 ;
  assign n46373 = ~n45902 & ~n45908 ;
  assign n46374 = n46372 & n46373 ;
  assign n46375 = ~n46372 & ~n46373 ;
  assign n46376 = ~n46374 & ~n46375 ;
  assign n46377 = x116 & n12506 ;
  assign n46378 = x114 & n13131 ;
  assign n46379 = x115 & n12501 ;
  assign n46380 = ~n46378 & ~n46379 ;
  assign n46381 = ~n46377 & n46380 ;
  assign n46382 = n12509 & n18336 ;
  assign n46383 = n46381 & ~n46382 ;
  assign n46384 = x44 & ~n46383 ;
  assign n46385 = x44 & ~n46384 ;
  assign n46386 = ~n46383 & ~n46384 ;
  assign n46387 = ~n46385 & ~n46386 ;
  assign n46388 = n46376 & ~n46387 ;
  assign n46389 = n46376 & ~n46388 ;
  assign n46390 = ~n46387 & ~n46388 ;
  assign n46391 = ~n46389 & ~n46390 ;
  assign n46392 = ~n45926 & n46391 ;
  assign n46393 = n45926 & ~n46391 ;
  assign n46394 = ~n46392 & ~n46393 ;
  assign n46395 = x119 & n10905 ;
  assign n46396 = x117 & n11466 ;
  assign n46397 = x118 & n10900 ;
  assign n46398 = ~n46396 & ~n46397 ;
  assign n46399 = ~n46395 & n46398 ;
  assign n46400 = n10908 & n20423 ;
  assign n46401 = n46399 & ~n46400 ;
  assign n46402 = x41 & ~n46401 ;
  assign n46403 = x41 & ~n46402 ;
  assign n46404 = ~n46401 & ~n46402 ;
  assign n46405 = ~n46403 & ~n46404 ;
  assign n46406 = ~n46394 & ~n46405 ;
  assign n46407 = n46394 & n46405 ;
  assign n46408 = ~n46406 & ~n46407 ;
  assign n46409 = ~n46252 & n46408 ;
  assign n46410 = n46252 & ~n46408 ;
  assign n46411 = ~n46409 & ~n46410 ;
  assign n46412 = x122 & n9433 ;
  assign n46413 = x120 & n9915 ;
  assign n46414 = x121 & n9428 ;
  assign n46415 = ~n46413 & ~n46414 ;
  assign n46416 = ~n46412 & n46415 ;
  assign n46417 = n9436 & n22622 ;
  assign n46418 = n46416 & ~n46417 ;
  assign n46419 = x38 & ~n46418 ;
  assign n46420 = x38 & ~n46419 ;
  assign n46421 = ~n46418 & ~n46419 ;
  assign n46422 = ~n46420 & ~n46421 ;
  assign n46423 = n46411 & ~n46422 ;
  assign n46424 = n46411 & ~n46423 ;
  assign n46425 = ~n46422 & ~n46423 ;
  assign n46426 = ~n46424 & ~n46425 ;
  assign n46427 = ~n45957 & ~n45963 ;
  assign n46428 = n46426 & n46427 ;
  assign n46429 = ~n46426 & ~n46427 ;
  assign n46430 = ~n46428 & ~n46429 ;
  assign n46431 = x125 & n8006 ;
  assign n46432 = x123 & n8474 ;
  assign n46433 = x124 & n8001 ;
  assign n46434 = ~n46432 & ~n46433 ;
  assign n46435 = ~n46431 & n46434 ;
  assign n46436 = n8009 & n24935 ;
  assign n46437 = n46435 & ~n46436 ;
  assign n46438 = x35 & ~n46437 ;
  assign n46439 = x35 & ~n46438 ;
  assign n46440 = ~n46437 & ~n46438 ;
  assign n46441 = ~n46439 & ~n46440 ;
  assign n46442 = n46430 & ~n46441 ;
  assign n46443 = ~n46430 & n46441 ;
  assign n46444 = n46251 & ~n46443 ;
  assign n46445 = ~n46442 & n46444 ;
  assign n46446 = n46251 & ~n46445 ;
  assign n46447 = ~n46443 & ~n46445 ;
  assign n46448 = ~n46442 & n46447 ;
  assign n46449 = ~n46446 & ~n46448 ;
  assign n46450 = ~n45996 & ~n46001 ;
  assign n46451 = ~n46449 & ~n46450 ;
  assign n46452 = ~n46449 & ~n46451 ;
  assign n46453 = ~n46450 & ~n46451 ;
  assign n46454 = ~n46452 & ~n46453 ;
  assign n46455 = ~n46003 & ~n46006 ;
  assign n46456 = ~n46454 & ~n46455 ;
  assign n46457 = n46454 & n46455 ;
  assign n46458 = ~n46456 & ~n46457 ;
  assign n46680 = n46458 & x222 ;
  assign n46459 = ~n46202 & ~n46208 ;
  assign n46460 = ~x126 & n7129 ;
  assign n46461 = ~x127 & n6720 ;
  assign n46462 = ~n46460 & ~n46461 ;
  assign n46463 = ~n6728 & n46462 ;
  assign n46464 = n27368 & n46462 ;
  assign n46465 = ~n46463 & ~n46464 ;
  assign n46466 = ~x32 & ~n46465 ;
  assign n46467 = x32 & n46465 ;
  assign n46468 = ~n46466 & ~n46467 ;
  assign n46469 = ~n46459 & ~n46468 ;
  assign n46470 = n46459 & n46468 ;
  assign n46471 = ~n46469 & ~n46470 ;
  assign n46472 = ~n46167 & ~n46169 ;
  assign n46473 = ~n46074 & ~n46080 ;
  assign n46474 = ~x104 & n20143 ;
  assign n46475 = ~x102 & n20854 ;
  assign n46476 = ~x103 & n20138 ;
  assign n46477 = ~n46475 & ~n46476 ;
  assign n46478 = ~n46474 & n46477 ;
  assign n46479 = n11380 & n20146 ;
  assign n46480 = n46478 & ~n46479 ;
  assign n46481 = ~x56 & ~n46480 ;
  assign n46482 = ~x56 & ~n46481 ;
  assign n46483 = ~n46480 & ~n46481 ;
  assign n46484 = ~n46482 & ~n46483 ;
  assign n46485 = ~n46057 & ~n46060 ;
  assign n46486 = ~x101 & n22325 ;
  assign n46487 = ~x99 & n23066 ;
  assign n46488 = ~x100 & n22320 ;
  assign n46489 = ~n46487 & ~n46488 ;
  assign n46490 = ~n46486 & n46489 ;
  assign n46491 = n9844 & n22328 ;
  assign n46492 = n46490 & ~n46491 ;
  assign n46493 = ~x59 & ~n46492 ;
  assign n46494 = ~x59 & ~n46493 ;
  assign n46495 = ~n46492 & ~n46493 ;
  assign n46496 = ~n46494 & ~n46495 ;
  assign n46497 = ~n46031 & ~n46042 ;
  assign n46498 = ~n46028 & ~n46497 ;
  assign n46499 = ~x94 & n27427 ;
  assign n46500 = ~x95 & ~n26217 ;
  assign n46501 = ~n46499 & ~n46500 ;
  assign n46502 = ~n46021 & ~n46024 ;
  assign n46503 = ~n46501 & n46502 ;
  assign n46504 = n46501 & ~n46502 ;
  assign n46505 = ~n46503 & ~n46504 ;
  assign n46506 = ~x98 & n24612 ;
  assign n46507 = ~x96 & n25390 ;
  assign n46508 = ~x97 & n24607 ;
  assign n46509 = ~n46507 & ~n46508 ;
  assign n46510 = ~n46506 & n46509 ;
  assign n46511 = n8426 & n24615 ;
  assign n46512 = n46510 & ~n46511 ;
  assign n46513 = ~x62 & ~n46512 ;
  assign n46514 = ~x62 & ~n46513 ;
  assign n46515 = ~n46512 & ~n46513 ;
  assign n46516 = ~n46514 & ~n46515 ;
  assign n46517 = ~n46505 & n46516 ;
  assign n46518 = n46505 & ~n46516 ;
  assign n46519 = ~n46517 & ~n46518 ;
  assign n46520 = ~n46498 & n46519 ;
  assign n46521 = ~n46498 & ~n46520 ;
  assign n46522 = n46519 & ~n46520 ;
  assign n46523 = ~n46521 & ~n46522 ;
  assign n46524 = ~n46496 & ~n46523 ;
  assign n46525 = n46496 & ~n46522 ;
  assign n46526 = ~n46521 & n46525 ;
  assign n46527 = ~n46524 & ~n46526 ;
  assign n46528 = ~n46485 & n46527 ;
  assign n46529 = ~n46485 & ~n46528 ;
  assign n46530 = n46527 & ~n46528 ;
  assign n46531 = ~n46529 & ~n46530 ;
  assign n46532 = ~n46484 & ~n46531 ;
  assign n46533 = n46484 & ~n46530 ;
  assign n46534 = ~n46529 & n46533 ;
  assign n46535 = ~n46532 & ~n46534 ;
  assign n46536 = ~n46473 & n46535 ;
  assign n46537 = n46473 & ~n46535 ;
  assign n46538 = ~n46536 & ~n46537 ;
  assign n46539 = ~x107 & n18025 ;
  assign n46540 = ~x105 & n18764 ;
  assign n46541 = ~x106 & n18020 ;
  assign n46542 = ~n46540 & ~n46541 ;
  assign n46543 = ~n46539 & n46542 ;
  assign n46544 = n13034 & n18028 ;
  assign n46545 = n46543 & ~n46544 ;
  assign n46546 = ~x53 & ~n46545 ;
  assign n46547 = ~x53 & ~n46546 ;
  assign n46548 = ~n46545 & ~n46546 ;
  assign n46549 = ~n46547 & ~n46548 ;
  assign n46550 = n46538 & ~n46549 ;
  assign n46551 = n46538 & ~n46550 ;
  assign n46552 = ~n46549 & ~n46550 ;
  assign n46553 = ~n46551 & ~n46552 ;
  assign n46554 = ~n46015 & ~n46096 ;
  assign n46555 = ~n46093 & ~n46554 ;
  assign n46556 = n46553 & n46555 ;
  assign n46557 = ~n46553 & ~n46555 ;
  assign n46558 = ~n46556 & ~n46557 ;
  assign n46559 = ~x110 & n16076 ;
  assign n46560 = ~x108 & n16756 ;
  assign n46561 = ~x109 & n16071 ;
  assign n46562 = ~n46560 & ~n46561 ;
  assign n46563 = ~n46559 & n46562 ;
  assign n46564 = n14802 & n16079 ;
  assign n46565 = n46563 & ~n46564 ;
  assign n46566 = ~x50 & ~n46565 ;
  assign n46567 = ~x50 & ~n46566 ;
  assign n46568 = ~n46565 & ~n46566 ;
  assign n46569 = ~n46567 & ~n46568 ;
  assign n46570 = n46558 & ~n46569 ;
  assign n46571 = n46558 & ~n46570 ;
  assign n46572 = ~n46569 & ~n46570 ;
  assign n46573 = ~n46571 & ~n46572 ;
  assign n46574 = ~n46111 & ~n46115 ;
  assign n46575 = n46573 & n46574 ;
  assign n46576 = ~n46573 & ~n46574 ;
  assign n46577 = ~n46575 & ~n46576 ;
  assign n46578 = ~x113 & n14233 ;
  assign n46579 = ~x111 & n14876 ;
  assign n46580 = ~x112 & n14228 ;
  assign n46581 = ~n46579 & ~n46580 ;
  assign n46582 = ~n46578 & n46581 ;
  assign n46583 = n14236 & n16684 ;
  assign n46584 = n46582 & ~n46583 ;
  assign n46585 = ~x47 & ~n46584 ;
  assign n46586 = ~x47 & ~n46585 ;
  assign n46587 = ~n46584 & ~n46585 ;
  assign n46588 = ~n46586 & ~n46587 ;
  assign n46589 = n46577 & ~n46588 ;
  assign n46590 = n46577 & ~n46589 ;
  assign n46591 = ~n46588 & ~n46589 ;
  assign n46592 = ~n46590 & ~n46591 ;
  assign n46593 = ~n46128 & ~n46134 ;
  assign n46594 = n46592 & n46593 ;
  assign n46595 = ~n46592 & ~n46593 ;
  assign n46596 = ~n46594 & ~n46595 ;
  assign n46597 = ~x116 & n12506 ;
  assign n46598 = ~x114 & n13131 ;
  assign n46599 = ~x115 & n12501 ;
  assign n46600 = ~n46598 & ~n46599 ;
  assign n46601 = ~n46597 & n46600 ;
  assign n46602 = n12509 & n18678 ;
  assign n46603 = n46601 & ~n46602 ;
  assign n46604 = ~x44 & ~n46603 ;
  assign n46605 = ~x44 & ~n46604 ;
  assign n46606 = ~n46603 & ~n46604 ;
  assign n46607 = ~n46605 & ~n46606 ;
  assign n46608 = n46596 & ~n46607 ;
  assign n46609 = n46596 & ~n46608 ;
  assign n46610 = ~n46607 & ~n46608 ;
  assign n46611 = ~n46609 & ~n46610 ;
  assign n46612 = ~n46152 & n46611 ;
  assign n46613 = n46152 & ~n46611 ;
  assign n46614 = ~n46612 & ~n46613 ;
  assign n46615 = ~x119 & n10905 ;
  assign n46616 = ~x117 & n11466 ;
  assign n46617 = ~x118 & n10900 ;
  assign n46618 = ~n46616 & ~n46617 ;
  assign n46619 = ~n46615 & n46618 ;
  assign n46620 = n10908 & n20778 ;
  assign n46621 = n46619 & ~n46620 ;
  assign n46622 = ~x41 & ~n46621 ;
  assign n46623 = ~x41 & ~n46622 ;
  assign n46624 = ~n46621 & ~n46622 ;
  assign n46625 = ~n46623 & ~n46624 ;
  assign n46626 = ~n46614 & ~n46625 ;
  assign n46627 = n46614 & n46625 ;
  assign n46628 = ~n46626 & ~n46627 ;
  assign n46629 = ~n46472 & n46628 ;
  assign n46630 = n46472 & ~n46628 ;
  assign n46631 = ~n46629 & ~n46630 ;
  assign n46632 = ~x122 & n9433 ;
  assign n46633 = ~x120 & n9915 ;
  assign n46634 = ~x121 & n9428 ;
  assign n46635 = ~n46633 & ~n46634 ;
  assign n46636 = ~n46632 & n46635 ;
  assign n46637 = n9436 & n22998 ;
  assign n46638 = n46636 & ~n46637 ;
  assign n46639 = ~x38 & ~n46638 ;
  assign n46640 = ~x38 & ~n46639 ;
  assign n46641 = ~n46638 & ~n46639 ;
  assign n46642 = ~n46640 & ~n46641 ;
  assign n46643 = n46631 & ~n46642 ;
  assign n46644 = n46631 & ~n46643 ;
  assign n46645 = ~n46642 & ~n46643 ;
  assign n46646 = ~n46644 & ~n46645 ;
  assign n46647 = ~n46183 & ~n46189 ;
  assign n46648 = n46646 & n46647 ;
  assign n46649 = ~n46646 & ~n46647 ;
  assign n46650 = ~n46648 & ~n46649 ;
  assign n46651 = ~x125 & n8006 ;
  assign n46652 = ~x123 & n8474 ;
  assign n46653 = ~x124 & n8001 ;
  assign n46654 = ~n46652 & ~n46653 ;
  assign n46655 = ~n46651 & n46654 ;
  assign n46656 = n8009 & n25330 ;
  assign n46657 = n46655 & ~n46656 ;
  assign n46658 = ~x35 & ~n46657 ;
  assign n46659 = ~x35 & ~n46658 ;
  assign n46660 = ~n46657 & ~n46658 ;
  assign n46661 = ~n46659 & ~n46660 ;
  assign n46662 = n46650 & ~n46661 ;
  assign n46663 = ~n46650 & n46661 ;
  assign n46664 = n46471 & ~n46663 ;
  assign n46665 = ~n46662 & n46664 ;
  assign n46666 = n46471 & ~n46665 ;
  assign n46667 = ~n46663 & ~n46665 ;
  assign n46668 = ~n46662 & n46667 ;
  assign n46669 = ~n46666 & ~n46668 ;
  assign n46670 = ~n46222 & ~n46227 ;
  assign n46671 = ~n46669 & ~n46670 ;
  assign n46672 = ~n46669 & ~n46671 ;
  assign n46673 = ~n46670 & ~n46671 ;
  assign n46674 = ~n46672 & ~n46673 ;
  assign n46675 = ~n46229 & ~n46232 ;
  assign n46676 = ~n46674 & ~n46675 ;
  assign n46677 = n46674 & n46675 ;
  assign n46678 = ~n46676 & ~n46677 ;
  assign n46681 = ~n46678 & ~x222 ;
  assign n46682 = ~n46680 & ~n46681 ;
  assign n46683 = ~n46451 & ~n46456 ;
  assign n46684 = ~n46249 & ~n46445 ;
  assign n46685 = ~n46429 & ~n46442 ;
  assign n46686 = x127 & n7129 ;
  assign n46687 = n6728 & n26962 ;
  assign n46688 = ~n46686 & ~n46687 ;
  assign n46689 = x32 & ~n46688 ;
  assign n46690 = x32 & ~n46689 ;
  assign n46691 = ~n46688 & ~n46689 ;
  assign n46692 = ~n46690 & ~n46691 ;
  assign n46693 = ~n46685 & ~n46692 ;
  assign n46694 = ~n46685 & ~n46693 ;
  assign n46695 = ~n46692 & ~n46693 ;
  assign n46696 = ~n46694 & ~n46695 ;
  assign n46697 = ~n45926 & ~n46391 ;
  assign n46698 = ~n46406 & ~n46697 ;
  assign n46699 = x120 & n10905 ;
  assign n46700 = x118 & n11466 ;
  assign n46701 = x119 & n10900 ;
  assign n46702 = ~n46700 & ~n46701 ;
  assign n46703 = ~n46699 & n46702 ;
  assign n46704 = n10908 & n21143 ;
  assign n46705 = n46703 & ~n46704 ;
  assign n46706 = x41 & ~n46705 ;
  assign n46707 = x41 & ~n46706 ;
  assign n46708 = ~n46705 & ~n46706 ;
  assign n46709 = ~n46707 & ~n46708 ;
  assign n46710 = ~n46375 & ~n46388 ;
  assign n46711 = x117 & n12506 ;
  assign n46712 = x115 & n13131 ;
  assign n46713 = x116 & n12501 ;
  assign n46714 = ~n46712 & ~n46713 ;
  assign n46715 = ~n46711 & n46714 ;
  assign n46716 = n12509 & n19026 ;
  assign n46717 = n46715 & ~n46716 ;
  assign n46718 = x44 & ~n46717 ;
  assign n46719 = x44 & ~n46718 ;
  assign n46720 = ~n46717 & ~n46718 ;
  assign n46721 = ~n46719 & ~n46720 ;
  assign n46722 = ~n46356 & ~n46369 ;
  assign n46723 = ~n46316 & ~n46330 ;
  assign n46724 = x108 & n18025 ;
  assign n46725 = x106 & n18764 ;
  assign n46726 = x107 & n18020 ;
  assign n46727 = ~n46725 & ~n46726 ;
  assign n46728 = ~n46724 & n46727 ;
  assign n46729 = n13323 & n18028 ;
  assign n46730 = n46728 & ~n46729 ;
  assign n46731 = x53 & ~n46730 ;
  assign n46732 = x53 & ~n46731 ;
  assign n46733 = ~n46730 & ~n46731 ;
  assign n46734 = ~n46732 & ~n46733 ;
  assign n46735 = ~n46308 & ~n46312 ;
  assign n46736 = x105 & n20143 ;
  assign n46737 = x103 & n20854 ;
  assign n46738 = x104 & n20138 ;
  assign n46739 = ~n46737 & ~n46738 ;
  assign n46740 = ~n46736 & n46739 ;
  assign n46741 = n11648 & n20146 ;
  assign n46742 = n46740 & ~n46741 ;
  assign n46743 = x56 & ~n46742 ;
  assign n46744 = x56 & ~n46743 ;
  assign n46745 = ~n46742 & ~n46743 ;
  assign n46746 = ~n46744 & ~n46745 ;
  assign n46747 = ~n46300 & ~n46304 ;
  assign n46748 = ~n46284 & ~n46298 ;
  assign n46749 = x95 & n27024 ;
  assign n46750 = x96 & ~n26217 ;
  assign n46751 = ~n46749 & ~n46750 ;
  assign n46752 = ~n46281 & n46751 ;
  assign n46753 = n46281 & ~n46751 ;
  assign n46754 = ~n46748 & ~n46753 ;
  assign n46755 = ~n46752 & n46754 ;
  assign n46756 = ~n46748 & ~n46755 ;
  assign n46757 = ~n46752 & ~n46755 ;
  assign n46758 = ~n46753 & n46757 ;
  assign n46759 = ~n46756 & ~n46758 ;
  assign n46760 = x99 & n24612 ;
  assign n46761 = x97 & n25390 ;
  assign n46762 = x98 & n24607 ;
  assign n46763 = ~n46761 & ~n46762 ;
  assign n46764 = ~n46760 & n46763 ;
  assign n46765 = n8660 & n24615 ;
  assign n46766 = n46764 & ~n46765 ;
  assign n46767 = x62 & ~n46766 ;
  assign n46768 = x62 & ~n46767 ;
  assign n46769 = ~n46766 & ~n46767 ;
  assign n46770 = ~n46768 & ~n46769 ;
  assign n46771 = ~n46759 & ~n46770 ;
  assign n46772 = ~n46759 & ~n46771 ;
  assign n46773 = ~n46770 & ~n46771 ;
  assign n46774 = ~n46772 & ~n46773 ;
  assign n46775 = x102 & n22325 ;
  assign n46776 = x100 & n23066 ;
  assign n46777 = x101 & n22320 ;
  assign n46778 = ~n46776 & ~n46777 ;
  assign n46779 = ~n46775 & n46778 ;
  assign n46780 = n10092 & n22328 ;
  assign n46781 = n46779 & ~n46780 ;
  assign n46782 = x59 & ~n46781 ;
  assign n46783 = x59 & ~n46782 ;
  assign n46784 = ~n46781 & ~n46782 ;
  assign n46785 = ~n46783 & ~n46784 ;
  assign n46786 = ~n46774 & n46785 ;
  assign n46787 = n46774 & ~n46785 ;
  assign n46788 = ~n46786 & ~n46787 ;
  assign n46789 = ~n46747 & ~n46788 ;
  assign n46790 = n46747 & n46788 ;
  assign n46791 = ~n46789 & ~n46790 ;
  assign n46792 = ~n46746 & n46791 ;
  assign n46793 = n46746 & ~n46791 ;
  assign n46794 = ~n46792 & ~n46793 ;
  assign n46795 = ~n46735 & n46794 ;
  assign n46796 = n46735 & ~n46794 ;
  assign n46797 = ~n46795 & ~n46796 ;
  assign n46798 = ~n46734 & n46797 ;
  assign n46799 = n46734 & ~n46797 ;
  assign n46800 = ~n46798 & ~n46799 ;
  assign n46801 = ~n46723 & n46800 ;
  assign n46802 = n46723 & ~n46800 ;
  assign n46803 = ~n46801 & ~n46802 ;
  assign n46804 = x111 & n16076 ;
  assign n46805 = x109 & n16756 ;
  assign n46806 = x110 & n16071 ;
  assign n46807 = ~n46805 & ~n46806 ;
  assign n46808 = ~n46804 & n46807 ;
  assign n46809 = n15111 & n16079 ;
  assign n46810 = n46808 & ~n46809 ;
  assign n46811 = x50 & ~n46810 ;
  assign n46812 = x50 & ~n46811 ;
  assign n46813 = ~n46810 & ~n46811 ;
  assign n46814 = ~n46812 & ~n46813 ;
  assign n46815 = n46803 & ~n46814 ;
  assign n46816 = n46803 & ~n46815 ;
  assign n46817 = ~n46814 & ~n46815 ;
  assign n46818 = ~n46816 & ~n46817 ;
  assign n46819 = ~n46337 & ~n46350 ;
  assign n46820 = n46818 & n46819 ;
  assign n46821 = ~n46818 & ~n46819 ;
  assign n46822 = ~n46820 & ~n46821 ;
  assign n46823 = x114 & n14233 ;
  assign n46824 = x112 & n14876 ;
  assign n46825 = x113 & n14228 ;
  assign n46826 = ~n46824 & ~n46825 ;
  assign n46827 = ~n46823 & n46826 ;
  assign n46828 = n14236 & n17012 ;
  assign n46829 = n46827 & ~n46828 ;
  assign n46830 = x47 & ~n46829 ;
  assign n46831 = x47 & ~n46830 ;
  assign n46832 = ~n46829 & ~n46830 ;
  assign n46833 = ~n46831 & ~n46832 ;
  assign n46834 = ~n46822 & n46833 ;
  assign n46835 = n46822 & ~n46833 ;
  assign n46836 = ~n46834 & ~n46835 ;
  assign n46837 = ~n46722 & n46836 ;
  assign n46838 = ~n46722 & ~n46837 ;
  assign n46839 = n46836 & ~n46837 ;
  assign n46840 = ~n46838 & ~n46839 ;
  assign n46841 = ~n46721 & ~n46840 ;
  assign n46842 = n46721 & ~n46839 ;
  assign n46843 = ~n46838 & n46842 ;
  assign n46844 = ~n46841 & ~n46843 ;
  assign n46845 = ~n46710 & n46844 ;
  assign n46846 = n46710 & ~n46844 ;
  assign n46847 = ~n46845 & ~n46846 ;
  assign n46848 = ~n46709 & n46847 ;
  assign n46849 = n46709 & ~n46847 ;
  assign n46850 = ~n46848 & ~n46849 ;
  assign n46851 = ~n46698 & n46850 ;
  assign n46852 = n46698 & ~n46850 ;
  assign n46853 = ~n46851 & ~n46852 ;
  assign n46854 = x123 & n9433 ;
  assign n46855 = x121 & n9915 ;
  assign n46856 = x122 & n9428 ;
  assign n46857 = ~n46855 & ~n46856 ;
  assign n46858 = ~n46854 & n46857 ;
  assign n46859 = n9436 & n23382 ;
  assign n46860 = n46858 & ~n46859 ;
  assign n46861 = x38 & ~n46860 ;
  assign n46862 = x38 & ~n46861 ;
  assign n46863 = ~n46860 & ~n46861 ;
  assign n46864 = ~n46862 & ~n46863 ;
  assign n46865 = n46853 & ~n46864 ;
  assign n46866 = n46853 & ~n46865 ;
  assign n46867 = ~n46864 & ~n46865 ;
  assign n46868 = ~n46866 & ~n46867 ;
  assign n46869 = ~n46409 & ~n46423 ;
  assign n46870 = n46868 & n46869 ;
  assign n46871 = ~n46868 & ~n46869 ;
  assign n46872 = ~n46870 & ~n46871 ;
  assign n46873 = x126 & n8006 ;
  assign n46874 = x124 & n8474 ;
  assign n46875 = x125 & n8001 ;
  assign n46876 = ~n46874 & ~n46875 ;
  assign n46877 = ~n46873 & n46876 ;
  assign n46878 = n8009 & n25735 ;
  assign n46879 = n46877 & ~n46878 ;
  assign n46880 = x35 & ~n46879 ;
  assign n46881 = x35 & ~n46880 ;
  assign n46882 = ~n46879 & ~n46880 ;
  assign n46883 = ~n46881 & ~n46882 ;
  assign n46884 = n46872 & ~n46883 ;
  assign n46885 = n46872 & ~n46884 ;
  assign n46886 = ~n46883 & ~n46884 ;
  assign n46887 = ~n46885 & ~n46886 ;
  assign n46888 = ~n46696 & n46887 ;
  assign n46889 = n46696 & ~n46887 ;
  assign n46890 = ~n46888 & ~n46889 ;
  assign n46891 = ~n46684 & ~n46890 ;
  assign n46892 = ~n46684 & ~n46891 ;
  assign n46893 = ~n46890 & ~n46891 ;
  assign n46894 = ~n46892 & ~n46893 ;
  assign n46895 = ~n46683 & ~n46894 ;
  assign n46896 = n46683 & ~n46893 ;
  assign n46897 = ~n46892 & n46896 ;
  assign n46898 = ~n46895 & ~n46897 ;
  assign n47116 = n46898 & x223 ;
  assign n46899 = ~n46671 & ~n46676 ;
  assign n46900 = ~n46469 & ~n46665 ;
  assign n46901 = ~n46649 & ~n46662 ;
  assign n46902 = ~x127 & n7129 ;
  assign n46903 = n6728 & n27365 ;
  assign n46904 = ~n46902 & ~n46903 ;
  assign n46905 = ~x32 & ~n46904 ;
  assign n46906 = ~x32 & ~n46905 ;
  assign n46907 = ~n46904 & ~n46905 ;
  assign n46908 = ~n46906 & ~n46907 ;
  assign n46909 = ~n46901 & ~n46908 ;
  assign n46910 = ~n46901 & ~n46909 ;
  assign n46911 = ~n46908 & ~n46909 ;
  assign n46912 = ~n46910 & ~n46911 ;
  assign n46913 = ~n46152 & ~n46611 ;
  assign n46914 = ~n46626 & ~n46913 ;
  assign n46915 = ~x120 & n10905 ;
  assign n46916 = ~x118 & n11466 ;
  assign n46917 = ~x119 & n10900 ;
  assign n46918 = ~n46916 & ~n46917 ;
  assign n46919 = ~n46915 & n46918 ;
  assign n46920 = n10908 & n21501 ;
  assign n46921 = n46919 & ~n46920 ;
  assign n46922 = ~x41 & ~n46921 ;
  assign n46923 = ~x41 & ~n46922 ;
  assign n46924 = ~n46921 & ~n46922 ;
  assign n46925 = ~n46923 & ~n46924 ;
  assign n46926 = ~n46595 & ~n46608 ;
  assign n46927 = ~x117 & n12506 ;
  assign n46928 = ~x115 & n13131 ;
  assign n46929 = ~x116 & n12501 ;
  assign n46930 = ~n46928 & ~n46929 ;
  assign n46931 = ~n46927 & n46930 ;
  assign n46932 = n12509 & n19365 ;
  assign n46933 = n46931 & ~n46932 ;
  assign n46934 = ~x44 & ~n46933 ;
  assign n46935 = ~x44 & ~n46934 ;
  assign n46936 = ~n46933 & ~n46934 ;
  assign n46937 = ~n46935 & ~n46936 ;
  assign n46938 = ~n46576 & ~n46589 ;
  assign n46939 = ~n46536 & ~n46550 ;
  assign n46940 = ~x108 & n18025 ;
  assign n46941 = ~x106 & n18764 ;
  assign n46942 = ~x107 & n18020 ;
  assign n46943 = ~n46941 & ~n46942 ;
  assign n46944 = ~n46940 & n46943 ;
  assign n46945 = n13601 & n18028 ;
  assign n46946 = n46944 & ~n46945 ;
  assign n46947 = ~x53 & ~n46946 ;
  assign n46948 = ~x53 & ~n46947 ;
  assign n46949 = ~n46946 & ~n46947 ;
  assign n46950 = ~n46948 & ~n46949 ;
  assign n46951 = ~n46528 & ~n46532 ;
  assign n46952 = ~x105 & n20143 ;
  assign n46953 = ~x103 & n20854 ;
  assign n46954 = ~x104 & n20138 ;
  assign n46955 = ~n46953 & ~n46954 ;
  assign n46956 = ~n46952 & n46955 ;
  assign n46957 = n11907 & n20146 ;
  assign n46958 = n46956 & ~n46957 ;
  assign n46959 = ~x56 & ~n46958 ;
  assign n46960 = ~x56 & ~n46959 ;
  assign n46961 = ~n46958 & ~n46959 ;
  assign n46962 = ~n46960 & ~n46961 ;
  assign n46963 = ~n46520 & ~n46524 ;
  assign n46964 = ~n46504 & ~n46518 ;
  assign n46965 = ~x95 & n27427 ;
  assign n46966 = ~x96 & ~n26217 ;
  assign n46967 = ~n46965 & ~n46966 ;
  assign n46968 = ~n46501 & n46967 ;
  assign n46969 = n46501 & ~n46967 ;
  assign n46970 = ~n46964 & ~n46969 ;
  assign n46971 = ~n46968 & n46970 ;
  assign n46972 = ~n46964 & ~n46971 ;
  assign n46973 = ~n46968 & ~n46971 ;
  assign n46974 = ~n46969 & n46973 ;
  assign n46975 = ~n46972 & ~n46974 ;
  assign n46976 = ~x99 & n24612 ;
  assign n46977 = ~x97 & n25390 ;
  assign n46978 = ~x98 & n24607 ;
  assign n46979 = ~n46977 & ~n46978 ;
  assign n46980 = ~n46976 & n46979 ;
  assign n46981 = n8885 & n24615 ;
  assign n46982 = n46980 & ~n46981 ;
  assign n46983 = ~x62 & ~n46982 ;
  assign n46984 = ~x62 & ~n46983 ;
  assign n46985 = ~n46982 & ~n46983 ;
  assign n46986 = ~n46984 & ~n46985 ;
  assign n46987 = ~n46975 & ~n46986 ;
  assign n46988 = ~n46975 & ~n46987 ;
  assign n46989 = ~n46986 & ~n46987 ;
  assign n46990 = ~n46988 & ~n46989 ;
  assign n46991 = ~x102 & n22325 ;
  assign n46992 = ~x100 & n23066 ;
  assign n46993 = ~x101 & n22320 ;
  assign n46994 = ~n46992 & ~n46993 ;
  assign n46995 = ~n46991 & n46994 ;
  assign n46996 = n10333 & n22328 ;
  assign n46997 = n46995 & ~n46996 ;
  assign n46998 = ~x59 & ~n46997 ;
  assign n46999 = ~x59 & ~n46998 ;
  assign n47000 = ~n46997 & ~n46998 ;
  assign n47001 = ~n46999 & ~n47000 ;
  assign n47002 = ~n46990 & n47001 ;
  assign n47003 = n46990 & ~n47001 ;
  assign n47004 = ~n47002 & ~n47003 ;
  assign n47005 = ~n46963 & ~n47004 ;
  assign n47006 = n46963 & n47004 ;
  assign n47007 = ~n47005 & ~n47006 ;
  assign n47008 = ~n46962 & n47007 ;
  assign n47009 = n46962 & ~n47007 ;
  assign n47010 = ~n47008 & ~n47009 ;
  assign n47011 = ~n46951 & n47010 ;
  assign n47012 = n46951 & ~n47010 ;
  assign n47013 = ~n47011 & ~n47012 ;
  assign n47014 = ~n46950 & n47013 ;
  assign n47015 = n46950 & ~n47013 ;
  assign n47016 = ~n47014 & ~n47015 ;
  assign n47017 = ~n46939 & n47016 ;
  assign n47018 = n46939 & ~n47016 ;
  assign n47019 = ~n47017 & ~n47018 ;
  assign n47020 = ~x111 & n16076 ;
  assign n47021 = ~x109 & n16756 ;
  assign n47022 = ~x110 & n16071 ;
  assign n47023 = ~n47021 & ~n47022 ;
  assign n47024 = ~n47020 & n47023 ;
  assign n47025 = n15411 & n16079 ;
  assign n47026 = n47024 & ~n47025 ;
  assign n47027 = ~x50 & ~n47026 ;
  assign n47028 = ~x50 & ~n47027 ;
  assign n47029 = ~n47026 & ~n47027 ;
  assign n47030 = ~n47028 & ~n47029 ;
  assign n47031 = n47019 & ~n47030 ;
  assign n47032 = n47019 & ~n47031 ;
  assign n47033 = ~n47030 & ~n47031 ;
  assign n47034 = ~n47032 & ~n47033 ;
  assign n47035 = ~n46557 & ~n46570 ;
  assign n47036 = n47034 & n47035 ;
  assign n47037 = ~n47034 & ~n47035 ;
  assign n47038 = ~n47036 & ~n47037 ;
  assign n47039 = ~x114 & n14233 ;
  assign n47040 = ~x112 & n14876 ;
  assign n47041 = ~x113 & n14228 ;
  assign n47042 = ~n47040 & ~n47041 ;
  assign n47043 = ~n47039 & n47042 ;
  assign n47044 = n14236 & n17333 ;
  assign n47045 = n47043 & ~n47044 ;
  assign n47046 = ~x47 & ~n47045 ;
  assign n47047 = ~x47 & ~n47046 ;
  assign n47048 = ~n47045 & ~n47046 ;
  assign n47049 = ~n47047 & ~n47048 ;
  assign n47050 = ~n47038 & n47049 ;
  assign n47051 = n47038 & ~n47049 ;
  assign n47052 = ~n47050 & ~n47051 ;
  assign n47053 = ~n46938 & n47052 ;
  assign n47054 = ~n46938 & ~n47053 ;
  assign n47055 = n47052 & ~n47053 ;
  assign n47056 = ~n47054 & ~n47055 ;
  assign n47057 = ~n46937 & ~n47056 ;
  assign n47058 = n46937 & ~n47055 ;
  assign n47059 = ~n47054 & n47058 ;
  assign n47060 = ~n47057 & ~n47059 ;
  assign n47061 = ~n46926 & n47060 ;
  assign n47062 = n46926 & ~n47060 ;
  assign n47063 = ~n47061 & ~n47062 ;
  assign n47064 = ~n46925 & n47063 ;
  assign n47065 = n46925 & ~n47063 ;
  assign n47066 = ~n47064 & ~n47065 ;
  assign n47067 = ~n46914 & n47066 ;
  assign n47068 = n46914 & ~n47066 ;
  assign n47069 = ~n47067 & ~n47068 ;
  assign n47070 = ~x123 & n9433 ;
  assign n47071 = ~x121 & n9915 ;
  assign n47072 = ~x122 & n9428 ;
  assign n47073 = ~n47071 & ~n47072 ;
  assign n47074 = ~n47070 & n47073 ;
  assign n47075 = n9436 & n23760 ;
  assign n47076 = n47074 & ~n47075 ;
  assign n47077 = ~x38 & ~n47076 ;
  assign n47078 = ~x38 & ~n47077 ;
  assign n47079 = ~n47076 & ~n47077 ;
  assign n47080 = ~n47078 & ~n47079 ;
  assign n47081 = n47069 & ~n47080 ;
  assign n47082 = n47069 & ~n47081 ;
  assign n47083 = ~n47080 & ~n47081 ;
  assign n47084 = ~n47082 & ~n47083 ;
  assign n47085 = ~n46629 & ~n46643 ;
  assign n47086 = n47084 & n47085 ;
  assign n47087 = ~n47084 & ~n47085 ;
  assign n47088 = ~n47086 & ~n47087 ;
  assign n47089 = ~x126 & n8006 ;
  assign n47090 = ~x124 & n8474 ;
  assign n47091 = ~x125 & n8001 ;
  assign n47092 = ~n47090 & ~n47091 ;
  assign n47093 = ~n47089 & n47092 ;
  assign n47094 = n8009 & n26128 ;
  assign n47095 = n47093 & ~n47094 ;
  assign n47096 = ~x35 & ~n47095 ;
  assign n47097 = ~x35 & ~n47096 ;
  assign n47098 = ~n47095 & ~n47096 ;
  assign n47099 = ~n47097 & ~n47098 ;
  assign n47100 = n47088 & ~n47099 ;
  assign n47101 = n47088 & ~n47100 ;
  assign n47102 = ~n47099 & ~n47100 ;
  assign n47103 = ~n47101 & ~n47102 ;
  assign n47104 = ~n46912 & n47103 ;
  assign n47105 = n46912 & ~n47103 ;
  assign n47106 = ~n47104 & ~n47105 ;
  assign n47107 = ~n46900 & ~n47106 ;
  assign n47108 = ~n46900 & ~n47107 ;
  assign n47109 = ~n47106 & ~n47107 ;
  assign n47110 = ~n47108 & ~n47109 ;
  assign n47111 = ~n46899 & ~n47110 ;
  assign n47112 = n46899 & ~n47109 ;
  assign n47113 = ~n47108 & n47112 ;
  assign n47114 = ~n47111 & ~n47113 ;
  assign n47117 = ~n47114 & ~x223 ;
  assign n47118 = ~n47116 & ~n47117 ;
  assign n47119 = ~n46891 & ~n46895 ;
  assign n47120 = ~n46696 & ~n46887 ;
  assign n47121 = ~n46693 & ~n47120 ;
  assign n47122 = ~n46837 & ~n46841 ;
  assign n47123 = ~n46821 & ~n46835 ;
  assign n47124 = ~n46774 & ~n46785 ;
  assign n47125 = ~n46771 & ~n47124 ;
  assign n47126 = x96 & n27024 ;
  assign n47127 = x97 & ~n26217 ;
  assign n47128 = ~n47126 & ~n47127 ;
  assign n47129 = ~x32 & ~n47128 ;
  assign n47130 = x32 & n47128 ;
  assign n47131 = ~n47129 & ~n47130 ;
  assign n47132 = ~n46751 & n47131 ;
  assign n47133 = ~n46751 & ~n47132 ;
  assign n47134 = n47131 & ~n47132 ;
  assign n47135 = ~n47133 & ~n47134 ;
  assign n47136 = ~n46757 & ~n47135 ;
  assign n47137 = ~n46757 & ~n47136 ;
  assign n47138 = ~n47135 & ~n47136 ;
  assign n47139 = ~n47137 & ~n47138 ;
  assign n47140 = x100 & n24612 ;
  assign n47141 = x98 & n25390 ;
  assign n47142 = x99 & n24607 ;
  assign n47143 = ~n47141 & ~n47142 ;
  assign n47144 = ~n47140 & n47143 ;
  assign n47145 = n9115 & n24615 ;
  assign n47146 = n47144 & ~n47145 ;
  assign n47147 = x62 & ~n47146 ;
  assign n47148 = x62 & ~n47147 ;
  assign n47149 = ~n47146 & ~n47147 ;
  assign n47150 = ~n47148 & ~n47149 ;
  assign n47151 = ~n47139 & n47150 ;
  assign n47152 = n47139 & ~n47150 ;
  assign n47153 = ~n47151 & ~n47152 ;
  assign n47154 = x103 & n22325 ;
  assign n47155 = x101 & n23066 ;
  assign n47156 = x102 & n22320 ;
  assign n47157 = ~n47155 & ~n47156 ;
  assign n47158 = ~n47154 & n47157 ;
  assign n47159 = n10588 & n22328 ;
  assign n47160 = n47158 & ~n47159 ;
  assign n47161 = x59 & ~n47160 ;
  assign n47162 = x59 & ~n47161 ;
  assign n47163 = ~n47160 & ~n47161 ;
  assign n47164 = ~n47162 & ~n47163 ;
  assign n47165 = ~n47153 & ~n47164 ;
  assign n47166 = n47153 & n47164 ;
  assign n47167 = ~n47165 & ~n47166 ;
  assign n47168 = ~n47125 & n47167 ;
  assign n47169 = n47125 & ~n47167 ;
  assign n47170 = ~n47168 & ~n47169 ;
  assign n47171 = x106 & n20143 ;
  assign n47172 = x104 & n20854 ;
  assign n47173 = x105 & n20138 ;
  assign n47174 = ~n47172 & ~n47173 ;
  assign n47175 = ~n47171 & n47174 ;
  assign n47176 = n12181 & n20146 ;
  assign n47177 = n47175 & ~n47176 ;
  assign n47178 = x56 & ~n47177 ;
  assign n47179 = x56 & ~n47178 ;
  assign n47180 = ~n47177 & ~n47178 ;
  assign n47181 = ~n47179 & ~n47180 ;
  assign n47182 = n47170 & ~n47181 ;
  assign n47183 = n47170 & ~n47182 ;
  assign n47184 = ~n47181 & ~n47182 ;
  assign n47185 = ~n47183 & ~n47184 ;
  assign n47186 = ~n46789 & ~n46792 ;
  assign n47187 = n47185 & n47186 ;
  assign n47188 = ~n47185 & ~n47186 ;
  assign n47189 = ~n47187 & ~n47188 ;
  assign n47190 = x109 & n18025 ;
  assign n47191 = x107 & n18764 ;
  assign n47192 = x108 & n18020 ;
  assign n47193 = ~n47191 & ~n47192 ;
  assign n47194 = ~n47190 & n47193 ;
  assign n47195 = n13894 & n18028 ;
  assign n47196 = n47194 & ~n47195 ;
  assign n47197 = x53 & ~n47196 ;
  assign n47198 = x53 & ~n47197 ;
  assign n47199 = ~n47196 & ~n47197 ;
  assign n47200 = ~n47198 & ~n47199 ;
  assign n47201 = n47189 & ~n47200 ;
  assign n47202 = n47189 & ~n47201 ;
  assign n47203 = ~n47200 & ~n47201 ;
  assign n47204 = ~n47202 & ~n47203 ;
  assign n47205 = ~n46795 & ~n46798 ;
  assign n47206 = n47204 & n47205 ;
  assign n47207 = ~n47204 & ~n47205 ;
  assign n47208 = ~n47206 & ~n47207 ;
  assign n47209 = x112 & n16076 ;
  assign n47210 = x110 & n16756 ;
  assign n47211 = x111 & n16071 ;
  assign n47212 = ~n47210 & ~n47211 ;
  assign n47213 = ~n47209 & n47212 ;
  assign n47214 = n15442 & n16079 ;
  assign n47215 = n47213 & ~n47214 ;
  assign n47216 = x50 & ~n47215 ;
  assign n47217 = x50 & ~n47216 ;
  assign n47218 = ~n47215 & ~n47216 ;
  assign n47219 = ~n47217 & ~n47218 ;
  assign n47220 = n47208 & ~n47219 ;
  assign n47221 = n47208 & ~n47220 ;
  assign n47222 = ~n47219 & ~n47220 ;
  assign n47223 = ~n47221 & ~n47222 ;
  assign n47224 = ~n46801 & ~n46815 ;
  assign n47225 = n47223 & n47224 ;
  assign n47226 = ~n47223 & ~n47224 ;
  assign n47227 = ~n47225 & ~n47226 ;
  assign n47228 = x115 & n14233 ;
  assign n47229 = x113 & n14876 ;
  assign n47230 = x114 & n14228 ;
  assign n47231 = ~n47229 & ~n47230 ;
  assign n47232 = ~n47228 & n47231 ;
  assign n47233 = n14236 & n17364 ;
  assign n47234 = n47232 & ~n47233 ;
  assign n47235 = x47 & ~n47234 ;
  assign n47236 = x47 & ~n47235 ;
  assign n47237 = ~n47234 & ~n47235 ;
  assign n47238 = ~n47236 & ~n47237 ;
  assign n47239 = n47227 & ~n47238 ;
  assign n47240 = ~n47227 & n47238 ;
  assign n47241 = ~n47123 & ~n47240 ;
  assign n47242 = ~n47239 & n47241 ;
  assign n47243 = ~n47123 & ~n47242 ;
  assign n47244 = ~n47239 & ~n47242 ;
  assign n47245 = ~n47240 & n47244 ;
  assign n47246 = ~n47243 & ~n47245 ;
  assign n47247 = x118 & n12506 ;
  assign n47248 = x116 & n13131 ;
  assign n47249 = x117 & n12501 ;
  assign n47250 = ~n47248 & ~n47249 ;
  assign n47251 = ~n47247 & n47250 ;
  assign n47252 = n12509 & n19395 ;
  assign n47253 = n47251 & ~n47252 ;
  assign n47254 = x44 & ~n47253 ;
  assign n47255 = x44 & ~n47254 ;
  assign n47256 = ~n47253 & ~n47254 ;
  assign n47257 = ~n47255 & ~n47256 ;
  assign n47258 = n47246 & n47257 ;
  assign n47259 = ~n47246 & ~n47257 ;
  assign n47260 = ~n47258 & ~n47259 ;
  assign n47261 = ~n47122 & n47260 ;
  assign n47262 = n47122 & ~n47260 ;
  assign n47263 = ~n47261 & ~n47262 ;
  assign n47264 = x121 & n10905 ;
  assign n47265 = x119 & n11466 ;
  assign n47266 = x120 & n10900 ;
  assign n47267 = ~n47265 & ~n47266 ;
  assign n47268 = ~n47264 & n47267 ;
  assign n47269 = n10908 & n21870 ;
  assign n47270 = n47268 & ~n47269 ;
  assign n47271 = x41 & ~n47270 ;
  assign n47272 = x41 & ~n47271 ;
  assign n47273 = ~n47270 & ~n47271 ;
  assign n47274 = ~n47272 & ~n47273 ;
  assign n47275 = n47263 & ~n47274 ;
  assign n47276 = n47263 & ~n47275 ;
  assign n47277 = ~n47274 & ~n47275 ;
  assign n47278 = ~n47276 & ~n47277 ;
  assign n47279 = ~n46845 & ~n46848 ;
  assign n47280 = n47278 & n47279 ;
  assign n47281 = ~n47278 & ~n47279 ;
  assign n47282 = ~n47280 & ~n47281 ;
  assign n47283 = x124 & n9433 ;
  assign n47284 = x122 & n9915 ;
  assign n47285 = x123 & n9428 ;
  assign n47286 = ~n47284 & ~n47285 ;
  assign n47287 = ~n47283 & n47286 ;
  assign n47288 = n9436 & n23796 ;
  assign n47289 = n47287 & ~n47288 ;
  assign n47290 = x38 & ~n47289 ;
  assign n47291 = x38 & ~n47290 ;
  assign n47292 = ~n47289 & ~n47290 ;
  assign n47293 = ~n47291 & ~n47292 ;
  assign n47294 = n47282 & ~n47293 ;
  assign n47295 = n47282 & ~n47294 ;
  assign n47296 = ~n47293 & ~n47294 ;
  assign n47297 = ~n47295 & ~n47296 ;
  assign n47298 = ~n46851 & ~n46865 ;
  assign n47299 = n47297 & n47298 ;
  assign n47300 = ~n47297 & ~n47298 ;
  assign n47301 = ~n47299 & ~n47300 ;
  assign n47302 = ~n46871 & ~n46884 ;
  assign n47303 = x127 & n8006 ;
  assign n47304 = x125 & n8474 ;
  assign n47305 = x126 & n8001 ;
  assign n47306 = ~n47304 & ~n47305 ;
  assign n47307 = ~n47303 & n47306 ;
  assign n47308 = n8009 & n26533 ;
  assign n47309 = n47307 & ~n47308 ;
  assign n47310 = x35 & ~n47309 ;
  assign n47311 = x35 & ~n47310 ;
  assign n47312 = ~n47309 & ~n47310 ;
  assign n47313 = ~n47311 & ~n47312 ;
  assign n47314 = ~n47302 & ~n47313 ;
  assign n47315 = ~n47302 & ~n47314 ;
  assign n47316 = ~n47313 & ~n47314 ;
  assign n47317 = ~n47315 & ~n47316 ;
  assign n47318 = ~n47301 & n47317 ;
  assign n47319 = n47301 & ~n47317 ;
  assign n47320 = ~n47318 & ~n47319 ;
  assign n47321 = ~n47121 & n47320 ;
  assign n47322 = n47121 & ~n47320 ;
  assign n47323 = ~n47321 & ~n47322 ;
  assign n47324 = ~n47119 & n47323 ;
  assign n47325 = n47119 & ~n47323 ;
  assign n47326 = ~n47324 & ~n47325 ;
  assign n47536 = n47326 & x224 ;
  assign n47327 = ~n47107 & ~n47111 ;
  assign n47328 = ~n46912 & ~n47103 ;
  assign n47329 = ~n46909 & ~n47328 ;
  assign n47330 = ~n47053 & ~n47057 ;
  assign n47331 = ~n47037 & ~n47051 ;
  assign n47332 = ~n46990 & ~n47001 ;
  assign n47333 = ~n46987 & ~n47332 ;
  assign n47334 = ~x96 & n27427 ;
  assign n47335 = ~x97 & ~n26217 ;
  assign n47336 = ~n47334 & ~n47335 ;
  assign n47337 = x32 & ~n47336 ;
  assign n47338 = ~x32 & n47336 ;
  assign n47339 = ~n47337 & ~n47338 ;
  assign n47340 = ~n46967 & n47339 ;
  assign n47341 = ~n46967 & ~n47340 ;
  assign n47342 = n47339 & ~n47340 ;
  assign n47343 = ~n47341 & ~n47342 ;
  assign n47344 = ~n46973 & ~n47343 ;
  assign n47345 = ~n46973 & ~n47344 ;
  assign n47346 = ~n47343 & ~n47344 ;
  assign n47347 = ~n47345 & ~n47346 ;
  assign n47348 = ~x100 & n24612 ;
  assign n47349 = ~x98 & n25390 ;
  assign n47350 = ~x99 & n24607 ;
  assign n47351 = ~n47349 & ~n47350 ;
  assign n47352 = ~n47348 & n47351 ;
  assign n47353 = n9338 & n24615 ;
  assign n47354 = n47352 & ~n47353 ;
  assign n47355 = ~x62 & ~n47354 ;
  assign n47356 = ~x62 & ~n47355 ;
  assign n47357 = ~n47354 & ~n47355 ;
  assign n47358 = ~n47356 & ~n47357 ;
  assign n47359 = ~n47347 & n47358 ;
  assign n47360 = n47347 & ~n47358 ;
  assign n47361 = ~n47359 & ~n47360 ;
  assign n47362 = ~x103 & n22325 ;
  assign n47363 = ~x101 & n23066 ;
  assign n47364 = ~x102 & n22320 ;
  assign n47365 = ~n47363 & ~n47364 ;
  assign n47366 = ~n47362 & n47365 ;
  assign n47367 = n10833 & n22328 ;
  assign n47368 = n47366 & ~n47367 ;
  assign n47369 = ~x59 & ~n47368 ;
  assign n47370 = ~x59 & ~n47369 ;
  assign n47371 = ~n47368 & ~n47369 ;
  assign n47372 = ~n47370 & ~n47371 ;
  assign n47373 = ~n47361 & ~n47372 ;
  assign n47374 = n47361 & n47372 ;
  assign n47375 = ~n47373 & ~n47374 ;
  assign n47376 = ~n47333 & n47375 ;
  assign n47377 = n47333 & ~n47375 ;
  assign n47378 = ~n47376 & ~n47377 ;
  assign n47379 = ~x106 & n20143 ;
  assign n47380 = ~x104 & n20854 ;
  assign n47381 = ~x105 & n20138 ;
  assign n47382 = ~n47380 & ~n47381 ;
  assign n47383 = ~n47379 & n47382 ;
  assign n47384 = n12447 & n20146 ;
  assign n47385 = n47383 & ~n47384 ;
  assign n47386 = ~x56 & ~n47385 ;
  assign n47387 = ~x56 & ~n47386 ;
  assign n47388 = ~n47385 & ~n47386 ;
  assign n47389 = ~n47387 & ~n47388 ;
  assign n47390 = n47378 & ~n47389 ;
  assign n47391 = n47378 & ~n47390 ;
  assign n47392 = ~n47389 & ~n47390 ;
  assign n47393 = ~n47391 & ~n47392 ;
  assign n47394 = ~n47005 & ~n47008 ;
  assign n47395 = n47393 & n47394 ;
  assign n47396 = ~n47393 & ~n47394 ;
  assign n47397 = ~n47395 & ~n47396 ;
  assign n47398 = ~x109 & n18025 ;
  assign n47399 = ~x107 & n18764 ;
  assign n47400 = ~x108 & n18020 ;
  assign n47401 = ~n47399 & ~n47400 ;
  assign n47402 = ~n47398 & n47401 ;
  assign n47403 = n14177 & n18028 ;
  assign n47404 = n47402 & ~n47403 ;
  assign n47405 = ~x53 & ~n47404 ;
  assign n47406 = ~x53 & ~n47405 ;
  assign n47407 = ~n47404 & ~n47405 ;
  assign n47408 = ~n47406 & ~n47407 ;
  assign n47409 = n47397 & ~n47408 ;
  assign n47410 = n47397 & ~n47409 ;
  assign n47411 = ~n47408 & ~n47409 ;
  assign n47412 = ~n47410 & ~n47411 ;
  assign n47413 = ~n47011 & ~n47014 ;
  assign n47414 = n47412 & n47413 ;
  assign n47415 = ~n47412 & ~n47413 ;
  assign n47416 = ~n47414 & ~n47415 ;
  assign n47417 = ~x112 & n16076 ;
  assign n47418 = ~x110 & n16756 ;
  assign n47419 = ~x111 & n16071 ;
  assign n47420 = ~n47418 & ~n47419 ;
  assign n47421 = ~n47417 & n47420 ;
  assign n47422 = n15744 & n16079 ;
  assign n47423 = n47421 & ~n47422 ;
  assign n47424 = ~x50 & ~n47423 ;
  assign n47425 = ~x50 & ~n47424 ;
  assign n47426 = ~n47423 & ~n47424 ;
  assign n47427 = ~n47425 & ~n47426 ;
  assign n47428 = n47416 & ~n47427 ;
  assign n47429 = n47416 & ~n47428 ;
  assign n47430 = ~n47427 & ~n47428 ;
  assign n47431 = ~n47429 & ~n47430 ;
  assign n47432 = ~n47017 & ~n47031 ;
  assign n47433 = n47431 & n47432 ;
  assign n47434 = ~n47431 & ~n47432 ;
  assign n47435 = ~n47433 & ~n47434 ;
  assign n47436 = ~x115 & n14233 ;
  assign n47437 = ~x113 & n14876 ;
  assign n47438 = ~x114 & n14228 ;
  assign n47439 = ~n47437 & ~n47438 ;
  assign n47440 = ~n47436 & n47439 ;
  assign n47441 = n14236 & n17683 ;
  assign n47442 = n47440 & ~n47441 ;
  assign n47443 = ~x47 & ~n47442 ;
  assign n47444 = ~x47 & ~n47443 ;
  assign n47445 = ~n47442 & ~n47443 ;
  assign n47446 = ~n47444 & ~n47445 ;
  assign n47447 = n47435 & ~n47446 ;
  assign n47448 = ~n47435 & n47446 ;
  assign n47449 = ~n47331 & ~n47448 ;
  assign n47450 = ~n47447 & n47449 ;
  assign n47451 = ~n47331 & ~n47450 ;
  assign n47452 = ~n47447 & ~n47450 ;
  assign n47453 = ~n47448 & n47452 ;
  assign n47454 = ~n47451 & ~n47453 ;
  assign n47455 = ~x118 & n12506 ;
  assign n47456 = ~x116 & n13131 ;
  assign n47457 = ~x117 & n12501 ;
  assign n47458 = ~n47456 & ~n47457 ;
  assign n47459 = ~n47455 & n47458 ;
  assign n47460 = n12509 & n19736 ;
  assign n47461 = n47459 & ~n47460 ;
  assign n47462 = ~x44 & ~n47461 ;
  assign n47463 = ~x44 & ~n47462 ;
  assign n47464 = ~n47461 & ~n47462 ;
  assign n47465 = ~n47463 & ~n47464 ;
  assign n47466 = n47454 & n47465 ;
  assign n47467 = ~n47454 & ~n47465 ;
  assign n47468 = ~n47466 & ~n47467 ;
  assign n47469 = ~n47330 & n47468 ;
  assign n47470 = n47330 & ~n47468 ;
  assign n47471 = ~n47469 & ~n47470 ;
  assign n47472 = ~x121 & n10905 ;
  assign n47473 = ~x119 & n11466 ;
  assign n47474 = ~x120 & n10900 ;
  assign n47475 = ~n47473 & ~n47474 ;
  assign n47476 = ~n47472 & n47475 ;
  assign n47477 = n10908 & n22229 ;
  assign n47478 = n47476 & ~n47477 ;
  assign n47479 = ~x41 & ~n47478 ;
  assign n47480 = ~x41 & ~n47479 ;
  assign n47481 = ~n47478 & ~n47479 ;
  assign n47482 = ~n47480 & ~n47481 ;
  assign n47483 = n47471 & ~n47482 ;
  assign n47484 = n47471 & ~n47483 ;
  assign n47485 = ~n47482 & ~n47483 ;
  assign n47486 = ~n47484 & ~n47485 ;
  assign n47487 = ~n47061 & ~n47064 ;
  assign n47488 = n47486 & n47487 ;
  assign n47489 = ~n47486 & ~n47487 ;
  assign n47490 = ~n47488 & ~n47489 ;
  assign n47491 = ~x124 & n9433 ;
  assign n47492 = ~x122 & n9915 ;
  assign n47493 = ~x123 & n9428 ;
  assign n47494 = ~n47492 & ~n47493 ;
  assign n47495 = ~n47491 & n47494 ;
  assign n47496 = n9436 & n24176 ;
  assign n47497 = n47495 & ~n47496 ;
  assign n47498 = ~x38 & ~n47497 ;
  assign n47499 = ~x38 & ~n47498 ;
  assign n47500 = ~n47497 & ~n47498 ;
  assign n47501 = ~n47499 & ~n47500 ;
  assign n47502 = n47490 & ~n47501 ;
  assign n47503 = n47490 & ~n47502 ;
  assign n47504 = ~n47501 & ~n47502 ;
  assign n47505 = ~n47503 & ~n47504 ;
  assign n47506 = ~n47067 & ~n47081 ;
  assign n47507 = n47505 & n47506 ;
  assign n47508 = ~n47505 & ~n47506 ;
  assign n47509 = ~n47507 & ~n47508 ;
  assign n47510 = ~n47087 & ~n47100 ;
  assign n47511 = ~x127 & n8006 ;
  assign n47512 = ~x125 & n8474 ;
  assign n47513 = ~x126 & n8001 ;
  assign n47514 = ~n47512 & ~n47513 ;
  assign n47515 = ~n47511 & n47514 ;
  assign n47516 = n8009 & n26932 ;
  assign n47517 = n47515 & ~n47516 ;
  assign n47518 = ~x35 & ~n47517 ;
  assign n47519 = ~x35 & ~n47518 ;
  assign n47520 = ~n47517 & ~n47518 ;
  assign n47521 = ~n47519 & ~n47520 ;
  assign n47522 = ~n47510 & ~n47521 ;
  assign n47523 = ~n47510 & ~n47522 ;
  assign n47524 = ~n47521 & ~n47522 ;
  assign n47525 = ~n47523 & ~n47524 ;
  assign n47526 = ~n47509 & n47525 ;
  assign n47527 = n47509 & ~n47525 ;
  assign n47528 = ~n47526 & ~n47527 ;
  assign n47529 = ~n47329 & n47528 ;
  assign n47530 = n47329 & ~n47528 ;
  assign n47531 = ~n47529 & ~n47530 ;
  assign n47532 = ~n47327 & n47531 ;
  assign n47533 = n47327 & ~n47531 ;
  assign n47534 = ~n47532 & ~n47533 ;
  assign n47537 = ~n47534 & ~x224 ;
  assign n47538 = ~n47536 & ~n47537 ;
  assign n47539 = ~n47294 & ~n47300 ;
  assign n47540 = x126 & n8474 ;
  assign n47541 = x127 & n8001 ;
  assign n47542 = ~n47540 & ~n47541 ;
  assign n47543 = ~n8009 & n47542 ;
  assign n47544 = n26965 & n47542 ;
  assign n47545 = ~n47543 & ~n47544 ;
  assign n47546 = x35 & ~n47545 ;
  assign n47547 = ~x35 & n47545 ;
  assign n47548 = ~n47546 & ~n47547 ;
  assign n47549 = ~n47539 & ~n47548 ;
  assign n47550 = n47539 & n47548 ;
  assign n47551 = ~n47549 & ~n47550 ;
  assign n47552 = ~n47259 & ~n47261 ;
  assign n47553 = ~n47165 & ~n47168 ;
  assign n47554 = x104 & n22325 ;
  assign n47555 = x102 & n23066 ;
  assign n47556 = x103 & n22320 ;
  assign n47557 = ~n47555 & ~n47556 ;
  assign n47558 = ~n47554 & n47557 ;
  assign n47559 = n11116 & n22328 ;
  assign n47560 = n47558 & ~n47559 ;
  assign n47561 = x59 & ~n47560 ;
  assign n47562 = x59 & ~n47561 ;
  assign n47563 = ~n47560 & ~n47561 ;
  assign n47564 = ~n47562 & ~n47563 ;
  assign n47565 = ~n47139 & ~n47150 ;
  assign n47566 = ~n47136 & ~n47565 ;
  assign n47567 = x97 & n27024 ;
  assign n47568 = x98 & ~n26217 ;
  assign n47569 = ~n47567 & ~n47568 ;
  assign n47570 = ~n47129 & ~n47132 ;
  assign n47571 = ~n47569 & n47570 ;
  assign n47572 = n47569 & ~n47570 ;
  assign n47573 = ~n47571 & ~n47572 ;
  assign n47574 = x101 & n24612 ;
  assign n47575 = x99 & n25390 ;
  assign n47576 = x100 & n24607 ;
  assign n47577 = ~n47575 & ~n47576 ;
  assign n47578 = ~n47574 & n47577 ;
  assign n47579 = n9601 & n24615 ;
  assign n47580 = n47578 & ~n47579 ;
  assign n47581 = x62 & ~n47580 ;
  assign n47582 = x62 & ~n47581 ;
  assign n47583 = ~n47580 & ~n47581 ;
  assign n47584 = ~n47582 & ~n47583 ;
  assign n47585 = ~n47573 & n47584 ;
  assign n47586 = n47573 & ~n47584 ;
  assign n47587 = ~n47585 & ~n47586 ;
  assign n47588 = ~n47566 & n47587 ;
  assign n47589 = ~n47566 & ~n47588 ;
  assign n47590 = n47587 & ~n47588 ;
  assign n47591 = ~n47589 & ~n47590 ;
  assign n47592 = ~n47564 & ~n47591 ;
  assign n47593 = n47564 & ~n47590 ;
  assign n47594 = ~n47589 & n47593 ;
  assign n47595 = ~n47592 & ~n47594 ;
  assign n47596 = ~n47553 & n47595 ;
  assign n47597 = n47553 & ~n47595 ;
  assign n47598 = ~n47596 & ~n47597 ;
  assign n47599 = x107 & n20143 ;
  assign n47600 = x105 & n20854 ;
  assign n47601 = x106 & n20138 ;
  assign n47602 = ~n47600 & ~n47601 ;
  assign n47603 = ~n47599 & n47602 ;
  assign n47604 = n12749 & n20146 ;
  assign n47605 = n47603 & ~n47604 ;
  assign n47606 = x56 & ~n47605 ;
  assign n47607 = x56 & ~n47606 ;
  assign n47608 = ~n47605 & ~n47606 ;
  assign n47609 = ~n47607 & ~n47608 ;
  assign n47610 = n47598 & ~n47609 ;
  assign n47611 = n47598 & ~n47610 ;
  assign n47612 = ~n47609 & ~n47610 ;
  assign n47613 = ~n47611 & ~n47612 ;
  assign n47614 = ~n47182 & ~n47188 ;
  assign n47615 = n47613 & n47614 ;
  assign n47616 = ~n47613 & ~n47614 ;
  assign n47617 = ~n47615 & ~n47616 ;
  assign n47618 = x110 & n18025 ;
  assign n47619 = x108 & n18764 ;
  assign n47620 = x109 & n18020 ;
  assign n47621 = ~n47619 & ~n47620 ;
  assign n47622 = ~n47618 & n47621 ;
  assign n47623 = n14497 & n18028 ;
  assign n47624 = n47622 & ~n47623 ;
  assign n47625 = x53 & ~n47624 ;
  assign n47626 = x53 & ~n47625 ;
  assign n47627 = ~n47624 & ~n47625 ;
  assign n47628 = ~n47626 & ~n47627 ;
  assign n47629 = n47617 & ~n47628 ;
  assign n47630 = n47617 & ~n47629 ;
  assign n47631 = ~n47628 & ~n47629 ;
  assign n47632 = ~n47630 & ~n47631 ;
  assign n47633 = ~n47201 & ~n47207 ;
  assign n47634 = n47632 & n47633 ;
  assign n47635 = ~n47632 & ~n47633 ;
  assign n47636 = ~n47634 & ~n47635 ;
  assign n47637 = x113 & n16076 ;
  assign n47638 = x111 & n16756 ;
  assign n47639 = x112 & n16071 ;
  assign n47640 = ~n47638 & ~n47639 ;
  assign n47641 = ~n47637 & n47640 ;
  assign n47642 = n16079 & n16361 ;
  assign n47643 = n47641 & ~n47642 ;
  assign n47644 = x50 & ~n47643 ;
  assign n47645 = x50 & ~n47644 ;
  assign n47646 = ~n47643 & ~n47644 ;
  assign n47647 = ~n47645 & ~n47646 ;
  assign n47648 = n47636 & ~n47647 ;
  assign n47649 = n47636 & ~n47648 ;
  assign n47650 = ~n47647 & ~n47648 ;
  assign n47651 = ~n47649 & ~n47650 ;
  assign n47652 = ~n47220 & ~n47226 ;
  assign n47653 = n47651 & n47652 ;
  assign n47654 = ~n47651 & ~n47652 ;
  assign n47655 = ~n47653 & ~n47654 ;
  assign n47656 = x116 & n14233 ;
  assign n47657 = x114 & n14876 ;
  assign n47658 = x115 & n14228 ;
  assign n47659 = ~n47657 & ~n47658 ;
  assign n47660 = ~n47656 & n47659 ;
  assign n47661 = n14236 & n18336 ;
  assign n47662 = n47660 & ~n47661 ;
  assign n47663 = x47 & ~n47662 ;
  assign n47664 = x47 & ~n47663 ;
  assign n47665 = ~n47662 & ~n47663 ;
  assign n47666 = ~n47664 & ~n47665 ;
  assign n47667 = n47655 & ~n47666 ;
  assign n47668 = n47655 & ~n47667 ;
  assign n47669 = ~n47666 & ~n47667 ;
  assign n47670 = ~n47668 & ~n47669 ;
  assign n47671 = ~n47244 & n47670 ;
  assign n47672 = n47244 & ~n47670 ;
  assign n47673 = ~n47671 & ~n47672 ;
  assign n47674 = x119 & n12506 ;
  assign n47675 = x117 & n13131 ;
  assign n47676 = x118 & n12501 ;
  assign n47677 = ~n47675 & ~n47676 ;
  assign n47678 = ~n47674 & n47677 ;
  assign n47679 = n12509 & n20423 ;
  assign n47680 = n47678 & ~n47679 ;
  assign n47681 = x44 & ~n47680 ;
  assign n47682 = x44 & ~n47681 ;
  assign n47683 = ~n47680 & ~n47681 ;
  assign n47684 = ~n47682 & ~n47683 ;
  assign n47685 = ~n47673 & ~n47684 ;
  assign n47686 = n47673 & n47684 ;
  assign n47687 = ~n47685 & ~n47686 ;
  assign n47688 = ~n47552 & n47687 ;
  assign n47689 = n47552 & ~n47687 ;
  assign n47690 = ~n47688 & ~n47689 ;
  assign n47691 = x122 & n10905 ;
  assign n47692 = x120 & n11466 ;
  assign n47693 = x121 & n10900 ;
  assign n47694 = ~n47692 & ~n47693 ;
  assign n47695 = ~n47691 & n47694 ;
  assign n47696 = n10908 & n22622 ;
  assign n47697 = n47695 & ~n47696 ;
  assign n47698 = x41 & ~n47697 ;
  assign n47699 = x41 & ~n47698 ;
  assign n47700 = ~n47697 & ~n47698 ;
  assign n47701 = ~n47699 & ~n47700 ;
  assign n47702 = n47690 & ~n47701 ;
  assign n47703 = n47690 & ~n47702 ;
  assign n47704 = ~n47701 & ~n47702 ;
  assign n47705 = ~n47703 & ~n47704 ;
  assign n47706 = ~n47275 & ~n47281 ;
  assign n47707 = n47705 & n47706 ;
  assign n47708 = ~n47705 & ~n47706 ;
  assign n47709 = ~n47707 & ~n47708 ;
  assign n47710 = x125 & n9433 ;
  assign n47711 = x123 & n9915 ;
  assign n47712 = x124 & n9428 ;
  assign n47713 = ~n47711 & ~n47712 ;
  assign n47714 = ~n47710 & n47713 ;
  assign n47715 = n9436 & n24935 ;
  assign n47716 = n47714 & ~n47715 ;
  assign n47717 = x38 & ~n47716 ;
  assign n47718 = x38 & ~n47717 ;
  assign n47719 = ~n47716 & ~n47717 ;
  assign n47720 = ~n47718 & ~n47719 ;
  assign n47721 = n47709 & ~n47720 ;
  assign n47722 = ~n47709 & n47720 ;
  assign n47723 = n47551 & ~n47722 ;
  assign n47724 = ~n47721 & n47723 ;
  assign n47725 = n47551 & ~n47724 ;
  assign n47726 = ~n47722 & ~n47724 ;
  assign n47727 = ~n47721 & n47726 ;
  assign n47728 = ~n47725 & ~n47727 ;
  assign n47729 = ~n47314 & ~n47319 ;
  assign n47730 = ~n47728 & ~n47729 ;
  assign n47731 = ~n47728 & ~n47730 ;
  assign n47732 = ~n47729 & ~n47730 ;
  assign n47733 = ~n47731 & ~n47732 ;
  assign n47734 = ~n47321 & ~n47324 ;
  assign n47735 = ~n47733 & ~n47734 ;
  assign n47736 = n47733 & n47734 ;
  assign n47737 = ~n47735 & ~n47736 ;
  assign n47938 = n47737 & x225 ;
  assign n47738 = ~n47502 & ~n47508 ;
  assign n47739 = ~x126 & n8474 ;
  assign n47740 = ~x127 & n8001 ;
  assign n47741 = ~n47739 & ~n47740 ;
  assign n47742 = ~n8009 & n47741 ;
  assign n47743 = n27368 & n47741 ;
  assign n47744 = ~n47742 & ~n47743 ;
  assign n47745 = ~x35 & ~n47744 ;
  assign n47746 = x35 & n47744 ;
  assign n47747 = ~n47745 & ~n47746 ;
  assign n47748 = ~n47738 & ~n47747 ;
  assign n47749 = n47738 & n47747 ;
  assign n47750 = ~n47748 & ~n47749 ;
  assign n47751 = ~n47467 & ~n47469 ;
  assign n47752 = ~n47373 & ~n47376 ;
  assign n47753 = ~x104 & n22325 ;
  assign n47754 = ~x102 & n23066 ;
  assign n47755 = ~x103 & n22320 ;
  assign n47756 = ~n47754 & ~n47755 ;
  assign n47757 = ~n47753 & n47756 ;
  assign n47758 = n11380 & n22328 ;
  assign n47759 = n47757 & ~n47758 ;
  assign n47760 = ~x59 & ~n47759 ;
  assign n47761 = ~x59 & ~n47760 ;
  assign n47762 = ~n47759 & ~n47760 ;
  assign n47763 = ~n47761 & ~n47762 ;
  assign n47764 = ~n47347 & ~n47358 ;
  assign n47765 = ~n47344 & ~n47764 ;
  assign n47766 = ~x97 & n27427 ;
  assign n47767 = ~x98 & ~n26217 ;
  assign n47768 = ~n47766 & ~n47767 ;
  assign n47769 = ~n47337 & ~n47340 ;
  assign n47770 = ~n47768 & n47769 ;
  assign n47771 = n47768 & ~n47769 ;
  assign n47772 = ~n47770 & ~n47771 ;
  assign n47773 = ~x101 & n24612 ;
  assign n47774 = ~x99 & n25390 ;
  assign n47775 = ~x100 & n24607 ;
  assign n47776 = ~n47774 & ~n47775 ;
  assign n47777 = ~n47773 & n47776 ;
  assign n47778 = n9844 & n24615 ;
  assign n47779 = n47777 & ~n47778 ;
  assign n47780 = ~x62 & ~n47779 ;
  assign n47781 = ~x62 & ~n47780 ;
  assign n47782 = ~n47779 & ~n47780 ;
  assign n47783 = ~n47781 & ~n47782 ;
  assign n47784 = ~n47772 & n47783 ;
  assign n47785 = n47772 & ~n47783 ;
  assign n47786 = ~n47784 & ~n47785 ;
  assign n47787 = ~n47765 & n47786 ;
  assign n47788 = ~n47765 & ~n47787 ;
  assign n47789 = n47786 & ~n47787 ;
  assign n47790 = ~n47788 & ~n47789 ;
  assign n47791 = ~n47763 & ~n47790 ;
  assign n47792 = n47763 & ~n47789 ;
  assign n47793 = ~n47788 & n47792 ;
  assign n47794 = ~n47791 & ~n47793 ;
  assign n47795 = ~n47752 & n47794 ;
  assign n47796 = n47752 & ~n47794 ;
  assign n47797 = ~n47795 & ~n47796 ;
  assign n47798 = ~x107 & n20143 ;
  assign n47799 = ~x105 & n20854 ;
  assign n47800 = ~x106 & n20138 ;
  assign n47801 = ~n47799 & ~n47800 ;
  assign n47802 = ~n47798 & n47801 ;
  assign n47803 = n13034 & n20146 ;
  assign n47804 = n47802 & ~n47803 ;
  assign n47805 = ~x56 & ~n47804 ;
  assign n47806 = ~x56 & ~n47805 ;
  assign n47807 = ~n47804 & ~n47805 ;
  assign n47808 = ~n47806 & ~n47807 ;
  assign n47809 = n47797 & ~n47808 ;
  assign n47810 = n47797 & ~n47809 ;
  assign n47811 = ~n47808 & ~n47809 ;
  assign n47812 = ~n47810 & ~n47811 ;
  assign n47813 = ~n47390 & ~n47396 ;
  assign n47814 = n47812 & n47813 ;
  assign n47815 = ~n47812 & ~n47813 ;
  assign n47816 = ~n47814 & ~n47815 ;
  assign n47817 = ~x110 & n18025 ;
  assign n47818 = ~x108 & n18764 ;
  assign n47819 = ~x109 & n18020 ;
  assign n47820 = ~n47818 & ~n47819 ;
  assign n47821 = ~n47817 & n47820 ;
  assign n47822 = n14802 & n18028 ;
  assign n47823 = n47821 & ~n47822 ;
  assign n47824 = ~x53 & ~n47823 ;
  assign n47825 = ~x53 & ~n47824 ;
  assign n47826 = ~n47823 & ~n47824 ;
  assign n47827 = ~n47825 & ~n47826 ;
  assign n47828 = n47816 & ~n47827 ;
  assign n47829 = n47816 & ~n47828 ;
  assign n47830 = ~n47827 & ~n47828 ;
  assign n47831 = ~n47829 & ~n47830 ;
  assign n47832 = ~n47409 & ~n47415 ;
  assign n47833 = n47831 & n47832 ;
  assign n47834 = ~n47831 & ~n47832 ;
  assign n47835 = ~n47833 & ~n47834 ;
  assign n47836 = ~x113 & n16076 ;
  assign n47837 = ~x111 & n16756 ;
  assign n47838 = ~x112 & n16071 ;
  assign n47839 = ~n47837 & ~n47838 ;
  assign n47840 = ~n47836 & n47839 ;
  assign n47841 = n16079 & n16684 ;
  assign n47842 = n47840 & ~n47841 ;
  assign n47843 = ~x50 & ~n47842 ;
  assign n47844 = ~x50 & ~n47843 ;
  assign n47845 = ~n47842 & ~n47843 ;
  assign n47846 = ~n47844 & ~n47845 ;
  assign n47847 = n47835 & ~n47846 ;
  assign n47848 = n47835 & ~n47847 ;
  assign n47849 = ~n47846 & ~n47847 ;
  assign n47850 = ~n47848 & ~n47849 ;
  assign n47851 = ~n47428 & ~n47434 ;
  assign n47852 = n47850 & n47851 ;
  assign n47853 = ~n47850 & ~n47851 ;
  assign n47854 = ~n47852 & ~n47853 ;
  assign n47855 = ~x116 & n14233 ;
  assign n47856 = ~x114 & n14876 ;
  assign n47857 = ~x115 & n14228 ;
  assign n47858 = ~n47856 & ~n47857 ;
  assign n47859 = ~n47855 & n47858 ;
  assign n47860 = n14236 & n18678 ;
  assign n47861 = n47859 & ~n47860 ;
  assign n47862 = ~x47 & ~n47861 ;
  assign n47863 = ~x47 & ~n47862 ;
  assign n47864 = ~n47861 & ~n47862 ;
  assign n47865 = ~n47863 & ~n47864 ;
  assign n47866 = n47854 & ~n47865 ;
  assign n47867 = n47854 & ~n47866 ;
  assign n47868 = ~n47865 & ~n47866 ;
  assign n47869 = ~n47867 & ~n47868 ;
  assign n47870 = ~n47452 & n47869 ;
  assign n47871 = n47452 & ~n47869 ;
  assign n47872 = ~n47870 & ~n47871 ;
  assign n47873 = ~x119 & n12506 ;
  assign n47874 = ~x117 & n13131 ;
  assign n47875 = ~x118 & n12501 ;
  assign n47876 = ~n47874 & ~n47875 ;
  assign n47877 = ~n47873 & n47876 ;
  assign n47878 = n12509 & n20778 ;
  assign n47879 = n47877 & ~n47878 ;
  assign n47880 = ~x44 & ~n47879 ;
  assign n47881 = ~x44 & ~n47880 ;
  assign n47882 = ~n47879 & ~n47880 ;
  assign n47883 = ~n47881 & ~n47882 ;
  assign n47884 = ~n47872 & ~n47883 ;
  assign n47885 = n47872 & n47883 ;
  assign n47886 = ~n47884 & ~n47885 ;
  assign n47887 = ~n47751 & n47886 ;
  assign n47888 = n47751 & ~n47886 ;
  assign n47889 = ~n47887 & ~n47888 ;
  assign n47890 = ~x122 & n10905 ;
  assign n47891 = ~x120 & n11466 ;
  assign n47892 = ~x121 & n10900 ;
  assign n47893 = ~n47891 & ~n47892 ;
  assign n47894 = ~n47890 & n47893 ;
  assign n47895 = n10908 & n22998 ;
  assign n47896 = n47894 & ~n47895 ;
  assign n47897 = ~x41 & ~n47896 ;
  assign n47898 = ~x41 & ~n47897 ;
  assign n47899 = ~n47896 & ~n47897 ;
  assign n47900 = ~n47898 & ~n47899 ;
  assign n47901 = n47889 & ~n47900 ;
  assign n47902 = n47889 & ~n47901 ;
  assign n47903 = ~n47900 & ~n47901 ;
  assign n47904 = ~n47902 & ~n47903 ;
  assign n47905 = ~n47483 & ~n47489 ;
  assign n47906 = n47904 & n47905 ;
  assign n47907 = ~n47904 & ~n47905 ;
  assign n47908 = ~n47906 & ~n47907 ;
  assign n47909 = ~x125 & n9433 ;
  assign n47910 = ~x123 & n9915 ;
  assign n47911 = ~x124 & n9428 ;
  assign n47912 = ~n47910 & ~n47911 ;
  assign n47913 = ~n47909 & n47912 ;
  assign n47914 = n9436 & n25330 ;
  assign n47915 = n47913 & ~n47914 ;
  assign n47916 = ~x38 & ~n47915 ;
  assign n47917 = ~x38 & ~n47916 ;
  assign n47918 = ~n47915 & ~n47916 ;
  assign n47919 = ~n47917 & ~n47918 ;
  assign n47920 = n47908 & ~n47919 ;
  assign n47921 = ~n47908 & n47919 ;
  assign n47922 = n47750 & ~n47921 ;
  assign n47923 = ~n47920 & n47922 ;
  assign n47924 = n47750 & ~n47923 ;
  assign n47925 = ~n47921 & ~n47923 ;
  assign n47926 = ~n47920 & n47925 ;
  assign n47927 = ~n47924 & ~n47926 ;
  assign n47928 = ~n47522 & ~n47527 ;
  assign n47929 = ~n47927 & ~n47928 ;
  assign n47930 = ~n47927 & ~n47929 ;
  assign n47931 = ~n47928 & ~n47929 ;
  assign n47932 = ~n47930 & ~n47931 ;
  assign n47933 = ~n47529 & ~n47532 ;
  assign n47934 = ~n47932 & ~n47933 ;
  assign n47935 = n47932 & n47933 ;
  assign n47936 = ~n47934 & ~n47935 ;
  assign n47939 = ~n47936 & ~x225 ;
  assign n47940 = ~n47938 & ~n47939 ;
  assign n47941 = ~n47730 & ~n47735 ;
  assign n47942 = ~n47549 & ~n47724 ;
  assign n47943 = ~n47708 & ~n47721 ;
  assign n47944 = x127 & n8474 ;
  assign n47945 = n8009 & n26962 ;
  assign n47946 = ~n47944 & ~n47945 ;
  assign n47947 = x35 & ~n47946 ;
  assign n47948 = x35 & ~n47947 ;
  assign n47949 = ~n47946 & ~n47947 ;
  assign n47950 = ~n47948 & ~n47949 ;
  assign n47951 = ~n47943 & ~n47950 ;
  assign n47952 = ~n47943 & ~n47951 ;
  assign n47953 = ~n47950 & ~n47951 ;
  assign n47954 = ~n47952 & ~n47953 ;
  assign n47955 = ~n47244 & ~n47670 ;
  assign n47956 = ~n47685 & ~n47955 ;
  assign n47957 = x120 & n12506 ;
  assign n47958 = x118 & n13131 ;
  assign n47959 = x119 & n12501 ;
  assign n47960 = ~n47958 & ~n47959 ;
  assign n47961 = ~n47957 & n47960 ;
  assign n47962 = n12509 & n21143 ;
  assign n47963 = n47961 & ~n47962 ;
  assign n47964 = x44 & ~n47963 ;
  assign n47965 = x44 & ~n47964 ;
  assign n47966 = ~n47963 & ~n47964 ;
  assign n47967 = ~n47965 & ~n47966 ;
  assign n47968 = ~n47654 & ~n47667 ;
  assign n47969 = x117 & n14233 ;
  assign n47970 = x115 & n14876 ;
  assign n47971 = x116 & n14228 ;
  assign n47972 = ~n47970 & ~n47971 ;
  assign n47973 = ~n47969 & n47972 ;
  assign n47974 = n14236 & n19026 ;
  assign n47975 = n47973 & ~n47974 ;
  assign n47976 = x47 & ~n47975 ;
  assign n47977 = x47 & ~n47976 ;
  assign n47978 = ~n47975 & ~n47976 ;
  assign n47979 = ~n47977 & ~n47978 ;
  assign n47980 = ~n47635 & ~n47648 ;
  assign n47981 = ~n47596 & ~n47610 ;
  assign n47982 = x108 & n20143 ;
  assign n47983 = x106 & n20854 ;
  assign n47984 = x107 & n20138 ;
  assign n47985 = ~n47983 & ~n47984 ;
  assign n47986 = ~n47982 & n47985 ;
  assign n47987 = n13323 & n20146 ;
  assign n47988 = n47986 & ~n47987 ;
  assign n47989 = x56 & ~n47988 ;
  assign n47990 = x56 & ~n47989 ;
  assign n47991 = ~n47988 & ~n47989 ;
  assign n47992 = ~n47990 & ~n47991 ;
  assign n47993 = ~n47588 & ~n47592 ;
  assign n47994 = ~n47572 & ~n47586 ;
  assign n47995 = x98 & n27024 ;
  assign n47996 = x99 & ~n26217 ;
  assign n47997 = ~n47995 & ~n47996 ;
  assign n47998 = ~n47569 & n47997 ;
  assign n47999 = n47569 & ~n47997 ;
  assign n48000 = ~n47994 & ~n47999 ;
  assign n48001 = ~n47998 & n48000 ;
  assign n48002 = ~n47994 & ~n48001 ;
  assign n48003 = ~n47998 & ~n48001 ;
  assign n48004 = ~n47999 & n48003 ;
  assign n48005 = ~n48002 & ~n48004 ;
  assign n48006 = x102 & n24612 ;
  assign n48007 = x100 & n25390 ;
  assign n48008 = x101 & n24607 ;
  assign n48009 = ~n48007 & ~n48008 ;
  assign n48010 = ~n48006 & n48009 ;
  assign n48011 = n10092 & n24615 ;
  assign n48012 = n48010 & ~n48011 ;
  assign n48013 = x62 & ~n48012 ;
  assign n48014 = x62 & ~n48013 ;
  assign n48015 = ~n48012 & ~n48013 ;
  assign n48016 = ~n48014 & ~n48015 ;
  assign n48017 = ~n48005 & ~n48016 ;
  assign n48018 = ~n48005 & ~n48017 ;
  assign n48019 = ~n48016 & ~n48017 ;
  assign n48020 = ~n48018 & ~n48019 ;
  assign n48021 = x105 & n22325 ;
  assign n48022 = x103 & n23066 ;
  assign n48023 = x104 & n22320 ;
  assign n48024 = ~n48022 & ~n48023 ;
  assign n48025 = ~n48021 & n48024 ;
  assign n48026 = n11648 & n22328 ;
  assign n48027 = n48025 & ~n48026 ;
  assign n48028 = x59 & ~n48027 ;
  assign n48029 = x59 & ~n48028 ;
  assign n48030 = ~n48027 & ~n48028 ;
  assign n48031 = ~n48029 & ~n48030 ;
  assign n48032 = ~n48020 & n48031 ;
  assign n48033 = n48020 & ~n48031 ;
  assign n48034 = ~n48032 & ~n48033 ;
  assign n48035 = ~n47993 & ~n48034 ;
  assign n48036 = n47993 & n48034 ;
  assign n48037 = ~n48035 & ~n48036 ;
  assign n48038 = ~n47992 & n48037 ;
  assign n48039 = n47992 & ~n48037 ;
  assign n48040 = ~n48038 & ~n48039 ;
  assign n48041 = ~n47981 & n48040 ;
  assign n48042 = n47981 & ~n48040 ;
  assign n48043 = ~n48041 & ~n48042 ;
  assign n48044 = x111 & n18025 ;
  assign n48045 = x109 & n18764 ;
  assign n48046 = x110 & n18020 ;
  assign n48047 = ~n48045 & ~n48046 ;
  assign n48048 = ~n48044 & n48047 ;
  assign n48049 = n15111 & n18028 ;
  assign n48050 = n48048 & ~n48049 ;
  assign n48051 = x53 & ~n48050 ;
  assign n48052 = x53 & ~n48051 ;
  assign n48053 = ~n48050 & ~n48051 ;
  assign n48054 = ~n48052 & ~n48053 ;
  assign n48055 = n48043 & ~n48054 ;
  assign n48056 = n48043 & ~n48055 ;
  assign n48057 = ~n48054 & ~n48055 ;
  assign n48058 = ~n48056 & ~n48057 ;
  assign n48059 = ~n47616 & ~n47629 ;
  assign n48060 = n48058 & n48059 ;
  assign n48061 = ~n48058 & ~n48059 ;
  assign n48062 = ~n48060 & ~n48061 ;
  assign n48063 = x114 & n16076 ;
  assign n48064 = x112 & n16756 ;
  assign n48065 = x113 & n16071 ;
  assign n48066 = ~n48064 & ~n48065 ;
  assign n48067 = ~n48063 & n48066 ;
  assign n48068 = n16079 & n17012 ;
  assign n48069 = n48067 & ~n48068 ;
  assign n48070 = x50 & ~n48069 ;
  assign n48071 = x50 & ~n48070 ;
  assign n48072 = ~n48069 & ~n48070 ;
  assign n48073 = ~n48071 & ~n48072 ;
  assign n48074 = ~n48062 & n48073 ;
  assign n48075 = n48062 & ~n48073 ;
  assign n48076 = ~n48074 & ~n48075 ;
  assign n48077 = ~n47980 & n48076 ;
  assign n48078 = ~n47980 & ~n48077 ;
  assign n48079 = n48076 & ~n48077 ;
  assign n48080 = ~n48078 & ~n48079 ;
  assign n48081 = ~n47979 & ~n48080 ;
  assign n48082 = n47979 & ~n48079 ;
  assign n48083 = ~n48078 & n48082 ;
  assign n48084 = ~n48081 & ~n48083 ;
  assign n48085 = ~n47968 & n48084 ;
  assign n48086 = n47968 & ~n48084 ;
  assign n48087 = ~n48085 & ~n48086 ;
  assign n48088 = ~n47967 & n48087 ;
  assign n48089 = n47967 & ~n48087 ;
  assign n48090 = ~n48088 & ~n48089 ;
  assign n48091 = ~n47956 & n48090 ;
  assign n48092 = n47956 & ~n48090 ;
  assign n48093 = ~n48091 & ~n48092 ;
  assign n48094 = x123 & n10905 ;
  assign n48095 = x121 & n11466 ;
  assign n48096 = x122 & n10900 ;
  assign n48097 = ~n48095 & ~n48096 ;
  assign n48098 = ~n48094 & n48097 ;
  assign n48099 = n10908 & n23382 ;
  assign n48100 = n48098 & ~n48099 ;
  assign n48101 = x41 & ~n48100 ;
  assign n48102 = x41 & ~n48101 ;
  assign n48103 = ~n48100 & ~n48101 ;
  assign n48104 = ~n48102 & ~n48103 ;
  assign n48105 = n48093 & ~n48104 ;
  assign n48106 = n48093 & ~n48105 ;
  assign n48107 = ~n48104 & ~n48105 ;
  assign n48108 = ~n48106 & ~n48107 ;
  assign n48109 = ~n47688 & ~n47702 ;
  assign n48110 = n48108 & n48109 ;
  assign n48111 = ~n48108 & ~n48109 ;
  assign n48112 = ~n48110 & ~n48111 ;
  assign n48113 = x126 & n9433 ;
  assign n48114 = x124 & n9915 ;
  assign n48115 = x125 & n9428 ;
  assign n48116 = ~n48114 & ~n48115 ;
  assign n48117 = ~n48113 & n48116 ;
  assign n48118 = n9436 & n25735 ;
  assign n48119 = n48117 & ~n48118 ;
  assign n48120 = x38 & ~n48119 ;
  assign n48121 = x38 & ~n48120 ;
  assign n48122 = ~n48119 & ~n48120 ;
  assign n48123 = ~n48121 & ~n48122 ;
  assign n48124 = n48112 & ~n48123 ;
  assign n48125 = n48112 & ~n48124 ;
  assign n48126 = ~n48123 & ~n48124 ;
  assign n48127 = ~n48125 & ~n48126 ;
  assign n48128 = ~n47954 & n48127 ;
  assign n48129 = n47954 & ~n48127 ;
  assign n48130 = ~n48128 & ~n48129 ;
  assign n48131 = ~n47942 & ~n48130 ;
  assign n48132 = n47942 & n48130 ;
  assign n48133 = ~n48131 & ~n48132 ;
  assign n48134 = ~n47941 & n48133 ;
  assign n48135 = n47941 & ~n48133 ;
  assign n48136 = ~n48134 & ~n48135 ;
  assign n48334 = n48136 & x226 ;
  assign n48137 = ~n47929 & ~n47934 ;
  assign n48138 = ~n47748 & ~n47923 ;
  assign n48139 = ~n47907 & ~n47920 ;
  assign n48140 = ~x127 & n8474 ;
  assign n48141 = n8009 & n27365 ;
  assign n48142 = ~n48140 & ~n48141 ;
  assign n48143 = ~x35 & ~n48142 ;
  assign n48144 = ~x35 & ~n48143 ;
  assign n48145 = ~n48142 & ~n48143 ;
  assign n48146 = ~n48144 & ~n48145 ;
  assign n48147 = ~n48139 & ~n48146 ;
  assign n48148 = ~n48139 & ~n48147 ;
  assign n48149 = ~n48146 & ~n48147 ;
  assign n48150 = ~n48148 & ~n48149 ;
  assign n48151 = ~n47452 & ~n47869 ;
  assign n48152 = ~n47884 & ~n48151 ;
  assign n48153 = ~x120 & n12506 ;
  assign n48154 = ~x118 & n13131 ;
  assign n48155 = ~x119 & n12501 ;
  assign n48156 = ~n48154 & ~n48155 ;
  assign n48157 = ~n48153 & n48156 ;
  assign n48158 = n12509 & n21501 ;
  assign n48159 = n48157 & ~n48158 ;
  assign n48160 = ~x44 & ~n48159 ;
  assign n48161 = ~x44 & ~n48160 ;
  assign n48162 = ~n48159 & ~n48160 ;
  assign n48163 = ~n48161 & ~n48162 ;
  assign n48164 = ~n47853 & ~n47866 ;
  assign n48165 = ~x117 & n14233 ;
  assign n48166 = ~x115 & n14876 ;
  assign n48167 = ~x116 & n14228 ;
  assign n48168 = ~n48166 & ~n48167 ;
  assign n48169 = ~n48165 & n48168 ;
  assign n48170 = n14236 & n19365 ;
  assign n48171 = n48169 & ~n48170 ;
  assign n48172 = ~x47 & ~n48171 ;
  assign n48173 = ~x47 & ~n48172 ;
  assign n48174 = ~n48171 & ~n48172 ;
  assign n48175 = ~n48173 & ~n48174 ;
  assign n48176 = ~n47834 & ~n47847 ;
  assign n48177 = ~n47795 & ~n47809 ;
  assign n48178 = ~x108 & n20143 ;
  assign n48179 = ~x106 & n20854 ;
  assign n48180 = ~x107 & n20138 ;
  assign n48181 = ~n48179 & ~n48180 ;
  assign n48182 = ~n48178 & n48181 ;
  assign n48183 = n13601 & n20146 ;
  assign n48184 = n48182 & ~n48183 ;
  assign n48185 = ~x56 & ~n48184 ;
  assign n48186 = ~x56 & ~n48185 ;
  assign n48187 = ~n48184 & ~n48185 ;
  assign n48188 = ~n48186 & ~n48187 ;
  assign n48189 = ~n47787 & ~n47791 ;
  assign n48190 = ~n47771 & ~n47785 ;
  assign n48191 = ~x98 & n27427 ;
  assign n48192 = ~x99 & ~n26217 ;
  assign n48193 = ~n48191 & ~n48192 ;
  assign n48194 = ~n47768 & n48193 ;
  assign n48195 = n47768 & ~n48193 ;
  assign n48196 = ~n48190 & ~n48195 ;
  assign n48197 = ~n48194 & n48196 ;
  assign n48198 = ~n48190 & ~n48197 ;
  assign n48199 = ~n48194 & ~n48197 ;
  assign n48200 = ~n48195 & n48199 ;
  assign n48201 = ~n48198 & ~n48200 ;
  assign n48202 = ~x102 & n24612 ;
  assign n48203 = ~x100 & n25390 ;
  assign n48204 = ~x101 & n24607 ;
  assign n48205 = ~n48203 & ~n48204 ;
  assign n48206 = ~n48202 & n48205 ;
  assign n48207 = n10333 & n24615 ;
  assign n48208 = n48206 & ~n48207 ;
  assign n48209 = ~x62 & ~n48208 ;
  assign n48210 = ~x62 & ~n48209 ;
  assign n48211 = ~n48208 & ~n48209 ;
  assign n48212 = ~n48210 & ~n48211 ;
  assign n48213 = ~n48201 & ~n48212 ;
  assign n48214 = ~n48201 & ~n48213 ;
  assign n48215 = ~n48212 & ~n48213 ;
  assign n48216 = ~n48214 & ~n48215 ;
  assign n48217 = ~x105 & n22325 ;
  assign n48218 = ~x103 & n23066 ;
  assign n48219 = ~x104 & n22320 ;
  assign n48220 = ~n48218 & ~n48219 ;
  assign n48221 = ~n48217 & n48220 ;
  assign n48222 = n11907 & n22328 ;
  assign n48223 = n48221 & ~n48222 ;
  assign n48224 = ~x59 & ~n48223 ;
  assign n48225 = ~x59 & ~n48224 ;
  assign n48226 = ~n48223 & ~n48224 ;
  assign n48227 = ~n48225 & ~n48226 ;
  assign n48228 = ~n48216 & n48227 ;
  assign n48229 = n48216 & ~n48227 ;
  assign n48230 = ~n48228 & ~n48229 ;
  assign n48231 = ~n48189 & ~n48230 ;
  assign n48232 = n48189 & n48230 ;
  assign n48233 = ~n48231 & ~n48232 ;
  assign n48234 = ~n48188 & n48233 ;
  assign n48235 = n48188 & ~n48233 ;
  assign n48236 = ~n48234 & ~n48235 ;
  assign n48237 = ~n48177 & n48236 ;
  assign n48238 = n48177 & ~n48236 ;
  assign n48239 = ~n48237 & ~n48238 ;
  assign n48240 = ~x111 & n18025 ;
  assign n48241 = ~x109 & n18764 ;
  assign n48242 = ~x110 & n18020 ;
  assign n48243 = ~n48241 & ~n48242 ;
  assign n48244 = ~n48240 & n48243 ;
  assign n48245 = n15411 & n18028 ;
  assign n48246 = n48244 & ~n48245 ;
  assign n48247 = ~x53 & ~n48246 ;
  assign n48248 = ~x53 & ~n48247 ;
  assign n48249 = ~n48246 & ~n48247 ;
  assign n48250 = ~n48248 & ~n48249 ;
  assign n48251 = n48239 & ~n48250 ;
  assign n48252 = n48239 & ~n48251 ;
  assign n48253 = ~n48250 & ~n48251 ;
  assign n48254 = ~n48252 & ~n48253 ;
  assign n48255 = ~n47815 & ~n47828 ;
  assign n48256 = n48254 & n48255 ;
  assign n48257 = ~n48254 & ~n48255 ;
  assign n48258 = ~n48256 & ~n48257 ;
  assign n48259 = ~x114 & n16076 ;
  assign n48260 = ~x112 & n16756 ;
  assign n48261 = ~x113 & n16071 ;
  assign n48262 = ~n48260 & ~n48261 ;
  assign n48263 = ~n48259 & n48262 ;
  assign n48264 = n16079 & n17333 ;
  assign n48265 = n48263 & ~n48264 ;
  assign n48266 = ~x50 & ~n48265 ;
  assign n48267 = ~x50 & ~n48266 ;
  assign n48268 = ~n48265 & ~n48266 ;
  assign n48269 = ~n48267 & ~n48268 ;
  assign n48270 = ~n48258 & n48269 ;
  assign n48271 = n48258 & ~n48269 ;
  assign n48272 = ~n48270 & ~n48271 ;
  assign n48273 = ~n48176 & n48272 ;
  assign n48274 = ~n48176 & ~n48273 ;
  assign n48275 = n48272 & ~n48273 ;
  assign n48276 = ~n48274 & ~n48275 ;
  assign n48277 = ~n48175 & ~n48276 ;
  assign n48278 = n48175 & ~n48275 ;
  assign n48279 = ~n48274 & n48278 ;
  assign n48280 = ~n48277 & ~n48279 ;
  assign n48281 = ~n48164 & n48280 ;
  assign n48282 = n48164 & ~n48280 ;
  assign n48283 = ~n48281 & ~n48282 ;
  assign n48284 = ~n48163 & n48283 ;
  assign n48285 = n48163 & ~n48283 ;
  assign n48286 = ~n48284 & ~n48285 ;
  assign n48287 = ~n48152 & n48286 ;
  assign n48288 = n48152 & ~n48286 ;
  assign n48289 = ~n48287 & ~n48288 ;
  assign n48290 = ~x123 & n10905 ;
  assign n48291 = ~x121 & n11466 ;
  assign n48292 = ~x122 & n10900 ;
  assign n48293 = ~n48291 & ~n48292 ;
  assign n48294 = ~n48290 & n48293 ;
  assign n48295 = n10908 & n23760 ;
  assign n48296 = n48294 & ~n48295 ;
  assign n48297 = ~x41 & ~n48296 ;
  assign n48298 = ~x41 & ~n48297 ;
  assign n48299 = ~n48296 & ~n48297 ;
  assign n48300 = ~n48298 & ~n48299 ;
  assign n48301 = n48289 & ~n48300 ;
  assign n48302 = n48289 & ~n48301 ;
  assign n48303 = ~n48300 & ~n48301 ;
  assign n48304 = ~n48302 & ~n48303 ;
  assign n48305 = ~n47887 & ~n47901 ;
  assign n48306 = n48304 & n48305 ;
  assign n48307 = ~n48304 & ~n48305 ;
  assign n48308 = ~n48306 & ~n48307 ;
  assign n48309 = ~x126 & n9433 ;
  assign n48310 = ~x124 & n9915 ;
  assign n48311 = ~x125 & n9428 ;
  assign n48312 = ~n48310 & ~n48311 ;
  assign n48313 = ~n48309 & n48312 ;
  assign n48314 = n9436 & n26128 ;
  assign n48315 = n48313 & ~n48314 ;
  assign n48316 = ~x38 & ~n48315 ;
  assign n48317 = ~x38 & ~n48316 ;
  assign n48318 = ~n48315 & ~n48316 ;
  assign n48319 = ~n48317 & ~n48318 ;
  assign n48320 = n48308 & ~n48319 ;
  assign n48321 = n48308 & ~n48320 ;
  assign n48322 = ~n48319 & ~n48320 ;
  assign n48323 = ~n48321 & ~n48322 ;
  assign n48324 = ~n48150 & n48323 ;
  assign n48325 = n48150 & ~n48323 ;
  assign n48326 = ~n48324 & ~n48325 ;
  assign n48327 = ~n48138 & ~n48326 ;
  assign n48328 = n48138 & n48326 ;
  assign n48329 = ~n48327 & ~n48328 ;
  assign n48330 = ~n48137 & n48329 ;
  assign n48331 = n48137 & ~n48329 ;
  assign n48332 = ~n48330 & ~n48331 ;
  assign n48335 = ~n48332 & ~x226 ;
  assign n48336 = ~n48334 & ~n48335 ;
  assign n48337 = ~n48131 & ~n48134 ;
  assign n48338 = ~n48077 & ~n48081 ;
  assign n48339 = x118 & n14233 ;
  assign n48340 = x116 & n14876 ;
  assign n48341 = x117 & n14228 ;
  assign n48342 = ~n48340 & ~n48341 ;
  assign n48343 = ~n48339 & n48342 ;
  assign n48344 = n14236 & n19395 ;
  assign n48345 = n48343 & ~n48344 ;
  assign n48346 = x47 & ~n48345 ;
  assign n48347 = x47 & ~n48346 ;
  assign n48348 = ~n48345 & ~n48346 ;
  assign n48349 = ~n48347 & ~n48348 ;
  assign n48350 = ~n48061 & ~n48075 ;
  assign n48351 = x99 & n27024 ;
  assign n48352 = x100 & ~n26217 ;
  assign n48353 = ~n48351 & ~n48352 ;
  assign n48354 = x35 & ~n47997 ;
  assign n48355 = ~x35 & n47997 ;
  assign n48356 = ~n48354 & ~n48355 ;
  assign n48357 = ~n48353 & ~n48356 ;
  assign n48358 = n48353 & n48356 ;
  assign n48359 = ~n48357 & ~n48358 ;
  assign n48360 = ~n48003 & n48359 ;
  assign n48361 = n48003 & ~n48359 ;
  assign n48362 = ~n48360 & ~n48361 ;
  assign n48363 = x103 & n24612 ;
  assign n48364 = x101 & n25390 ;
  assign n48365 = x102 & n24607 ;
  assign n48366 = ~n48364 & ~n48365 ;
  assign n48367 = ~n48363 & n48366 ;
  assign n48368 = n10588 & n24615 ;
  assign n48369 = n48367 & ~n48368 ;
  assign n48370 = x62 & ~n48369 ;
  assign n48371 = x62 & ~n48370 ;
  assign n48372 = ~n48369 & ~n48370 ;
  assign n48373 = ~n48371 & ~n48372 ;
  assign n48374 = ~n48362 & n48373 ;
  assign n48375 = n48362 & ~n48373 ;
  assign n48376 = ~n48374 & ~n48375 ;
  assign n48377 = x106 & n22325 ;
  assign n48378 = x104 & n23066 ;
  assign n48379 = x105 & n22320 ;
  assign n48380 = ~n48378 & ~n48379 ;
  assign n48381 = ~n48377 & n48380 ;
  assign n48382 = n12181 & n22328 ;
  assign n48383 = n48381 & ~n48382 ;
  assign n48384 = x59 & ~n48383 ;
  assign n48385 = x59 & ~n48384 ;
  assign n48386 = ~n48383 & ~n48384 ;
  assign n48387 = ~n48385 & ~n48386 ;
  assign n48388 = n48376 & ~n48387 ;
  assign n48389 = n48376 & ~n48388 ;
  assign n48390 = ~n48387 & ~n48388 ;
  assign n48391 = ~n48389 & ~n48390 ;
  assign n48392 = ~n48020 & ~n48031 ;
  assign n48393 = ~n48017 & ~n48392 ;
  assign n48394 = ~n48391 & ~n48393 ;
  assign n48395 = ~n48391 & ~n48394 ;
  assign n48396 = ~n48393 & ~n48394 ;
  assign n48397 = ~n48395 & ~n48396 ;
  assign n48398 = x109 & n20143 ;
  assign n48399 = x107 & n20854 ;
  assign n48400 = x108 & n20138 ;
  assign n48401 = ~n48399 & ~n48400 ;
  assign n48402 = ~n48398 & n48401 ;
  assign n48403 = n13894 & n20146 ;
  assign n48404 = n48402 & ~n48403 ;
  assign n48405 = x56 & ~n48404 ;
  assign n48406 = x56 & ~n48405 ;
  assign n48407 = ~n48404 & ~n48405 ;
  assign n48408 = ~n48406 & ~n48407 ;
  assign n48409 = ~n48397 & ~n48408 ;
  assign n48410 = ~n48397 & ~n48409 ;
  assign n48411 = ~n48408 & ~n48409 ;
  assign n48412 = ~n48410 & ~n48411 ;
  assign n48413 = ~n48035 & ~n48038 ;
  assign n48414 = n48412 & n48413 ;
  assign n48415 = ~n48412 & ~n48413 ;
  assign n48416 = ~n48414 & ~n48415 ;
  assign n48417 = x112 & n18025 ;
  assign n48418 = x110 & n18764 ;
  assign n48419 = x111 & n18020 ;
  assign n48420 = ~n48418 & ~n48419 ;
  assign n48421 = ~n48417 & n48420 ;
  assign n48422 = n15442 & n18028 ;
  assign n48423 = n48421 & ~n48422 ;
  assign n48424 = x53 & ~n48423 ;
  assign n48425 = x53 & ~n48424 ;
  assign n48426 = ~n48423 & ~n48424 ;
  assign n48427 = ~n48425 & ~n48426 ;
  assign n48428 = n48416 & ~n48427 ;
  assign n48429 = n48416 & ~n48428 ;
  assign n48430 = ~n48427 & ~n48428 ;
  assign n48431 = ~n48429 & ~n48430 ;
  assign n48432 = ~n48041 & ~n48055 ;
  assign n48433 = n48431 & n48432 ;
  assign n48434 = ~n48431 & ~n48432 ;
  assign n48435 = ~n48433 & ~n48434 ;
  assign n48436 = x115 & n16076 ;
  assign n48437 = x113 & n16756 ;
  assign n48438 = x114 & n16071 ;
  assign n48439 = ~n48437 & ~n48438 ;
  assign n48440 = ~n48436 & n48439 ;
  assign n48441 = n16079 & n17364 ;
  assign n48442 = n48440 & ~n48441 ;
  assign n48443 = x50 & ~n48442 ;
  assign n48444 = x50 & ~n48443 ;
  assign n48445 = ~n48442 & ~n48443 ;
  assign n48446 = ~n48444 & ~n48445 ;
  assign n48447 = ~n48435 & n48446 ;
  assign n48448 = n48435 & ~n48446 ;
  assign n48449 = ~n48447 & ~n48448 ;
  assign n48450 = ~n48350 & n48449 ;
  assign n48451 = n48350 & ~n48449 ;
  assign n48452 = ~n48450 & ~n48451 ;
  assign n48453 = ~n48349 & n48452 ;
  assign n48454 = n48349 & ~n48452 ;
  assign n48455 = ~n48453 & ~n48454 ;
  assign n48456 = ~n48338 & n48455 ;
  assign n48457 = n48338 & ~n48455 ;
  assign n48458 = ~n48456 & ~n48457 ;
  assign n48459 = x121 & n12506 ;
  assign n48460 = x119 & n13131 ;
  assign n48461 = x120 & n12501 ;
  assign n48462 = ~n48460 & ~n48461 ;
  assign n48463 = ~n48459 & n48462 ;
  assign n48464 = n12509 & n21870 ;
  assign n48465 = n48463 & ~n48464 ;
  assign n48466 = x44 & ~n48465 ;
  assign n48467 = x44 & ~n48466 ;
  assign n48468 = ~n48465 & ~n48466 ;
  assign n48469 = ~n48467 & ~n48468 ;
  assign n48470 = n48458 & ~n48469 ;
  assign n48471 = n48458 & ~n48470 ;
  assign n48472 = ~n48469 & ~n48470 ;
  assign n48473 = ~n48471 & ~n48472 ;
  assign n48474 = ~n48085 & ~n48088 ;
  assign n48475 = n48473 & n48474 ;
  assign n48476 = ~n48473 & ~n48474 ;
  assign n48477 = ~n48475 & ~n48476 ;
  assign n48478 = x124 & n10905 ;
  assign n48479 = x122 & n11466 ;
  assign n48480 = x123 & n10900 ;
  assign n48481 = ~n48479 & ~n48480 ;
  assign n48482 = ~n48478 & n48481 ;
  assign n48483 = n10908 & n23796 ;
  assign n48484 = n48482 & ~n48483 ;
  assign n48485 = x41 & ~n48484 ;
  assign n48486 = x41 & ~n48485 ;
  assign n48487 = ~n48484 & ~n48485 ;
  assign n48488 = ~n48486 & ~n48487 ;
  assign n48489 = n48477 & ~n48488 ;
  assign n48490 = n48477 & ~n48489 ;
  assign n48491 = ~n48488 & ~n48489 ;
  assign n48492 = ~n48490 & ~n48491 ;
  assign n48493 = ~n48091 & ~n48105 ;
  assign n48494 = n48492 & n48493 ;
  assign n48495 = ~n48492 & ~n48493 ;
  assign n48496 = ~n48494 & ~n48495 ;
  assign n48497 = x127 & n9433 ;
  assign n48498 = x125 & n9915 ;
  assign n48499 = x126 & n9428 ;
  assign n48500 = ~n48498 & ~n48499 ;
  assign n48501 = ~n48497 & n48500 ;
  assign n48502 = n9436 & n26533 ;
  assign n48503 = n48501 & ~n48502 ;
  assign n48504 = x38 & ~n48503 ;
  assign n48505 = x38 & ~n48504 ;
  assign n48506 = ~n48503 & ~n48504 ;
  assign n48507 = ~n48505 & ~n48506 ;
  assign n48508 = n48496 & ~n48507 ;
  assign n48509 = n48496 & ~n48508 ;
  assign n48510 = ~n48507 & ~n48508 ;
  assign n48511 = ~n48509 & ~n48510 ;
  assign n48512 = ~n48111 & ~n48124 ;
  assign n48513 = n48511 & n48512 ;
  assign n48514 = ~n48511 & ~n48512 ;
  assign n48515 = ~n48513 & ~n48514 ;
  assign n48516 = ~n47954 & ~n48127 ;
  assign n48517 = ~n47951 & ~n48516 ;
  assign n48518 = n48515 & ~n48517 ;
  assign n48519 = ~n48515 & n48517 ;
  assign n48520 = ~n48518 & ~n48519 ;
  assign n48521 = ~n48337 & n48520 ;
  assign n48522 = n48337 & ~n48520 ;
  assign n48523 = ~n48521 & ~n48522 ;
  assign n48712 = n48523 & x227 ;
  assign n48524 = ~n48327 & ~n48330 ;
  assign n48525 = ~n48273 & ~n48277 ;
  assign n48526 = ~x118 & n14233 ;
  assign n48527 = ~x116 & n14876 ;
  assign n48528 = ~x117 & n14228 ;
  assign n48529 = ~n48527 & ~n48528 ;
  assign n48530 = ~n48526 & n48529 ;
  assign n48531 = n14236 & n19736 ;
  assign n48532 = n48530 & ~n48531 ;
  assign n48533 = ~x47 & ~n48532 ;
  assign n48534 = ~x47 & ~n48533 ;
  assign n48535 = ~n48532 & ~n48533 ;
  assign n48536 = ~n48534 & ~n48535 ;
  assign n48537 = ~n48257 & ~n48271 ;
  assign n48538 = ~x99 & n27427 ;
  assign n48539 = ~x100 & ~n26217 ;
  assign n48540 = ~n48538 & ~n48539 ;
  assign n48541 = ~x35 & ~n48193 ;
  assign n48542 = x35 & n48193 ;
  assign n48543 = ~n48541 & ~n48542 ;
  assign n48544 = ~n48540 & ~n48543 ;
  assign n48545 = n48540 & n48543 ;
  assign n48546 = ~n48544 & ~n48545 ;
  assign n48547 = ~n48199 & n48546 ;
  assign n48548 = n48199 & ~n48546 ;
  assign n48549 = ~n48547 & ~n48548 ;
  assign n48550 = ~x103 & n24612 ;
  assign n48551 = ~x101 & n25390 ;
  assign n48552 = ~x102 & n24607 ;
  assign n48553 = ~n48551 & ~n48552 ;
  assign n48554 = ~n48550 & n48553 ;
  assign n48555 = n10833 & n24615 ;
  assign n48556 = n48554 & ~n48555 ;
  assign n48557 = ~x62 & ~n48556 ;
  assign n48558 = ~x62 & ~n48557 ;
  assign n48559 = ~n48556 & ~n48557 ;
  assign n48560 = ~n48558 & ~n48559 ;
  assign n48561 = ~n48549 & n48560 ;
  assign n48562 = n48549 & ~n48560 ;
  assign n48563 = ~n48561 & ~n48562 ;
  assign n48564 = ~x106 & n22325 ;
  assign n48565 = ~x104 & n23066 ;
  assign n48566 = ~x105 & n22320 ;
  assign n48567 = ~n48565 & ~n48566 ;
  assign n48568 = ~n48564 & n48567 ;
  assign n48569 = n12447 & n22328 ;
  assign n48570 = n48568 & ~n48569 ;
  assign n48571 = ~x59 & ~n48570 ;
  assign n48572 = ~x59 & ~n48571 ;
  assign n48573 = ~n48570 & ~n48571 ;
  assign n48574 = ~n48572 & ~n48573 ;
  assign n48575 = n48563 & ~n48574 ;
  assign n48576 = n48563 & ~n48575 ;
  assign n48577 = ~n48574 & ~n48575 ;
  assign n48578 = ~n48576 & ~n48577 ;
  assign n48579 = ~n48216 & ~n48227 ;
  assign n48580 = ~n48213 & ~n48579 ;
  assign n48581 = ~n48578 & ~n48580 ;
  assign n48582 = ~n48578 & ~n48581 ;
  assign n48583 = ~n48580 & ~n48581 ;
  assign n48584 = ~n48582 & ~n48583 ;
  assign n48585 = ~x109 & n20143 ;
  assign n48586 = ~x107 & n20854 ;
  assign n48587 = ~x108 & n20138 ;
  assign n48588 = ~n48586 & ~n48587 ;
  assign n48589 = ~n48585 & n48588 ;
  assign n48590 = n14177 & n20146 ;
  assign n48591 = n48589 & ~n48590 ;
  assign n48592 = ~x56 & ~n48591 ;
  assign n48593 = ~x56 & ~n48592 ;
  assign n48594 = ~n48591 & ~n48592 ;
  assign n48595 = ~n48593 & ~n48594 ;
  assign n48596 = ~n48584 & ~n48595 ;
  assign n48597 = ~n48584 & ~n48596 ;
  assign n48598 = ~n48595 & ~n48596 ;
  assign n48599 = ~n48597 & ~n48598 ;
  assign n48600 = ~n48231 & ~n48234 ;
  assign n48601 = n48599 & n48600 ;
  assign n48602 = ~n48599 & ~n48600 ;
  assign n48603 = ~n48601 & ~n48602 ;
  assign n48604 = ~x112 & n18025 ;
  assign n48605 = ~x110 & n18764 ;
  assign n48606 = ~x111 & n18020 ;
  assign n48607 = ~n48605 & ~n48606 ;
  assign n48608 = ~n48604 & n48607 ;
  assign n48609 = n15744 & n18028 ;
  assign n48610 = n48608 & ~n48609 ;
  assign n48611 = ~x53 & ~n48610 ;
  assign n48612 = ~x53 & ~n48611 ;
  assign n48613 = ~n48610 & ~n48611 ;
  assign n48614 = ~n48612 & ~n48613 ;
  assign n48615 = n48603 & ~n48614 ;
  assign n48616 = n48603 & ~n48615 ;
  assign n48617 = ~n48614 & ~n48615 ;
  assign n48618 = ~n48616 & ~n48617 ;
  assign n48619 = ~n48237 & ~n48251 ;
  assign n48620 = n48618 & n48619 ;
  assign n48621 = ~n48618 & ~n48619 ;
  assign n48622 = ~n48620 & ~n48621 ;
  assign n48623 = ~x115 & n16076 ;
  assign n48624 = ~x113 & n16756 ;
  assign n48625 = ~x114 & n16071 ;
  assign n48626 = ~n48624 & ~n48625 ;
  assign n48627 = ~n48623 & n48626 ;
  assign n48628 = n16079 & n17683 ;
  assign n48629 = n48627 & ~n48628 ;
  assign n48630 = ~x50 & ~n48629 ;
  assign n48631 = ~x50 & ~n48630 ;
  assign n48632 = ~n48629 & ~n48630 ;
  assign n48633 = ~n48631 & ~n48632 ;
  assign n48634 = ~n48622 & n48633 ;
  assign n48635 = n48622 & ~n48633 ;
  assign n48636 = ~n48634 & ~n48635 ;
  assign n48637 = ~n48537 & n48636 ;
  assign n48638 = n48537 & ~n48636 ;
  assign n48639 = ~n48637 & ~n48638 ;
  assign n48640 = ~n48536 & n48639 ;
  assign n48641 = n48536 & ~n48639 ;
  assign n48642 = ~n48640 & ~n48641 ;
  assign n48643 = ~n48525 & n48642 ;
  assign n48644 = n48525 & ~n48642 ;
  assign n48645 = ~n48643 & ~n48644 ;
  assign n48646 = ~x121 & n12506 ;
  assign n48647 = ~x119 & n13131 ;
  assign n48648 = ~x120 & n12501 ;
  assign n48649 = ~n48647 & ~n48648 ;
  assign n48650 = ~n48646 & n48649 ;
  assign n48651 = n12509 & n22229 ;
  assign n48652 = n48650 & ~n48651 ;
  assign n48653 = ~x44 & ~n48652 ;
  assign n48654 = ~x44 & ~n48653 ;
  assign n48655 = ~n48652 & ~n48653 ;
  assign n48656 = ~n48654 & ~n48655 ;
  assign n48657 = n48645 & ~n48656 ;
  assign n48658 = n48645 & ~n48657 ;
  assign n48659 = ~n48656 & ~n48657 ;
  assign n48660 = ~n48658 & ~n48659 ;
  assign n48661 = ~n48281 & ~n48284 ;
  assign n48662 = n48660 & n48661 ;
  assign n48663 = ~n48660 & ~n48661 ;
  assign n48664 = ~n48662 & ~n48663 ;
  assign n48665 = ~x124 & n10905 ;
  assign n48666 = ~x122 & n11466 ;
  assign n48667 = ~x123 & n10900 ;
  assign n48668 = ~n48666 & ~n48667 ;
  assign n48669 = ~n48665 & n48668 ;
  assign n48670 = n10908 & n24176 ;
  assign n48671 = n48669 & ~n48670 ;
  assign n48672 = ~x41 & ~n48671 ;
  assign n48673 = ~x41 & ~n48672 ;
  assign n48674 = ~n48671 & ~n48672 ;
  assign n48675 = ~n48673 & ~n48674 ;
  assign n48676 = n48664 & ~n48675 ;
  assign n48677 = n48664 & ~n48676 ;
  assign n48678 = ~n48675 & ~n48676 ;
  assign n48679 = ~n48677 & ~n48678 ;
  assign n48680 = ~n48287 & ~n48301 ;
  assign n48681 = n48679 & n48680 ;
  assign n48682 = ~n48679 & ~n48680 ;
  assign n48683 = ~n48681 & ~n48682 ;
  assign n48684 = ~x127 & n9433 ;
  assign n48685 = ~x125 & n9915 ;
  assign n48686 = ~x126 & n9428 ;
  assign n48687 = ~n48685 & ~n48686 ;
  assign n48688 = ~n48684 & n48687 ;
  assign n48689 = n9436 & n26932 ;
  assign n48690 = n48688 & ~n48689 ;
  assign n48691 = ~x38 & ~n48690 ;
  assign n48692 = ~x38 & ~n48691 ;
  assign n48693 = ~n48690 & ~n48691 ;
  assign n48694 = ~n48692 & ~n48693 ;
  assign n48695 = n48683 & ~n48694 ;
  assign n48696 = n48683 & ~n48695 ;
  assign n48697 = ~n48694 & ~n48695 ;
  assign n48698 = ~n48696 & ~n48697 ;
  assign n48699 = ~n48307 & ~n48320 ;
  assign n48700 = n48698 & n48699 ;
  assign n48701 = ~n48698 & ~n48699 ;
  assign n48702 = ~n48700 & ~n48701 ;
  assign n48703 = ~n48150 & ~n48323 ;
  assign n48704 = ~n48147 & ~n48703 ;
  assign n48705 = n48702 & ~n48704 ;
  assign n48706 = ~n48702 & n48704 ;
  assign n48707 = ~n48705 & ~n48706 ;
  assign n48708 = ~n48524 & n48707 ;
  assign n48709 = n48524 & ~n48707 ;
  assign n48710 = ~n48708 & ~n48709 ;
  assign n48713 = ~n48710 & ~x227 ;
  assign n48714 = ~n48712 & ~n48713 ;
  assign n48715 = ~n48489 & ~n48495 ;
  assign n48716 = x126 & n9915 ;
  assign n48717 = x127 & n9428 ;
  assign n48718 = ~n48716 & ~n48717 ;
  assign n48719 = ~n9436 & n48718 ;
  assign n48720 = n26965 & n48718 ;
  assign n48721 = ~n48719 & ~n48720 ;
  assign n48722 = x38 & ~n48721 ;
  assign n48723 = ~x38 & n48721 ;
  assign n48724 = ~n48722 & ~n48723 ;
  assign n48725 = ~n48715 & ~n48724 ;
  assign n48726 = n48715 & n48724 ;
  assign n48727 = ~n48725 & ~n48726 ;
  assign n48728 = x104 & n24612 ;
  assign n48729 = x102 & n25390 ;
  assign n48730 = x103 & n24607 ;
  assign n48731 = ~n48729 & ~n48730 ;
  assign n48732 = ~n48728 & n48731 ;
  assign n48733 = n11116 & n24615 ;
  assign n48734 = n48732 & ~n48733 ;
  assign n48735 = x62 & ~n48734 ;
  assign n48736 = x62 & ~n48735 ;
  assign n48737 = ~n48734 & ~n48735 ;
  assign n48738 = ~n48736 & ~n48737 ;
  assign n48739 = x100 & n27024 ;
  assign n48740 = x101 & ~n26217 ;
  assign n48741 = ~n48739 & ~n48740 ;
  assign n48742 = ~x35 & ~n47997 ;
  assign n48743 = ~n48357 & ~n48742 ;
  assign n48744 = n48741 & ~n48743 ;
  assign n48745 = n48741 & ~n48744 ;
  assign n48746 = ~n48743 & ~n48744 ;
  assign n48747 = ~n48745 & ~n48746 ;
  assign n48748 = ~n48738 & ~n48747 ;
  assign n48749 = ~n48738 & ~n48748 ;
  assign n48750 = ~n48747 & ~n48748 ;
  assign n48751 = ~n48749 & ~n48750 ;
  assign n48752 = ~n48360 & ~n48375 ;
  assign n48753 = n48751 & n48752 ;
  assign n48754 = ~n48751 & ~n48752 ;
  assign n48755 = ~n48753 & ~n48754 ;
  assign n48756 = x107 & n22325 ;
  assign n48757 = x105 & n23066 ;
  assign n48758 = x106 & n22320 ;
  assign n48759 = ~n48757 & ~n48758 ;
  assign n48760 = ~n48756 & n48759 ;
  assign n48761 = n12749 & n22328 ;
  assign n48762 = n48760 & ~n48761 ;
  assign n48763 = x59 & ~n48762 ;
  assign n48764 = x59 & ~n48763 ;
  assign n48765 = ~n48762 & ~n48763 ;
  assign n48766 = ~n48764 & ~n48765 ;
  assign n48767 = n48755 & ~n48766 ;
  assign n48768 = n48755 & ~n48767 ;
  assign n48769 = ~n48766 & ~n48767 ;
  assign n48770 = ~n48768 & ~n48769 ;
  assign n48771 = ~n48388 & ~n48394 ;
  assign n48772 = n48770 & n48771 ;
  assign n48773 = ~n48770 & ~n48771 ;
  assign n48774 = ~n48772 & ~n48773 ;
  assign n48775 = x110 & n20143 ;
  assign n48776 = x108 & n20854 ;
  assign n48777 = x109 & n20138 ;
  assign n48778 = ~n48776 & ~n48777 ;
  assign n48779 = ~n48775 & n48778 ;
  assign n48780 = n14497 & n20146 ;
  assign n48781 = n48779 & ~n48780 ;
  assign n48782 = x56 & ~n48781 ;
  assign n48783 = x56 & ~n48782 ;
  assign n48784 = ~n48781 & ~n48782 ;
  assign n48785 = ~n48783 & ~n48784 ;
  assign n48786 = n48774 & ~n48785 ;
  assign n48787 = n48774 & ~n48786 ;
  assign n48788 = ~n48785 & ~n48786 ;
  assign n48789 = ~n48787 & ~n48788 ;
  assign n48790 = ~n48409 & ~n48415 ;
  assign n48791 = n48789 & n48790 ;
  assign n48792 = ~n48789 & ~n48790 ;
  assign n48793 = ~n48791 & ~n48792 ;
  assign n48794 = x113 & n18025 ;
  assign n48795 = x111 & n18764 ;
  assign n48796 = x112 & n18020 ;
  assign n48797 = ~n48795 & ~n48796 ;
  assign n48798 = ~n48794 & n48797 ;
  assign n48799 = n16361 & n18028 ;
  assign n48800 = n48798 & ~n48799 ;
  assign n48801 = x53 & ~n48800 ;
  assign n48802 = x53 & ~n48801 ;
  assign n48803 = ~n48800 & ~n48801 ;
  assign n48804 = ~n48802 & ~n48803 ;
  assign n48805 = n48793 & ~n48804 ;
  assign n48806 = n48793 & ~n48805 ;
  assign n48807 = ~n48804 & ~n48805 ;
  assign n48808 = ~n48806 & ~n48807 ;
  assign n48809 = ~n48428 & ~n48434 ;
  assign n48810 = n48808 & n48809 ;
  assign n48811 = ~n48808 & ~n48809 ;
  assign n48812 = ~n48810 & ~n48811 ;
  assign n48813 = x116 & n16076 ;
  assign n48814 = x114 & n16756 ;
  assign n48815 = x115 & n16071 ;
  assign n48816 = ~n48814 & ~n48815 ;
  assign n48817 = ~n48813 & n48816 ;
  assign n48818 = n16079 & n18336 ;
  assign n48819 = n48817 & ~n48818 ;
  assign n48820 = x50 & ~n48819 ;
  assign n48821 = x50 & ~n48820 ;
  assign n48822 = ~n48819 & ~n48820 ;
  assign n48823 = ~n48821 & ~n48822 ;
  assign n48824 = n48812 & ~n48823 ;
  assign n48825 = n48812 & ~n48824 ;
  assign n48826 = ~n48823 & ~n48824 ;
  assign n48827 = ~n48825 & ~n48826 ;
  assign n48828 = ~n48448 & ~n48450 ;
  assign n48829 = ~n48827 & ~n48828 ;
  assign n48830 = ~n48827 & ~n48829 ;
  assign n48831 = ~n48828 & ~n48829 ;
  assign n48832 = ~n48830 & ~n48831 ;
  assign n48833 = x119 & n14233 ;
  assign n48834 = x117 & n14876 ;
  assign n48835 = x118 & n14228 ;
  assign n48836 = ~n48834 & ~n48835 ;
  assign n48837 = ~n48833 & n48836 ;
  assign n48838 = n14236 & n20423 ;
  assign n48839 = n48837 & ~n48838 ;
  assign n48840 = x47 & ~n48839 ;
  assign n48841 = x47 & ~n48840 ;
  assign n48842 = ~n48839 & ~n48840 ;
  assign n48843 = ~n48841 & ~n48842 ;
  assign n48844 = ~n48832 & ~n48843 ;
  assign n48845 = ~n48832 & ~n48844 ;
  assign n48846 = ~n48843 & ~n48844 ;
  assign n48847 = ~n48845 & ~n48846 ;
  assign n48848 = ~n48453 & ~n48456 ;
  assign n48849 = n48847 & n48848 ;
  assign n48850 = ~n48847 & ~n48848 ;
  assign n48851 = ~n48849 & ~n48850 ;
  assign n48852 = x122 & n12506 ;
  assign n48853 = x120 & n13131 ;
  assign n48854 = x121 & n12501 ;
  assign n48855 = ~n48853 & ~n48854 ;
  assign n48856 = ~n48852 & n48855 ;
  assign n48857 = n12509 & n22622 ;
  assign n48858 = n48856 & ~n48857 ;
  assign n48859 = x44 & ~n48858 ;
  assign n48860 = x44 & ~n48859 ;
  assign n48861 = ~n48858 & ~n48859 ;
  assign n48862 = ~n48860 & ~n48861 ;
  assign n48863 = n48851 & ~n48862 ;
  assign n48864 = n48851 & ~n48863 ;
  assign n48865 = ~n48862 & ~n48863 ;
  assign n48866 = ~n48864 & ~n48865 ;
  assign n48867 = ~n48470 & ~n48476 ;
  assign n48868 = n48866 & n48867 ;
  assign n48869 = ~n48866 & ~n48867 ;
  assign n48870 = ~n48868 & ~n48869 ;
  assign n48871 = x125 & n10905 ;
  assign n48872 = x123 & n11466 ;
  assign n48873 = x124 & n10900 ;
  assign n48874 = ~n48872 & ~n48873 ;
  assign n48875 = ~n48871 & n48874 ;
  assign n48876 = n10908 & n24935 ;
  assign n48877 = n48875 & ~n48876 ;
  assign n48878 = x41 & ~n48877 ;
  assign n48879 = x41 & ~n48878 ;
  assign n48880 = ~n48877 & ~n48878 ;
  assign n48881 = ~n48879 & ~n48880 ;
  assign n48882 = n48870 & ~n48881 ;
  assign n48883 = ~n48870 & n48881 ;
  assign n48884 = n48727 & ~n48883 ;
  assign n48885 = ~n48882 & n48884 ;
  assign n48886 = n48727 & ~n48885 ;
  assign n48887 = ~n48883 & ~n48885 ;
  assign n48888 = ~n48882 & n48887 ;
  assign n48889 = ~n48886 & ~n48888 ;
  assign n48890 = ~n48508 & ~n48514 ;
  assign n48891 = n48889 & n48890 ;
  assign n48892 = ~n48889 & ~n48890 ;
  assign n48893 = ~n48891 & ~n48892 ;
  assign n48894 = ~n48518 & ~n48521 ;
  assign n48895 = n48893 & ~n48894 ;
  assign n48896 = ~n48893 & n48894 ;
  assign n48897 = ~n48895 & ~n48896 ;
  assign n49082 = n48897 & x228 ;
  assign n48898 = ~n48676 & ~n48682 ;
  assign n48899 = ~x126 & n9915 ;
  assign n48900 = ~x127 & n9428 ;
  assign n48901 = ~n48899 & ~n48900 ;
  assign n48902 = ~n9436 & n48901 ;
  assign n48903 = n27368 & n48901 ;
  assign n48904 = ~n48902 & ~n48903 ;
  assign n48905 = ~x38 & ~n48904 ;
  assign n48906 = x38 & n48904 ;
  assign n48907 = ~n48905 & ~n48906 ;
  assign n48908 = ~n48898 & ~n48907 ;
  assign n48909 = n48898 & n48907 ;
  assign n48910 = ~n48908 & ~n48909 ;
  assign n48911 = ~x104 & n24612 ;
  assign n48912 = ~x102 & n25390 ;
  assign n48913 = ~x103 & n24607 ;
  assign n48914 = ~n48912 & ~n48913 ;
  assign n48915 = ~n48911 & n48914 ;
  assign n48916 = n11380 & n24615 ;
  assign n48917 = n48915 & ~n48916 ;
  assign n48918 = ~x62 & ~n48917 ;
  assign n48919 = ~x62 & ~n48918 ;
  assign n48920 = ~n48917 & ~n48918 ;
  assign n48921 = ~n48919 & ~n48920 ;
  assign n48922 = ~x100 & n27427 ;
  assign n48923 = ~x101 & ~n26217 ;
  assign n48924 = ~n48922 & ~n48923 ;
  assign n48925 = x35 & ~n48193 ;
  assign n48926 = ~n48544 & ~n48925 ;
  assign n48927 = n48924 & ~n48926 ;
  assign n48928 = n48924 & ~n48927 ;
  assign n48929 = ~n48926 & ~n48927 ;
  assign n48930 = ~n48928 & ~n48929 ;
  assign n48931 = ~n48921 & ~n48930 ;
  assign n48932 = ~n48921 & ~n48931 ;
  assign n48933 = ~n48930 & ~n48931 ;
  assign n48934 = ~n48932 & ~n48933 ;
  assign n48935 = ~n48547 & ~n48562 ;
  assign n48936 = n48934 & n48935 ;
  assign n48937 = ~n48934 & ~n48935 ;
  assign n48938 = ~n48936 & ~n48937 ;
  assign n48939 = ~x107 & n22325 ;
  assign n48940 = ~x105 & n23066 ;
  assign n48941 = ~x106 & n22320 ;
  assign n48942 = ~n48940 & ~n48941 ;
  assign n48943 = ~n48939 & n48942 ;
  assign n48944 = n13034 & n22328 ;
  assign n48945 = n48943 & ~n48944 ;
  assign n48946 = ~x59 & ~n48945 ;
  assign n48947 = ~x59 & ~n48946 ;
  assign n48948 = ~n48945 & ~n48946 ;
  assign n48949 = ~n48947 & ~n48948 ;
  assign n48950 = n48938 & ~n48949 ;
  assign n48951 = n48938 & ~n48950 ;
  assign n48952 = ~n48949 & ~n48950 ;
  assign n48953 = ~n48951 & ~n48952 ;
  assign n48954 = ~n48575 & ~n48581 ;
  assign n48955 = n48953 & n48954 ;
  assign n48956 = ~n48953 & ~n48954 ;
  assign n48957 = ~n48955 & ~n48956 ;
  assign n48958 = ~x110 & n20143 ;
  assign n48959 = ~x108 & n20854 ;
  assign n48960 = ~x109 & n20138 ;
  assign n48961 = ~n48959 & ~n48960 ;
  assign n48962 = ~n48958 & n48961 ;
  assign n48963 = n14802 & n20146 ;
  assign n48964 = n48962 & ~n48963 ;
  assign n48965 = ~x56 & ~n48964 ;
  assign n48966 = ~x56 & ~n48965 ;
  assign n48967 = ~n48964 & ~n48965 ;
  assign n48968 = ~n48966 & ~n48967 ;
  assign n48969 = n48957 & ~n48968 ;
  assign n48970 = n48957 & ~n48969 ;
  assign n48971 = ~n48968 & ~n48969 ;
  assign n48972 = ~n48970 & ~n48971 ;
  assign n48973 = ~n48596 & ~n48602 ;
  assign n48974 = n48972 & n48973 ;
  assign n48975 = ~n48972 & ~n48973 ;
  assign n48976 = ~n48974 & ~n48975 ;
  assign n48977 = ~x113 & n18025 ;
  assign n48978 = ~x111 & n18764 ;
  assign n48979 = ~x112 & n18020 ;
  assign n48980 = ~n48978 & ~n48979 ;
  assign n48981 = ~n48977 & n48980 ;
  assign n48982 = n16684 & n18028 ;
  assign n48983 = n48981 & ~n48982 ;
  assign n48984 = ~x53 & ~n48983 ;
  assign n48985 = ~x53 & ~n48984 ;
  assign n48986 = ~n48983 & ~n48984 ;
  assign n48987 = ~n48985 & ~n48986 ;
  assign n48988 = n48976 & ~n48987 ;
  assign n48989 = n48976 & ~n48988 ;
  assign n48990 = ~n48987 & ~n48988 ;
  assign n48991 = ~n48989 & ~n48990 ;
  assign n48992 = ~n48615 & ~n48621 ;
  assign n48993 = n48991 & n48992 ;
  assign n48994 = ~n48991 & ~n48992 ;
  assign n48995 = ~n48993 & ~n48994 ;
  assign n48996 = ~x116 & n16076 ;
  assign n48997 = ~x114 & n16756 ;
  assign n48998 = ~x115 & n16071 ;
  assign n48999 = ~n48997 & ~n48998 ;
  assign n49000 = ~n48996 & n48999 ;
  assign n49001 = n16079 & n18678 ;
  assign n49002 = n49000 & ~n49001 ;
  assign n49003 = ~x50 & ~n49002 ;
  assign n49004 = ~x50 & ~n49003 ;
  assign n49005 = ~n49002 & ~n49003 ;
  assign n49006 = ~n49004 & ~n49005 ;
  assign n49007 = n48995 & ~n49006 ;
  assign n49008 = n48995 & ~n49007 ;
  assign n49009 = ~n49006 & ~n49007 ;
  assign n49010 = ~n49008 & ~n49009 ;
  assign n49011 = ~n48635 & ~n48637 ;
  assign n49012 = ~n49010 & ~n49011 ;
  assign n49013 = ~n49010 & ~n49012 ;
  assign n49014 = ~n49011 & ~n49012 ;
  assign n49015 = ~n49013 & ~n49014 ;
  assign n49016 = ~x119 & n14233 ;
  assign n49017 = ~x117 & n14876 ;
  assign n49018 = ~x118 & n14228 ;
  assign n49019 = ~n49017 & ~n49018 ;
  assign n49020 = ~n49016 & n49019 ;
  assign n49021 = n14236 & n20778 ;
  assign n49022 = n49020 & ~n49021 ;
  assign n49023 = ~x47 & ~n49022 ;
  assign n49024 = ~x47 & ~n49023 ;
  assign n49025 = ~n49022 & ~n49023 ;
  assign n49026 = ~n49024 & ~n49025 ;
  assign n49027 = ~n49015 & ~n49026 ;
  assign n49028 = ~n49015 & ~n49027 ;
  assign n49029 = ~n49026 & ~n49027 ;
  assign n49030 = ~n49028 & ~n49029 ;
  assign n49031 = ~n48640 & ~n48643 ;
  assign n49032 = n49030 & n49031 ;
  assign n49033 = ~n49030 & ~n49031 ;
  assign n49034 = ~n49032 & ~n49033 ;
  assign n49035 = ~x122 & n12506 ;
  assign n49036 = ~x120 & n13131 ;
  assign n49037 = ~x121 & n12501 ;
  assign n49038 = ~n49036 & ~n49037 ;
  assign n49039 = ~n49035 & n49038 ;
  assign n49040 = n12509 & n22998 ;
  assign n49041 = n49039 & ~n49040 ;
  assign n49042 = ~x44 & ~n49041 ;
  assign n49043 = ~x44 & ~n49042 ;
  assign n49044 = ~n49041 & ~n49042 ;
  assign n49045 = ~n49043 & ~n49044 ;
  assign n49046 = n49034 & ~n49045 ;
  assign n49047 = n49034 & ~n49046 ;
  assign n49048 = ~n49045 & ~n49046 ;
  assign n49049 = ~n49047 & ~n49048 ;
  assign n49050 = ~n48657 & ~n48663 ;
  assign n49051 = n49049 & n49050 ;
  assign n49052 = ~n49049 & ~n49050 ;
  assign n49053 = ~n49051 & ~n49052 ;
  assign n49054 = ~x125 & n10905 ;
  assign n49055 = ~x123 & n11466 ;
  assign n49056 = ~x124 & n10900 ;
  assign n49057 = ~n49055 & ~n49056 ;
  assign n49058 = ~n49054 & n49057 ;
  assign n49059 = n10908 & n25330 ;
  assign n49060 = n49058 & ~n49059 ;
  assign n49061 = ~x41 & ~n49060 ;
  assign n49062 = ~x41 & ~n49061 ;
  assign n49063 = ~n49060 & ~n49061 ;
  assign n49064 = ~n49062 & ~n49063 ;
  assign n49065 = n49053 & ~n49064 ;
  assign n49066 = ~n49053 & n49064 ;
  assign n49067 = n48910 & ~n49066 ;
  assign n49068 = ~n49065 & n49067 ;
  assign n49069 = n48910 & ~n49068 ;
  assign n49070 = ~n49066 & ~n49068 ;
  assign n49071 = ~n49065 & n49070 ;
  assign n49072 = ~n49069 & ~n49071 ;
  assign n49073 = ~n48695 & ~n48701 ;
  assign n49074 = n49072 & n49073 ;
  assign n49075 = ~n49072 & ~n49073 ;
  assign n49076 = ~n49074 & ~n49075 ;
  assign n49077 = ~n48705 & ~n48708 ;
  assign n49078 = n49076 & ~n49077 ;
  assign n49079 = ~n49076 & n49077 ;
  assign n49080 = ~n49078 & ~n49079 ;
  assign n49083 = ~n49080 & ~x228 ;
  assign n49084 = ~n49082 & ~n49083 ;
  assign n49085 = ~n48892 & ~n48895 ;
  assign n49086 = ~n48725 & ~n48885 ;
  assign n49087 = ~n48869 & ~n48882 ;
  assign n49088 = x127 & n9915 ;
  assign n49089 = n9436 & n26962 ;
  assign n49090 = ~n49088 & ~n49089 ;
  assign n49091 = x38 & ~n49090 ;
  assign n49092 = x38 & ~n49091 ;
  assign n49093 = ~n49090 & ~n49091 ;
  assign n49094 = ~n49092 & ~n49093 ;
  assign n49095 = ~n49087 & ~n49094 ;
  assign n49096 = ~n49087 & ~n49095 ;
  assign n49097 = ~n49094 & ~n49095 ;
  assign n49098 = ~n49096 & ~n49097 ;
  assign n49099 = ~n48829 & ~n48844 ;
  assign n49100 = x120 & n14233 ;
  assign n49101 = x118 & n14876 ;
  assign n49102 = x119 & n14228 ;
  assign n49103 = ~n49101 & ~n49102 ;
  assign n49104 = ~n49100 & n49103 ;
  assign n49105 = n14236 & n21143 ;
  assign n49106 = n49104 & ~n49105 ;
  assign n49107 = x47 & ~n49106 ;
  assign n49108 = x47 & ~n49107 ;
  assign n49109 = ~n49106 & ~n49107 ;
  assign n49110 = ~n49108 & ~n49109 ;
  assign n49111 = ~n48811 & ~n48824 ;
  assign n49112 = x117 & n16076 ;
  assign n49113 = x115 & n16756 ;
  assign n49114 = x116 & n16071 ;
  assign n49115 = ~n49113 & ~n49114 ;
  assign n49116 = ~n49112 & n49115 ;
  assign n49117 = n16079 & n19026 ;
  assign n49118 = n49116 & ~n49117 ;
  assign n49119 = x50 & ~n49118 ;
  assign n49120 = x50 & ~n49119 ;
  assign n49121 = ~n49118 & ~n49119 ;
  assign n49122 = ~n49120 & ~n49121 ;
  assign n49123 = ~n48792 & ~n48805 ;
  assign n49124 = ~n48744 & ~n48748 ;
  assign n49125 = x101 & n27024 ;
  assign n49126 = x102 & ~n26217 ;
  assign n49127 = ~n49125 & ~n49126 ;
  assign n49128 = n48741 & ~n49127 ;
  assign n49129 = n48741 & ~n49128 ;
  assign n49130 = ~n49127 & ~n49128 ;
  assign n49131 = ~n49129 & ~n49130 ;
  assign n49132 = ~n49124 & ~n49131 ;
  assign n49133 = ~n49124 & ~n49132 ;
  assign n49134 = ~n49131 & ~n49132 ;
  assign n49135 = ~n49133 & ~n49134 ;
  assign n49136 = x105 & n24612 ;
  assign n49137 = x103 & n25390 ;
  assign n49138 = x104 & n24607 ;
  assign n49139 = ~n49137 & ~n49138 ;
  assign n49140 = ~n49136 & n49139 ;
  assign n49141 = n11648 & n24615 ;
  assign n49142 = n49140 & ~n49141 ;
  assign n49143 = x62 & ~n49142 ;
  assign n49144 = x62 & ~n49143 ;
  assign n49145 = ~n49142 & ~n49143 ;
  assign n49146 = ~n49144 & ~n49145 ;
  assign n49147 = ~n49135 & ~n49146 ;
  assign n49148 = ~n49135 & ~n49147 ;
  assign n49149 = ~n49146 & ~n49147 ;
  assign n49150 = ~n49148 & ~n49149 ;
  assign n49151 = x108 & n22325 ;
  assign n49152 = x106 & n23066 ;
  assign n49153 = x107 & n22320 ;
  assign n49154 = ~n49152 & ~n49153 ;
  assign n49155 = ~n49151 & n49154 ;
  assign n49156 = n13323 & n22328 ;
  assign n49157 = n49155 & ~n49156 ;
  assign n49158 = x59 & ~n49157 ;
  assign n49159 = x59 & ~n49158 ;
  assign n49160 = ~n49157 & ~n49158 ;
  assign n49161 = ~n49159 & ~n49160 ;
  assign n49162 = ~n49150 & n49161 ;
  assign n49163 = n49150 & ~n49161 ;
  assign n49164 = ~n49162 & ~n49163 ;
  assign n49165 = ~n48754 & ~n48767 ;
  assign n49166 = n49164 & n49165 ;
  assign n49167 = ~n49164 & ~n49165 ;
  assign n49168 = ~n49166 & ~n49167 ;
  assign n49169 = x111 & n20143 ;
  assign n49170 = x109 & n20854 ;
  assign n49171 = x110 & n20138 ;
  assign n49172 = ~n49170 & ~n49171 ;
  assign n49173 = ~n49169 & n49172 ;
  assign n49174 = n15111 & n20146 ;
  assign n49175 = n49173 & ~n49174 ;
  assign n49176 = x56 & ~n49175 ;
  assign n49177 = x56 & ~n49176 ;
  assign n49178 = ~n49175 & ~n49176 ;
  assign n49179 = ~n49177 & ~n49178 ;
  assign n49180 = n49168 & ~n49179 ;
  assign n49181 = n49168 & ~n49180 ;
  assign n49182 = ~n49179 & ~n49180 ;
  assign n49183 = ~n49181 & ~n49182 ;
  assign n49184 = ~n48773 & ~n48786 ;
  assign n49185 = n49183 & n49184 ;
  assign n49186 = ~n49183 & ~n49184 ;
  assign n49187 = ~n49185 & ~n49186 ;
  assign n49188 = x114 & n18025 ;
  assign n49189 = x112 & n18764 ;
  assign n49190 = x113 & n18020 ;
  assign n49191 = ~n49189 & ~n49190 ;
  assign n49192 = ~n49188 & n49191 ;
  assign n49193 = n17012 & n18028 ;
  assign n49194 = n49192 & ~n49193 ;
  assign n49195 = x53 & ~n49194 ;
  assign n49196 = x53 & ~n49195 ;
  assign n49197 = ~n49194 & ~n49195 ;
  assign n49198 = ~n49196 & ~n49197 ;
  assign n49199 = ~n49187 & n49198 ;
  assign n49200 = n49187 & ~n49198 ;
  assign n49201 = ~n49199 & ~n49200 ;
  assign n49202 = ~n49123 & n49201 ;
  assign n49203 = ~n49123 & ~n49202 ;
  assign n49204 = n49201 & ~n49202 ;
  assign n49205 = ~n49203 & ~n49204 ;
  assign n49206 = ~n49122 & ~n49205 ;
  assign n49207 = n49122 & ~n49204 ;
  assign n49208 = ~n49203 & n49207 ;
  assign n49209 = ~n49206 & ~n49208 ;
  assign n49210 = ~n49111 & n49209 ;
  assign n49211 = n49111 & ~n49209 ;
  assign n49212 = ~n49210 & ~n49211 ;
  assign n49213 = ~n49110 & n49212 ;
  assign n49214 = n49110 & ~n49212 ;
  assign n49215 = ~n49213 & ~n49214 ;
  assign n49216 = ~n49099 & n49215 ;
  assign n49217 = n49099 & ~n49215 ;
  assign n49218 = ~n49216 & ~n49217 ;
  assign n49219 = x123 & n12506 ;
  assign n49220 = x121 & n13131 ;
  assign n49221 = x122 & n12501 ;
  assign n49222 = ~n49220 & ~n49221 ;
  assign n49223 = ~n49219 & n49222 ;
  assign n49224 = n12509 & n23382 ;
  assign n49225 = n49223 & ~n49224 ;
  assign n49226 = x44 & ~n49225 ;
  assign n49227 = x44 & ~n49226 ;
  assign n49228 = ~n49225 & ~n49226 ;
  assign n49229 = ~n49227 & ~n49228 ;
  assign n49230 = n49218 & ~n49229 ;
  assign n49231 = n49218 & ~n49230 ;
  assign n49232 = ~n49229 & ~n49230 ;
  assign n49233 = ~n49231 & ~n49232 ;
  assign n49234 = ~n48850 & ~n48863 ;
  assign n49235 = n49233 & n49234 ;
  assign n49236 = ~n49233 & ~n49234 ;
  assign n49237 = ~n49235 & ~n49236 ;
  assign n49238 = x126 & n10905 ;
  assign n49239 = x124 & n11466 ;
  assign n49240 = x125 & n10900 ;
  assign n49241 = ~n49239 & ~n49240 ;
  assign n49242 = ~n49238 & n49241 ;
  assign n49243 = n10908 & n25735 ;
  assign n49244 = n49242 & ~n49243 ;
  assign n49245 = x41 & ~n49244 ;
  assign n49246 = x41 & ~n49245 ;
  assign n49247 = ~n49244 & ~n49245 ;
  assign n49248 = ~n49246 & ~n49247 ;
  assign n49249 = n49237 & ~n49248 ;
  assign n49250 = n49237 & ~n49249 ;
  assign n49251 = ~n49248 & ~n49249 ;
  assign n49252 = ~n49250 & ~n49251 ;
  assign n49253 = ~n49098 & n49252 ;
  assign n49254 = n49098 & ~n49252 ;
  assign n49255 = ~n49253 & ~n49254 ;
  assign n49256 = ~n49086 & ~n49255 ;
  assign n49257 = n49086 & n49255 ;
  assign n49258 = ~n49256 & ~n49257 ;
  assign n49259 = ~n49085 & n49258 ;
  assign n49260 = n49085 & ~n49258 ;
  assign n49261 = ~n49259 & ~n49260 ;
  assign n49440 = n49261 & x229 ;
  assign n49262 = ~n49075 & ~n49078 ;
  assign n49263 = ~n48908 & ~n49068 ;
  assign n49264 = ~n49052 & ~n49065 ;
  assign n49265 = ~x127 & n9915 ;
  assign n49266 = n9436 & n27365 ;
  assign n49267 = ~n49265 & ~n49266 ;
  assign n49268 = ~x38 & ~n49267 ;
  assign n49269 = ~x38 & ~n49268 ;
  assign n49270 = ~n49267 & ~n49268 ;
  assign n49271 = ~n49269 & ~n49270 ;
  assign n49272 = ~n49264 & ~n49271 ;
  assign n49273 = ~n49264 & ~n49272 ;
  assign n49274 = ~n49271 & ~n49272 ;
  assign n49275 = ~n49273 & ~n49274 ;
  assign n49276 = ~n49012 & ~n49027 ;
  assign n49277 = ~x120 & n14233 ;
  assign n49278 = ~x118 & n14876 ;
  assign n49279 = ~x119 & n14228 ;
  assign n49280 = ~n49278 & ~n49279 ;
  assign n49281 = ~n49277 & n49280 ;
  assign n49282 = n14236 & n21501 ;
  assign n49283 = n49281 & ~n49282 ;
  assign n49284 = ~x47 & ~n49283 ;
  assign n49285 = ~x47 & ~n49284 ;
  assign n49286 = ~n49283 & ~n49284 ;
  assign n49287 = ~n49285 & ~n49286 ;
  assign n49288 = ~n48994 & ~n49007 ;
  assign n49289 = ~x117 & n16076 ;
  assign n49290 = ~x115 & n16756 ;
  assign n49291 = ~x116 & n16071 ;
  assign n49292 = ~n49290 & ~n49291 ;
  assign n49293 = ~n49289 & n49292 ;
  assign n49294 = n16079 & n19365 ;
  assign n49295 = n49293 & ~n49294 ;
  assign n49296 = ~x50 & ~n49295 ;
  assign n49297 = ~x50 & ~n49296 ;
  assign n49298 = ~n49295 & ~n49296 ;
  assign n49299 = ~n49297 & ~n49298 ;
  assign n49300 = ~n48975 & ~n48988 ;
  assign n49301 = ~n48927 & ~n48931 ;
  assign n49302 = ~x101 & n27427 ;
  assign n49303 = ~x102 & ~n26217 ;
  assign n49304 = ~n49302 & ~n49303 ;
  assign n49305 = n48924 & ~n49304 ;
  assign n49306 = n48924 & ~n49305 ;
  assign n49307 = ~n49304 & ~n49305 ;
  assign n49308 = ~n49306 & ~n49307 ;
  assign n49309 = ~n49301 & ~n49308 ;
  assign n49310 = ~n49301 & ~n49309 ;
  assign n49311 = ~n49308 & ~n49309 ;
  assign n49312 = ~n49310 & ~n49311 ;
  assign n49313 = ~x105 & n24612 ;
  assign n49314 = ~x103 & n25390 ;
  assign n49315 = ~x104 & n24607 ;
  assign n49316 = ~n49314 & ~n49315 ;
  assign n49317 = ~n49313 & n49316 ;
  assign n49318 = n11907 & n24615 ;
  assign n49319 = n49317 & ~n49318 ;
  assign n49320 = ~x62 & ~n49319 ;
  assign n49321 = ~x62 & ~n49320 ;
  assign n49322 = ~n49319 & ~n49320 ;
  assign n49323 = ~n49321 & ~n49322 ;
  assign n49324 = ~n49312 & ~n49323 ;
  assign n49325 = ~n49312 & ~n49324 ;
  assign n49326 = ~n49323 & ~n49324 ;
  assign n49327 = ~n49325 & ~n49326 ;
  assign n49328 = ~x108 & n22325 ;
  assign n49329 = ~x106 & n23066 ;
  assign n49330 = ~x107 & n22320 ;
  assign n49331 = ~n49329 & ~n49330 ;
  assign n49332 = ~n49328 & n49331 ;
  assign n49333 = n13601 & n22328 ;
  assign n49334 = n49332 & ~n49333 ;
  assign n49335 = ~x59 & ~n49334 ;
  assign n49336 = ~x59 & ~n49335 ;
  assign n49337 = ~n49334 & ~n49335 ;
  assign n49338 = ~n49336 & ~n49337 ;
  assign n49339 = ~n49327 & n49338 ;
  assign n49340 = n49327 & ~n49338 ;
  assign n49341 = ~n49339 & ~n49340 ;
  assign n49342 = ~n48937 & ~n48950 ;
  assign n49343 = n49341 & n49342 ;
  assign n49344 = ~n49341 & ~n49342 ;
  assign n49345 = ~n49343 & ~n49344 ;
  assign n49346 = ~x111 & n20143 ;
  assign n49347 = ~x109 & n20854 ;
  assign n49348 = ~x110 & n20138 ;
  assign n49349 = ~n49347 & ~n49348 ;
  assign n49350 = ~n49346 & n49349 ;
  assign n49351 = n15411 & n20146 ;
  assign n49352 = n49350 & ~n49351 ;
  assign n49353 = ~x56 & ~n49352 ;
  assign n49354 = ~x56 & ~n49353 ;
  assign n49355 = ~n49352 & ~n49353 ;
  assign n49356 = ~n49354 & ~n49355 ;
  assign n49357 = n49345 & ~n49356 ;
  assign n49358 = n49345 & ~n49357 ;
  assign n49359 = ~n49356 & ~n49357 ;
  assign n49360 = ~n49358 & ~n49359 ;
  assign n49361 = ~n48956 & ~n48969 ;
  assign n49362 = n49360 & n49361 ;
  assign n49363 = ~n49360 & ~n49361 ;
  assign n49364 = ~n49362 & ~n49363 ;
  assign n49365 = ~x114 & n18025 ;
  assign n49366 = ~x112 & n18764 ;
  assign n49367 = ~x113 & n18020 ;
  assign n49368 = ~n49366 & ~n49367 ;
  assign n49369 = ~n49365 & n49368 ;
  assign n49370 = n17333 & n18028 ;
  assign n49371 = n49369 & ~n49370 ;
  assign n49372 = ~x53 & ~n49371 ;
  assign n49373 = ~x53 & ~n49372 ;
  assign n49374 = ~n49371 & ~n49372 ;
  assign n49375 = ~n49373 & ~n49374 ;
  assign n49376 = ~n49364 & n49375 ;
  assign n49377 = n49364 & ~n49375 ;
  assign n49378 = ~n49376 & ~n49377 ;
  assign n49379 = ~n49300 & n49378 ;
  assign n49380 = ~n49300 & ~n49379 ;
  assign n49381 = n49378 & ~n49379 ;
  assign n49382 = ~n49380 & ~n49381 ;
  assign n49383 = ~n49299 & ~n49382 ;
  assign n49384 = n49299 & ~n49381 ;
  assign n49385 = ~n49380 & n49384 ;
  assign n49386 = ~n49383 & ~n49385 ;
  assign n49387 = ~n49288 & n49386 ;
  assign n49388 = n49288 & ~n49386 ;
  assign n49389 = ~n49387 & ~n49388 ;
  assign n49390 = ~n49287 & n49389 ;
  assign n49391 = n49287 & ~n49389 ;
  assign n49392 = ~n49390 & ~n49391 ;
  assign n49393 = ~n49276 & n49392 ;
  assign n49394 = n49276 & ~n49392 ;
  assign n49395 = ~n49393 & ~n49394 ;
  assign n49396 = ~x123 & n12506 ;
  assign n49397 = ~x121 & n13131 ;
  assign n49398 = ~x122 & n12501 ;
  assign n49399 = ~n49397 & ~n49398 ;
  assign n49400 = ~n49396 & n49399 ;
  assign n49401 = n12509 & n23760 ;
  assign n49402 = n49400 & ~n49401 ;
  assign n49403 = ~x44 & ~n49402 ;
  assign n49404 = ~x44 & ~n49403 ;
  assign n49405 = ~n49402 & ~n49403 ;
  assign n49406 = ~n49404 & ~n49405 ;
  assign n49407 = n49395 & ~n49406 ;
  assign n49408 = n49395 & ~n49407 ;
  assign n49409 = ~n49406 & ~n49407 ;
  assign n49410 = ~n49408 & ~n49409 ;
  assign n49411 = ~n49033 & ~n49046 ;
  assign n49412 = n49410 & n49411 ;
  assign n49413 = ~n49410 & ~n49411 ;
  assign n49414 = ~n49412 & ~n49413 ;
  assign n49415 = ~x126 & n10905 ;
  assign n49416 = ~x124 & n11466 ;
  assign n49417 = ~x125 & n10900 ;
  assign n49418 = ~n49416 & ~n49417 ;
  assign n49419 = ~n49415 & n49418 ;
  assign n49420 = n10908 & n26128 ;
  assign n49421 = n49419 & ~n49420 ;
  assign n49422 = ~x41 & ~n49421 ;
  assign n49423 = ~x41 & ~n49422 ;
  assign n49424 = ~n49421 & ~n49422 ;
  assign n49425 = ~n49423 & ~n49424 ;
  assign n49426 = n49414 & ~n49425 ;
  assign n49427 = n49414 & ~n49426 ;
  assign n49428 = ~n49425 & ~n49426 ;
  assign n49429 = ~n49427 & ~n49428 ;
  assign n49430 = ~n49275 & n49429 ;
  assign n49431 = n49275 & ~n49429 ;
  assign n49432 = ~n49430 & ~n49431 ;
  assign n49433 = ~n49263 & ~n49432 ;
  assign n49434 = n49263 & n49432 ;
  assign n49435 = ~n49433 & ~n49434 ;
  assign n49436 = ~n49262 & n49435 ;
  assign n49437 = n49262 & ~n49435 ;
  assign n49438 = ~n49436 & ~n49437 ;
  assign n49441 = ~n49438 & ~x229 ;
  assign n49442 = ~n49440 & ~n49441 ;
  assign n49443 = ~n49256 & ~n49259 ;
  assign n49444 = ~n49202 & ~n49206 ;
  assign n49445 = x118 & n16076 ;
  assign n49446 = x116 & n16756 ;
  assign n49447 = x117 & n16071 ;
  assign n49448 = ~n49446 & ~n49447 ;
  assign n49449 = ~n49445 & n49448 ;
  assign n49450 = n16079 & n19395 ;
  assign n49451 = n49449 & ~n49450 ;
  assign n49452 = x50 & ~n49451 ;
  assign n49453 = x50 & ~n49452 ;
  assign n49454 = ~n49451 & ~n49452 ;
  assign n49455 = ~n49453 & ~n49454 ;
  assign n49456 = ~n49186 & ~n49200 ;
  assign n49457 = ~n49128 & ~n49132 ;
  assign n49458 = x102 & n27024 ;
  assign n49459 = x103 & ~n26217 ;
  assign n49460 = ~n49458 & ~n49459 ;
  assign n49461 = x38 & ~n48741 ;
  assign n49462 = ~x38 & n48741 ;
  assign n49463 = ~n49461 & ~n49462 ;
  assign n49464 = ~n49460 & ~n49463 ;
  assign n49465 = n49460 & n49463 ;
  assign n49466 = ~n49464 & ~n49465 ;
  assign n49467 = ~n49457 & n49466 ;
  assign n49468 = n49457 & ~n49466 ;
  assign n49469 = ~n49467 & ~n49468 ;
  assign n49470 = x106 & n24612 ;
  assign n49471 = x104 & n25390 ;
  assign n49472 = x105 & n24607 ;
  assign n49473 = ~n49471 & ~n49472 ;
  assign n49474 = ~n49470 & n49473 ;
  assign n49475 = n12181 & n24615 ;
  assign n49476 = n49474 & ~n49475 ;
  assign n49477 = x62 & ~n49476 ;
  assign n49478 = x62 & ~n49477 ;
  assign n49479 = ~n49476 & ~n49477 ;
  assign n49480 = ~n49478 & ~n49479 ;
  assign n49481 = n49469 & ~n49480 ;
  assign n49482 = n49469 & ~n49481 ;
  assign n49483 = ~n49480 & ~n49481 ;
  assign n49484 = ~n49482 & ~n49483 ;
  assign n49485 = x109 & n22325 ;
  assign n49486 = x107 & n23066 ;
  assign n49487 = x108 & n22320 ;
  assign n49488 = ~n49486 & ~n49487 ;
  assign n49489 = ~n49485 & n49488 ;
  assign n49490 = n13894 & n22328 ;
  assign n49491 = n49489 & ~n49490 ;
  assign n49492 = x59 & ~n49491 ;
  assign n49493 = x59 & ~n49492 ;
  assign n49494 = ~n49491 & ~n49492 ;
  assign n49495 = ~n49493 & ~n49494 ;
  assign n49496 = ~n49484 & ~n49495 ;
  assign n49497 = ~n49484 & ~n49496 ;
  assign n49498 = ~n49495 & ~n49496 ;
  assign n49499 = ~n49497 & ~n49498 ;
  assign n49500 = ~n49150 & ~n49161 ;
  assign n49501 = ~n49147 & ~n49500 ;
  assign n49502 = ~n49499 & ~n49501 ;
  assign n49503 = ~n49499 & ~n49502 ;
  assign n49504 = ~n49501 & ~n49502 ;
  assign n49505 = ~n49503 & ~n49504 ;
  assign n49506 = x112 & n20143 ;
  assign n49507 = x110 & n20854 ;
  assign n49508 = x111 & n20138 ;
  assign n49509 = ~n49507 & ~n49508 ;
  assign n49510 = ~n49506 & n49509 ;
  assign n49511 = n15442 & n20146 ;
  assign n49512 = n49510 & ~n49511 ;
  assign n49513 = x56 & ~n49512 ;
  assign n49514 = x56 & ~n49513 ;
  assign n49515 = ~n49512 & ~n49513 ;
  assign n49516 = ~n49514 & ~n49515 ;
  assign n49517 = ~n49505 & ~n49516 ;
  assign n49518 = ~n49505 & ~n49517 ;
  assign n49519 = ~n49516 & ~n49517 ;
  assign n49520 = ~n49518 & ~n49519 ;
  assign n49521 = ~n49167 & ~n49180 ;
  assign n49522 = n49520 & n49521 ;
  assign n49523 = ~n49520 & ~n49521 ;
  assign n49524 = ~n49522 & ~n49523 ;
  assign n49525 = x115 & n18025 ;
  assign n49526 = x113 & n18764 ;
  assign n49527 = x114 & n18020 ;
  assign n49528 = ~n49526 & ~n49527 ;
  assign n49529 = ~n49525 & n49528 ;
  assign n49530 = n17364 & n18028 ;
  assign n49531 = n49529 & ~n49530 ;
  assign n49532 = x53 & ~n49531 ;
  assign n49533 = x53 & ~n49532 ;
  assign n49534 = ~n49531 & ~n49532 ;
  assign n49535 = ~n49533 & ~n49534 ;
  assign n49536 = ~n49524 & n49535 ;
  assign n49537 = n49524 & ~n49535 ;
  assign n49538 = ~n49536 & ~n49537 ;
  assign n49539 = ~n49456 & n49538 ;
  assign n49540 = n49456 & ~n49538 ;
  assign n49541 = ~n49539 & ~n49540 ;
  assign n49542 = ~n49455 & n49541 ;
  assign n49543 = n49455 & ~n49541 ;
  assign n49544 = ~n49542 & ~n49543 ;
  assign n49545 = ~n49444 & n49544 ;
  assign n49546 = n49444 & ~n49544 ;
  assign n49547 = ~n49545 & ~n49546 ;
  assign n49548 = x121 & n14233 ;
  assign n49549 = x119 & n14876 ;
  assign n49550 = x120 & n14228 ;
  assign n49551 = ~n49549 & ~n49550 ;
  assign n49552 = ~n49548 & n49551 ;
  assign n49553 = n14236 & n21870 ;
  assign n49554 = n49552 & ~n49553 ;
  assign n49555 = x47 & ~n49554 ;
  assign n49556 = x47 & ~n49555 ;
  assign n49557 = ~n49554 & ~n49555 ;
  assign n49558 = ~n49556 & ~n49557 ;
  assign n49559 = n49547 & ~n49558 ;
  assign n49560 = n49547 & ~n49559 ;
  assign n49561 = ~n49558 & ~n49559 ;
  assign n49562 = ~n49560 & ~n49561 ;
  assign n49563 = ~n49210 & ~n49213 ;
  assign n49564 = n49562 & n49563 ;
  assign n49565 = ~n49562 & ~n49563 ;
  assign n49566 = ~n49564 & ~n49565 ;
  assign n49567 = x124 & n12506 ;
  assign n49568 = x122 & n13131 ;
  assign n49569 = x123 & n12501 ;
  assign n49570 = ~n49568 & ~n49569 ;
  assign n49571 = ~n49567 & n49570 ;
  assign n49572 = n12509 & n23796 ;
  assign n49573 = n49571 & ~n49572 ;
  assign n49574 = x44 & ~n49573 ;
  assign n49575 = x44 & ~n49574 ;
  assign n49576 = ~n49573 & ~n49574 ;
  assign n49577 = ~n49575 & ~n49576 ;
  assign n49578 = n49566 & ~n49577 ;
  assign n49579 = n49566 & ~n49578 ;
  assign n49580 = ~n49577 & ~n49578 ;
  assign n49581 = ~n49579 & ~n49580 ;
  assign n49582 = ~n49216 & ~n49230 ;
  assign n49583 = n49581 & n49582 ;
  assign n49584 = ~n49581 & ~n49582 ;
  assign n49585 = ~n49583 & ~n49584 ;
  assign n49586 = x127 & n10905 ;
  assign n49587 = x125 & n11466 ;
  assign n49588 = x126 & n10900 ;
  assign n49589 = ~n49587 & ~n49588 ;
  assign n49590 = ~n49586 & n49589 ;
  assign n49591 = n10908 & n26533 ;
  assign n49592 = n49590 & ~n49591 ;
  assign n49593 = x41 & ~n49592 ;
  assign n49594 = x41 & ~n49593 ;
  assign n49595 = ~n49592 & ~n49593 ;
  assign n49596 = ~n49594 & ~n49595 ;
  assign n49597 = n49585 & ~n49596 ;
  assign n49598 = n49585 & ~n49597 ;
  assign n49599 = ~n49596 & ~n49597 ;
  assign n49600 = ~n49598 & ~n49599 ;
  assign n49601 = ~n49236 & ~n49249 ;
  assign n49602 = n49600 & n49601 ;
  assign n49603 = ~n49600 & ~n49601 ;
  assign n49604 = ~n49602 & ~n49603 ;
  assign n49605 = ~n49098 & ~n49252 ;
  assign n49606 = ~n49095 & ~n49605 ;
  assign n49607 = n49604 & ~n49606 ;
  assign n49608 = ~n49604 & n49606 ;
  assign n49609 = ~n49607 & ~n49608 ;
  assign n49610 = ~n49443 & n49609 ;
  assign n49611 = n49443 & ~n49609 ;
  assign n49612 = ~n49610 & ~n49611 ;
  assign n49784 = n49612 & x230 ;
  assign n49613 = ~n49433 & ~n49436 ;
  assign n49614 = ~n49379 & ~n49383 ;
  assign n49615 = ~x118 & n16076 ;
  assign n49616 = ~x116 & n16756 ;
  assign n49617 = ~x117 & n16071 ;
  assign n49618 = ~n49616 & ~n49617 ;
  assign n49619 = ~n49615 & n49618 ;
  assign n49620 = n16079 & n19736 ;
  assign n49621 = n49619 & ~n49620 ;
  assign n49622 = ~x50 & ~n49621 ;
  assign n49623 = ~x50 & ~n49622 ;
  assign n49624 = ~n49621 & ~n49622 ;
  assign n49625 = ~n49623 & ~n49624 ;
  assign n49626 = ~n49363 & ~n49377 ;
  assign n49627 = ~n49305 & ~n49309 ;
  assign n49628 = ~x102 & n27427 ;
  assign n49629 = ~x103 & ~n26217 ;
  assign n49630 = ~n49628 & ~n49629 ;
  assign n49631 = ~x38 & ~n48924 ;
  assign n49632 = x38 & n48924 ;
  assign n49633 = ~n49631 & ~n49632 ;
  assign n49634 = ~n49630 & ~n49633 ;
  assign n49635 = n49630 & n49633 ;
  assign n49636 = ~n49634 & ~n49635 ;
  assign n49637 = ~n49627 & n49636 ;
  assign n49638 = n49627 & ~n49636 ;
  assign n49639 = ~n49637 & ~n49638 ;
  assign n49640 = ~x106 & n24612 ;
  assign n49641 = ~x104 & n25390 ;
  assign n49642 = ~x105 & n24607 ;
  assign n49643 = ~n49641 & ~n49642 ;
  assign n49644 = ~n49640 & n49643 ;
  assign n49645 = n12447 & n24615 ;
  assign n49646 = n49644 & ~n49645 ;
  assign n49647 = ~x62 & ~n49646 ;
  assign n49648 = ~x62 & ~n49647 ;
  assign n49649 = ~n49646 & ~n49647 ;
  assign n49650 = ~n49648 & ~n49649 ;
  assign n49651 = n49639 & ~n49650 ;
  assign n49652 = n49639 & ~n49651 ;
  assign n49653 = ~n49650 & ~n49651 ;
  assign n49654 = ~n49652 & ~n49653 ;
  assign n49655 = ~x109 & n22325 ;
  assign n49656 = ~x107 & n23066 ;
  assign n49657 = ~x108 & n22320 ;
  assign n49658 = ~n49656 & ~n49657 ;
  assign n49659 = ~n49655 & n49658 ;
  assign n49660 = n14177 & n22328 ;
  assign n49661 = n49659 & ~n49660 ;
  assign n49662 = ~x59 & ~n49661 ;
  assign n49663 = ~x59 & ~n49662 ;
  assign n49664 = ~n49661 & ~n49662 ;
  assign n49665 = ~n49663 & ~n49664 ;
  assign n49666 = ~n49654 & ~n49665 ;
  assign n49667 = ~n49654 & ~n49666 ;
  assign n49668 = ~n49665 & ~n49666 ;
  assign n49669 = ~n49667 & ~n49668 ;
  assign n49670 = ~n49327 & ~n49338 ;
  assign n49671 = ~n49324 & ~n49670 ;
  assign n49672 = ~n49669 & ~n49671 ;
  assign n49673 = ~n49669 & ~n49672 ;
  assign n49674 = ~n49671 & ~n49672 ;
  assign n49675 = ~n49673 & ~n49674 ;
  assign n49676 = ~x112 & n20143 ;
  assign n49677 = ~x110 & n20854 ;
  assign n49678 = ~x111 & n20138 ;
  assign n49679 = ~n49677 & ~n49678 ;
  assign n49680 = ~n49676 & n49679 ;
  assign n49681 = n15744 & n20146 ;
  assign n49682 = n49680 & ~n49681 ;
  assign n49683 = ~x56 & ~n49682 ;
  assign n49684 = ~x56 & ~n49683 ;
  assign n49685 = ~n49682 & ~n49683 ;
  assign n49686 = ~n49684 & ~n49685 ;
  assign n49687 = ~n49675 & ~n49686 ;
  assign n49688 = ~n49675 & ~n49687 ;
  assign n49689 = ~n49686 & ~n49687 ;
  assign n49690 = ~n49688 & ~n49689 ;
  assign n49691 = ~n49344 & ~n49357 ;
  assign n49692 = n49690 & n49691 ;
  assign n49693 = ~n49690 & ~n49691 ;
  assign n49694 = ~n49692 & ~n49693 ;
  assign n49695 = ~x115 & n18025 ;
  assign n49696 = ~x113 & n18764 ;
  assign n49697 = ~x114 & n18020 ;
  assign n49698 = ~n49696 & ~n49697 ;
  assign n49699 = ~n49695 & n49698 ;
  assign n49700 = n17683 & n18028 ;
  assign n49701 = n49699 & ~n49700 ;
  assign n49702 = ~x53 & ~n49701 ;
  assign n49703 = ~x53 & ~n49702 ;
  assign n49704 = ~n49701 & ~n49702 ;
  assign n49705 = ~n49703 & ~n49704 ;
  assign n49706 = ~n49694 & n49705 ;
  assign n49707 = n49694 & ~n49705 ;
  assign n49708 = ~n49706 & ~n49707 ;
  assign n49709 = ~n49626 & n49708 ;
  assign n49710 = n49626 & ~n49708 ;
  assign n49711 = ~n49709 & ~n49710 ;
  assign n49712 = ~n49625 & n49711 ;
  assign n49713 = n49625 & ~n49711 ;
  assign n49714 = ~n49712 & ~n49713 ;
  assign n49715 = ~n49614 & n49714 ;
  assign n49716 = n49614 & ~n49714 ;
  assign n49717 = ~n49715 & ~n49716 ;
  assign n49718 = ~x121 & n14233 ;
  assign n49719 = ~x119 & n14876 ;
  assign n49720 = ~x120 & n14228 ;
  assign n49721 = ~n49719 & ~n49720 ;
  assign n49722 = ~n49718 & n49721 ;
  assign n49723 = n14236 & n22229 ;
  assign n49724 = n49722 & ~n49723 ;
  assign n49725 = ~x47 & ~n49724 ;
  assign n49726 = ~x47 & ~n49725 ;
  assign n49727 = ~n49724 & ~n49725 ;
  assign n49728 = ~n49726 & ~n49727 ;
  assign n49729 = n49717 & ~n49728 ;
  assign n49730 = n49717 & ~n49729 ;
  assign n49731 = ~n49728 & ~n49729 ;
  assign n49732 = ~n49730 & ~n49731 ;
  assign n49733 = ~n49387 & ~n49390 ;
  assign n49734 = n49732 & n49733 ;
  assign n49735 = ~n49732 & ~n49733 ;
  assign n49736 = ~n49734 & ~n49735 ;
  assign n49737 = ~x124 & n12506 ;
  assign n49738 = ~x122 & n13131 ;
  assign n49739 = ~x123 & n12501 ;
  assign n49740 = ~n49738 & ~n49739 ;
  assign n49741 = ~n49737 & n49740 ;
  assign n49742 = n12509 & n24176 ;
  assign n49743 = n49741 & ~n49742 ;
  assign n49744 = ~x44 & ~n49743 ;
  assign n49745 = ~x44 & ~n49744 ;
  assign n49746 = ~n49743 & ~n49744 ;
  assign n49747 = ~n49745 & ~n49746 ;
  assign n49748 = n49736 & ~n49747 ;
  assign n49749 = n49736 & ~n49748 ;
  assign n49750 = ~n49747 & ~n49748 ;
  assign n49751 = ~n49749 & ~n49750 ;
  assign n49752 = ~n49393 & ~n49407 ;
  assign n49753 = n49751 & n49752 ;
  assign n49754 = ~n49751 & ~n49752 ;
  assign n49755 = ~n49753 & ~n49754 ;
  assign n49756 = ~x127 & n10905 ;
  assign n49757 = ~x125 & n11466 ;
  assign n49758 = ~x126 & n10900 ;
  assign n49759 = ~n49757 & ~n49758 ;
  assign n49760 = ~n49756 & n49759 ;
  assign n49761 = n10908 & n26932 ;
  assign n49762 = n49760 & ~n49761 ;
  assign n49763 = ~x41 & ~n49762 ;
  assign n49764 = ~x41 & ~n49763 ;
  assign n49765 = ~n49762 & ~n49763 ;
  assign n49766 = ~n49764 & ~n49765 ;
  assign n49767 = n49755 & ~n49766 ;
  assign n49768 = n49755 & ~n49767 ;
  assign n49769 = ~n49766 & ~n49767 ;
  assign n49770 = ~n49768 & ~n49769 ;
  assign n49771 = ~n49413 & ~n49426 ;
  assign n49772 = n49770 & n49771 ;
  assign n49773 = ~n49770 & ~n49771 ;
  assign n49774 = ~n49772 & ~n49773 ;
  assign n49775 = ~n49275 & ~n49429 ;
  assign n49776 = ~n49272 & ~n49775 ;
  assign n49777 = n49774 & ~n49776 ;
  assign n49778 = ~n49774 & n49776 ;
  assign n49779 = ~n49777 & ~n49778 ;
  assign n49780 = ~n49613 & n49779 ;
  assign n49781 = n49613 & ~n49779 ;
  assign n49782 = ~n49780 & ~n49781 ;
  assign n49785 = ~n49782 & ~x230 ;
  assign n49786 = ~n49784 & ~n49785 ;
  assign n49787 = ~n49578 & ~n49584 ;
  assign n49788 = x126 & n11466 ;
  assign n49789 = x127 & n10900 ;
  assign n49790 = ~n49788 & ~n49789 ;
  assign n49791 = ~n10908 & n49790 ;
  assign n49792 = n26965 & n49790 ;
  assign n49793 = ~n49791 & ~n49792 ;
  assign n49794 = x41 & ~n49793 ;
  assign n49795 = ~x41 & n49793 ;
  assign n49796 = ~n49794 & ~n49795 ;
  assign n49797 = ~n49787 & ~n49796 ;
  assign n49798 = n49787 & n49796 ;
  assign n49799 = ~n49797 & ~n49798 ;
  assign n49800 = ~n49467 & ~n49481 ;
  assign n49801 = x103 & n27024 ;
  assign n49802 = x104 & ~n26217 ;
  assign n49803 = ~n49801 & ~n49802 ;
  assign n49804 = ~x38 & ~n48741 ;
  assign n49805 = ~n49464 & ~n49804 ;
  assign n49806 = n49803 & ~n49805 ;
  assign n49807 = ~n49803 & n49805 ;
  assign n49808 = ~n49806 & ~n49807 ;
  assign n49809 = x107 & n24612 ;
  assign n49810 = x105 & n25390 ;
  assign n49811 = x106 & n24607 ;
  assign n49812 = ~n49810 & ~n49811 ;
  assign n49813 = ~n49809 & n49812 ;
  assign n49814 = ~n24615 & n49813 ;
  assign n49815 = ~n12749 & n49813 ;
  assign n49816 = ~n49814 & ~n49815 ;
  assign n49817 = x62 & ~n49816 ;
  assign n49818 = ~x62 & n49816 ;
  assign n49819 = ~n49817 & ~n49818 ;
  assign n49820 = n49808 & ~n49819 ;
  assign n49821 = ~n49808 & n49819 ;
  assign n49822 = ~n49820 & ~n49821 ;
  assign n49823 = ~n49800 & n49822 ;
  assign n49824 = n49800 & ~n49822 ;
  assign n49825 = ~n49823 & ~n49824 ;
  assign n49826 = x110 & n22325 ;
  assign n49827 = x108 & n23066 ;
  assign n49828 = x109 & n22320 ;
  assign n49829 = ~n49827 & ~n49828 ;
  assign n49830 = ~n49826 & n49829 ;
  assign n49831 = n14497 & n22328 ;
  assign n49832 = n49830 & ~n49831 ;
  assign n49833 = x59 & ~n49832 ;
  assign n49834 = x59 & ~n49833 ;
  assign n49835 = ~n49832 & ~n49833 ;
  assign n49836 = ~n49834 & ~n49835 ;
  assign n49837 = n49825 & ~n49836 ;
  assign n49838 = n49825 & ~n49837 ;
  assign n49839 = ~n49836 & ~n49837 ;
  assign n49840 = ~n49838 & ~n49839 ;
  assign n49841 = ~n49496 & ~n49502 ;
  assign n49842 = n49840 & n49841 ;
  assign n49843 = ~n49840 & ~n49841 ;
  assign n49844 = ~n49842 & ~n49843 ;
  assign n49845 = x113 & n20143 ;
  assign n49846 = x111 & n20854 ;
  assign n49847 = x112 & n20138 ;
  assign n49848 = ~n49846 & ~n49847 ;
  assign n49849 = ~n49845 & n49848 ;
  assign n49850 = n16361 & n20146 ;
  assign n49851 = n49849 & ~n49850 ;
  assign n49852 = x56 & ~n49851 ;
  assign n49853 = x56 & ~n49852 ;
  assign n49854 = ~n49851 & ~n49852 ;
  assign n49855 = ~n49853 & ~n49854 ;
  assign n49856 = n49844 & ~n49855 ;
  assign n49857 = n49844 & ~n49856 ;
  assign n49858 = ~n49855 & ~n49856 ;
  assign n49859 = ~n49857 & ~n49858 ;
  assign n49860 = ~n49517 & ~n49523 ;
  assign n49861 = n49859 & n49860 ;
  assign n49862 = ~n49859 & ~n49860 ;
  assign n49863 = ~n49861 & ~n49862 ;
  assign n49864 = x116 & n18025 ;
  assign n49865 = x114 & n18764 ;
  assign n49866 = x115 & n18020 ;
  assign n49867 = ~n49865 & ~n49866 ;
  assign n49868 = ~n49864 & n49867 ;
  assign n49869 = n18028 & n18336 ;
  assign n49870 = n49868 & ~n49869 ;
  assign n49871 = x53 & ~n49870 ;
  assign n49872 = x53 & ~n49871 ;
  assign n49873 = ~n49870 & ~n49871 ;
  assign n49874 = ~n49872 & ~n49873 ;
  assign n49875 = n49863 & ~n49874 ;
  assign n49876 = n49863 & ~n49875 ;
  assign n49877 = ~n49874 & ~n49875 ;
  assign n49878 = ~n49876 & ~n49877 ;
  assign n49879 = ~n49537 & ~n49539 ;
  assign n49880 = ~n49878 & ~n49879 ;
  assign n49881 = ~n49878 & ~n49880 ;
  assign n49882 = ~n49879 & ~n49880 ;
  assign n49883 = ~n49881 & ~n49882 ;
  assign n49884 = x119 & n16076 ;
  assign n49885 = x117 & n16756 ;
  assign n49886 = x118 & n16071 ;
  assign n49887 = ~n49885 & ~n49886 ;
  assign n49888 = ~n49884 & n49887 ;
  assign n49889 = n16079 & n20423 ;
  assign n49890 = n49888 & ~n49889 ;
  assign n49891 = x50 & ~n49890 ;
  assign n49892 = x50 & ~n49891 ;
  assign n49893 = ~n49890 & ~n49891 ;
  assign n49894 = ~n49892 & ~n49893 ;
  assign n49895 = ~n49883 & ~n49894 ;
  assign n49896 = ~n49883 & ~n49895 ;
  assign n49897 = ~n49894 & ~n49895 ;
  assign n49898 = ~n49896 & ~n49897 ;
  assign n49899 = ~n49542 & ~n49545 ;
  assign n49900 = n49898 & n49899 ;
  assign n49901 = ~n49898 & ~n49899 ;
  assign n49902 = ~n49900 & ~n49901 ;
  assign n49903 = x122 & n14233 ;
  assign n49904 = x120 & n14876 ;
  assign n49905 = x121 & n14228 ;
  assign n49906 = ~n49904 & ~n49905 ;
  assign n49907 = ~n49903 & n49906 ;
  assign n49908 = n14236 & n22622 ;
  assign n49909 = n49907 & ~n49908 ;
  assign n49910 = x47 & ~n49909 ;
  assign n49911 = x47 & ~n49910 ;
  assign n49912 = ~n49909 & ~n49910 ;
  assign n49913 = ~n49911 & ~n49912 ;
  assign n49914 = n49902 & ~n49913 ;
  assign n49915 = n49902 & ~n49914 ;
  assign n49916 = ~n49913 & ~n49914 ;
  assign n49917 = ~n49915 & ~n49916 ;
  assign n49918 = ~n49559 & ~n49565 ;
  assign n49919 = n49917 & n49918 ;
  assign n49920 = ~n49917 & ~n49918 ;
  assign n49921 = ~n49919 & ~n49920 ;
  assign n49922 = x125 & n12506 ;
  assign n49923 = x123 & n13131 ;
  assign n49924 = x124 & n12501 ;
  assign n49925 = ~n49923 & ~n49924 ;
  assign n49926 = ~n49922 & n49925 ;
  assign n49927 = n12509 & n24935 ;
  assign n49928 = n49926 & ~n49927 ;
  assign n49929 = x44 & ~n49928 ;
  assign n49930 = x44 & ~n49929 ;
  assign n49931 = ~n49928 & ~n49929 ;
  assign n49932 = ~n49930 & ~n49931 ;
  assign n49933 = n49921 & ~n49932 ;
  assign n49934 = ~n49921 & n49932 ;
  assign n49935 = n49799 & ~n49934 ;
  assign n49936 = ~n49933 & n49935 ;
  assign n49937 = n49799 & ~n49936 ;
  assign n49938 = ~n49934 & ~n49936 ;
  assign n49939 = ~n49933 & n49938 ;
  assign n49940 = ~n49937 & ~n49939 ;
  assign n49941 = ~n49597 & ~n49603 ;
  assign n49942 = n49940 & n49941 ;
  assign n49943 = ~n49940 & ~n49941 ;
  assign n49944 = ~n49942 & ~n49943 ;
  assign n49945 = ~n49607 & ~n49610 ;
  assign n49946 = n49944 & ~n49945 ;
  assign n49947 = ~n49944 & n49945 ;
  assign n49948 = ~n49946 & ~n49947 ;
  assign n50112 = n49948 & x231 ;
  assign n49949 = ~n49748 & ~n49754 ;
  assign n49950 = ~x126 & n11466 ;
  assign n49951 = ~x127 & n10900 ;
  assign n49952 = ~n49950 & ~n49951 ;
  assign n49953 = ~n10908 & n49952 ;
  assign n49954 = n27368 & n49952 ;
  assign n49955 = ~n49953 & ~n49954 ;
  assign n49956 = ~x41 & ~n49955 ;
  assign n49957 = x41 & n49955 ;
  assign n49958 = ~n49956 & ~n49957 ;
  assign n49959 = ~n49949 & ~n49958 ;
  assign n49960 = n49949 & n49958 ;
  assign n49961 = ~n49959 & ~n49960 ;
  assign n49962 = ~n49637 & ~n49651 ;
  assign n49963 = ~x103 & n27427 ;
  assign n49964 = ~x104 & ~n26217 ;
  assign n49965 = ~n49963 & ~n49964 ;
  assign n49966 = x38 & ~n48924 ;
  assign n49967 = ~n49634 & ~n49966 ;
  assign n49968 = n49965 & ~n49967 ;
  assign n49969 = ~n49965 & n49967 ;
  assign n49970 = ~n49968 & ~n49969 ;
  assign n49971 = ~x107 & n24612 ;
  assign n49972 = ~x105 & n25390 ;
  assign n49973 = ~x106 & n24607 ;
  assign n49974 = ~n49972 & ~n49973 ;
  assign n49975 = ~n49971 & n49974 ;
  assign n49976 = ~n24615 & n49975 ;
  assign n49977 = ~n13034 & n49975 ;
  assign n49978 = ~n49976 & ~n49977 ;
  assign n49979 = ~x62 & ~n49978 ;
  assign n49980 = x62 & n49978 ;
  assign n49981 = ~n49979 & ~n49980 ;
  assign n49982 = n49970 & ~n49981 ;
  assign n49983 = ~n49970 & n49981 ;
  assign n49984 = ~n49982 & ~n49983 ;
  assign n49985 = ~n49962 & n49984 ;
  assign n49986 = n49962 & ~n49984 ;
  assign n49987 = ~n49985 & ~n49986 ;
  assign n49988 = ~x110 & n22325 ;
  assign n49989 = ~x108 & n23066 ;
  assign n49990 = ~x109 & n22320 ;
  assign n49991 = ~n49989 & ~n49990 ;
  assign n49992 = ~n49988 & n49991 ;
  assign n49993 = n14802 & n22328 ;
  assign n49994 = n49992 & ~n49993 ;
  assign n49995 = ~x59 & ~n49994 ;
  assign n49996 = ~x59 & ~n49995 ;
  assign n49997 = ~n49994 & ~n49995 ;
  assign n49998 = ~n49996 & ~n49997 ;
  assign n49999 = n49987 & ~n49998 ;
  assign n50000 = n49987 & ~n49999 ;
  assign n50001 = ~n49998 & ~n49999 ;
  assign n50002 = ~n50000 & ~n50001 ;
  assign n50003 = ~n49666 & ~n49672 ;
  assign n50004 = n50002 & n50003 ;
  assign n50005 = ~n50002 & ~n50003 ;
  assign n50006 = ~n50004 & ~n50005 ;
  assign n50007 = ~x113 & n20143 ;
  assign n50008 = ~x111 & n20854 ;
  assign n50009 = ~x112 & n20138 ;
  assign n50010 = ~n50008 & ~n50009 ;
  assign n50011 = ~n50007 & n50010 ;
  assign n50012 = n16684 & n20146 ;
  assign n50013 = n50011 & ~n50012 ;
  assign n50014 = ~x56 & ~n50013 ;
  assign n50015 = ~x56 & ~n50014 ;
  assign n50016 = ~n50013 & ~n50014 ;
  assign n50017 = ~n50015 & ~n50016 ;
  assign n50018 = n50006 & ~n50017 ;
  assign n50019 = n50006 & ~n50018 ;
  assign n50020 = ~n50017 & ~n50018 ;
  assign n50021 = ~n50019 & ~n50020 ;
  assign n50022 = ~n49687 & ~n49693 ;
  assign n50023 = n50021 & n50022 ;
  assign n50024 = ~n50021 & ~n50022 ;
  assign n50025 = ~n50023 & ~n50024 ;
  assign n50026 = ~x116 & n18025 ;
  assign n50027 = ~x114 & n18764 ;
  assign n50028 = ~x115 & n18020 ;
  assign n50029 = ~n50027 & ~n50028 ;
  assign n50030 = ~n50026 & n50029 ;
  assign n50031 = n18028 & n18678 ;
  assign n50032 = n50030 & ~n50031 ;
  assign n50033 = ~x53 & ~n50032 ;
  assign n50034 = ~x53 & ~n50033 ;
  assign n50035 = ~n50032 & ~n50033 ;
  assign n50036 = ~n50034 & ~n50035 ;
  assign n50037 = n50025 & ~n50036 ;
  assign n50038 = n50025 & ~n50037 ;
  assign n50039 = ~n50036 & ~n50037 ;
  assign n50040 = ~n50038 & ~n50039 ;
  assign n50041 = ~n49707 & ~n49709 ;
  assign n50042 = ~n50040 & ~n50041 ;
  assign n50043 = ~n50040 & ~n50042 ;
  assign n50044 = ~n50041 & ~n50042 ;
  assign n50045 = ~n50043 & ~n50044 ;
  assign n50046 = ~x119 & n16076 ;
  assign n50047 = ~x117 & n16756 ;
  assign n50048 = ~x118 & n16071 ;
  assign n50049 = ~n50047 & ~n50048 ;
  assign n50050 = ~n50046 & n50049 ;
  assign n50051 = n16079 & n20778 ;
  assign n50052 = n50050 & ~n50051 ;
  assign n50053 = ~x50 & ~n50052 ;
  assign n50054 = ~x50 & ~n50053 ;
  assign n50055 = ~n50052 & ~n50053 ;
  assign n50056 = ~n50054 & ~n50055 ;
  assign n50057 = ~n50045 & ~n50056 ;
  assign n50058 = ~n50045 & ~n50057 ;
  assign n50059 = ~n50056 & ~n50057 ;
  assign n50060 = ~n50058 & ~n50059 ;
  assign n50061 = ~n49712 & ~n49715 ;
  assign n50062 = n50060 & n50061 ;
  assign n50063 = ~n50060 & ~n50061 ;
  assign n50064 = ~n50062 & ~n50063 ;
  assign n50065 = ~x122 & n14233 ;
  assign n50066 = ~x120 & n14876 ;
  assign n50067 = ~x121 & n14228 ;
  assign n50068 = ~n50066 & ~n50067 ;
  assign n50069 = ~n50065 & n50068 ;
  assign n50070 = n14236 & n22998 ;
  assign n50071 = n50069 & ~n50070 ;
  assign n50072 = ~x47 & ~n50071 ;
  assign n50073 = ~x47 & ~n50072 ;
  assign n50074 = ~n50071 & ~n50072 ;
  assign n50075 = ~n50073 & ~n50074 ;
  assign n50076 = n50064 & ~n50075 ;
  assign n50077 = n50064 & ~n50076 ;
  assign n50078 = ~n50075 & ~n50076 ;
  assign n50079 = ~n50077 & ~n50078 ;
  assign n50080 = ~n49729 & ~n49735 ;
  assign n50081 = n50079 & n50080 ;
  assign n50082 = ~n50079 & ~n50080 ;
  assign n50083 = ~n50081 & ~n50082 ;
  assign n50084 = ~x125 & n12506 ;
  assign n50085 = ~x123 & n13131 ;
  assign n50086 = ~x124 & n12501 ;
  assign n50087 = ~n50085 & ~n50086 ;
  assign n50088 = ~n50084 & n50087 ;
  assign n50089 = n12509 & n25330 ;
  assign n50090 = n50088 & ~n50089 ;
  assign n50091 = ~x44 & ~n50090 ;
  assign n50092 = ~x44 & ~n50091 ;
  assign n50093 = ~n50090 & ~n50091 ;
  assign n50094 = ~n50092 & ~n50093 ;
  assign n50095 = n50083 & ~n50094 ;
  assign n50096 = ~n50083 & n50094 ;
  assign n50097 = n49961 & ~n50096 ;
  assign n50098 = ~n50095 & n50097 ;
  assign n50099 = n49961 & ~n50098 ;
  assign n50100 = ~n50096 & ~n50098 ;
  assign n50101 = ~n50095 & n50100 ;
  assign n50102 = ~n50099 & ~n50101 ;
  assign n50103 = ~n49767 & ~n49773 ;
  assign n50104 = n50102 & n50103 ;
  assign n50105 = ~n50102 & ~n50103 ;
  assign n50106 = ~n50104 & ~n50105 ;
  assign n50107 = ~n49777 & ~n49780 ;
  assign n50108 = n50106 & ~n50107 ;
  assign n50109 = ~n50106 & n50107 ;
  assign n50110 = ~n50108 & ~n50109 ;
  assign n50113 = ~n50110 & ~x231 ;
  assign n50114 = ~n50112 & ~n50113 ;
  assign n50115 = ~n49943 & ~n49946 ;
  assign n50116 = ~n49797 & ~n49936 ;
  assign n50117 = ~n49920 & ~n49933 ;
  assign n50118 = x127 & n11466 ;
  assign n50119 = n10908 & n26962 ;
  assign n50120 = ~n50118 & ~n50119 ;
  assign n50121 = x41 & ~n50120 ;
  assign n50122 = x41 & ~n50121 ;
  assign n50123 = ~n50120 & ~n50121 ;
  assign n50124 = ~n50122 & ~n50123 ;
  assign n50125 = ~n50117 & ~n50124 ;
  assign n50126 = ~n50117 & ~n50125 ;
  assign n50127 = ~n50124 & ~n50125 ;
  assign n50128 = ~n50126 & ~n50127 ;
  assign n50129 = ~n49880 & ~n49895 ;
  assign n50130 = x120 & n16076 ;
  assign n50131 = x118 & n16756 ;
  assign n50132 = x119 & n16071 ;
  assign n50133 = ~n50131 & ~n50132 ;
  assign n50134 = ~n50130 & n50133 ;
  assign n50135 = n16079 & n21143 ;
  assign n50136 = n50134 & ~n50135 ;
  assign n50137 = x50 & ~n50136 ;
  assign n50138 = x50 & ~n50137 ;
  assign n50139 = ~n50136 & ~n50137 ;
  assign n50140 = ~n50138 & ~n50139 ;
  assign n50141 = ~n49862 & ~n49875 ;
  assign n50142 = x117 & n18025 ;
  assign n50143 = x115 & n18764 ;
  assign n50144 = x116 & n18020 ;
  assign n50145 = ~n50143 & ~n50144 ;
  assign n50146 = ~n50142 & n50145 ;
  assign n50147 = n18028 & n19026 ;
  assign n50148 = n50146 & ~n50147 ;
  assign n50149 = x53 & ~n50148 ;
  assign n50150 = x53 & ~n50149 ;
  assign n50151 = ~n50148 & ~n50149 ;
  assign n50152 = ~n50150 & ~n50151 ;
  assign n50153 = ~n49843 & ~n49856 ;
  assign n50154 = ~n49823 & ~n49837 ;
  assign n50155 = ~n49806 & ~n49820 ;
  assign n50156 = x104 & n27024 ;
  assign n50157 = x105 & ~n26217 ;
  assign n50158 = ~n50156 & ~n50157 ;
  assign n50159 = n49803 & ~n50158 ;
  assign n50160 = n49803 & ~n50159 ;
  assign n50161 = ~n50158 & ~n50159 ;
  assign n50162 = ~n50160 & ~n50161 ;
  assign n50163 = ~n50155 & ~n50162 ;
  assign n50164 = ~n50155 & ~n50163 ;
  assign n50165 = ~n50162 & ~n50163 ;
  assign n50166 = ~n50164 & ~n50165 ;
  assign n50167 = x108 & n24612 ;
  assign n50168 = x106 & n25390 ;
  assign n50169 = x107 & n24607 ;
  assign n50170 = ~n50168 & ~n50169 ;
  assign n50171 = ~n50167 & n50170 ;
  assign n50172 = n13323 & n24615 ;
  assign n50173 = n50171 & ~n50172 ;
  assign n50174 = x62 & ~n50173 ;
  assign n50175 = x62 & ~n50174 ;
  assign n50176 = ~n50173 & ~n50174 ;
  assign n50177 = ~n50175 & ~n50176 ;
  assign n50178 = ~n50166 & n50177 ;
  assign n50179 = n50166 & ~n50177 ;
  assign n50180 = ~n50178 & ~n50179 ;
  assign n50181 = x111 & n22325 ;
  assign n50182 = x109 & n23066 ;
  assign n50183 = x110 & n22320 ;
  assign n50184 = ~n50182 & ~n50183 ;
  assign n50185 = ~n50181 & n50184 ;
  assign n50186 = n15111 & n22328 ;
  assign n50187 = n50185 & ~n50186 ;
  assign n50188 = x59 & ~n50187 ;
  assign n50189 = x59 & ~n50188 ;
  assign n50190 = ~n50187 & ~n50188 ;
  assign n50191 = ~n50189 & ~n50190 ;
  assign n50192 = ~n50180 & ~n50191 ;
  assign n50193 = n50180 & n50191 ;
  assign n50194 = ~n50192 & ~n50193 ;
  assign n50195 = n50154 & ~n50194 ;
  assign n50196 = ~n50154 & n50194 ;
  assign n50197 = ~n50195 & ~n50196 ;
  assign n50198 = x114 & n20143 ;
  assign n50199 = x112 & n20854 ;
  assign n50200 = x113 & n20138 ;
  assign n50201 = ~n50199 & ~n50200 ;
  assign n50202 = ~n50198 & n50201 ;
  assign n50203 = n17012 & n20146 ;
  assign n50204 = n50202 & ~n50203 ;
  assign n50205 = x56 & ~n50204 ;
  assign n50206 = x56 & ~n50205 ;
  assign n50207 = ~n50204 & ~n50205 ;
  assign n50208 = ~n50206 & ~n50207 ;
  assign n50209 = ~n50197 & n50208 ;
  assign n50210 = n50197 & ~n50208 ;
  assign n50211 = ~n50209 & ~n50210 ;
  assign n50212 = ~n50153 & n50211 ;
  assign n50213 = ~n50153 & ~n50212 ;
  assign n50214 = n50211 & ~n50212 ;
  assign n50215 = ~n50213 & ~n50214 ;
  assign n50216 = ~n50152 & ~n50215 ;
  assign n50217 = n50152 & ~n50214 ;
  assign n50218 = ~n50213 & n50217 ;
  assign n50219 = ~n50216 & ~n50218 ;
  assign n50220 = ~n50141 & n50219 ;
  assign n50221 = ~n50141 & ~n50220 ;
  assign n50222 = n50219 & ~n50220 ;
  assign n50223 = ~n50221 & ~n50222 ;
  assign n50224 = ~n50140 & ~n50223 ;
  assign n50225 = n50140 & ~n50222 ;
  assign n50226 = ~n50221 & n50225 ;
  assign n50227 = ~n50224 & ~n50226 ;
  assign n50228 = ~n50129 & n50227 ;
  assign n50229 = n50129 & ~n50227 ;
  assign n50230 = ~n50228 & ~n50229 ;
  assign n50231 = x123 & n14233 ;
  assign n50232 = x121 & n14876 ;
  assign n50233 = x122 & n14228 ;
  assign n50234 = ~n50232 & ~n50233 ;
  assign n50235 = ~n50231 & n50234 ;
  assign n50236 = n14236 & n23382 ;
  assign n50237 = n50235 & ~n50236 ;
  assign n50238 = x47 & ~n50237 ;
  assign n50239 = x47 & ~n50238 ;
  assign n50240 = ~n50237 & ~n50238 ;
  assign n50241 = ~n50239 & ~n50240 ;
  assign n50242 = n50230 & ~n50241 ;
  assign n50243 = n50230 & ~n50242 ;
  assign n50244 = ~n50241 & ~n50242 ;
  assign n50245 = ~n50243 & ~n50244 ;
  assign n50246 = ~n49901 & ~n49914 ;
  assign n50247 = n50245 & n50246 ;
  assign n50248 = ~n50245 & ~n50246 ;
  assign n50249 = ~n50247 & ~n50248 ;
  assign n50250 = x126 & n12506 ;
  assign n50251 = x124 & n13131 ;
  assign n50252 = x125 & n12501 ;
  assign n50253 = ~n50251 & ~n50252 ;
  assign n50254 = ~n50250 & n50253 ;
  assign n50255 = n12509 & n25735 ;
  assign n50256 = n50254 & ~n50255 ;
  assign n50257 = x44 & ~n50256 ;
  assign n50258 = x44 & ~n50257 ;
  assign n50259 = ~n50256 & ~n50257 ;
  assign n50260 = ~n50258 & ~n50259 ;
  assign n50261 = n50249 & ~n50260 ;
  assign n50262 = n50249 & ~n50261 ;
  assign n50263 = ~n50260 & ~n50261 ;
  assign n50264 = ~n50262 & ~n50263 ;
  assign n50265 = ~n50128 & n50264 ;
  assign n50266 = n50128 & ~n50264 ;
  assign n50267 = ~n50265 & ~n50266 ;
  assign n50268 = ~n50116 & ~n50267 ;
  assign n50269 = n50116 & n50267 ;
  assign n50270 = ~n50268 & ~n50269 ;
  assign n50271 = ~n50115 & n50270 ;
  assign n50272 = n50115 & ~n50270 ;
  assign n50273 = ~n50271 & ~n50272 ;
  assign n50434 = n50273 & x232 ;
  assign n50274 = ~n50105 & ~n50108 ;
  assign n50275 = ~n49959 & ~n50098 ;
  assign n50276 = ~n50082 & ~n50095 ;
  assign n50277 = ~x127 & n11466 ;
  assign n50278 = n10908 & n27365 ;
  assign n50279 = ~n50277 & ~n50278 ;
  assign n50280 = ~x41 & ~n50279 ;
  assign n50281 = ~x41 & ~n50280 ;
  assign n50282 = ~n50279 & ~n50280 ;
  assign n50283 = ~n50281 & ~n50282 ;
  assign n50284 = ~n50276 & ~n50283 ;
  assign n50285 = ~n50276 & ~n50284 ;
  assign n50286 = ~n50283 & ~n50284 ;
  assign n50287 = ~n50285 & ~n50286 ;
  assign n50288 = ~n50042 & ~n50057 ;
  assign n50289 = ~x120 & n16076 ;
  assign n50290 = ~x118 & n16756 ;
  assign n50291 = ~x119 & n16071 ;
  assign n50292 = ~n50290 & ~n50291 ;
  assign n50293 = ~n50289 & n50292 ;
  assign n50294 = n16079 & n21501 ;
  assign n50295 = n50293 & ~n50294 ;
  assign n50296 = ~x50 & ~n50295 ;
  assign n50297 = ~x50 & ~n50296 ;
  assign n50298 = ~n50295 & ~n50296 ;
  assign n50299 = ~n50297 & ~n50298 ;
  assign n50300 = ~n50024 & ~n50037 ;
  assign n50301 = ~x117 & n18025 ;
  assign n50302 = ~x115 & n18764 ;
  assign n50303 = ~x116 & n18020 ;
  assign n50304 = ~n50302 & ~n50303 ;
  assign n50305 = ~n50301 & n50304 ;
  assign n50306 = n18028 & n19365 ;
  assign n50307 = n50305 & ~n50306 ;
  assign n50308 = ~x53 & ~n50307 ;
  assign n50309 = ~x53 & ~n50308 ;
  assign n50310 = ~n50307 & ~n50308 ;
  assign n50311 = ~n50309 & ~n50310 ;
  assign n50312 = ~n50005 & ~n50018 ;
  assign n50313 = ~n49985 & ~n49999 ;
  assign n50314 = ~n49968 & ~n49982 ;
  assign n50315 = ~x104 & n27427 ;
  assign n50316 = ~x105 & ~n26217 ;
  assign n50317 = ~n50315 & ~n50316 ;
  assign n50318 = n49965 & ~n50317 ;
  assign n50319 = n49965 & ~n50318 ;
  assign n50320 = ~n50317 & ~n50318 ;
  assign n50321 = ~n50319 & ~n50320 ;
  assign n50322 = ~n50314 & ~n50321 ;
  assign n50323 = ~n50314 & ~n50322 ;
  assign n50324 = ~n50321 & ~n50322 ;
  assign n50325 = ~n50323 & ~n50324 ;
  assign n50326 = ~x108 & n24612 ;
  assign n50327 = ~x106 & n25390 ;
  assign n50328 = ~x107 & n24607 ;
  assign n50329 = ~n50327 & ~n50328 ;
  assign n50330 = ~n50326 & n50329 ;
  assign n50331 = n13601 & n24615 ;
  assign n50332 = n50330 & ~n50331 ;
  assign n50333 = ~x62 & ~n50332 ;
  assign n50334 = ~x62 & ~n50333 ;
  assign n50335 = ~n50332 & ~n50333 ;
  assign n50336 = ~n50334 & ~n50335 ;
  assign n50337 = ~n50325 & n50336 ;
  assign n50338 = n50325 & ~n50336 ;
  assign n50339 = ~n50337 & ~n50338 ;
  assign n50340 = ~x111 & n22325 ;
  assign n50341 = ~x109 & n23066 ;
  assign n50342 = ~x110 & n22320 ;
  assign n50343 = ~n50341 & ~n50342 ;
  assign n50344 = ~n50340 & n50343 ;
  assign n50345 = n15411 & n22328 ;
  assign n50346 = n50344 & ~n50345 ;
  assign n50347 = ~x59 & ~n50346 ;
  assign n50348 = ~x59 & ~n50347 ;
  assign n50349 = ~n50346 & ~n50347 ;
  assign n50350 = ~n50348 & ~n50349 ;
  assign n50351 = ~n50339 & ~n50350 ;
  assign n50352 = n50339 & n50350 ;
  assign n50353 = ~n50351 & ~n50352 ;
  assign n50354 = n50313 & ~n50353 ;
  assign n50355 = ~n50313 & n50353 ;
  assign n50356 = ~n50354 & ~n50355 ;
  assign n50357 = ~x114 & n20143 ;
  assign n50358 = ~x112 & n20854 ;
  assign n50359 = ~x113 & n20138 ;
  assign n50360 = ~n50358 & ~n50359 ;
  assign n50361 = ~n50357 & n50360 ;
  assign n50362 = n17333 & n20146 ;
  assign n50363 = n50361 & ~n50362 ;
  assign n50364 = ~x56 & ~n50363 ;
  assign n50365 = ~x56 & ~n50364 ;
  assign n50366 = ~n50363 & ~n50364 ;
  assign n50367 = ~n50365 & ~n50366 ;
  assign n50368 = ~n50356 & n50367 ;
  assign n50369 = n50356 & ~n50367 ;
  assign n50370 = ~n50368 & ~n50369 ;
  assign n50371 = ~n50312 & n50370 ;
  assign n50372 = ~n50312 & ~n50371 ;
  assign n50373 = n50370 & ~n50371 ;
  assign n50374 = ~n50372 & ~n50373 ;
  assign n50375 = ~n50311 & ~n50374 ;
  assign n50376 = n50311 & ~n50373 ;
  assign n50377 = ~n50372 & n50376 ;
  assign n50378 = ~n50375 & ~n50377 ;
  assign n50379 = ~n50300 & n50378 ;
  assign n50380 = ~n50300 & ~n50379 ;
  assign n50381 = n50378 & ~n50379 ;
  assign n50382 = ~n50380 & ~n50381 ;
  assign n50383 = ~n50299 & ~n50382 ;
  assign n50384 = n50299 & ~n50381 ;
  assign n50385 = ~n50380 & n50384 ;
  assign n50386 = ~n50383 & ~n50385 ;
  assign n50387 = ~n50288 & n50386 ;
  assign n50388 = n50288 & ~n50386 ;
  assign n50389 = ~n50387 & ~n50388 ;
  assign n50390 = ~x123 & n14233 ;
  assign n50391 = ~x121 & n14876 ;
  assign n50392 = ~x122 & n14228 ;
  assign n50393 = ~n50391 & ~n50392 ;
  assign n50394 = ~n50390 & n50393 ;
  assign n50395 = n14236 & n23760 ;
  assign n50396 = n50394 & ~n50395 ;
  assign n50397 = ~x47 & ~n50396 ;
  assign n50398 = ~x47 & ~n50397 ;
  assign n50399 = ~n50396 & ~n50397 ;
  assign n50400 = ~n50398 & ~n50399 ;
  assign n50401 = n50389 & ~n50400 ;
  assign n50402 = n50389 & ~n50401 ;
  assign n50403 = ~n50400 & ~n50401 ;
  assign n50404 = ~n50402 & ~n50403 ;
  assign n50405 = ~n50063 & ~n50076 ;
  assign n50406 = n50404 & n50405 ;
  assign n50407 = ~n50404 & ~n50405 ;
  assign n50408 = ~n50406 & ~n50407 ;
  assign n50409 = ~x126 & n12506 ;
  assign n50410 = ~x124 & n13131 ;
  assign n50411 = ~x125 & n12501 ;
  assign n50412 = ~n50410 & ~n50411 ;
  assign n50413 = ~n50409 & n50412 ;
  assign n50414 = n12509 & n26128 ;
  assign n50415 = n50413 & ~n50414 ;
  assign n50416 = ~x44 & ~n50415 ;
  assign n50417 = ~x44 & ~n50416 ;
  assign n50418 = ~n50415 & ~n50416 ;
  assign n50419 = ~n50417 & ~n50418 ;
  assign n50420 = n50408 & ~n50419 ;
  assign n50421 = n50408 & ~n50420 ;
  assign n50422 = ~n50419 & ~n50420 ;
  assign n50423 = ~n50421 & ~n50422 ;
  assign n50424 = ~n50287 & n50423 ;
  assign n50425 = n50287 & ~n50423 ;
  assign n50426 = ~n50424 & ~n50425 ;
  assign n50427 = ~n50275 & ~n50426 ;
  assign n50428 = n50275 & n50426 ;
  assign n50429 = ~n50427 & ~n50428 ;
  assign n50430 = ~n50274 & n50429 ;
  assign n50431 = n50274 & ~n50429 ;
  assign n50432 = ~n50430 & ~n50431 ;
  assign n50435 = ~n50432 & ~x232 ;
  assign n50436 = ~n50434 & ~n50435 ;
  assign n50437 = ~n50268 & ~n50271 ;
  assign n50438 = ~n50220 & ~n50224 ;
  assign n50439 = x121 & n16076 ;
  assign n50440 = x119 & n16756 ;
  assign n50441 = x120 & n16071 ;
  assign n50442 = ~n50440 & ~n50441 ;
  assign n50443 = ~n50439 & n50442 ;
  assign n50444 = n16079 & n21870 ;
  assign n50445 = n50443 & ~n50444 ;
  assign n50446 = x50 & ~n50445 ;
  assign n50447 = x50 & ~n50446 ;
  assign n50448 = ~n50445 & ~n50446 ;
  assign n50449 = ~n50447 & ~n50448 ;
  assign n50450 = ~n50212 & ~n50216 ;
  assign n50451 = ~n50196 & ~n50210 ;
  assign n50452 = x115 & n20143 ;
  assign n50453 = x113 & n20854 ;
  assign n50454 = x114 & n20138 ;
  assign n50455 = ~n50453 & ~n50454 ;
  assign n50456 = ~n50452 & n50455 ;
  assign n50457 = n17364 & n20146 ;
  assign n50458 = n50456 & ~n50457 ;
  assign n50459 = x56 & ~n50458 ;
  assign n50460 = x56 & ~n50459 ;
  assign n50461 = ~n50458 & ~n50459 ;
  assign n50462 = ~n50460 & ~n50461 ;
  assign n50463 = x41 & ~n49803 ;
  assign n50464 = ~x41 & n49803 ;
  assign n50465 = ~n50463 & ~n50464 ;
  assign n50466 = x105 & n27024 ;
  assign n50467 = x106 & ~n26217 ;
  assign n50468 = ~n50466 & ~n50467 ;
  assign n50469 = n50465 & n50468 ;
  assign n50470 = ~n50465 & ~n50468 ;
  assign n50471 = ~n50469 & ~n50470 ;
  assign n50472 = x109 & n24612 ;
  assign n50473 = x107 & n25390 ;
  assign n50474 = x108 & n24607 ;
  assign n50475 = ~n50473 & ~n50474 ;
  assign n50476 = ~n50472 & n50475 ;
  assign n50477 = n13894 & n24615 ;
  assign n50478 = n50476 & ~n50477 ;
  assign n50479 = x62 & ~n50478 ;
  assign n50480 = x62 & ~n50479 ;
  assign n50481 = ~n50478 & ~n50479 ;
  assign n50482 = ~n50480 & ~n50481 ;
  assign n50483 = n50471 & ~n50482 ;
  assign n50484 = n50471 & ~n50483 ;
  assign n50485 = ~n50482 & ~n50483 ;
  assign n50486 = ~n50484 & ~n50485 ;
  assign n50487 = ~n50159 & ~n50163 ;
  assign n50488 = n50486 & n50487 ;
  assign n50489 = ~n50486 & ~n50487 ;
  assign n50490 = ~n50488 & ~n50489 ;
  assign n50491 = x112 & n22325 ;
  assign n50492 = x110 & n23066 ;
  assign n50493 = x111 & n22320 ;
  assign n50494 = ~n50492 & ~n50493 ;
  assign n50495 = ~n50491 & n50494 ;
  assign n50496 = n15442 & n22328 ;
  assign n50497 = n50495 & ~n50496 ;
  assign n50498 = x59 & ~n50497 ;
  assign n50499 = x59 & ~n50498 ;
  assign n50500 = ~n50497 & ~n50498 ;
  assign n50501 = ~n50499 & ~n50500 ;
  assign n50502 = n50490 & ~n50501 ;
  assign n50503 = n50490 & ~n50502 ;
  assign n50504 = ~n50501 & ~n50502 ;
  assign n50505 = ~n50503 & ~n50504 ;
  assign n50506 = ~n50166 & ~n50177 ;
  assign n50507 = ~n50192 & ~n50506 ;
  assign n50508 = ~n50505 & ~n50507 ;
  assign n50509 = n50505 & n50507 ;
  assign n50510 = ~n50508 & ~n50509 ;
  assign n50511 = ~n50462 & n50510 ;
  assign n50512 = ~n50462 & ~n50511 ;
  assign n50513 = n50510 & ~n50511 ;
  assign n50514 = ~n50512 & ~n50513 ;
  assign n50515 = ~n50451 & ~n50514 ;
  assign n50516 = ~n50451 & ~n50515 ;
  assign n50517 = ~n50514 & ~n50515 ;
  assign n50518 = ~n50516 & ~n50517 ;
  assign n50519 = x118 & n18025 ;
  assign n50520 = x116 & n18764 ;
  assign n50521 = x117 & n18020 ;
  assign n50522 = ~n50520 & ~n50521 ;
  assign n50523 = ~n50519 & n50522 ;
  assign n50524 = n18028 & n19395 ;
  assign n50525 = n50523 & ~n50524 ;
  assign n50526 = x53 & ~n50525 ;
  assign n50527 = x53 & ~n50526 ;
  assign n50528 = ~n50525 & ~n50526 ;
  assign n50529 = ~n50527 & ~n50528 ;
  assign n50530 = n50518 & n50529 ;
  assign n50531 = ~n50518 & ~n50529 ;
  assign n50532 = ~n50530 & ~n50531 ;
  assign n50533 = ~n50450 & n50532 ;
  assign n50534 = n50450 & ~n50532 ;
  assign n50535 = ~n50533 & ~n50534 ;
  assign n50536 = n50449 & ~n50535 ;
  assign n50537 = ~n50449 & n50535 ;
  assign n50538 = ~n50536 & ~n50537 ;
  assign n50539 = ~n50438 & n50538 ;
  assign n50540 = n50438 & ~n50538 ;
  assign n50541 = ~n50539 & ~n50540 ;
  assign n50542 = x124 & n14233 ;
  assign n50543 = x122 & n14876 ;
  assign n50544 = x123 & n14228 ;
  assign n50545 = ~n50543 & ~n50544 ;
  assign n50546 = ~n50542 & n50545 ;
  assign n50547 = n14236 & n23796 ;
  assign n50548 = n50546 & ~n50547 ;
  assign n50549 = x47 & ~n50548 ;
  assign n50550 = x47 & ~n50549 ;
  assign n50551 = ~n50548 & ~n50549 ;
  assign n50552 = ~n50550 & ~n50551 ;
  assign n50553 = n50541 & ~n50552 ;
  assign n50554 = n50541 & ~n50553 ;
  assign n50555 = ~n50552 & ~n50553 ;
  assign n50556 = ~n50554 & ~n50555 ;
  assign n50557 = ~n50228 & ~n50242 ;
  assign n50558 = n50556 & n50557 ;
  assign n50559 = ~n50556 & ~n50557 ;
  assign n50560 = ~n50558 & ~n50559 ;
  assign n50561 = x127 & n12506 ;
  assign n50562 = x125 & n13131 ;
  assign n50563 = x126 & n12501 ;
  assign n50564 = ~n50562 & ~n50563 ;
  assign n50565 = ~n50561 & n50564 ;
  assign n50566 = n12509 & n26533 ;
  assign n50567 = n50565 & ~n50566 ;
  assign n50568 = x44 & ~n50567 ;
  assign n50569 = x44 & ~n50568 ;
  assign n50570 = ~n50567 & ~n50568 ;
  assign n50571 = ~n50569 & ~n50570 ;
  assign n50572 = n50560 & ~n50571 ;
  assign n50573 = n50560 & ~n50572 ;
  assign n50574 = ~n50571 & ~n50572 ;
  assign n50575 = ~n50573 & ~n50574 ;
  assign n50576 = ~n50248 & ~n50261 ;
  assign n50577 = n50575 & n50576 ;
  assign n50578 = ~n50575 & ~n50576 ;
  assign n50579 = ~n50577 & ~n50578 ;
  assign n50580 = ~n50128 & ~n50264 ;
  assign n50581 = ~n50125 & ~n50580 ;
  assign n50582 = n50579 & ~n50581 ;
  assign n50583 = ~n50579 & n50581 ;
  assign n50584 = ~n50582 & ~n50583 ;
  assign n50585 = ~n50437 & n50584 ;
  assign n50586 = n50437 & ~n50584 ;
  assign n50587 = ~n50585 & ~n50586 ;
  assign n50740 = n50587 & x233 ;
  assign n50588 = ~n50427 & ~n50430 ;
  assign n50589 = ~n50379 & ~n50383 ;
  assign n50590 = ~x121 & n16076 ;
  assign n50591 = ~x119 & n16756 ;
  assign n50592 = ~x120 & n16071 ;
  assign n50593 = ~n50591 & ~n50592 ;
  assign n50594 = ~n50590 & n50593 ;
  assign n50595 = n16079 & n22229 ;
  assign n50596 = n50594 & ~n50595 ;
  assign n50597 = ~x50 & ~n50596 ;
  assign n50598 = ~x50 & ~n50597 ;
  assign n50599 = ~n50596 & ~n50597 ;
  assign n50600 = ~n50598 & ~n50599 ;
  assign n50601 = ~n50371 & ~n50375 ;
  assign n50602 = ~n50355 & ~n50369 ;
  assign n50603 = ~x115 & n20143 ;
  assign n50604 = ~x113 & n20854 ;
  assign n50605 = ~x114 & n20138 ;
  assign n50606 = ~n50604 & ~n50605 ;
  assign n50607 = ~n50603 & n50606 ;
  assign n50608 = n17683 & n20146 ;
  assign n50609 = n50607 & ~n50608 ;
  assign n50610 = ~x56 & ~n50609 ;
  assign n50611 = ~x56 & ~n50610 ;
  assign n50612 = ~n50609 & ~n50610 ;
  assign n50613 = ~n50611 & ~n50612 ;
  assign n50614 = ~x41 & ~n49965 ;
  assign n50615 = x41 & n49965 ;
  assign n50616 = ~n50614 & ~n50615 ;
  assign n50617 = ~x105 & n27427 ;
  assign n50618 = ~x106 & ~n26217 ;
  assign n50619 = ~n50617 & ~n50618 ;
  assign n50620 = n50616 & n50619 ;
  assign n50621 = ~n50616 & ~n50619 ;
  assign n50622 = ~n50620 & ~n50621 ;
  assign n50623 = ~x109 & n24612 ;
  assign n50624 = ~x107 & n25390 ;
  assign n50625 = ~x108 & n24607 ;
  assign n50626 = ~n50624 & ~n50625 ;
  assign n50627 = ~n50623 & n50626 ;
  assign n50628 = n14177 & n24615 ;
  assign n50629 = n50627 & ~n50628 ;
  assign n50630 = ~x62 & ~n50629 ;
  assign n50631 = ~x62 & ~n50630 ;
  assign n50632 = ~n50629 & ~n50630 ;
  assign n50633 = ~n50631 & ~n50632 ;
  assign n50634 = n50622 & ~n50633 ;
  assign n50635 = n50622 & ~n50634 ;
  assign n50636 = ~n50633 & ~n50634 ;
  assign n50637 = ~n50635 & ~n50636 ;
  assign n50638 = ~n50318 & ~n50322 ;
  assign n50639 = n50637 & n50638 ;
  assign n50640 = ~n50637 & ~n50638 ;
  assign n50641 = ~n50639 & ~n50640 ;
  assign n50642 = ~x112 & n22325 ;
  assign n50643 = ~x110 & n23066 ;
  assign n50644 = ~x111 & n22320 ;
  assign n50645 = ~n50643 & ~n50644 ;
  assign n50646 = ~n50642 & n50645 ;
  assign n50647 = n15744 & n22328 ;
  assign n50648 = n50646 & ~n50647 ;
  assign n50649 = ~x59 & ~n50648 ;
  assign n50650 = ~x59 & ~n50649 ;
  assign n50651 = ~n50648 & ~n50649 ;
  assign n50652 = ~n50650 & ~n50651 ;
  assign n50653 = n50641 & ~n50652 ;
  assign n50654 = n50641 & ~n50653 ;
  assign n50655 = ~n50652 & ~n50653 ;
  assign n50656 = ~n50654 & ~n50655 ;
  assign n50657 = ~n50325 & ~n50336 ;
  assign n50658 = ~n50351 & ~n50657 ;
  assign n50659 = ~n50656 & ~n50658 ;
  assign n50660 = n50656 & n50658 ;
  assign n50661 = ~n50659 & ~n50660 ;
  assign n50662 = ~n50613 & n50661 ;
  assign n50663 = ~n50613 & ~n50662 ;
  assign n50664 = n50661 & ~n50662 ;
  assign n50665 = ~n50663 & ~n50664 ;
  assign n50666 = ~n50602 & ~n50665 ;
  assign n50667 = ~n50602 & ~n50666 ;
  assign n50668 = ~n50665 & ~n50666 ;
  assign n50669 = ~n50667 & ~n50668 ;
  assign n50670 = ~x118 & n18025 ;
  assign n50671 = ~x116 & n18764 ;
  assign n50672 = ~x117 & n18020 ;
  assign n50673 = ~n50671 & ~n50672 ;
  assign n50674 = ~n50670 & n50673 ;
  assign n50675 = n18028 & n19736 ;
  assign n50676 = n50674 & ~n50675 ;
  assign n50677 = ~x53 & ~n50676 ;
  assign n50678 = ~x53 & ~n50677 ;
  assign n50679 = ~n50676 & ~n50677 ;
  assign n50680 = ~n50678 & ~n50679 ;
  assign n50681 = n50669 & n50680 ;
  assign n50682 = ~n50669 & ~n50680 ;
  assign n50683 = ~n50681 & ~n50682 ;
  assign n50684 = ~n50601 & n50683 ;
  assign n50685 = n50601 & ~n50683 ;
  assign n50686 = ~n50684 & ~n50685 ;
  assign n50687 = n50600 & ~n50686 ;
  assign n50688 = ~n50600 & n50686 ;
  assign n50689 = ~n50687 & ~n50688 ;
  assign n50690 = ~n50589 & n50689 ;
  assign n50691 = n50589 & ~n50689 ;
  assign n50692 = ~n50690 & ~n50691 ;
  assign n50693 = ~x124 & n14233 ;
  assign n50694 = ~x122 & n14876 ;
  assign n50695 = ~x123 & n14228 ;
  assign n50696 = ~n50694 & ~n50695 ;
  assign n50697 = ~n50693 & n50696 ;
  assign n50698 = n14236 & n24176 ;
  assign n50699 = n50697 & ~n50698 ;
  assign n50700 = ~x47 & ~n50699 ;
  assign n50701 = ~x47 & ~n50700 ;
  assign n50702 = ~n50699 & ~n50700 ;
  assign n50703 = ~n50701 & ~n50702 ;
  assign n50704 = n50692 & ~n50703 ;
  assign n50705 = n50692 & ~n50704 ;
  assign n50706 = ~n50703 & ~n50704 ;
  assign n50707 = ~n50705 & ~n50706 ;
  assign n50708 = ~n50387 & ~n50401 ;
  assign n50709 = n50707 & n50708 ;
  assign n50710 = ~n50707 & ~n50708 ;
  assign n50711 = ~n50709 & ~n50710 ;
  assign n50712 = ~x127 & n12506 ;
  assign n50713 = ~x125 & n13131 ;
  assign n50714 = ~x126 & n12501 ;
  assign n50715 = ~n50713 & ~n50714 ;
  assign n50716 = ~n50712 & n50715 ;
  assign n50717 = n12509 & n26932 ;
  assign n50718 = n50716 & ~n50717 ;
  assign n50719 = ~x44 & ~n50718 ;
  assign n50720 = ~x44 & ~n50719 ;
  assign n50721 = ~n50718 & ~n50719 ;
  assign n50722 = ~n50720 & ~n50721 ;
  assign n50723 = n50711 & ~n50722 ;
  assign n50724 = n50711 & ~n50723 ;
  assign n50725 = ~n50722 & ~n50723 ;
  assign n50726 = ~n50724 & ~n50725 ;
  assign n50727 = ~n50407 & ~n50420 ;
  assign n50728 = n50726 & n50727 ;
  assign n50729 = ~n50726 & ~n50727 ;
  assign n50730 = ~n50728 & ~n50729 ;
  assign n50731 = ~n50287 & ~n50423 ;
  assign n50732 = ~n50284 & ~n50731 ;
  assign n50733 = n50730 & ~n50732 ;
  assign n50734 = ~n50730 & n50732 ;
  assign n50735 = ~n50733 & ~n50734 ;
  assign n50736 = ~n50588 & n50735 ;
  assign n50737 = n50588 & ~n50735 ;
  assign n50738 = ~n50736 & ~n50737 ;
  assign n50741 = ~n50738 & ~x233 ;
  assign n50742 = ~n50740 & ~n50741 ;
  assign n50743 = ~n50553 & ~n50559 ;
  assign n50744 = x126 & n13131 ;
  assign n50745 = x127 & n12501 ;
  assign n50746 = ~n50744 & ~n50745 ;
  assign n50747 = ~n12509 & n50746 ;
  assign n50748 = n26965 & n50746 ;
  assign n50749 = ~n50747 & ~n50748 ;
  assign n50750 = x44 & ~n50749 ;
  assign n50751 = ~x44 & n50749 ;
  assign n50752 = ~n50750 & ~n50751 ;
  assign n50753 = ~n50743 & ~n50752 ;
  assign n50754 = n50743 & n50752 ;
  assign n50755 = ~n50753 & ~n50754 ;
  assign n50756 = x125 & n14233 ;
  assign n50757 = x123 & n14876 ;
  assign n50758 = x124 & n14228 ;
  assign n50759 = ~n50757 & ~n50758 ;
  assign n50760 = ~n50756 & n50759 ;
  assign n50761 = n14236 & n24935 ;
  assign n50762 = n50760 & ~n50761 ;
  assign n50763 = x47 & ~n50762 ;
  assign n50764 = x47 & ~n50763 ;
  assign n50765 = ~n50762 & ~n50763 ;
  assign n50766 = ~n50764 & ~n50765 ;
  assign n50767 = ~n50537 & ~n50539 ;
  assign n50768 = ~n50531 & ~n50533 ;
  assign n50769 = ~n50483 & ~n50489 ;
  assign n50770 = x106 & n27024 ;
  assign n50771 = x107 & ~n26217 ;
  assign n50772 = ~n50770 & ~n50771 ;
  assign n50773 = ~x41 & ~n49803 ;
  assign n50774 = ~n50470 & ~n50773 ;
  assign n50775 = n50772 & ~n50774 ;
  assign n50776 = n50772 & ~n50775 ;
  assign n50777 = ~n50774 & ~n50775 ;
  assign n50778 = ~n50776 & ~n50777 ;
  assign n50779 = x110 & n24612 ;
  assign n50780 = x108 & n25390 ;
  assign n50781 = x109 & n24607 ;
  assign n50782 = ~n50780 & ~n50781 ;
  assign n50783 = ~n50779 & n50782 ;
  assign n50784 = ~n24615 & n50783 ;
  assign n50785 = ~n14497 & n50783 ;
  assign n50786 = ~n50784 & ~n50785 ;
  assign n50787 = x62 & ~n50786 ;
  assign n50788 = ~x62 & n50786 ;
  assign n50789 = ~n50787 & ~n50788 ;
  assign n50790 = ~n50778 & ~n50789 ;
  assign n50791 = n50778 & n50789 ;
  assign n50792 = ~n50790 & ~n50791 ;
  assign n50793 = ~n50769 & n50792 ;
  assign n50794 = n50769 & ~n50792 ;
  assign n50795 = ~n50793 & ~n50794 ;
  assign n50796 = x113 & n22325 ;
  assign n50797 = x111 & n23066 ;
  assign n50798 = x112 & n22320 ;
  assign n50799 = ~n50797 & ~n50798 ;
  assign n50800 = ~n50796 & n50799 ;
  assign n50801 = n16361 & n22328 ;
  assign n50802 = n50800 & ~n50801 ;
  assign n50803 = x59 & ~n50802 ;
  assign n50804 = x59 & ~n50803 ;
  assign n50805 = ~n50802 & ~n50803 ;
  assign n50806 = ~n50804 & ~n50805 ;
  assign n50807 = n50795 & ~n50806 ;
  assign n50808 = n50795 & ~n50807 ;
  assign n50809 = ~n50806 & ~n50807 ;
  assign n50810 = ~n50808 & ~n50809 ;
  assign n50811 = ~n50502 & ~n50508 ;
  assign n50812 = n50810 & n50811 ;
  assign n50813 = ~n50810 & ~n50811 ;
  assign n50814 = ~n50812 & ~n50813 ;
  assign n50815 = x116 & n20143 ;
  assign n50816 = x114 & n20854 ;
  assign n50817 = x115 & n20138 ;
  assign n50818 = ~n50816 & ~n50817 ;
  assign n50819 = ~n50815 & n50818 ;
  assign n50820 = n18336 & n20146 ;
  assign n50821 = n50819 & ~n50820 ;
  assign n50822 = x56 & ~n50821 ;
  assign n50823 = x56 & ~n50822 ;
  assign n50824 = ~n50821 & ~n50822 ;
  assign n50825 = ~n50823 & ~n50824 ;
  assign n50826 = n50814 & ~n50825 ;
  assign n50827 = n50814 & ~n50826 ;
  assign n50828 = ~n50825 & ~n50826 ;
  assign n50829 = ~n50827 & ~n50828 ;
  assign n50830 = ~n50511 & ~n50515 ;
  assign n50831 = n50829 & n50830 ;
  assign n50832 = ~n50829 & ~n50830 ;
  assign n50833 = ~n50831 & ~n50832 ;
  assign n50834 = x119 & n18025 ;
  assign n50835 = x117 & n18764 ;
  assign n50836 = x118 & n18020 ;
  assign n50837 = ~n50835 & ~n50836 ;
  assign n50838 = ~n50834 & n50837 ;
  assign n50839 = n18028 & n20423 ;
  assign n50840 = n50838 & ~n50839 ;
  assign n50841 = x53 & ~n50840 ;
  assign n50842 = x53 & ~n50841 ;
  assign n50843 = ~n50840 & ~n50841 ;
  assign n50844 = ~n50842 & ~n50843 ;
  assign n50845 = n50833 & ~n50844 ;
  assign n50846 = n50833 & ~n50845 ;
  assign n50847 = ~n50844 & ~n50845 ;
  assign n50848 = ~n50846 & ~n50847 ;
  assign n50849 = ~n50768 & n50848 ;
  assign n50850 = n50768 & ~n50848 ;
  assign n50851 = ~n50849 & ~n50850 ;
  assign n50852 = x122 & n16076 ;
  assign n50853 = x120 & n16756 ;
  assign n50854 = x121 & n16071 ;
  assign n50855 = ~n50853 & ~n50854 ;
  assign n50856 = ~n50852 & n50855 ;
  assign n50857 = n16079 & n22622 ;
  assign n50858 = n50856 & ~n50857 ;
  assign n50859 = x50 & ~n50858 ;
  assign n50860 = x50 & ~n50859 ;
  assign n50861 = ~n50858 & ~n50859 ;
  assign n50862 = ~n50860 & ~n50861 ;
  assign n50863 = n50851 & n50862 ;
  assign n50864 = ~n50851 & ~n50862 ;
  assign n50865 = ~n50863 & ~n50864 ;
  assign n50866 = ~n50767 & n50865 ;
  assign n50867 = ~n50767 & ~n50866 ;
  assign n50868 = n50865 & ~n50866 ;
  assign n50869 = ~n50867 & ~n50868 ;
  assign n50870 = ~n50766 & ~n50869 ;
  assign n50871 = ~n50766 & ~n50870 ;
  assign n50872 = ~n50869 & ~n50870 ;
  assign n50873 = ~n50871 & ~n50872 ;
  assign n50874 = n50755 & ~n50873 ;
  assign n50875 = n50755 & ~n50874 ;
  assign n50876 = ~n50873 & ~n50874 ;
  assign n50877 = ~n50875 & ~n50876 ;
  assign n50878 = ~n50572 & ~n50578 ;
  assign n50879 = n50877 & n50878 ;
  assign n50880 = ~n50877 & ~n50878 ;
  assign n50881 = ~n50879 & ~n50880 ;
  assign n50882 = ~n50582 & ~n50585 ;
  assign n50883 = n50881 & ~n50882 ;
  assign n50884 = ~n50881 & n50882 ;
  assign n50885 = ~n50883 & ~n50884 ;
  assign n51030 = n50885 & x234 ;
  assign n50886 = ~n50704 & ~n50710 ;
  assign n50887 = ~x126 & n13131 ;
  assign n50888 = ~x127 & n12501 ;
  assign n50889 = ~n50887 & ~n50888 ;
  assign n50890 = ~n12509 & n50889 ;
  assign n50891 = n27368 & n50889 ;
  assign n50892 = ~n50890 & ~n50891 ;
  assign n50893 = ~x44 & ~n50892 ;
  assign n50894 = x44 & n50892 ;
  assign n50895 = ~n50893 & ~n50894 ;
  assign n50896 = ~n50886 & ~n50895 ;
  assign n50897 = n50886 & n50895 ;
  assign n50898 = ~n50896 & ~n50897 ;
  assign n50899 = ~x125 & n14233 ;
  assign n50900 = ~x123 & n14876 ;
  assign n50901 = ~x124 & n14228 ;
  assign n50902 = ~n50900 & ~n50901 ;
  assign n50903 = ~n50899 & n50902 ;
  assign n50904 = n14236 & n25330 ;
  assign n50905 = n50903 & ~n50904 ;
  assign n50906 = ~x47 & ~n50905 ;
  assign n50907 = ~x47 & ~n50906 ;
  assign n50908 = ~n50905 & ~n50906 ;
  assign n50909 = ~n50907 & ~n50908 ;
  assign n50910 = ~n50688 & ~n50690 ;
  assign n50911 = ~n50682 & ~n50684 ;
  assign n50912 = ~n50634 & ~n50640 ;
  assign n50913 = ~x106 & n27427 ;
  assign n50914 = ~x107 & ~n26217 ;
  assign n50915 = ~n50913 & ~n50914 ;
  assign n50916 = x41 & ~n49965 ;
  assign n50917 = ~n50621 & ~n50916 ;
  assign n50918 = n50915 & ~n50917 ;
  assign n50919 = n50915 & ~n50918 ;
  assign n50920 = ~n50917 & ~n50918 ;
  assign n50921 = ~n50919 & ~n50920 ;
  assign n50922 = ~x110 & n24612 ;
  assign n50923 = ~x108 & n25390 ;
  assign n50924 = ~x109 & n24607 ;
  assign n50925 = ~n50923 & ~n50924 ;
  assign n50926 = ~n50922 & n50925 ;
  assign n50927 = ~n24615 & n50926 ;
  assign n50928 = ~n14802 & n50926 ;
  assign n50929 = ~n50927 & ~n50928 ;
  assign n50930 = ~x62 & ~n50929 ;
  assign n50931 = x62 & n50929 ;
  assign n50932 = ~n50930 & ~n50931 ;
  assign n50933 = ~n50921 & ~n50932 ;
  assign n50934 = n50921 & n50932 ;
  assign n50935 = ~n50933 & ~n50934 ;
  assign n50936 = ~n50912 & n50935 ;
  assign n50937 = n50912 & ~n50935 ;
  assign n50938 = ~n50936 & ~n50937 ;
  assign n50939 = ~x113 & n22325 ;
  assign n50940 = ~x111 & n23066 ;
  assign n50941 = ~x112 & n22320 ;
  assign n50942 = ~n50940 & ~n50941 ;
  assign n50943 = ~n50939 & n50942 ;
  assign n50944 = n16684 & n22328 ;
  assign n50945 = n50943 & ~n50944 ;
  assign n50946 = ~x59 & ~n50945 ;
  assign n50947 = ~x59 & ~n50946 ;
  assign n50948 = ~n50945 & ~n50946 ;
  assign n50949 = ~n50947 & ~n50948 ;
  assign n50950 = n50938 & ~n50949 ;
  assign n50951 = n50938 & ~n50950 ;
  assign n50952 = ~n50949 & ~n50950 ;
  assign n50953 = ~n50951 & ~n50952 ;
  assign n50954 = ~n50653 & ~n50659 ;
  assign n50955 = n50953 & n50954 ;
  assign n50956 = ~n50953 & ~n50954 ;
  assign n50957 = ~n50955 & ~n50956 ;
  assign n50958 = ~x116 & n20143 ;
  assign n50959 = ~x114 & n20854 ;
  assign n50960 = ~x115 & n20138 ;
  assign n50961 = ~n50959 & ~n50960 ;
  assign n50962 = ~n50958 & n50961 ;
  assign n50963 = n18678 & n20146 ;
  assign n50964 = n50962 & ~n50963 ;
  assign n50965 = ~x56 & ~n50964 ;
  assign n50966 = ~x56 & ~n50965 ;
  assign n50967 = ~n50964 & ~n50965 ;
  assign n50968 = ~n50966 & ~n50967 ;
  assign n50969 = n50957 & ~n50968 ;
  assign n50970 = n50957 & ~n50969 ;
  assign n50971 = ~n50968 & ~n50969 ;
  assign n50972 = ~n50970 & ~n50971 ;
  assign n50973 = ~n50662 & ~n50666 ;
  assign n50974 = n50972 & n50973 ;
  assign n50975 = ~n50972 & ~n50973 ;
  assign n50976 = ~n50974 & ~n50975 ;
  assign n50977 = ~x119 & n18025 ;
  assign n50978 = ~x117 & n18764 ;
  assign n50979 = ~x118 & n18020 ;
  assign n50980 = ~n50978 & ~n50979 ;
  assign n50981 = ~n50977 & n50980 ;
  assign n50982 = n18028 & n20778 ;
  assign n50983 = n50981 & ~n50982 ;
  assign n50984 = ~x53 & ~n50983 ;
  assign n50985 = ~x53 & ~n50984 ;
  assign n50986 = ~n50983 & ~n50984 ;
  assign n50987 = ~n50985 & ~n50986 ;
  assign n50988 = n50976 & ~n50987 ;
  assign n50989 = n50976 & ~n50988 ;
  assign n50990 = ~n50987 & ~n50988 ;
  assign n50991 = ~n50989 & ~n50990 ;
  assign n50992 = ~n50911 & n50991 ;
  assign n50993 = n50911 & ~n50991 ;
  assign n50994 = ~n50992 & ~n50993 ;
  assign n50995 = ~x122 & n16076 ;
  assign n50996 = ~x120 & n16756 ;
  assign n50997 = ~x121 & n16071 ;
  assign n50998 = ~n50996 & ~n50997 ;
  assign n50999 = ~n50995 & n50998 ;
  assign n51000 = n16079 & n22998 ;
  assign n51001 = n50999 & ~n51000 ;
  assign n51002 = ~x50 & ~n51001 ;
  assign n51003 = ~x50 & ~n51002 ;
  assign n51004 = ~n51001 & ~n51002 ;
  assign n51005 = ~n51003 & ~n51004 ;
  assign n51006 = n50994 & n51005 ;
  assign n51007 = ~n50994 & ~n51005 ;
  assign n51008 = ~n51006 & ~n51007 ;
  assign n51009 = ~n50910 & n51008 ;
  assign n51010 = ~n50910 & ~n51009 ;
  assign n51011 = n51008 & ~n51009 ;
  assign n51012 = ~n51010 & ~n51011 ;
  assign n51013 = ~n50909 & ~n51012 ;
  assign n51014 = ~n50909 & ~n51013 ;
  assign n51015 = ~n51012 & ~n51013 ;
  assign n51016 = ~n51014 & ~n51015 ;
  assign n51017 = n50898 & ~n51016 ;
  assign n51018 = n50898 & ~n51017 ;
  assign n51019 = ~n51016 & ~n51017 ;
  assign n51020 = ~n51018 & ~n51019 ;
  assign n51021 = ~n50723 & ~n50729 ;
  assign n51022 = n51020 & n51021 ;
  assign n51023 = ~n51020 & ~n51021 ;
  assign n51024 = ~n51022 & ~n51023 ;
  assign n51025 = ~n50733 & ~n50736 ;
  assign n51026 = n51024 & ~n51025 ;
  assign n51027 = ~n51024 & n51025 ;
  assign n51028 = ~n51026 & ~n51027 ;
  assign n51031 = ~n51028 & ~x234 ;
  assign n51032 = ~n51030 & ~n51031 ;
  assign n51033 = ~n50880 & ~n50883 ;
  assign n51034 = ~n50753 & ~n50874 ;
  assign n51035 = ~n50866 & ~n50870 ;
  assign n51036 = x127 & n13131 ;
  assign n51037 = n12509 & n26962 ;
  assign n51038 = ~n51036 & ~n51037 ;
  assign n51039 = x44 & ~n51038 ;
  assign n51040 = x44 & ~n51039 ;
  assign n51041 = ~n51038 & ~n51039 ;
  assign n51042 = ~n51040 & ~n51041 ;
  assign n51043 = ~n51035 & ~n51042 ;
  assign n51044 = ~n51035 & ~n51043 ;
  assign n51045 = ~n51042 & ~n51043 ;
  assign n51046 = ~n51044 & ~n51045 ;
  assign n51047 = ~n50832 & ~n50845 ;
  assign n51048 = x120 & n18025 ;
  assign n51049 = x118 & n18764 ;
  assign n51050 = x119 & n18020 ;
  assign n51051 = ~n51049 & ~n51050 ;
  assign n51052 = ~n51048 & n51051 ;
  assign n51053 = n18028 & n21143 ;
  assign n51054 = n51052 & ~n51053 ;
  assign n51055 = x53 & ~n51054 ;
  assign n51056 = x53 & ~n51055 ;
  assign n51057 = ~n51054 & ~n51055 ;
  assign n51058 = ~n51056 & ~n51057 ;
  assign n51059 = ~n50813 & ~n50826 ;
  assign n51060 = x117 & n20143 ;
  assign n51061 = x115 & n20854 ;
  assign n51062 = x116 & n20138 ;
  assign n51063 = ~n51061 & ~n51062 ;
  assign n51064 = ~n51060 & n51063 ;
  assign n51065 = n19026 & n20146 ;
  assign n51066 = n51064 & ~n51065 ;
  assign n51067 = x56 & ~n51066 ;
  assign n51068 = x56 & ~n51067 ;
  assign n51069 = ~n51066 & ~n51067 ;
  assign n51070 = ~n51068 & ~n51069 ;
  assign n51071 = ~n50793 & ~n50807 ;
  assign n51072 = x114 & n22325 ;
  assign n51073 = x112 & n23066 ;
  assign n51074 = x113 & n22320 ;
  assign n51075 = ~n51073 & ~n51074 ;
  assign n51076 = ~n51072 & n51075 ;
  assign n51077 = n17012 & n22328 ;
  assign n51078 = n51076 & ~n51077 ;
  assign n51079 = x59 & ~n51078 ;
  assign n51080 = x59 & ~n51079 ;
  assign n51081 = ~n51078 & ~n51079 ;
  assign n51082 = ~n51080 & ~n51081 ;
  assign n51083 = ~n50775 & ~n50790 ;
  assign n51084 = x107 & n27024 ;
  assign n51085 = x108 & ~n26217 ;
  assign n51086 = ~n51084 & ~n51085 ;
  assign n51087 = n50772 & ~n51086 ;
  assign n51088 = ~n50772 & n51086 ;
  assign n51089 = ~n51087 & ~n51088 ;
  assign n51090 = x111 & n24612 ;
  assign n51091 = x109 & n25390 ;
  assign n51092 = x110 & n24607 ;
  assign n51093 = ~n51091 & ~n51092 ;
  assign n51094 = ~n51090 & n51093 ;
  assign n51095 = ~n24615 & n51094 ;
  assign n51096 = ~n15111 & n51094 ;
  assign n51097 = ~n51095 & ~n51096 ;
  assign n51098 = x62 & ~n51097 ;
  assign n51099 = ~x62 & n51097 ;
  assign n51100 = ~n51098 & ~n51099 ;
  assign n51101 = n51089 & ~n51100 ;
  assign n51102 = ~n51089 & n51100 ;
  assign n51103 = ~n51101 & ~n51102 ;
  assign n51104 = ~n51083 & n51103 ;
  assign n51105 = ~n51083 & ~n51104 ;
  assign n51106 = n51103 & ~n51104 ;
  assign n51107 = ~n51105 & ~n51106 ;
  assign n51108 = ~n51082 & ~n51107 ;
  assign n51109 = n51082 & ~n51106 ;
  assign n51110 = ~n51105 & n51109 ;
  assign n51111 = ~n51108 & ~n51110 ;
  assign n51112 = ~n51071 & n51111 ;
  assign n51113 = ~n51071 & ~n51112 ;
  assign n51114 = n51111 & ~n51112 ;
  assign n51115 = ~n51113 & ~n51114 ;
  assign n51116 = ~n51070 & ~n51115 ;
  assign n51117 = n51070 & ~n51114 ;
  assign n51118 = ~n51113 & n51117 ;
  assign n51119 = ~n51116 & ~n51118 ;
  assign n51120 = ~n51059 & n51119 ;
  assign n51121 = ~n51059 & ~n51120 ;
  assign n51122 = n51119 & ~n51120 ;
  assign n51123 = ~n51121 & ~n51122 ;
  assign n51124 = ~n51058 & ~n51123 ;
  assign n51125 = n51058 & ~n51122 ;
  assign n51126 = ~n51121 & n51125 ;
  assign n51127 = ~n51124 & ~n51126 ;
  assign n51128 = ~n51047 & n51127 ;
  assign n51129 = n51047 & ~n51127 ;
  assign n51130 = ~n51128 & ~n51129 ;
  assign n51131 = x123 & n16076 ;
  assign n51132 = x121 & n16756 ;
  assign n51133 = x122 & n16071 ;
  assign n51134 = ~n51132 & ~n51133 ;
  assign n51135 = ~n51131 & n51134 ;
  assign n51136 = n16079 & n23382 ;
  assign n51137 = n51135 & ~n51136 ;
  assign n51138 = x50 & ~n51137 ;
  assign n51139 = x50 & ~n51138 ;
  assign n51140 = ~n51137 & ~n51138 ;
  assign n51141 = ~n51139 & ~n51140 ;
  assign n51142 = n51130 & ~n51141 ;
  assign n51143 = n51130 & ~n51142 ;
  assign n51144 = ~n51141 & ~n51142 ;
  assign n51145 = ~n51143 & ~n51144 ;
  assign n51146 = ~n50768 & ~n50848 ;
  assign n51147 = ~n50864 & ~n51146 ;
  assign n51148 = ~n51145 & ~n51147 ;
  assign n51149 = ~n51145 & ~n51148 ;
  assign n51150 = ~n51147 & ~n51148 ;
  assign n51151 = ~n51149 & ~n51150 ;
  assign n51152 = x126 & n14233 ;
  assign n51153 = x124 & n14876 ;
  assign n51154 = x125 & n14228 ;
  assign n51155 = ~n51153 & ~n51154 ;
  assign n51156 = ~n51152 & n51155 ;
  assign n51157 = n14236 & n25735 ;
  assign n51158 = n51156 & ~n51157 ;
  assign n51159 = x47 & ~n51158 ;
  assign n51160 = x47 & ~n51159 ;
  assign n51161 = ~n51158 & ~n51159 ;
  assign n51162 = ~n51160 & ~n51161 ;
  assign n51163 = ~n51151 & ~n51162 ;
  assign n51164 = ~n51151 & ~n51163 ;
  assign n51165 = ~n51162 & ~n51163 ;
  assign n51166 = ~n51164 & ~n51165 ;
  assign n51167 = ~n51046 & n51166 ;
  assign n51168 = n51046 & ~n51166 ;
  assign n51169 = ~n51167 & ~n51168 ;
  assign n51170 = ~n51034 & ~n51169 ;
  assign n51171 = n51034 & n51169 ;
  assign n51172 = ~n51170 & ~n51171 ;
  assign n51173 = ~n51033 & n51172 ;
  assign n51174 = n51033 & ~n51172 ;
  assign n51175 = ~n51173 & ~n51174 ;
  assign n51320 = n51175 & x235 ;
  assign n51176 = ~n51023 & ~n51026 ;
  assign n51177 = ~n50896 & ~n51017 ;
  assign n51178 = ~n51009 & ~n51013 ;
  assign n51179 = ~x127 & n13131 ;
  assign n51180 = n12509 & n27365 ;
  assign n51181 = ~n51179 & ~n51180 ;
  assign n51182 = ~x44 & ~n51181 ;
  assign n51183 = ~x44 & ~n51182 ;
  assign n51184 = ~n51181 & ~n51182 ;
  assign n51185 = ~n51183 & ~n51184 ;
  assign n51186 = ~n51178 & ~n51185 ;
  assign n51187 = ~n51178 & ~n51186 ;
  assign n51188 = ~n51185 & ~n51186 ;
  assign n51189 = ~n51187 & ~n51188 ;
  assign n51190 = ~n50975 & ~n50988 ;
  assign n51191 = ~x120 & n18025 ;
  assign n51192 = ~x118 & n18764 ;
  assign n51193 = ~x119 & n18020 ;
  assign n51194 = ~n51192 & ~n51193 ;
  assign n51195 = ~n51191 & n51194 ;
  assign n51196 = n18028 & n21501 ;
  assign n51197 = n51195 & ~n51196 ;
  assign n51198 = ~x53 & ~n51197 ;
  assign n51199 = ~x53 & ~n51198 ;
  assign n51200 = ~n51197 & ~n51198 ;
  assign n51201 = ~n51199 & ~n51200 ;
  assign n51202 = ~n50956 & ~n50969 ;
  assign n51203 = ~x117 & n20143 ;
  assign n51204 = ~x115 & n20854 ;
  assign n51205 = ~x116 & n20138 ;
  assign n51206 = ~n51204 & ~n51205 ;
  assign n51207 = ~n51203 & n51206 ;
  assign n51208 = n19365 & n20146 ;
  assign n51209 = n51207 & ~n51208 ;
  assign n51210 = ~x56 & ~n51209 ;
  assign n51211 = ~x56 & ~n51210 ;
  assign n51212 = ~n51209 & ~n51210 ;
  assign n51213 = ~n51211 & ~n51212 ;
  assign n51214 = ~n50936 & ~n50950 ;
  assign n51215 = ~x114 & n22325 ;
  assign n51216 = ~x112 & n23066 ;
  assign n51217 = ~x113 & n22320 ;
  assign n51218 = ~n51216 & ~n51217 ;
  assign n51219 = ~n51215 & n51218 ;
  assign n51220 = n17333 & n22328 ;
  assign n51221 = n51219 & ~n51220 ;
  assign n51222 = ~x59 & ~n51221 ;
  assign n51223 = ~x59 & ~n51222 ;
  assign n51224 = ~n51221 & ~n51222 ;
  assign n51225 = ~n51223 & ~n51224 ;
  assign n51226 = ~n50918 & ~n50933 ;
  assign n51227 = ~x107 & n27427 ;
  assign n51228 = ~x108 & ~n26217 ;
  assign n51229 = ~n51227 & ~n51228 ;
  assign n51230 = n50915 & ~n51229 ;
  assign n51231 = ~n50915 & n51229 ;
  assign n51232 = ~n51230 & ~n51231 ;
  assign n51233 = ~x111 & n24612 ;
  assign n51234 = ~x109 & n25390 ;
  assign n51235 = ~x110 & n24607 ;
  assign n51236 = ~n51234 & ~n51235 ;
  assign n51237 = ~n51233 & n51236 ;
  assign n51238 = ~n24615 & n51237 ;
  assign n51239 = ~n15411 & n51237 ;
  assign n51240 = ~n51238 & ~n51239 ;
  assign n51241 = ~x62 & ~n51240 ;
  assign n51242 = x62 & n51240 ;
  assign n51243 = ~n51241 & ~n51242 ;
  assign n51244 = n51232 & ~n51243 ;
  assign n51245 = ~n51232 & n51243 ;
  assign n51246 = ~n51244 & ~n51245 ;
  assign n51247 = ~n51226 & n51246 ;
  assign n51248 = ~n51226 & ~n51247 ;
  assign n51249 = n51246 & ~n51247 ;
  assign n51250 = ~n51248 & ~n51249 ;
  assign n51251 = ~n51225 & ~n51250 ;
  assign n51252 = n51225 & ~n51249 ;
  assign n51253 = ~n51248 & n51252 ;
  assign n51254 = ~n51251 & ~n51253 ;
  assign n51255 = ~n51214 & n51254 ;
  assign n51256 = ~n51214 & ~n51255 ;
  assign n51257 = n51254 & ~n51255 ;
  assign n51258 = ~n51256 & ~n51257 ;
  assign n51259 = ~n51213 & ~n51258 ;
  assign n51260 = n51213 & ~n51257 ;
  assign n51261 = ~n51256 & n51260 ;
  assign n51262 = ~n51259 & ~n51261 ;
  assign n51263 = ~n51202 & n51262 ;
  assign n51264 = ~n51202 & ~n51263 ;
  assign n51265 = n51262 & ~n51263 ;
  assign n51266 = ~n51264 & ~n51265 ;
  assign n51267 = ~n51201 & ~n51266 ;
  assign n51268 = n51201 & ~n51265 ;
  assign n51269 = ~n51264 & n51268 ;
  assign n51270 = ~n51267 & ~n51269 ;
  assign n51271 = ~n51190 & n51270 ;
  assign n51272 = n51190 & ~n51270 ;
  assign n51273 = ~n51271 & ~n51272 ;
  assign n51274 = ~x123 & n16076 ;
  assign n51275 = ~x121 & n16756 ;
  assign n51276 = ~x122 & n16071 ;
  assign n51277 = ~n51275 & ~n51276 ;
  assign n51278 = ~n51274 & n51277 ;
  assign n51279 = n16079 & n23760 ;
  assign n51280 = n51278 & ~n51279 ;
  assign n51281 = ~x50 & ~n51280 ;
  assign n51282 = ~x50 & ~n51281 ;
  assign n51283 = ~n51280 & ~n51281 ;
  assign n51284 = ~n51282 & ~n51283 ;
  assign n51285 = n51273 & ~n51284 ;
  assign n51286 = n51273 & ~n51285 ;
  assign n51287 = ~n51284 & ~n51285 ;
  assign n51288 = ~n51286 & ~n51287 ;
  assign n51289 = ~n50911 & ~n50991 ;
  assign n51290 = ~n51007 & ~n51289 ;
  assign n51291 = ~n51288 & ~n51290 ;
  assign n51292 = ~n51288 & ~n51291 ;
  assign n51293 = ~n51290 & ~n51291 ;
  assign n51294 = ~n51292 & ~n51293 ;
  assign n51295 = ~x126 & n14233 ;
  assign n51296 = ~x124 & n14876 ;
  assign n51297 = ~x125 & n14228 ;
  assign n51298 = ~n51296 & ~n51297 ;
  assign n51299 = ~n51295 & n51298 ;
  assign n51300 = n14236 & n26128 ;
  assign n51301 = n51299 & ~n51300 ;
  assign n51302 = ~x47 & ~n51301 ;
  assign n51303 = ~x47 & ~n51302 ;
  assign n51304 = ~n51301 & ~n51302 ;
  assign n51305 = ~n51303 & ~n51304 ;
  assign n51306 = ~n51294 & ~n51305 ;
  assign n51307 = ~n51294 & ~n51306 ;
  assign n51308 = ~n51305 & ~n51306 ;
  assign n51309 = ~n51307 & ~n51308 ;
  assign n51310 = ~n51189 & n51309 ;
  assign n51311 = n51189 & ~n51309 ;
  assign n51312 = ~n51310 & ~n51311 ;
  assign n51313 = ~n51177 & ~n51312 ;
  assign n51314 = n51177 & n51312 ;
  assign n51315 = ~n51313 & ~n51314 ;
  assign n51316 = ~n51176 & n51315 ;
  assign n51317 = n51176 & ~n51315 ;
  assign n51318 = ~n51316 & ~n51317 ;
  assign n51321 = ~n51318 & ~x235 ;
  assign n51322 = ~n51320 & ~n51321 ;
  assign n51323 = ~n51170 & ~n51173 ;
  assign n51324 = ~n51128 & ~n51142 ;
  assign n51325 = x124 & n16076 ;
  assign n51326 = x122 & n16756 ;
  assign n51327 = x123 & n16071 ;
  assign n51328 = ~n51326 & ~n51327 ;
  assign n51329 = ~n51325 & n51328 ;
  assign n51330 = n16079 & n23796 ;
  assign n51331 = n51329 & ~n51330 ;
  assign n51332 = x50 & ~n51331 ;
  assign n51333 = x50 & ~n51332 ;
  assign n51334 = ~n51331 & ~n51332 ;
  assign n51335 = ~n51333 & ~n51334 ;
  assign n51336 = ~n51120 & ~n51124 ;
  assign n51337 = x121 & n18025 ;
  assign n51338 = x119 & n18764 ;
  assign n51339 = x120 & n18020 ;
  assign n51340 = ~n51338 & ~n51339 ;
  assign n51341 = ~n51337 & n51340 ;
  assign n51342 = n18028 & n21870 ;
  assign n51343 = n51341 & ~n51342 ;
  assign n51344 = x53 & ~n51343 ;
  assign n51345 = x53 & ~n51344 ;
  assign n51346 = ~n51343 & ~n51344 ;
  assign n51347 = ~n51345 & ~n51346 ;
  assign n51348 = ~n51112 & ~n51116 ;
  assign n51349 = x118 & n20143 ;
  assign n51350 = x116 & n20854 ;
  assign n51351 = x117 & n20138 ;
  assign n51352 = ~n51350 & ~n51351 ;
  assign n51353 = ~n51349 & n51352 ;
  assign n51354 = n19395 & n20146 ;
  assign n51355 = n51353 & ~n51354 ;
  assign n51356 = x56 & ~n51355 ;
  assign n51357 = x56 & ~n51356 ;
  assign n51358 = ~n51355 & ~n51356 ;
  assign n51359 = ~n51357 & ~n51358 ;
  assign n51360 = ~n51104 & ~n51108 ;
  assign n51361 = ~n51087 & ~n51101 ;
  assign n51362 = x108 & n27024 ;
  assign n51363 = x109 & ~n26217 ;
  assign n51364 = ~n51362 & ~n51363 ;
  assign n51365 = ~x44 & ~n51364 ;
  assign n51366 = x44 & n51364 ;
  assign n51367 = ~n51365 & ~n51366 ;
  assign n51368 = ~n50772 & n51367 ;
  assign n51369 = ~n50772 & ~n51368 ;
  assign n51370 = n51367 & ~n51368 ;
  assign n51371 = ~n51369 & ~n51370 ;
  assign n51372 = ~n51361 & ~n51371 ;
  assign n51373 = ~n51361 & ~n51372 ;
  assign n51374 = ~n51371 & ~n51372 ;
  assign n51375 = ~n51373 & ~n51374 ;
  assign n51376 = x112 & n24612 ;
  assign n51377 = x110 & n25390 ;
  assign n51378 = x111 & n24607 ;
  assign n51379 = ~n51377 & ~n51378 ;
  assign n51380 = ~n51376 & n51379 ;
  assign n51381 = n15442 & n24615 ;
  assign n51382 = n51380 & ~n51381 ;
  assign n51383 = x62 & ~n51382 ;
  assign n51384 = x62 & ~n51383 ;
  assign n51385 = ~n51382 & ~n51383 ;
  assign n51386 = ~n51384 & ~n51385 ;
  assign n51387 = ~n51375 & ~n51386 ;
  assign n51388 = ~n51375 & ~n51387 ;
  assign n51389 = ~n51386 & ~n51387 ;
  assign n51390 = ~n51388 & ~n51389 ;
  assign n51391 = x115 & n22325 ;
  assign n51392 = x113 & n23066 ;
  assign n51393 = x114 & n22320 ;
  assign n51394 = ~n51392 & ~n51393 ;
  assign n51395 = ~n51391 & n51394 ;
  assign n51396 = n17364 & n22328 ;
  assign n51397 = n51395 & ~n51396 ;
  assign n51398 = x59 & ~n51397 ;
  assign n51399 = x59 & ~n51398 ;
  assign n51400 = ~n51397 & ~n51398 ;
  assign n51401 = ~n51399 & ~n51400 ;
  assign n51402 = n51390 & n51401 ;
  assign n51403 = ~n51390 & ~n51401 ;
  assign n51404 = ~n51402 & ~n51403 ;
  assign n51405 = ~n51360 & n51404 ;
  assign n51406 = n51360 & ~n51404 ;
  assign n51407 = ~n51405 & ~n51406 ;
  assign n51408 = n51359 & ~n51407 ;
  assign n51409 = ~n51359 & n51407 ;
  assign n51410 = ~n51408 & ~n51409 ;
  assign n51411 = ~n51348 & n51410 ;
  assign n51412 = n51348 & ~n51410 ;
  assign n51413 = ~n51411 & ~n51412 ;
  assign n51414 = n51347 & ~n51413 ;
  assign n51415 = ~n51347 & n51413 ;
  assign n51416 = ~n51414 & ~n51415 ;
  assign n51417 = ~n51336 & n51416 ;
  assign n51418 = n51336 & ~n51416 ;
  assign n51419 = ~n51417 & ~n51418 ;
  assign n51420 = n51335 & ~n51419 ;
  assign n51421 = ~n51335 & n51419 ;
  assign n51422 = ~n51420 & ~n51421 ;
  assign n51423 = ~n51324 & n51422 ;
  assign n51424 = n51324 & ~n51422 ;
  assign n51425 = ~n51423 & ~n51424 ;
  assign n51426 = x127 & n14233 ;
  assign n51427 = x125 & n14876 ;
  assign n51428 = x126 & n14228 ;
  assign n51429 = ~n51427 & ~n51428 ;
  assign n51430 = ~n51426 & n51429 ;
  assign n51431 = n14236 & n26533 ;
  assign n51432 = n51430 & ~n51431 ;
  assign n51433 = x47 & ~n51432 ;
  assign n51434 = x47 & ~n51433 ;
  assign n51435 = ~n51432 & ~n51433 ;
  assign n51436 = ~n51434 & ~n51435 ;
  assign n51437 = n51425 & ~n51436 ;
  assign n51438 = n51425 & ~n51437 ;
  assign n51439 = ~n51436 & ~n51437 ;
  assign n51440 = ~n51438 & ~n51439 ;
  assign n51441 = ~n51148 & ~n51163 ;
  assign n51442 = n51440 & n51441 ;
  assign n51443 = ~n51440 & ~n51441 ;
  assign n51444 = ~n51442 & ~n51443 ;
  assign n51445 = ~n51046 & ~n51166 ;
  assign n51446 = ~n51043 & ~n51445 ;
  assign n51447 = n51444 & ~n51446 ;
  assign n51448 = ~n51444 & n51446 ;
  assign n51449 = ~n51447 & ~n51448 ;
  assign n51450 = ~n51323 & n51449 ;
  assign n51451 = n51323 & ~n51449 ;
  assign n51452 = ~n51450 & ~n51451 ;
  assign n51584 = n51452 & x236 ;
  assign n51453 = ~n51313 & ~n51316 ;
  assign n51454 = ~n51271 & ~n51285 ;
  assign n51455 = ~x124 & n16076 ;
  assign n51456 = ~x122 & n16756 ;
  assign n51457 = ~x123 & n16071 ;
  assign n51458 = ~n51456 & ~n51457 ;
  assign n51459 = ~n51455 & n51458 ;
  assign n51460 = n16079 & n24176 ;
  assign n51461 = n51459 & ~n51460 ;
  assign n51462 = ~x50 & ~n51461 ;
  assign n51463 = ~x50 & ~n51462 ;
  assign n51464 = ~n51461 & ~n51462 ;
  assign n51465 = ~n51463 & ~n51464 ;
  assign n51466 = ~n51263 & ~n51267 ;
  assign n51467 = ~x121 & n18025 ;
  assign n51468 = ~x119 & n18764 ;
  assign n51469 = ~x120 & n18020 ;
  assign n51470 = ~n51468 & ~n51469 ;
  assign n51471 = ~n51467 & n51470 ;
  assign n51472 = n18028 & n22229 ;
  assign n51473 = n51471 & ~n51472 ;
  assign n51474 = ~x53 & ~n51473 ;
  assign n51475 = ~x53 & ~n51474 ;
  assign n51476 = ~n51473 & ~n51474 ;
  assign n51477 = ~n51475 & ~n51476 ;
  assign n51478 = ~n51255 & ~n51259 ;
  assign n51479 = ~x118 & n20143 ;
  assign n51480 = ~x116 & n20854 ;
  assign n51481 = ~x117 & n20138 ;
  assign n51482 = ~n51480 & ~n51481 ;
  assign n51483 = ~n51479 & n51482 ;
  assign n51484 = n19736 & n20146 ;
  assign n51485 = n51483 & ~n51484 ;
  assign n51486 = ~x56 & ~n51485 ;
  assign n51487 = ~x56 & ~n51486 ;
  assign n51488 = ~n51485 & ~n51486 ;
  assign n51489 = ~n51487 & ~n51488 ;
  assign n51490 = ~n51247 & ~n51251 ;
  assign n51491 = ~n51230 & ~n51244 ;
  assign n51492 = ~x108 & n27427 ;
  assign n51493 = ~x109 & ~n26217 ;
  assign n51494 = ~n51492 & ~n51493 ;
  assign n51495 = x44 & ~n51494 ;
  assign n51496 = ~x44 & n51494 ;
  assign n51497 = ~n51495 & ~n51496 ;
  assign n51498 = ~n50915 & n51497 ;
  assign n51499 = ~n50915 & ~n51498 ;
  assign n51500 = n51497 & ~n51498 ;
  assign n51501 = ~n51499 & ~n51500 ;
  assign n51502 = ~n51491 & ~n51501 ;
  assign n51503 = ~n51491 & ~n51502 ;
  assign n51504 = ~n51501 & ~n51502 ;
  assign n51505 = ~n51503 & ~n51504 ;
  assign n51506 = ~x112 & n24612 ;
  assign n51507 = ~x110 & n25390 ;
  assign n51508 = ~x111 & n24607 ;
  assign n51509 = ~n51507 & ~n51508 ;
  assign n51510 = ~n51506 & n51509 ;
  assign n51511 = n15744 & n24615 ;
  assign n51512 = n51510 & ~n51511 ;
  assign n51513 = ~x62 & ~n51512 ;
  assign n51514 = ~x62 & ~n51513 ;
  assign n51515 = ~n51512 & ~n51513 ;
  assign n51516 = ~n51514 & ~n51515 ;
  assign n51517 = ~n51505 & ~n51516 ;
  assign n51518 = ~n51505 & ~n51517 ;
  assign n51519 = ~n51516 & ~n51517 ;
  assign n51520 = ~n51518 & ~n51519 ;
  assign n51521 = ~x115 & n22325 ;
  assign n51522 = ~x113 & n23066 ;
  assign n51523 = ~x114 & n22320 ;
  assign n51524 = ~n51522 & ~n51523 ;
  assign n51525 = ~n51521 & n51524 ;
  assign n51526 = n17683 & n22328 ;
  assign n51527 = n51525 & ~n51526 ;
  assign n51528 = ~x59 & ~n51527 ;
  assign n51529 = ~x59 & ~n51528 ;
  assign n51530 = ~n51527 & ~n51528 ;
  assign n51531 = ~n51529 & ~n51530 ;
  assign n51532 = n51520 & n51531 ;
  assign n51533 = ~n51520 & ~n51531 ;
  assign n51534 = ~n51532 & ~n51533 ;
  assign n51535 = ~n51490 & n51534 ;
  assign n51536 = n51490 & ~n51534 ;
  assign n51537 = ~n51535 & ~n51536 ;
  assign n51538 = n51489 & ~n51537 ;
  assign n51539 = ~n51489 & n51537 ;
  assign n51540 = ~n51538 & ~n51539 ;
  assign n51541 = ~n51478 & n51540 ;
  assign n51542 = n51478 & ~n51540 ;
  assign n51543 = ~n51541 & ~n51542 ;
  assign n51544 = n51477 & ~n51543 ;
  assign n51545 = ~n51477 & n51543 ;
  assign n51546 = ~n51544 & ~n51545 ;
  assign n51547 = ~n51466 & n51546 ;
  assign n51548 = n51466 & ~n51546 ;
  assign n51549 = ~n51547 & ~n51548 ;
  assign n51550 = n51465 & ~n51549 ;
  assign n51551 = ~n51465 & n51549 ;
  assign n51552 = ~n51550 & ~n51551 ;
  assign n51553 = ~n51454 & n51552 ;
  assign n51554 = n51454 & ~n51552 ;
  assign n51555 = ~n51553 & ~n51554 ;
  assign n51556 = ~x127 & n14233 ;
  assign n51557 = ~x125 & n14876 ;
  assign n51558 = ~x126 & n14228 ;
  assign n51559 = ~n51557 & ~n51558 ;
  assign n51560 = ~n51556 & n51559 ;
  assign n51561 = n14236 & n26932 ;
  assign n51562 = n51560 & ~n51561 ;
  assign n51563 = ~x47 & ~n51562 ;
  assign n51564 = ~x47 & ~n51563 ;
  assign n51565 = ~n51562 & ~n51563 ;
  assign n51566 = ~n51564 & ~n51565 ;
  assign n51567 = n51555 & ~n51566 ;
  assign n51568 = n51555 & ~n51567 ;
  assign n51569 = ~n51566 & ~n51567 ;
  assign n51570 = ~n51568 & ~n51569 ;
  assign n51571 = ~n51291 & ~n51306 ;
  assign n51572 = n51570 & n51571 ;
  assign n51573 = ~n51570 & ~n51571 ;
  assign n51574 = ~n51572 & ~n51573 ;
  assign n51575 = ~n51189 & ~n51309 ;
  assign n51576 = ~n51186 & ~n51575 ;
  assign n51577 = n51574 & ~n51576 ;
  assign n51578 = ~n51574 & n51576 ;
  assign n51579 = ~n51577 & ~n51578 ;
  assign n51580 = ~n51453 & n51579 ;
  assign n51581 = n51453 & ~n51579 ;
  assign n51582 = ~n51580 & ~n51581 ;
  assign n51585 = ~n51582 & ~x236 ;
  assign n51586 = ~n51584 & ~n51585 ;
  assign n51587 = ~n51421 & ~n51423 ;
  assign n51588 = x126 & n14876 ;
  assign n51589 = x127 & n14228 ;
  assign n51590 = ~n51588 & ~n51589 ;
  assign n51591 = ~n14236 & n51590 ;
  assign n51592 = n26965 & n51590 ;
  assign n51593 = ~n51591 & ~n51592 ;
  assign n51594 = x47 & ~n51593 ;
  assign n51595 = ~x47 & n51593 ;
  assign n51596 = ~n51594 & ~n51595 ;
  assign n51597 = ~n51587 & ~n51596 ;
  assign n51598 = n51587 & n51596 ;
  assign n51599 = ~n51597 & ~n51598 ;
  assign n51600 = x125 & n16076 ;
  assign n51601 = x123 & n16756 ;
  assign n51602 = x124 & n16071 ;
  assign n51603 = ~n51601 & ~n51602 ;
  assign n51604 = ~n51600 & n51603 ;
  assign n51605 = n16079 & n24935 ;
  assign n51606 = n51604 & ~n51605 ;
  assign n51607 = x50 & ~n51606 ;
  assign n51608 = x50 & ~n51607 ;
  assign n51609 = ~n51606 & ~n51607 ;
  assign n51610 = ~n51608 & ~n51609 ;
  assign n51611 = ~n51415 & ~n51417 ;
  assign n51612 = ~n51409 & ~n51411 ;
  assign n51613 = ~n51403 & ~n51405 ;
  assign n51614 = x116 & n22325 ;
  assign n51615 = x114 & n23066 ;
  assign n51616 = x115 & n22320 ;
  assign n51617 = ~n51615 & ~n51616 ;
  assign n51618 = ~n51614 & n51617 ;
  assign n51619 = n18336 & n22328 ;
  assign n51620 = n51618 & ~n51619 ;
  assign n51621 = x59 & ~n51620 ;
  assign n51622 = x59 & ~n51621 ;
  assign n51623 = ~n51620 & ~n51621 ;
  assign n51624 = ~n51622 & ~n51623 ;
  assign n51625 = ~n51372 & ~n51387 ;
  assign n51626 = x109 & n27024 ;
  assign n51627 = x110 & ~n26217 ;
  assign n51628 = ~n51626 & ~n51627 ;
  assign n51629 = ~n51365 & ~n51368 ;
  assign n51630 = ~n51628 & n51629 ;
  assign n51631 = n51628 & ~n51629 ;
  assign n51632 = ~n51630 & ~n51631 ;
  assign n51633 = x113 & n24612 ;
  assign n51634 = x111 & n25390 ;
  assign n51635 = x112 & n24607 ;
  assign n51636 = ~n51634 & ~n51635 ;
  assign n51637 = ~n51633 & n51636 ;
  assign n51638 = n16361 & n24615 ;
  assign n51639 = n51637 & ~n51638 ;
  assign n51640 = x62 & ~n51639 ;
  assign n51641 = x62 & ~n51640 ;
  assign n51642 = ~n51639 & ~n51640 ;
  assign n51643 = ~n51641 & ~n51642 ;
  assign n51644 = ~n51632 & n51643 ;
  assign n51645 = n51632 & ~n51643 ;
  assign n51646 = ~n51644 & ~n51645 ;
  assign n51647 = ~n51625 & n51646 ;
  assign n51648 = ~n51625 & ~n51647 ;
  assign n51649 = n51646 & ~n51647 ;
  assign n51650 = ~n51648 & ~n51649 ;
  assign n51651 = ~n51624 & ~n51650 ;
  assign n51652 = n51624 & ~n51649 ;
  assign n51653 = ~n51648 & n51652 ;
  assign n51654 = ~n51651 & ~n51653 ;
  assign n51655 = ~n51613 & n51654 ;
  assign n51656 = n51613 & ~n51654 ;
  assign n51657 = ~n51655 & ~n51656 ;
  assign n51658 = x119 & n20143 ;
  assign n51659 = x117 & n20854 ;
  assign n51660 = x118 & n20138 ;
  assign n51661 = ~n51659 & ~n51660 ;
  assign n51662 = ~n51658 & n51661 ;
  assign n51663 = n20146 & n20423 ;
  assign n51664 = n51662 & ~n51663 ;
  assign n51665 = x56 & ~n51664 ;
  assign n51666 = x56 & ~n51665 ;
  assign n51667 = ~n51664 & ~n51665 ;
  assign n51668 = ~n51666 & ~n51667 ;
  assign n51669 = n51657 & ~n51668 ;
  assign n51670 = n51657 & ~n51669 ;
  assign n51671 = ~n51668 & ~n51669 ;
  assign n51672 = ~n51670 & ~n51671 ;
  assign n51673 = ~n51612 & n51672 ;
  assign n51674 = n51612 & ~n51672 ;
  assign n51675 = ~n51673 & ~n51674 ;
  assign n51676 = x122 & n18025 ;
  assign n51677 = x120 & n18764 ;
  assign n51678 = x121 & n18020 ;
  assign n51679 = ~n51677 & ~n51678 ;
  assign n51680 = ~n51676 & n51679 ;
  assign n51681 = n18028 & n22622 ;
  assign n51682 = n51680 & ~n51681 ;
  assign n51683 = x53 & ~n51682 ;
  assign n51684 = x53 & ~n51683 ;
  assign n51685 = ~n51682 & ~n51683 ;
  assign n51686 = ~n51684 & ~n51685 ;
  assign n51687 = n51675 & n51686 ;
  assign n51688 = ~n51675 & ~n51686 ;
  assign n51689 = ~n51687 & ~n51688 ;
  assign n51690 = ~n51611 & n51689 ;
  assign n51691 = ~n51611 & ~n51690 ;
  assign n51692 = n51689 & ~n51690 ;
  assign n51693 = ~n51691 & ~n51692 ;
  assign n51694 = ~n51610 & ~n51693 ;
  assign n51695 = ~n51610 & ~n51694 ;
  assign n51696 = ~n51693 & ~n51694 ;
  assign n51697 = ~n51695 & ~n51696 ;
  assign n51698 = n51599 & ~n51697 ;
  assign n51699 = n51599 & ~n51698 ;
  assign n51700 = ~n51697 & ~n51698 ;
  assign n51701 = ~n51699 & ~n51700 ;
  assign n51702 = ~n51437 & ~n51443 ;
  assign n51703 = n51701 & n51702 ;
  assign n51704 = ~n51701 & ~n51702 ;
  assign n51705 = ~n51703 & ~n51704 ;
  assign n51706 = ~n51447 & ~n51450 ;
  assign n51707 = n51705 & ~n51706 ;
  assign n51708 = ~n51705 & n51706 ;
  assign n51709 = ~n51707 & ~n51708 ;
  assign n51834 = n51709 & x237 ;
  assign n51710 = ~n51551 & ~n51553 ;
  assign n51711 = ~x126 & n14876 ;
  assign n51712 = ~x127 & n14228 ;
  assign n51713 = ~n51711 & ~n51712 ;
  assign n51714 = ~n14236 & n51713 ;
  assign n51715 = n27368 & n51713 ;
  assign n51716 = ~n51714 & ~n51715 ;
  assign n51717 = ~x47 & ~n51716 ;
  assign n51718 = x47 & n51716 ;
  assign n51719 = ~n51717 & ~n51718 ;
  assign n51720 = ~n51710 & ~n51719 ;
  assign n51721 = n51710 & n51719 ;
  assign n51722 = ~n51720 & ~n51721 ;
  assign n51723 = ~x125 & n16076 ;
  assign n51724 = ~x123 & n16756 ;
  assign n51725 = ~x124 & n16071 ;
  assign n51726 = ~n51724 & ~n51725 ;
  assign n51727 = ~n51723 & n51726 ;
  assign n51728 = n16079 & n25330 ;
  assign n51729 = n51727 & ~n51728 ;
  assign n51730 = ~x50 & ~n51729 ;
  assign n51731 = ~x50 & ~n51730 ;
  assign n51732 = ~n51729 & ~n51730 ;
  assign n51733 = ~n51731 & ~n51732 ;
  assign n51734 = ~n51545 & ~n51547 ;
  assign n51735 = ~n51539 & ~n51541 ;
  assign n51736 = ~n51533 & ~n51535 ;
  assign n51737 = ~x116 & n22325 ;
  assign n51738 = ~x114 & n23066 ;
  assign n51739 = ~x115 & n22320 ;
  assign n51740 = ~n51738 & ~n51739 ;
  assign n51741 = ~n51737 & n51740 ;
  assign n51742 = n18678 & n22328 ;
  assign n51743 = n51741 & ~n51742 ;
  assign n51744 = ~x59 & ~n51743 ;
  assign n51745 = ~x59 & ~n51744 ;
  assign n51746 = ~n51743 & ~n51744 ;
  assign n51747 = ~n51745 & ~n51746 ;
  assign n51748 = ~n51502 & ~n51517 ;
  assign n51749 = ~x109 & n27427 ;
  assign n51750 = ~x110 & ~n26217 ;
  assign n51751 = ~n51749 & ~n51750 ;
  assign n51752 = ~n51495 & ~n51498 ;
  assign n51753 = ~n51751 & n51752 ;
  assign n51754 = n51751 & ~n51752 ;
  assign n51755 = ~n51753 & ~n51754 ;
  assign n51756 = ~x113 & n24612 ;
  assign n51757 = ~x111 & n25390 ;
  assign n51758 = ~x112 & n24607 ;
  assign n51759 = ~n51757 & ~n51758 ;
  assign n51760 = ~n51756 & n51759 ;
  assign n51761 = n16684 & n24615 ;
  assign n51762 = n51760 & ~n51761 ;
  assign n51763 = ~x62 & ~n51762 ;
  assign n51764 = ~x62 & ~n51763 ;
  assign n51765 = ~n51762 & ~n51763 ;
  assign n51766 = ~n51764 & ~n51765 ;
  assign n51767 = ~n51755 & n51766 ;
  assign n51768 = n51755 & ~n51766 ;
  assign n51769 = ~n51767 & ~n51768 ;
  assign n51770 = ~n51748 & n51769 ;
  assign n51771 = ~n51748 & ~n51770 ;
  assign n51772 = n51769 & ~n51770 ;
  assign n51773 = ~n51771 & ~n51772 ;
  assign n51774 = ~n51747 & ~n51773 ;
  assign n51775 = n51747 & ~n51772 ;
  assign n51776 = ~n51771 & n51775 ;
  assign n51777 = ~n51774 & ~n51776 ;
  assign n51778 = ~n51736 & n51777 ;
  assign n51779 = n51736 & ~n51777 ;
  assign n51780 = ~n51778 & ~n51779 ;
  assign n51781 = ~x119 & n20143 ;
  assign n51782 = ~x117 & n20854 ;
  assign n51783 = ~x118 & n20138 ;
  assign n51784 = ~n51782 & ~n51783 ;
  assign n51785 = ~n51781 & n51784 ;
  assign n51786 = n20146 & n20778 ;
  assign n51787 = n51785 & ~n51786 ;
  assign n51788 = ~x56 & ~n51787 ;
  assign n51789 = ~x56 & ~n51788 ;
  assign n51790 = ~n51787 & ~n51788 ;
  assign n51791 = ~n51789 & ~n51790 ;
  assign n51792 = n51780 & ~n51791 ;
  assign n51793 = n51780 & ~n51792 ;
  assign n51794 = ~n51791 & ~n51792 ;
  assign n51795 = ~n51793 & ~n51794 ;
  assign n51796 = ~n51735 & n51795 ;
  assign n51797 = n51735 & ~n51795 ;
  assign n51798 = ~n51796 & ~n51797 ;
  assign n51799 = ~x122 & n18025 ;
  assign n51800 = ~x120 & n18764 ;
  assign n51801 = ~x121 & n18020 ;
  assign n51802 = ~n51800 & ~n51801 ;
  assign n51803 = ~n51799 & n51802 ;
  assign n51804 = n18028 & n22998 ;
  assign n51805 = n51803 & ~n51804 ;
  assign n51806 = ~x53 & ~n51805 ;
  assign n51807 = ~x53 & ~n51806 ;
  assign n51808 = ~n51805 & ~n51806 ;
  assign n51809 = ~n51807 & ~n51808 ;
  assign n51810 = n51798 & n51809 ;
  assign n51811 = ~n51798 & ~n51809 ;
  assign n51812 = ~n51810 & ~n51811 ;
  assign n51813 = ~n51734 & n51812 ;
  assign n51814 = ~n51734 & ~n51813 ;
  assign n51815 = n51812 & ~n51813 ;
  assign n51816 = ~n51814 & ~n51815 ;
  assign n51817 = ~n51733 & ~n51816 ;
  assign n51818 = ~n51733 & ~n51817 ;
  assign n51819 = ~n51816 & ~n51817 ;
  assign n51820 = ~n51818 & ~n51819 ;
  assign n51821 = n51722 & ~n51820 ;
  assign n51822 = n51722 & ~n51821 ;
  assign n51823 = ~n51820 & ~n51821 ;
  assign n51824 = ~n51822 & ~n51823 ;
  assign n51825 = ~n51567 & ~n51573 ;
  assign n51826 = n51824 & n51825 ;
  assign n51827 = ~n51824 & ~n51825 ;
  assign n51828 = ~n51826 & ~n51827 ;
  assign n51829 = ~n51577 & ~n51580 ;
  assign n51830 = n51828 & ~n51829 ;
  assign n51831 = ~n51828 & n51829 ;
  assign n51832 = ~n51830 & ~n51831 ;
  assign n51835 = ~n51832 & ~x237 ;
  assign n51836 = ~n51834 & ~n51835 ;
  assign n51837 = ~n51655 & ~n51669 ;
  assign n51838 = x120 & n20143 ;
  assign n51839 = x118 & n20854 ;
  assign n51840 = x119 & n20138 ;
  assign n51841 = ~n51839 & ~n51840 ;
  assign n51842 = ~n51838 & n51841 ;
  assign n51843 = n20146 & n21143 ;
  assign n51844 = n51842 & ~n51843 ;
  assign n51845 = x56 & ~n51844 ;
  assign n51846 = x56 & ~n51845 ;
  assign n51847 = ~n51844 & ~n51845 ;
  assign n51848 = ~n51846 & ~n51847 ;
  assign n51849 = ~n51647 & ~n51651 ;
  assign n51850 = x117 & n22325 ;
  assign n51851 = x115 & n23066 ;
  assign n51852 = x116 & n22320 ;
  assign n51853 = ~n51851 & ~n51852 ;
  assign n51854 = ~n51850 & n51853 ;
  assign n51855 = n19026 & n22328 ;
  assign n51856 = n51854 & ~n51855 ;
  assign n51857 = x59 & ~n51856 ;
  assign n51858 = x59 & ~n51857 ;
  assign n51859 = ~n51856 & ~n51857 ;
  assign n51860 = ~n51858 & ~n51859 ;
  assign n51861 = ~n51631 & ~n51645 ;
  assign n51862 = x110 & n27024 ;
  assign n51863 = x111 & ~n26217 ;
  assign n51864 = ~n51862 & ~n51863 ;
  assign n51865 = n51628 & ~n51864 ;
  assign n51866 = ~n51628 & n51864 ;
  assign n51867 = ~n51861 & ~n51866 ;
  assign n51868 = ~n51865 & n51867 ;
  assign n51869 = ~n51861 & ~n51868 ;
  assign n51870 = ~n51866 & ~n51868 ;
  assign n51871 = ~n51865 & n51870 ;
  assign n51872 = ~n51869 & ~n51871 ;
  assign n51873 = x114 & n24612 ;
  assign n51874 = x112 & n25390 ;
  assign n51875 = x113 & n24607 ;
  assign n51876 = ~n51874 & ~n51875 ;
  assign n51877 = ~n51873 & n51876 ;
  assign n51878 = n17012 & n24615 ;
  assign n51879 = n51877 & ~n51878 ;
  assign n51880 = x62 & ~n51879 ;
  assign n51881 = x62 & ~n51880 ;
  assign n51882 = ~n51879 & ~n51880 ;
  assign n51883 = ~n51881 & ~n51882 ;
  assign n51884 = ~n51872 & n51883 ;
  assign n51885 = n51872 & ~n51883 ;
  assign n51886 = ~n51884 & ~n51885 ;
  assign n51887 = ~n51860 & ~n51886 ;
  assign n51888 = n51860 & n51886 ;
  assign n51889 = ~n51887 & ~n51888 ;
  assign n51890 = ~n51849 & n51889 ;
  assign n51891 = ~n51849 & ~n51890 ;
  assign n51892 = n51889 & ~n51890 ;
  assign n51893 = ~n51891 & ~n51892 ;
  assign n51894 = ~n51848 & ~n51893 ;
  assign n51895 = n51848 & ~n51892 ;
  assign n51896 = ~n51891 & n51895 ;
  assign n51897 = ~n51894 & ~n51896 ;
  assign n51898 = ~n51837 & n51897 ;
  assign n51899 = n51837 & ~n51897 ;
  assign n51900 = ~n51898 & ~n51899 ;
  assign n51901 = x123 & n18025 ;
  assign n51902 = x121 & n18764 ;
  assign n51903 = x122 & n18020 ;
  assign n51904 = ~n51902 & ~n51903 ;
  assign n51905 = ~n51901 & n51904 ;
  assign n51906 = n18028 & n23382 ;
  assign n51907 = n51905 & ~n51906 ;
  assign n51908 = x53 & ~n51907 ;
  assign n51909 = x53 & ~n51908 ;
  assign n51910 = ~n51907 & ~n51908 ;
  assign n51911 = ~n51909 & ~n51910 ;
  assign n51912 = n51900 & ~n51911 ;
  assign n51913 = n51900 & ~n51912 ;
  assign n51914 = ~n51911 & ~n51912 ;
  assign n51915 = ~n51913 & ~n51914 ;
  assign n51916 = ~n51612 & ~n51672 ;
  assign n51917 = ~n51688 & ~n51916 ;
  assign n51918 = ~n51915 & ~n51917 ;
  assign n51919 = ~n51915 & ~n51918 ;
  assign n51920 = ~n51917 & ~n51918 ;
  assign n51921 = ~n51919 & ~n51920 ;
  assign n51922 = x126 & n16076 ;
  assign n51923 = x124 & n16756 ;
  assign n51924 = x125 & n16071 ;
  assign n51925 = ~n51923 & ~n51924 ;
  assign n51926 = ~n51922 & n51925 ;
  assign n51927 = n16079 & n25735 ;
  assign n51928 = n51926 & ~n51927 ;
  assign n51929 = x50 & ~n51928 ;
  assign n51930 = x50 & ~n51929 ;
  assign n51931 = ~n51928 & ~n51929 ;
  assign n51932 = ~n51930 & ~n51931 ;
  assign n51933 = ~n51921 & ~n51932 ;
  assign n51934 = ~n51921 & ~n51933 ;
  assign n51935 = ~n51932 & ~n51933 ;
  assign n51936 = ~n51934 & ~n51935 ;
  assign n51937 = ~n51690 & ~n51694 ;
  assign n51938 = x127 & n14876 ;
  assign n51939 = ~n14236 & ~n51938 ;
  assign n51940 = ~n26962 & ~n51938 ;
  assign n51941 = ~n51939 & ~n51940 ;
  assign n51942 = x47 & ~n51941 ;
  assign n51943 = ~x47 & n51941 ;
  assign n51944 = ~n51942 & ~n51943 ;
  assign n51945 = ~n51937 & ~n51944 ;
  assign n51946 = n51937 & n51944 ;
  assign n51947 = ~n51945 & ~n51946 ;
  assign n51948 = ~n51936 & n51947 ;
  assign n51949 = ~n51936 & ~n51948 ;
  assign n51950 = n51947 & ~n51948 ;
  assign n51951 = ~n51949 & ~n51950 ;
  assign n51952 = ~n51597 & ~n51698 ;
  assign n51953 = n51951 & n51952 ;
  assign n51954 = ~n51951 & ~n51952 ;
  assign n51955 = ~n51953 & ~n51954 ;
  assign n51956 = ~n51704 & ~n51707 ;
  assign n51957 = n51955 & ~n51956 ;
  assign n51958 = ~n51955 & n51956 ;
  assign n51959 = ~n51957 & ~n51958 ;
  assign n52084 = n51959 & x238 ;
  assign n51960 = ~n51778 & ~n51792 ;
  assign n51961 = ~x120 & n20143 ;
  assign n51962 = ~x118 & n20854 ;
  assign n51963 = ~x119 & n20138 ;
  assign n51964 = ~n51962 & ~n51963 ;
  assign n51965 = ~n51961 & n51964 ;
  assign n51966 = n20146 & n21501 ;
  assign n51967 = n51965 & ~n51966 ;
  assign n51968 = ~x56 & ~n51967 ;
  assign n51969 = ~x56 & ~n51968 ;
  assign n51970 = ~n51967 & ~n51968 ;
  assign n51971 = ~n51969 & ~n51970 ;
  assign n51972 = ~n51770 & ~n51774 ;
  assign n51973 = ~x117 & n22325 ;
  assign n51974 = ~x115 & n23066 ;
  assign n51975 = ~x116 & n22320 ;
  assign n51976 = ~n51974 & ~n51975 ;
  assign n51977 = ~n51973 & n51976 ;
  assign n51978 = n19365 & n22328 ;
  assign n51979 = n51977 & ~n51978 ;
  assign n51980 = ~x59 & ~n51979 ;
  assign n51981 = ~x59 & ~n51980 ;
  assign n51982 = ~n51979 & ~n51980 ;
  assign n51983 = ~n51981 & ~n51982 ;
  assign n51984 = ~n51754 & ~n51768 ;
  assign n51985 = ~x110 & n27427 ;
  assign n51986 = ~x111 & ~n26217 ;
  assign n51987 = ~n51985 & ~n51986 ;
  assign n51988 = n51751 & ~n51987 ;
  assign n51989 = ~n51751 & n51987 ;
  assign n51990 = ~n51984 & ~n51989 ;
  assign n51991 = ~n51988 & n51990 ;
  assign n51992 = ~n51984 & ~n51991 ;
  assign n51993 = ~n51989 & ~n51991 ;
  assign n51994 = ~n51988 & n51993 ;
  assign n51995 = ~n51992 & ~n51994 ;
  assign n51996 = ~x114 & n24612 ;
  assign n51997 = ~x112 & n25390 ;
  assign n51998 = ~x113 & n24607 ;
  assign n51999 = ~n51997 & ~n51998 ;
  assign n52000 = ~n51996 & n51999 ;
  assign n52001 = n17333 & n24615 ;
  assign n52002 = n52000 & ~n52001 ;
  assign n52003 = ~x62 & ~n52002 ;
  assign n52004 = ~x62 & ~n52003 ;
  assign n52005 = ~n52002 & ~n52003 ;
  assign n52006 = ~n52004 & ~n52005 ;
  assign n52007 = ~n51995 & n52006 ;
  assign n52008 = n51995 & ~n52006 ;
  assign n52009 = ~n52007 & ~n52008 ;
  assign n52010 = ~n51983 & ~n52009 ;
  assign n52011 = n51983 & n52009 ;
  assign n52012 = ~n52010 & ~n52011 ;
  assign n52013 = ~n51972 & n52012 ;
  assign n52014 = ~n51972 & ~n52013 ;
  assign n52015 = n52012 & ~n52013 ;
  assign n52016 = ~n52014 & ~n52015 ;
  assign n52017 = ~n51971 & ~n52016 ;
  assign n52018 = n51971 & ~n52015 ;
  assign n52019 = ~n52014 & n52018 ;
  assign n52020 = ~n52017 & ~n52019 ;
  assign n52021 = ~n51960 & n52020 ;
  assign n52022 = n51960 & ~n52020 ;
  assign n52023 = ~n52021 & ~n52022 ;
  assign n52024 = ~x123 & n18025 ;
  assign n52025 = ~x121 & n18764 ;
  assign n52026 = ~x122 & n18020 ;
  assign n52027 = ~n52025 & ~n52026 ;
  assign n52028 = ~n52024 & n52027 ;
  assign n52029 = n18028 & n23760 ;
  assign n52030 = n52028 & ~n52029 ;
  assign n52031 = ~x53 & ~n52030 ;
  assign n52032 = ~x53 & ~n52031 ;
  assign n52033 = ~n52030 & ~n52031 ;
  assign n52034 = ~n52032 & ~n52033 ;
  assign n52035 = n52023 & ~n52034 ;
  assign n52036 = n52023 & ~n52035 ;
  assign n52037 = ~n52034 & ~n52035 ;
  assign n52038 = ~n52036 & ~n52037 ;
  assign n52039 = ~n51735 & ~n51795 ;
  assign n52040 = ~n51811 & ~n52039 ;
  assign n52041 = ~n52038 & ~n52040 ;
  assign n52042 = ~n52038 & ~n52041 ;
  assign n52043 = ~n52040 & ~n52041 ;
  assign n52044 = ~n52042 & ~n52043 ;
  assign n52045 = ~x126 & n16076 ;
  assign n52046 = ~x124 & n16756 ;
  assign n52047 = ~x125 & n16071 ;
  assign n52048 = ~n52046 & ~n52047 ;
  assign n52049 = ~n52045 & n52048 ;
  assign n52050 = n16079 & n26128 ;
  assign n52051 = n52049 & ~n52050 ;
  assign n52052 = ~x50 & ~n52051 ;
  assign n52053 = ~x50 & ~n52052 ;
  assign n52054 = ~n52051 & ~n52052 ;
  assign n52055 = ~n52053 & ~n52054 ;
  assign n52056 = ~n52044 & ~n52055 ;
  assign n52057 = ~n52044 & ~n52056 ;
  assign n52058 = ~n52055 & ~n52056 ;
  assign n52059 = ~n52057 & ~n52058 ;
  assign n52060 = ~n51813 & ~n51817 ;
  assign n52061 = ~x127 & n14876 ;
  assign n52062 = ~n14236 & ~n52061 ;
  assign n52063 = ~n27365 & ~n52061 ;
  assign n52064 = ~n52062 & ~n52063 ;
  assign n52065 = ~x47 & ~n52064 ;
  assign n52066 = x47 & n52064 ;
  assign n52067 = ~n52065 & ~n52066 ;
  assign n52068 = ~n52060 & ~n52067 ;
  assign n52069 = n52060 & n52067 ;
  assign n52070 = ~n52068 & ~n52069 ;
  assign n52071 = ~n52059 & n52070 ;
  assign n52072 = ~n52059 & ~n52071 ;
  assign n52073 = n52070 & ~n52071 ;
  assign n52074 = ~n52072 & ~n52073 ;
  assign n52075 = ~n51720 & ~n51821 ;
  assign n52076 = n52074 & n52075 ;
  assign n52077 = ~n52074 & ~n52075 ;
  assign n52078 = ~n52076 & ~n52077 ;
  assign n52079 = ~n51827 & ~n51830 ;
  assign n52080 = n52078 & ~n52079 ;
  assign n52081 = ~n52078 & n52079 ;
  assign n52082 = ~n52080 & ~n52081 ;
  assign n52085 = ~n52082 & ~x238 ;
  assign n52086 = ~n52084 & ~n52085 ;
  assign n52087 = ~n51898 & ~n51912 ;
  assign n52088 = x124 & n18025 ;
  assign n52089 = x122 & n18764 ;
  assign n52090 = x123 & n18020 ;
  assign n52091 = ~n52089 & ~n52090 ;
  assign n52092 = ~n52088 & n52091 ;
  assign n52093 = n18028 & n23796 ;
  assign n52094 = n52092 & ~n52093 ;
  assign n52095 = x53 & ~n52094 ;
  assign n52096 = x53 & ~n52095 ;
  assign n52097 = ~n52094 & ~n52095 ;
  assign n52098 = ~n52096 & ~n52097 ;
  assign n52099 = ~n51890 & ~n51894 ;
  assign n52100 = x121 & n20143 ;
  assign n52101 = x119 & n20854 ;
  assign n52102 = x120 & n20138 ;
  assign n52103 = ~n52101 & ~n52102 ;
  assign n52104 = ~n52100 & n52103 ;
  assign n52105 = n20146 & n21870 ;
  assign n52106 = n52104 & ~n52105 ;
  assign n52107 = x56 & ~n52106 ;
  assign n52108 = x56 & ~n52107 ;
  assign n52109 = ~n52106 & ~n52107 ;
  assign n52110 = ~n52108 & ~n52109 ;
  assign n52111 = ~n51872 & ~n51883 ;
  assign n52112 = ~n51887 & ~n52111 ;
  assign n52113 = x115 & n24612 ;
  assign n52114 = x113 & n25390 ;
  assign n52115 = x114 & n24607 ;
  assign n52116 = ~n52114 & ~n52115 ;
  assign n52117 = ~n52113 & n52116 ;
  assign n52118 = n17364 & n24615 ;
  assign n52119 = n52117 & ~n52118 ;
  assign n52120 = x62 & ~n52119 ;
  assign n52121 = x62 & ~n52120 ;
  assign n52122 = ~n52119 & ~n52120 ;
  assign n52123 = ~n52121 & ~n52122 ;
  assign n52124 = x111 & n27024 ;
  assign n52125 = x112 & ~n26217 ;
  assign n52126 = ~n52124 & ~n52125 ;
  assign n52127 = x47 & ~n51864 ;
  assign n52128 = ~x47 & n51864 ;
  assign n52129 = ~n52127 & ~n52128 ;
  assign n52130 = ~n52126 & ~n52129 ;
  assign n52131 = n52126 & n52129 ;
  assign n52132 = ~n52130 & ~n52131 ;
  assign n52133 = ~n52123 & n52132 ;
  assign n52134 = ~n52123 & ~n52133 ;
  assign n52135 = n52132 & ~n52133 ;
  assign n52136 = ~n52134 & ~n52135 ;
  assign n52137 = ~n51870 & ~n52136 ;
  assign n52138 = ~n51870 & ~n52137 ;
  assign n52139 = ~n52136 & ~n52137 ;
  assign n52140 = ~n52138 & ~n52139 ;
  assign n52141 = x118 & n22325 ;
  assign n52142 = x116 & n23066 ;
  assign n52143 = x117 & n22320 ;
  assign n52144 = ~n52142 & ~n52143 ;
  assign n52145 = ~n52141 & n52144 ;
  assign n52146 = n19395 & n22328 ;
  assign n52147 = n52145 & ~n52146 ;
  assign n52148 = x59 & ~n52147 ;
  assign n52149 = x59 & ~n52148 ;
  assign n52150 = ~n52147 & ~n52148 ;
  assign n52151 = ~n52149 & ~n52150 ;
  assign n52152 = n52140 & n52151 ;
  assign n52153 = ~n52140 & ~n52151 ;
  assign n52154 = ~n52152 & ~n52153 ;
  assign n52155 = ~n52112 & n52154 ;
  assign n52156 = n52112 & ~n52154 ;
  assign n52157 = ~n52155 & ~n52156 ;
  assign n52158 = n52110 & ~n52157 ;
  assign n52159 = ~n52110 & n52157 ;
  assign n52160 = ~n52158 & ~n52159 ;
  assign n52161 = ~n52099 & n52160 ;
  assign n52162 = n52099 & ~n52160 ;
  assign n52163 = ~n52161 & ~n52162 ;
  assign n52164 = n52098 & ~n52163 ;
  assign n52165 = ~n52098 & n52163 ;
  assign n52166 = ~n52164 & ~n52165 ;
  assign n52167 = ~n52087 & n52166 ;
  assign n52168 = n52087 & ~n52166 ;
  assign n52169 = ~n52167 & ~n52168 ;
  assign n52170 = x127 & n16076 ;
  assign n52171 = x125 & n16756 ;
  assign n52172 = x126 & n16071 ;
  assign n52173 = ~n52171 & ~n52172 ;
  assign n52174 = ~n52170 & n52173 ;
  assign n52175 = n16079 & n26533 ;
  assign n52176 = n52174 & ~n52175 ;
  assign n52177 = x50 & ~n52176 ;
  assign n52178 = x50 & ~n52177 ;
  assign n52179 = ~n52176 & ~n52177 ;
  assign n52180 = ~n52178 & ~n52179 ;
  assign n52181 = n52169 & ~n52180 ;
  assign n52182 = n52169 & ~n52181 ;
  assign n52183 = ~n52180 & ~n52181 ;
  assign n52184 = ~n52182 & ~n52183 ;
  assign n52185 = ~n51918 & ~n51933 ;
  assign n52186 = n52184 & n52185 ;
  assign n52187 = ~n52184 & ~n52185 ;
  assign n52188 = ~n52186 & ~n52187 ;
  assign n52189 = ~n51945 & ~n51948 ;
  assign n52190 = ~n52188 & n52189 ;
  assign n52191 = n52188 & ~n52189 ;
  assign n52192 = ~n52190 & ~n52191 ;
  assign n52193 = ~n51954 & ~n51957 ;
  assign n52194 = n52192 & ~n52193 ;
  assign n52195 = ~n52192 & n52193 ;
  assign n52196 = ~n52194 & ~n52195 ;
  assign n52308 = n52196 & x239 ;
  assign n52197 = ~n52021 & ~n52035 ;
  assign n52198 = ~x124 & n18025 ;
  assign n52199 = ~x122 & n18764 ;
  assign n52200 = ~x123 & n18020 ;
  assign n52201 = ~n52199 & ~n52200 ;
  assign n52202 = ~n52198 & n52201 ;
  assign n52203 = n18028 & n24176 ;
  assign n52204 = n52202 & ~n52203 ;
  assign n52205 = ~x53 & ~n52204 ;
  assign n52206 = ~x53 & ~n52205 ;
  assign n52207 = ~n52204 & ~n52205 ;
  assign n52208 = ~n52206 & ~n52207 ;
  assign n52209 = ~n52013 & ~n52017 ;
  assign n52210 = ~x121 & n20143 ;
  assign n52211 = ~x119 & n20854 ;
  assign n52212 = ~x120 & n20138 ;
  assign n52213 = ~n52211 & ~n52212 ;
  assign n52214 = ~n52210 & n52213 ;
  assign n52215 = n20146 & n22229 ;
  assign n52216 = n52214 & ~n52215 ;
  assign n52217 = ~x56 & ~n52216 ;
  assign n52218 = ~x56 & ~n52217 ;
  assign n52219 = ~n52216 & ~n52217 ;
  assign n52220 = ~n52218 & ~n52219 ;
  assign n52221 = ~n51995 & ~n52006 ;
  assign n52222 = ~n52010 & ~n52221 ;
  assign n52223 = ~x115 & n24612 ;
  assign n52224 = ~x113 & n25390 ;
  assign n52225 = ~x114 & n24607 ;
  assign n52226 = ~n52224 & ~n52225 ;
  assign n52227 = ~n52223 & n52226 ;
  assign n52228 = n17683 & n24615 ;
  assign n52229 = n52227 & ~n52228 ;
  assign n52230 = ~x62 & ~n52229 ;
  assign n52231 = ~x62 & ~n52230 ;
  assign n52232 = ~n52229 & ~n52230 ;
  assign n52233 = ~n52231 & ~n52232 ;
  assign n52234 = ~x111 & n27427 ;
  assign n52235 = ~x112 & ~n26217 ;
  assign n52236 = ~n52234 & ~n52235 ;
  assign n52237 = ~x47 & ~n51987 ;
  assign n52238 = x47 & n51987 ;
  assign n52239 = ~n52237 & ~n52238 ;
  assign n52240 = ~n52236 & ~n52239 ;
  assign n52241 = n52236 & n52239 ;
  assign n52242 = ~n52240 & ~n52241 ;
  assign n52243 = ~n52233 & n52242 ;
  assign n52244 = ~n52233 & ~n52243 ;
  assign n52245 = n52242 & ~n52243 ;
  assign n52246 = ~n52244 & ~n52245 ;
  assign n52247 = ~n51993 & ~n52246 ;
  assign n52248 = ~n51993 & ~n52247 ;
  assign n52249 = ~n52246 & ~n52247 ;
  assign n52250 = ~n52248 & ~n52249 ;
  assign n52251 = ~x118 & n22325 ;
  assign n52252 = ~x116 & n23066 ;
  assign n52253 = ~x117 & n22320 ;
  assign n52254 = ~n52252 & ~n52253 ;
  assign n52255 = ~n52251 & n52254 ;
  assign n52256 = n19736 & n22328 ;
  assign n52257 = n52255 & ~n52256 ;
  assign n52258 = ~x59 & ~n52257 ;
  assign n52259 = ~x59 & ~n52258 ;
  assign n52260 = ~n52257 & ~n52258 ;
  assign n52261 = ~n52259 & ~n52260 ;
  assign n52262 = n52250 & n52261 ;
  assign n52263 = ~n52250 & ~n52261 ;
  assign n52264 = ~n52262 & ~n52263 ;
  assign n52265 = ~n52222 & n52264 ;
  assign n52266 = n52222 & ~n52264 ;
  assign n52267 = ~n52265 & ~n52266 ;
  assign n52268 = n52220 & ~n52267 ;
  assign n52269 = ~n52220 & n52267 ;
  assign n52270 = ~n52268 & ~n52269 ;
  assign n52271 = ~n52209 & n52270 ;
  assign n52272 = n52209 & ~n52270 ;
  assign n52273 = ~n52271 & ~n52272 ;
  assign n52274 = n52208 & ~n52273 ;
  assign n52275 = ~n52208 & n52273 ;
  assign n52276 = ~n52274 & ~n52275 ;
  assign n52277 = ~n52197 & n52276 ;
  assign n52278 = n52197 & ~n52276 ;
  assign n52279 = ~n52277 & ~n52278 ;
  assign n52280 = ~x127 & n16076 ;
  assign n52281 = ~x125 & n16756 ;
  assign n52282 = ~x126 & n16071 ;
  assign n52283 = ~n52281 & ~n52282 ;
  assign n52284 = ~n52280 & n52283 ;
  assign n52285 = n16079 & n26932 ;
  assign n52286 = n52284 & ~n52285 ;
  assign n52287 = ~x50 & ~n52286 ;
  assign n52288 = ~x50 & ~n52287 ;
  assign n52289 = ~n52286 & ~n52287 ;
  assign n52290 = ~n52288 & ~n52289 ;
  assign n52291 = n52279 & ~n52290 ;
  assign n52292 = n52279 & ~n52291 ;
  assign n52293 = ~n52290 & ~n52291 ;
  assign n52294 = ~n52292 & ~n52293 ;
  assign n52295 = ~n52041 & ~n52056 ;
  assign n52296 = n52294 & n52295 ;
  assign n52297 = ~n52294 & ~n52295 ;
  assign n52298 = ~n52296 & ~n52297 ;
  assign n52299 = ~n52068 & ~n52071 ;
  assign n52300 = ~n52298 & n52299 ;
  assign n52301 = n52298 & ~n52299 ;
  assign n52302 = ~n52300 & ~n52301 ;
  assign n52303 = ~n52077 & ~n52080 ;
  assign n52304 = n52302 & ~n52303 ;
  assign n52305 = ~n52302 & n52303 ;
  assign n52306 = ~n52304 & ~n52305 ;
  assign n52309 = ~n52306 & ~x239 ;
  assign n52310 = ~n52308 & ~n52309 ;
  assign n52311 = ~n52165 & ~n52167 ;
  assign n52312 = x125 & n18025 ;
  assign n52313 = x123 & n18764 ;
  assign n52314 = x124 & n18020 ;
  assign n52315 = ~n52313 & ~n52314 ;
  assign n52316 = ~n52312 & n52315 ;
  assign n52317 = n18028 & n24935 ;
  assign n52318 = n52316 & ~n52317 ;
  assign n52319 = x53 & ~n52318 ;
  assign n52320 = x53 & ~n52319 ;
  assign n52321 = ~n52318 & ~n52319 ;
  assign n52322 = ~n52320 & ~n52321 ;
  assign n52323 = ~n52159 & ~n52161 ;
  assign n52324 = x122 & n20143 ;
  assign n52325 = x120 & n20854 ;
  assign n52326 = x121 & n20138 ;
  assign n52327 = ~n52325 & ~n52326 ;
  assign n52328 = ~n52324 & n52327 ;
  assign n52329 = n20146 & n22622 ;
  assign n52330 = n52328 & ~n52329 ;
  assign n52331 = x56 & ~n52330 ;
  assign n52332 = x56 & ~n52331 ;
  assign n52333 = ~n52330 & ~n52331 ;
  assign n52334 = ~n52332 & ~n52333 ;
  assign n52335 = ~n52153 & ~n52155 ;
  assign n52336 = x119 & n22325 ;
  assign n52337 = x117 & n23066 ;
  assign n52338 = x118 & n22320 ;
  assign n52339 = ~n52337 & ~n52338 ;
  assign n52340 = ~n52336 & n52339 ;
  assign n52341 = n20423 & n22328 ;
  assign n52342 = n52340 & ~n52341 ;
  assign n52343 = x59 & ~n52342 ;
  assign n52344 = x59 & ~n52343 ;
  assign n52345 = ~n52342 & ~n52343 ;
  assign n52346 = ~n52344 & ~n52345 ;
  assign n52347 = ~n52133 & ~n52137 ;
  assign n52348 = x112 & n27024 ;
  assign n52349 = x113 & ~n26217 ;
  assign n52350 = ~n52348 & ~n52349 ;
  assign n52351 = ~x47 & ~n51864 ;
  assign n52352 = ~n52130 & ~n52351 ;
  assign n52353 = n52350 & ~n52352 ;
  assign n52354 = ~n52350 & n52352 ;
  assign n52355 = ~n52353 & ~n52354 ;
  assign n52356 = x116 & n24612 ;
  assign n52357 = x114 & n25390 ;
  assign n52358 = x115 & n24607 ;
  assign n52359 = ~n52357 & ~n52358 ;
  assign n52360 = ~n52356 & n52359 ;
  assign n52361 = ~n24615 & n52360 ;
  assign n52362 = ~n18336 & n52360 ;
  assign n52363 = ~n52361 & ~n52362 ;
  assign n52364 = x62 & ~n52363 ;
  assign n52365 = ~x62 & n52363 ;
  assign n52366 = ~n52364 & ~n52365 ;
  assign n52367 = n52355 & ~n52366 ;
  assign n52368 = ~n52355 & n52366 ;
  assign n52369 = ~n52367 & ~n52368 ;
  assign n52370 = ~n52347 & n52369 ;
  assign n52371 = ~n52347 & ~n52370 ;
  assign n52372 = n52369 & ~n52370 ;
  assign n52373 = ~n52371 & ~n52372 ;
  assign n52374 = ~n52346 & ~n52373 ;
  assign n52375 = n52346 & ~n52372 ;
  assign n52376 = ~n52371 & n52375 ;
  assign n52377 = ~n52374 & ~n52376 ;
  assign n52378 = ~n52335 & n52377 ;
  assign n52379 = n52335 & ~n52377 ;
  assign n52380 = ~n52378 & ~n52379 ;
  assign n52381 = ~n52334 & n52380 ;
  assign n52382 = n52334 & ~n52380 ;
  assign n52383 = ~n52381 & ~n52382 ;
  assign n52384 = ~n52323 & n52383 ;
  assign n52385 = ~n52323 & ~n52384 ;
  assign n52386 = n52383 & ~n52384 ;
  assign n52387 = ~n52385 & ~n52386 ;
  assign n52388 = ~n52322 & ~n52387 ;
  assign n52389 = n52322 & ~n52386 ;
  assign n52390 = ~n52385 & n52389 ;
  assign n52391 = ~n52388 & ~n52390 ;
  assign n52392 = ~n52311 & n52391 ;
  assign n52393 = n52311 & ~n52391 ;
  assign n52394 = ~n52392 & ~n52393 ;
  assign n52395 = x126 & n16756 ;
  assign n52396 = x127 & n16071 ;
  assign n52397 = ~n52395 & ~n52396 ;
  assign n52398 = n16079 & ~n26965 ;
  assign n52399 = n52397 & ~n52398 ;
  assign n52400 = x50 & ~n52399 ;
  assign n52401 = x50 & ~n52400 ;
  assign n52402 = ~n52399 & ~n52400 ;
  assign n52403 = ~n52401 & ~n52402 ;
  assign n52404 = n52394 & ~n52403 ;
  assign n52405 = n52394 & ~n52404 ;
  assign n52406 = ~n52403 & ~n52404 ;
  assign n52407 = ~n52405 & ~n52406 ;
  assign n52408 = ~n52181 & ~n52187 ;
  assign n52409 = n52407 & n52408 ;
  assign n52410 = ~n52407 & ~n52408 ;
  assign n52411 = ~n52409 & ~n52410 ;
  assign n52412 = ~n52191 & ~n52194 ;
  assign n52413 = n52411 & ~n52412 ;
  assign n52414 = ~n52411 & n52412 ;
  assign n52415 = ~n52413 & ~n52414 ;
  assign n52522 = n52415 & x240 ;
  assign n52416 = ~n52275 & ~n52277 ;
  assign n52417 = ~x125 & n18025 ;
  assign n52418 = ~x123 & n18764 ;
  assign n52419 = ~x124 & n18020 ;
  assign n52420 = ~n52418 & ~n52419 ;
  assign n52421 = ~n52417 & n52420 ;
  assign n52422 = n18028 & n25330 ;
  assign n52423 = n52421 & ~n52422 ;
  assign n52424 = ~x53 & ~n52423 ;
  assign n52425 = ~x53 & ~n52424 ;
  assign n52426 = ~n52423 & ~n52424 ;
  assign n52427 = ~n52425 & ~n52426 ;
  assign n52428 = ~n52269 & ~n52271 ;
  assign n52429 = ~x122 & n20143 ;
  assign n52430 = ~x120 & n20854 ;
  assign n52431 = ~x121 & n20138 ;
  assign n52432 = ~n52430 & ~n52431 ;
  assign n52433 = ~n52429 & n52432 ;
  assign n52434 = n20146 & n22998 ;
  assign n52435 = n52433 & ~n52434 ;
  assign n52436 = ~x56 & ~n52435 ;
  assign n52437 = ~x56 & ~n52436 ;
  assign n52438 = ~n52435 & ~n52436 ;
  assign n52439 = ~n52437 & ~n52438 ;
  assign n52440 = ~n52263 & ~n52265 ;
  assign n52441 = ~x119 & n22325 ;
  assign n52442 = ~x117 & n23066 ;
  assign n52443 = ~x118 & n22320 ;
  assign n52444 = ~n52442 & ~n52443 ;
  assign n52445 = ~n52441 & n52444 ;
  assign n52446 = n20778 & n22328 ;
  assign n52447 = n52445 & ~n52446 ;
  assign n52448 = ~x59 & ~n52447 ;
  assign n52449 = ~x59 & ~n52448 ;
  assign n52450 = ~n52447 & ~n52448 ;
  assign n52451 = ~n52449 & ~n52450 ;
  assign n52452 = ~n52243 & ~n52247 ;
  assign n52453 = ~x112 & n27427 ;
  assign n52454 = ~x113 & ~n26217 ;
  assign n52455 = ~n52453 & ~n52454 ;
  assign n52456 = x47 & ~n51987 ;
  assign n52457 = ~n52240 & ~n52456 ;
  assign n52458 = n52455 & ~n52457 ;
  assign n52459 = ~n52455 & n52457 ;
  assign n52460 = ~n52458 & ~n52459 ;
  assign n52461 = ~x116 & n24612 ;
  assign n52462 = ~x114 & n25390 ;
  assign n52463 = ~x115 & n24607 ;
  assign n52464 = ~n52462 & ~n52463 ;
  assign n52465 = ~n52461 & n52464 ;
  assign n52466 = ~n24615 & n52465 ;
  assign n52467 = ~n18678 & n52465 ;
  assign n52468 = ~n52466 & ~n52467 ;
  assign n52469 = ~x62 & ~n52468 ;
  assign n52470 = x62 & n52468 ;
  assign n52471 = ~n52469 & ~n52470 ;
  assign n52472 = n52460 & ~n52471 ;
  assign n52473 = ~n52460 & n52471 ;
  assign n52474 = ~n52472 & ~n52473 ;
  assign n52475 = ~n52452 & n52474 ;
  assign n52476 = ~n52452 & ~n52475 ;
  assign n52477 = n52474 & ~n52475 ;
  assign n52478 = ~n52476 & ~n52477 ;
  assign n52479 = ~n52451 & ~n52478 ;
  assign n52480 = n52451 & ~n52477 ;
  assign n52481 = ~n52476 & n52480 ;
  assign n52482 = ~n52479 & ~n52481 ;
  assign n52483 = ~n52440 & n52482 ;
  assign n52484 = n52440 & ~n52482 ;
  assign n52485 = ~n52483 & ~n52484 ;
  assign n52486 = ~n52439 & n52485 ;
  assign n52487 = n52439 & ~n52485 ;
  assign n52488 = ~n52486 & ~n52487 ;
  assign n52489 = ~n52428 & n52488 ;
  assign n52490 = ~n52428 & ~n52489 ;
  assign n52491 = n52488 & ~n52489 ;
  assign n52492 = ~n52490 & ~n52491 ;
  assign n52493 = ~n52427 & ~n52492 ;
  assign n52494 = n52427 & ~n52491 ;
  assign n52495 = ~n52490 & n52494 ;
  assign n52496 = ~n52493 & ~n52495 ;
  assign n52497 = ~n52416 & n52496 ;
  assign n52498 = n52416 & ~n52496 ;
  assign n52499 = ~n52497 & ~n52498 ;
  assign n52500 = ~x126 & n16756 ;
  assign n52501 = ~x127 & n16071 ;
  assign n52502 = ~n52500 & ~n52501 ;
  assign n52503 = n16079 & ~n27368 ;
  assign n52504 = n52502 & ~n52503 ;
  assign n52505 = ~x50 & ~n52504 ;
  assign n52506 = ~x50 & ~n52505 ;
  assign n52507 = ~n52504 & ~n52505 ;
  assign n52508 = ~n52506 & ~n52507 ;
  assign n52509 = n52499 & ~n52508 ;
  assign n52510 = n52499 & ~n52509 ;
  assign n52511 = ~n52508 & ~n52509 ;
  assign n52512 = ~n52510 & ~n52511 ;
  assign n52513 = ~n52291 & ~n52297 ;
  assign n52514 = n52512 & n52513 ;
  assign n52515 = ~n52512 & ~n52513 ;
  assign n52516 = ~n52514 & ~n52515 ;
  assign n52517 = ~n52301 & ~n52304 ;
  assign n52518 = n52516 & ~n52517 ;
  assign n52519 = ~n52516 & n52517 ;
  assign n52520 = ~n52518 & ~n52519 ;
  assign n52523 = ~n52520 & ~x240 ;
  assign n52524 = ~n52522 & ~n52523 ;
  assign n52525 = ~n52370 & ~n52374 ;
  assign n52526 = x117 & n24612 ;
  assign n52527 = x115 & n25390 ;
  assign n52528 = x116 & n24607 ;
  assign n52529 = ~n52527 & ~n52528 ;
  assign n52530 = ~n52526 & n52529 ;
  assign n52531 = n19026 & n24615 ;
  assign n52532 = n52530 & ~n52531 ;
  assign n52533 = x62 & ~n52532 ;
  assign n52534 = x62 & ~n52533 ;
  assign n52535 = ~n52532 & ~n52533 ;
  assign n52536 = ~n52534 & ~n52535 ;
  assign n52537 = x113 & n27024 ;
  assign n52538 = x114 & ~n26217 ;
  assign n52539 = ~n52537 & ~n52538 ;
  assign n52540 = n52350 & ~n52539 ;
  assign n52541 = n52350 & ~n52540 ;
  assign n52542 = ~n52539 & ~n52540 ;
  assign n52543 = ~n52541 & ~n52542 ;
  assign n52544 = ~n52536 & ~n52543 ;
  assign n52545 = ~n52536 & ~n52544 ;
  assign n52546 = ~n52543 & ~n52544 ;
  assign n52547 = ~n52545 & ~n52546 ;
  assign n52548 = ~n52353 & ~n52367 ;
  assign n52549 = n52547 & n52548 ;
  assign n52550 = ~n52547 & ~n52548 ;
  assign n52551 = ~n52549 & ~n52550 ;
  assign n52552 = x120 & n22325 ;
  assign n52553 = x118 & n23066 ;
  assign n52554 = x119 & n22320 ;
  assign n52555 = ~n52553 & ~n52554 ;
  assign n52556 = ~n52552 & n52555 ;
  assign n52557 = n21143 & n22328 ;
  assign n52558 = n52556 & ~n52557 ;
  assign n52559 = x59 & ~n52558 ;
  assign n52560 = x59 & ~n52559 ;
  assign n52561 = ~n52558 & ~n52559 ;
  assign n52562 = ~n52560 & ~n52561 ;
  assign n52563 = ~n52551 & n52562 ;
  assign n52564 = n52551 & ~n52562 ;
  assign n52565 = ~n52563 & ~n52564 ;
  assign n52566 = ~n52525 & n52565 ;
  assign n52567 = n52525 & ~n52565 ;
  assign n52568 = ~n52566 & ~n52567 ;
  assign n52569 = x123 & n20143 ;
  assign n52570 = x121 & n20854 ;
  assign n52571 = x122 & n20138 ;
  assign n52572 = ~n52570 & ~n52571 ;
  assign n52573 = ~n52569 & n52572 ;
  assign n52574 = n20146 & n23382 ;
  assign n52575 = n52573 & ~n52574 ;
  assign n52576 = x56 & ~n52575 ;
  assign n52577 = x56 & ~n52576 ;
  assign n52578 = ~n52575 & ~n52576 ;
  assign n52579 = ~n52577 & ~n52578 ;
  assign n52580 = n52568 & ~n52579 ;
  assign n52581 = n52568 & ~n52580 ;
  assign n52582 = ~n52579 & ~n52580 ;
  assign n52583 = ~n52581 & ~n52582 ;
  assign n52584 = ~n52378 & ~n52381 ;
  assign n52585 = n52583 & n52584 ;
  assign n52586 = ~n52583 & ~n52584 ;
  assign n52587 = ~n52585 & ~n52586 ;
  assign n52588 = x126 & n18025 ;
  assign n52589 = x124 & n18764 ;
  assign n52590 = x125 & n18020 ;
  assign n52591 = ~n52589 & ~n52590 ;
  assign n52592 = ~n52588 & n52591 ;
  assign n52593 = n18028 & n25735 ;
  assign n52594 = n52592 & ~n52593 ;
  assign n52595 = x53 & ~n52594 ;
  assign n52596 = x53 & ~n52595 ;
  assign n52597 = ~n52594 & ~n52595 ;
  assign n52598 = ~n52596 & ~n52597 ;
  assign n52599 = n52587 & ~n52598 ;
  assign n52600 = n52587 & ~n52599 ;
  assign n52601 = ~n52598 & ~n52599 ;
  assign n52602 = ~n52600 & ~n52601 ;
  assign n52603 = ~n52384 & ~n52388 ;
  assign n52604 = x127 & n16756 ;
  assign n52605 = ~n16079 & ~n52604 ;
  assign n52606 = ~n26962 & ~n52604 ;
  assign n52607 = ~n52605 & ~n52606 ;
  assign n52608 = x50 & ~n52607 ;
  assign n52609 = ~x50 & n52607 ;
  assign n52610 = ~n52608 & ~n52609 ;
  assign n52611 = ~n52603 & ~n52610 ;
  assign n52612 = n52603 & n52610 ;
  assign n52613 = ~n52611 & ~n52612 ;
  assign n52614 = ~n52602 & n52613 ;
  assign n52615 = ~n52602 & ~n52614 ;
  assign n52616 = n52613 & ~n52614 ;
  assign n52617 = ~n52615 & ~n52616 ;
  assign n52618 = ~n52392 & ~n52404 ;
  assign n52619 = n52617 & n52618 ;
  assign n52620 = ~n52617 & ~n52618 ;
  assign n52621 = ~n52619 & ~n52620 ;
  assign n52622 = ~n52410 & ~n52413 ;
  assign n52623 = n52621 & ~n52622 ;
  assign n52624 = ~n52621 & n52622 ;
  assign n52625 = ~n52623 & ~n52624 ;
  assign n52728 = n52625 & x241 ;
  assign n52626 = ~n52475 & ~n52479 ;
  assign n52627 = ~x117 & n24612 ;
  assign n52628 = ~x115 & n25390 ;
  assign n52629 = ~x116 & n24607 ;
  assign n52630 = ~n52628 & ~n52629 ;
  assign n52631 = ~n52627 & n52630 ;
  assign n52632 = n19365 & n24615 ;
  assign n52633 = n52631 & ~n52632 ;
  assign n52634 = ~x62 & ~n52633 ;
  assign n52635 = ~x62 & ~n52634 ;
  assign n52636 = ~n52633 & ~n52634 ;
  assign n52637 = ~n52635 & ~n52636 ;
  assign n52638 = ~x113 & n27427 ;
  assign n52639 = ~x114 & ~n26217 ;
  assign n52640 = ~n52638 & ~n52639 ;
  assign n52641 = n52455 & ~n52640 ;
  assign n52642 = n52455 & ~n52641 ;
  assign n52643 = ~n52640 & ~n52641 ;
  assign n52644 = ~n52642 & ~n52643 ;
  assign n52645 = ~n52637 & ~n52644 ;
  assign n52646 = ~n52637 & ~n52645 ;
  assign n52647 = ~n52644 & ~n52645 ;
  assign n52648 = ~n52646 & ~n52647 ;
  assign n52649 = ~n52458 & ~n52472 ;
  assign n52650 = n52648 & n52649 ;
  assign n52651 = ~n52648 & ~n52649 ;
  assign n52652 = ~n52650 & ~n52651 ;
  assign n52653 = ~x120 & n22325 ;
  assign n52654 = ~x118 & n23066 ;
  assign n52655 = ~x119 & n22320 ;
  assign n52656 = ~n52654 & ~n52655 ;
  assign n52657 = ~n52653 & n52656 ;
  assign n52658 = n21501 & n22328 ;
  assign n52659 = n52657 & ~n52658 ;
  assign n52660 = ~x59 & ~n52659 ;
  assign n52661 = ~x59 & ~n52660 ;
  assign n52662 = ~n52659 & ~n52660 ;
  assign n52663 = ~n52661 & ~n52662 ;
  assign n52664 = ~n52652 & n52663 ;
  assign n52665 = n52652 & ~n52663 ;
  assign n52666 = ~n52664 & ~n52665 ;
  assign n52667 = ~n52626 & n52666 ;
  assign n52668 = n52626 & ~n52666 ;
  assign n52669 = ~n52667 & ~n52668 ;
  assign n52670 = ~x123 & n20143 ;
  assign n52671 = ~x121 & n20854 ;
  assign n52672 = ~x122 & n20138 ;
  assign n52673 = ~n52671 & ~n52672 ;
  assign n52674 = ~n52670 & n52673 ;
  assign n52675 = n20146 & n23760 ;
  assign n52676 = n52674 & ~n52675 ;
  assign n52677 = ~x56 & ~n52676 ;
  assign n52678 = ~x56 & ~n52677 ;
  assign n52679 = ~n52676 & ~n52677 ;
  assign n52680 = ~n52678 & ~n52679 ;
  assign n52681 = n52669 & ~n52680 ;
  assign n52682 = n52669 & ~n52681 ;
  assign n52683 = ~n52680 & ~n52681 ;
  assign n52684 = ~n52682 & ~n52683 ;
  assign n52685 = ~n52483 & ~n52486 ;
  assign n52686 = n52684 & n52685 ;
  assign n52687 = ~n52684 & ~n52685 ;
  assign n52688 = ~n52686 & ~n52687 ;
  assign n52689 = ~x126 & n18025 ;
  assign n52690 = ~x124 & n18764 ;
  assign n52691 = ~x125 & n18020 ;
  assign n52692 = ~n52690 & ~n52691 ;
  assign n52693 = ~n52689 & n52692 ;
  assign n52694 = n18028 & n26128 ;
  assign n52695 = n52693 & ~n52694 ;
  assign n52696 = ~x53 & ~n52695 ;
  assign n52697 = ~x53 & ~n52696 ;
  assign n52698 = ~n52695 & ~n52696 ;
  assign n52699 = ~n52697 & ~n52698 ;
  assign n52700 = n52688 & ~n52699 ;
  assign n52701 = n52688 & ~n52700 ;
  assign n52702 = ~n52699 & ~n52700 ;
  assign n52703 = ~n52701 & ~n52702 ;
  assign n52704 = ~n52489 & ~n52493 ;
  assign n52705 = ~x127 & n16756 ;
  assign n52706 = ~n16079 & ~n52705 ;
  assign n52707 = ~n27365 & ~n52705 ;
  assign n52708 = ~n52706 & ~n52707 ;
  assign n52709 = ~x50 & ~n52708 ;
  assign n52710 = x50 & n52708 ;
  assign n52711 = ~n52709 & ~n52710 ;
  assign n52712 = ~n52704 & ~n52711 ;
  assign n52713 = n52704 & n52711 ;
  assign n52714 = ~n52712 & ~n52713 ;
  assign n52715 = ~n52703 & n52714 ;
  assign n52716 = ~n52703 & ~n52715 ;
  assign n52717 = n52714 & ~n52715 ;
  assign n52718 = ~n52716 & ~n52717 ;
  assign n52719 = ~n52497 & ~n52509 ;
  assign n52720 = n52718 & n52719 ;
  assign n52721 = ~n52718 & ~n52719 ;
  assign n52722 = ~n52720 & ~n52721 ;
  assign n52723 = ~n52515 & ~n52518 ;
  assign n52724 = n52722 & ~n52723 ;
  assign n52725 = ~n52722 & n52723 ;
  assign n52726 = ~n52724 & ~n52725 ;
  assign n52729 = ~n52726 & ~x241 ;
  assign n52730 = ~n52728 & ~n52729 ;
  assign n52731 = ~n52566 & ~n52580 ;
  assign n52732 = x124 & n20143 ;
  assign n52733 = x122 & n20854 ;
  assign n52734 = x123 & n20138 ;
  assign n52735 = ~n52733 & ~n52734 ;
  assign n52736 = ~n52732 & n52735 ;
  assign n52737 = n20146 & n23796 ;
  assign n52738 = n52736 & ~n52737 ;
  assign n52739 = x56 & ~n52738 ;
  assign n52740 = x56 & ~n52739 ;
  assign n52741 = ~n52738 & ~n52739 ;
  assign n52742 = ~n52740 & ~n52741 ;
  assign n52743 = ~n52550 & ~n52564 ;
  assign n52744 = x121 & n22325 ;
  assign n52745 = x119 & n23066 ;
  assign n52746 = x120 & n22320 ;
  assign n52747 = ~n52745 & ~n52746 ;
  assign n52748 = ~n52744 & n52747 ;
  assign n52749 = n21870 & n22328 ;
  assign n52750 = n52748 & ~n52749 ;
  assign n52751 = x59 & ~n52750 ;
  assign n52752 = x59 & ~n52751 ;
  assign n52753 = ~n52750 & ~n52751 ;
  assign n52754 = ~n52752 & ~n52753 ;
  assign n52755 = x118 & n24612 ;
  assign n52756 = x116 & n25390 ;
  assign n52757 = x117 & n24607 ;
  assign n52758 = ~n52756 & ~n52757 ;
  assign n52759 = ~n52755 & n52758 ;
  assign n52760 = n19395 & n24615 ;
  assign n52761 = n52759 & ~n52760 ;
  assign n52762 = x62 & ~n52761 ;
  assign n52763 = x62 & ~n52762 ;
  assign n52764 = ~n52761 & ~n52762 ;
  assign n52765 = ~n52763 & ~n52764 ;
  assign n52766 = ~n52540 & ~n52544 ;
  assign n52767 = x114 & n27024 ;
  assign n52768 = x115 & ~n26217 ;
  assign n52769 = ~n52767 & ~n52768 ;
  assign n52770 = ~x50 & ~n52769 ;
  assign n52771 = x50 & n52769 ;
  assign n52772 = ~n52770 & ~n52771 ;
  assign n52773 = ~n52350 & n52772 ;
  assign n52774 = n52350 & ~n52772 ;
  assign n52775 = ~n52773 & ~n52774 ;
  assign n52776 = ~n52766 & n52775 ;
  assign n52777 = ~n52766 & ~n52776 ;
  assign n52778 = n52775 & ~n52776 ;
  assign n52779 = ~n52777 & ~n52778 ;
  assign n52780 = ~n52765 & ~n52779 ;
  assign n52781 = n52765 & ~n52778 ;
  assign n52782 = ~n52777 & n52781 ;
  assign n52783 = ~n52780 & ~n52782 ;
  assign n52784 = ~n52754 & n52783 ;
  assign n52785 = ~n52754 & ~n52784 ;
  assign n52786 = n52783 & ~n52784 ;
  assign n52787 = ~n52785 & ~n52786 ;
  assign n52788 = ~n52743 & ~n52787 ;
  assign n52789 = n52743 & ~n52786 ;
  assign n52790 = ~n52785 & n52789 ;
  assign n52791 = ~n52788 & ~n52790 ;
  assign n52792 = ~n52742 & n52791 ;
  assign n52793 = n52742 & ~n52791 ;
  assign n52794 = ~n52792 & ~n52793 ;
  assign n52795 = ~n52731 & n52794 ;
  assign n52796 = n52731 & ~n52794 ;
  assign n52797 = ~n52795 & ~n52796 ;
  assign n52798 = x127 & n18025 ;
  assign n52799 = x125 & n18764 ;
  assign n52800 = x126 & n18020 ;
  assign n52801 = ~n52799 & ~n52800 ;
  assign n52802 = ~n52798 & n52801 ;
  assign n52803 = n18028 & n26533 ;
  assign n52804 = n52802 & ~n52803 ;
  assign n52805 = x53 & ~n52804 ;
  assign n52806 = x53 & ~n52805 ;
  assign n52807 = ~n52804 & ~n52805 ;
  assign n52808 = ~n52806 & ~n52807 ;
  assign n52809 = n52797 & ~n52808 ;
  assign n52810 = n52797 & ~n52809 ;
  assign n52811 = ~n52808 & ~n52809 ;
  assign n52812 = ~n52810 & ~n52811 ;
  assign n52813 = ~n52586 & ~n52599 ;
  assign n52814 = n52812 & n52813 ;
  assign n52815 = ~n52812 & ~n52813 ;
  assign n52816 = ~n52814 & ~n52815 ;
  assign n52817 = ~n52611 & ~n52614 ;
  assign n52818 = ~n52816 & n52817 ;
  assign n52819 = n52816 & ~n52817 ;
  assign n52820 = ~n52818 & ~n52819 ;
  assign n52821 = ~n52620 & ~n52623 ;
  assign n52822 = n52820 & ~n52821 ;
  assign n52823 = ~n52820 & n52821 ;
  assign n52824 = ~n52822 & ~n52823 ;
  assign n52920 = n52824 & x242 ;
  assign n52825 = ~n52667 & ~n52681 ;
  assign n52826 = ~x124 & n20143 ;
  assign n52827 = ~x122 & n20854 ;
  assign n52828 = ~x123 & n20138 ;
  assign n52829 = ~n52827 & ~n52828 ;
  assign n52830 = ~n52826 & n52829 ;
  assign n52831 = n20146 & n24176 ;
  assign n52832 = n52830 & ~n52831 ;
  assign n52833 = ~x56 & ~n52832 ;
  assign n52834 = ~x56 & ~n52833 ;
  assign n52835 = ~n52832 & ~n52833 ;
  assign n52836 = ~n52834 & ~n52835 ;
  assign n52837 = ~n52651 & ~n52665 ;
  assign n52838 = ~x121 & n22325 ;
  assign n52839 = ~x119 & n23066 ;
  assign n52840 = ~x120 & n22320 ;
  assign n52841 = ~n52839 & ~n52840 ;
  assign n52842 = ~n52838 & n52841 ;
  assign n52843 = n22229 & n22328 ;
  assign n52844 = n52842 & ~n52843 ;
  assign n52845 = ~x59 & ~n52844 ;
  assign n52846 = ~x59 & ~n52845 ;
  assign n52847 = ~n52844 & ~n52845 ;
  assign n52848 = ~n52846 & ~n52847 ;
  assign n52849 = ~x118 & n24612 ;
  assign n52850 = ~x116 & n25390 ;
  assign n52851 = ~x117 & n24607 ;
  assign n52852 = ~n52850 & ~n52851 ;
  assign n52853 = ~n52849 & n52852 ;
  assign n52854 = n19736 & n24615 ;
  assign n52855 = n52853 & ~n52854 ;
  assign n52856 = ~x62 & ~n52855 ;
  assign n52857 = ~x62 & ~n52856 ;
  assign n52858 = ~n52855 & ~n52856 ;
  assign n52859 = ~n52857 & ~n52858 ;
  assign n52860 = ~n52641 & ~n52645 ;
  assign n52861 = ~x114 & n27427 ;
  assign n52862 = ~x115 & ~n26217 ;
  assign n52863 = ~n52861 & ~n52862 ;
  assign n52864 = x50 & ~n52863 ;
  assign n52865 = ~x50 & n52863 ;
  assign n52866 = ~n52864 & ~n52865 ;
  assign n52867 = ~n52455 & n52866 ;
  assign n52868 = n52455 & ~n52866 ;
  assign n52869 = ~n52867 & ~n52868 ;
  assign n52870 = ~n52860 & n52869 ;
  assign n52871 = ~n52860 & ~n52870 ;
  assign n52872 = n52869 & ~n52870 ;
  assign n52873 = ~n52871 & ~n52872 ;
  assign n52874 = ~n52859 & ~n52873 ;
  assign n52875 = n52859 & ~n52872 ;
  assign n52876 = ~n52871 & n52875 ;
  assign n52877 = ~n52874 & ~n52876 ;
  assign n52878 = ~n52848 & n52877 ;
  assign n52879 = ~n52848 & ~n52878 ;
  assign n52880 = n52877 & ~n52878 ;
  assign n52881 = ~n52879 & ~n52880 ;
  assign n52882 = ~n52837 & ~n52881 ;
  assign n52883 = n52837 & ~n52880 ;
  assign n52884 = ~n52879 & n52883 ;
  assign n52885 = ~n52882 & ~n52884 ;
  assign n52886 = ~n52836 & n52885 ;
  assign n52887 = n52836 & ~n52885 ;
  assign n52888 = ~n52886 & ~n52887 ;
  assign n52889 = ~n52825 & n52888 ;
  assign n52890 = n52825 & ~n52888 ;
  assign n52891 = ~n52889 & ~n52890 ;
  assign n52892 = ~x127 & n18025 ;
  assign n52893 = ~x125 & n18764 ;
  assign n52894 = ~x126 & n18020 ;
  assign n52895 = ~n52893 & ~n52894 ;
  assign n52896 = ~n52892 & n52895 ;
  assign n52897 = n18028 & n26932 ;
  assign n52898 = n52896 & ~n52897 ;
  assign n52899 = ~x53 & ~n52898 ;
  assign n52900 = ~x53 & ~n52899 ;
  assign n52901 = ~n52898 & ~n52899 ;
  assign n52902 = ~n52900 & ~n52901 ;
  assign n52903 = n52891 & ~n52902 ;
  assign n52904 = n52891 & ~n52903 ;
  assign n52905 = ~n52902 & ~n52903 ;
  assign n52906 = ~n52904 & ~n52905 ;
  assign n52907 = ~n52687 & ~n52700 ;
  assign n52908 = n52906 & n52907 ;
  assign n52909 = ~n52906 & ~n52907 ;
  assign n52910 = ~n52908 & ~n52909 ;
  assign n52911 = ~n52712 & ~n52715 ;
  assign n52912 = ~n52910 & n52911 ;
  assign n52913 = n52910 & ~n52911 ;
  assign n52914 = ~n52912 & ~n52913 ;
  assign n52915 = ~n52721 & ~n52724 ;
  assign n52916 = n52914 & ~n52915 ;
  assign n52917 = ~n52914 & n52915 ;
  assign n52918 = ~n52916 & ~n52917 ;
  assign n52921 = ~n52918 & ~x242 ;
  assign n52922 = ~n52920 & ~n52921 ;
  assign n52923 = ~n52792 & ~n52795 ;
  assign n52924 = x125 & n20143 ;
  assign n52925 = x123 & n20854 ;
  assign n52926 = x124 & n20138 ;
  assign n52927 = ~n52925 & ~n52926 ;
  assign n52928 = ~n52924 & n52927 ;
  assign n52929 = n20146 & n24935 ;
  assign n52930 = n52928 & ~n52929 ;
  assign n52931 = x56 & ~n52930 ;
  assign n52932 = x56 & ~n52931 ;
  assign n52933 = ~n52930 & ~n52931 ;
  assign n52934 = ~n52932 & ~n52933 ;
  assign n52935 = ~n52784 & ~n52788 ;
  assign n52936 = x122 & n22325 ;
  assign n52937 = x120 & n23066 ;
  assign n52938 = x121 & n22320 ;
  assign n52939 = ~n52937 & ~n52938 ;
  assign n52940 = ~n52936 & n52939 ;
  assign n52941 = n22328 & n22622 ;
  assign n52942 = n52940 & ~n52941 ;
  assign n52943 = x59 & ~n52942 ;
  assign n52944 = x59 & ~n52943 ;
  assign n52945 = ~n52942 & ~n52943 ;
  assign n52946 = ~n52944 & ~n52945 ;
  assign n52947 = ~n52776 & ~n52780 ;
  assign n52948 = x115 & n27024 ;
  assign n52949 = x116 & ~n26217 ;
  assign n52950 = ~n52948 & ~n52949 ;
  assign n52951 = ~n52770 & ~n52773 ;
  assign n52952 = ~n52950 & n52951 ;
  assign n52953 = n52950 & ~n52951 ;
  assign n52954 = ~n52952 & ~n52953 ;
  assign n52955 = x119 & n24612 ;
  assign n52956 = x117 & n25390 ;
  assign n52957 = x118 & n24607 ;
  assign n52958 = ~n52956 & ~n52957 ;
  assign n52959 = ~n52955 & n52958 ;
  assign n52960 = n20423 & n24615 ;
  assign n52961 = n52959 & ~n52960 ;
  assign n52962 = x62 & ~n52961 ;
  assign n52963 = x62 & ~n52962 ;
  assign n52964 = ~n52961 & ~n52962 ;
  assign n52965 = ~n52963 & ~n52964 ;
  assign n52966 = ~n52954 & n52965 ;
  assign n52967 = n52954 & ~n52965 ;
  assign n52968 = ~n52966 & ~n52967 ;
  assign n52969 = ~n52947 & n52968 ;
  assign n52970 = n52947 & ~n52968 ;
  assign n52971 = ~n52969 & ~n52970 ;
  assign n52972 = ~n52946 & n52971 ;
  assign n52973 = n52946 & ~n52971 ;
  assign n52974 = ~n52972 & ~n52973 ;
  assign n52975 = ~n52935 & n52974 ;
  assign n52976 = ~n52935 & ~n52975 ;
  assign n52977 = n52974 & ~n52975 ;
  assign n52978 = ~n52976 & ~n52977 ;
  assign n52979 = ~n52934 & ~n52978 ;
  assign n52980 = n52934 & ~n52977 ;
  assign n52981 = ~n52976 & n52980 ;
  assign n52982 = ~n52979 & ~n52981 ;
  assign n52983 = ~n52923 & n52982 ;
  assign n52984 = n52923 & ~n52982 ;
  assign n52985 = ~n52983 & ~n52984 ;
  assign n52986 = x126 & n18764 ;
  assign n52987 = x127 & n18020 ;
  assign n52988 = ~n52986 & ~n52987 ;
  assign n52989 = n18028 & ~n26965 ;
  assign n52990 = n52988 & ~n52989 ;
  assign n52991 = x53 & ~n52990 ;
  assign n52992 = x53 & ~n52991 ;
  assign n52993 = ~n52990 & ~n52991 ;
  assign n52994 = ~n52992 & ~n52993 ;
  assign n52995 = n52985 & ~n52994 ;
  assign n52996 = n52985 & ~n52995 ;
  assign n52997 = ~n52994 & ~n52995 ;
  assign n52998 = ~n52996 & ~n52997 ;
  assign n52999 = ~n52809 & ~n52815 ;
  assign n53000 = n52998 & n52999 ;
  assign n53001 = ~n52998 & ~n52999 ;
  assign n53002 = ~n53000 & ~n53001 ;
  assign n53003 = ~n52819 & ~n52822 ;
  assign n53004 = n53002 & ~n53003 ;
  assign n53005 = ~n53002 & n53003 ;
  assign n53006 = ~n53004 & ~n53005 ;
  assign n53092 = n53006 & x243 ;
  assign n53007 = ~n52886 & ~n52889 ;
  assign n53008 = ~x125 & n20143 ;
  assign n53009 = ~x123 & n20854 ;
  assign n53010 = ~x124 & n20138 ;
  assign n53011 = ~n53009 & ~n53010 ;
  assign n53012 = ~n53008 & n53011 ;
  assign n53013 = n20146 & n25330 ;
  assign n53014 = n53012 & ~n53013 ;
  assign n53015 = ~x56 & ~n53014 ;
  assign n53016 = ~x56 & ~n53015 ;
  assign n53017 = ~n53014 & ~n53015 ;
  assign n53018 = ~n53016 & ~n53017 ;
  assign n53019 = ~n52878 & ~n52882 ;
  assign n53020 = ~x122 & n22325 ;
  assign n53021 = ~x120 & n23066 ;
  assign n53022 = ~x121 & n22320 ;
  assign n53023 = ~n53021 & ~n53022 ;
  assign n53024 = ~n53020 & n53023 ;
  assign n53025 = n22328 & n22998 ;
  assign n53026 = n53024 & ~n53025 ;
  assign n53027 = ~x59 & ~n53026 ;
  assign n53028 = ~x59 & ~n53027 ;
  assign n53029 = ~n53026 & ~n53027 ;
  assign n53030 = ~n53028 & ~n53029 ;
  assign n53031 = ~n52870 & ~n52874 ;
  assign n53032 = ~x115 & n27427 ;
  assign n53033 = ~x116 & ~n26217 ;
  assign n53034 = ~n53032 & ~n53033 ;
  assign n53035 = ~n52864 & ~n52867 ;
  assign n53036 = ~n53034 & n53035 ;
  assign n53037 = n53034 & ~n53035 ;
  assign n53038 = ~n53036 & ~n53037 ;
  assign n53039 = ~x119 & n24612 ;
  assign n53040 = ~x117 & n25390 ;
  assign n53041 = ~x118 & n24607 ;
  assign n53042 = ~n53040 & ~n53041 ;
  assign n53043 = ~n53039 & n53042 ;
  assign n53044 = n20778 & n24615 ;
  assign n53045 = n53043 & ~n53044 ;
  assign n53046 = ~x62 & ~n53045 ;
  assign n53047 = ~x62 & ~n53046 ;
  assign n53048 = ~n53045 & ~n53046 ;
  assign n53049 = ~n53047 & ~n53048 ;
  assign n53050 = ~n53038 & n53049 ;
  assign n53051 = n53038 & ~n53049 ;
  assign n53052 = ~n53050 & ~n53051 ;
  assign n53053 = ~n53031 & n53052 ;
  assign n53054 = n53031 & ~n53052 ;
  assign n53055 = ~n53053 & ~n53054 ;
  assign n53056 = ~n53030 & n53055 ;
  assign n53057 = n53030 & ~n53055 ;
  assign n53058 = ~n53056 & ~n53057 ;
  assign n53059 = ~n53019 & n53058 ;
  assign n53060 = ~n53019 & ~n53059 ;
  assign n53061 = n53058 & ~n53059 ;
  assign n53062 = ~n53060 & ~n53061 ;
  assign n53063 = ~n53018 & ~n53062 ;
  assign n53064 = n53018 & ~n53061 ;
  assign n53065 = ~n53060 & n53064 ;
  assign n53066 = ~n53063 & ~n53065 ;
  assign n53067 = ~n53007 & n53066 ;
  assign n53068 = n53007 & ~n53066 ;
  assign n53069 = ~n53067 & ~n53068 ;
  assign n53070 = ~x126 & n18764 ;
  assign n53071 = ~x127 & n18020 ;
  assign n53072 = ~n53070 & ~n53071 ;
  assign n53073 = n18028 & ~n27368 ;
  assign n53074 = n53072 & ~n53073 ;
  assign n53075 = ~x53 & ~n53074 ;
  assign n53076 = ~x53 & ~n53075 ;
  assign n53077 = ~n53074 & ~n53075 ;
  assign n53078 = ~n53076 & ~n53077 ;
  assign n53079 = n53069 & ~n53078 ;
  assign n53080 = n53069 & ~n53079 ;
  assign n53081 = ~n53078 & ~n53079 ;
  assign n53082 = ~n53080 & ~n53081 ;
  assign n53083 = ~n52903 & ~n52909 ;
  assign n53084 = n53082 & n53083 ;
  assign n53085 = ~n53082 & ~n53083 ;
  assign n53086 = ~n53084 & ~n53085 ;
  assign n53087 = ~n52913 & ~n52916 ;
  assign n53088 = n53086 & ~n53087 ;
  assign n53089 = ~n53086 & n53087 ;
  assign n53090 = ~n53088 & ~n53089 ;
  assign n53093 = ~n53090 & ~x243 ;
  assign n53094 = ~n53092 & ~n53093 ;
  assign n53095 = ~n52969 & ~n52972 ;
  assign n53096 = ~n52953 & ~n52967 ;
  assign n53097 = x116 & n27024 ;
  assign n53098 = x117 & ~n26217 ;
  assign n53099 = ~n53097 & ~n53098 ;
  assign n53100 = n52950 & ~n53099 ;
  assign n53101 = ~n52950 & n53099 ;
  assign n53102 = ~n53096 & ~n53101 ;
  assign n53103 = ~n53100 & n53102 ;
  assign n53104 = ~n53096 & ~n53103 ;
  assign n53105 = ~n53101 & ~n53103 ;
  assign n53106 = ~n53100 & n53105 ;
  assign n53107 = ~n53104 & ~n53106 ;
  assign n53108 = x120 & n24612 ;
  assign n53109 = x118 & n25390 ;
  assign n53110 = x119 & n24607 ;
  assign n53111 = ~n53109 & ~n53110 ;
  assign n53112 = ~n53108 & n53111 ;
  assign n53113 = n21143 & n24615 ;
  assign n53114 = n53112 & ~n53113 ;
  assign n53115 = x62 & ~n53114 ;
  assign n53116 = x62 & ~n53115 ;
  assign n53117 = ~n53114 & ~n53115 ;
  assign n53118 = ~n53116 & ~n53117 ;
  assign n53119 = ~n53107 & n53118 ;
  assign n53120 = n53107 & ~n53118 ;
  assign n53121 = ~n53119 & ~n53120 ;
  assign n53122 = x123 & n22325 ;
  assign n53123 = x121 & n23066 ;
  assign n53124 = x122 & n22320 ;
  assign n53125 = ~n53123 & ~n53124 ;
  assign n53126 = ~n53122 & n53125 ;
  assign n53127 = n22328 & n23382 ;
  assign n53128 = n53126 & ~n53127 ;
  assign n53129 = x59 & ~n53128 ;
  assign n53130 = x59 & ~n53129 ;
  assign n53131 = ~n53128 & ~n53129 ;
  assign n53132 = ~n53130 & ~n53131 ;
  assign n53133 = ~n53121 & ~n53132 ;
  assign n53134 = n53121 & n53132 ;
  assign n53135 = ~n53133 & ~n53134 ;
  assign n53136 = n53095 & ~n53135 ;
  assign n53137 = ~n53095 & n53135 ;
  assign n53138 = ~n53136 & ~n53137 ;
  assign n53139 = x126 & n20143 ;
  assign n53140 = x124 & n20854 ;
  assign n53141 = x125 & n20138 ;
  assign n53142 = ~n53140 & ~n53141 ;
  assign n53143 = ~n53139 & n53142 ;
  assign n53144 = n20146 & n25735 ;
  assign n53145 = n53143 & ~n53144 ;
  assign n53146 = x56 & ~n53145 ;
  assign n53147 = x56 & ~n53146 ;
  assign n53148 = ~n53145 & ~n53146 ;
  assign n53149 = ~n53147 & ~n53148 ;
  assign n53150 = n53138 & ~n53149 ;
  assign n53151 = n53138 & ~n53150 ;
  assign n53152 = ~n53149 & ~n53150 ;
  assign n53153 = ~n53151 & ~n53152 ;
  assign n53154 = ~n52975 & ~n52979 ;
  assign n53155 = x127 & n18764 ;
  assign n53156 = ~n18028 & ~n53155 ;
  assign n53157 = ~n26962 & ~n53155 ;
  assign n53158 = ~n53156 & ~n53157 ;
  assign n53159 = x53 & ~n53158 ;
  assign n53160 = ~x53 & n53158 ;
  assign n53161 = ~n53159 & ~n53160 ;
  assign n53162 = ~n53154 & ~n53161 ;
  assign n53163 = n53154 & n53161 ;
  assign n53164 = ~n53162 & ~n53163 ;
  assign n53165 = ~n53153 & n53164 ;
  assign n53166 = ~n53153 & ~n53165 ;
  assign n53167 = n53164 & ~n53165 ;
  assign n53168 = ~n53166 & ~n53167 ;
  assign n53169 = ~n52983 & ~n52995 ;
  assign n53170 = n53168 & n53169 ;
  assign n53171 = ~n53168 & ~n53169 ;
  assign n53172 = ~n53170 & ~n53171 ;
  assign n53173 = ~n53001 & ~n53004 ;
  assign n53174 = n53172 & ~n53173 ;
  assign n53175 = ~n53172 & n53173 ;
  assign n53176 = ~n53174 & ~n53175 ;
  assign n53260 = n53176 & x244 ;
  assign n53177 = ~n53053 & ~n53056 ;
  assign n53178 = ~n53037 & ~n53051 ;
  assign n53179 = ~x116 & n27427 ;
  assign n53180 = ~x117 & ~n26217 ;
  assign n53181 = ~n53179 & ~n53180 ;
  assign n53182 = n53034 & ~n53181 ;
  assign n53183 = ~n53034 & n53181 ;
  assign n53184 = ~n53178 & ~n53183 ;
  assign n53185 = ~n53182 & n53184 ;
  assign n53186 = ~n53178 & ~n53185 ;
  assign n53187 = ~n53183 & ~n53185 ;
  assign n53188 = ~n53182 & n53187 ;
  assign n53189 = ~n53186 & ~n53188 ;
  assign n53190 = ~x120 & n24612 ;
  assign n53191 = ~x118 & n25390 ;
  assign n53192 = ~x119 & n24607 ;
  assign n53193 = ~n53191 & ~n53192 ;
  assign n53194 = ~n53190 & n53193 ;
  assign n53195 = n21501 & n24615 ;
  assign n53196 = n53194 & ~n53195 ;
  assign n53197 = ~x62 & ~n53196 ;
  assign n53198 = ~x62 & ~n53197 ;
  assign n53199 = ~n53196 & ~n53197 ;
  assign n53200 = ~n53198 & ~n53199 ;
  assign n53201 = ~n53189 & n53200 ;
  assign n53202 = n53189 & ~n53200 ;
  assign n53203 = ~n53201 & ~n53202 ;
  assign n53204 = ~x123 & n22325 ;
  assign n53205 = ~x121 & n23066 ;
  assign n53206 = ~x122 & n22320 ;
  assign n53207 = ~n53205 & ~n53206 ;
  assign n53208 = ~n53204 & n53207 ;
  assign n53209 = n22328 & n23760 ;
  assign n53210 = n53208 & ~n53209 ;
  assign n53211 = ~x59 & ~n53210 ;
  assign n53212 = ~x59 & ~n53211 ;
  assign n53213 = ~n53210 & ~n53211 ;
  assign n53214 = ~n53212 & ~n53213 ;
  assign n53215 = ~n53203 & ~n53214 ;
  assign n53216 = n53203 & n53214 ;
  assign n53217 = ~n53215 & ~n53216 ;
  assign n53218 = n53177 & ~n53217 ;
  assign n53219 = ~n53177 & n53217 ;
  assign n53220 = ~n53218 & ~n53219 ;
  assign n53221 = ~x126 & n20143 ;
  assign n53222 = ~x124 & n20854 ;
  assign n53223 = ~x125 & n20138 ;
  assign n53224 = ~n53222 & ~n53223 ;
  assign n53225 = ~n53221 & n53224 ;
  assign n53226 = n20146 & n26128 ;
  assign n53227 = n53225 & ~n53226 ;
  assign n53228 = ~x56 & ~n53227 ;
  assign n53229 = ~x56 & ~n53228 ;
  assign n53230 = ~n53227 & ~n53228 ;
  assign n53231 = ~n53229 & ~n53230 ;
  assign n53232 = n53220 & ~n53231 ;
  assign n53233 = n53220 & ~n53232 ;
  assign n53234 = ~n53231 & ~n53232 ;
  assign n53235 = ~n53233 & ~n53234 ;
  assign n53236 = ~n53059 & ~n53063 ;
  assign n53237 = ~x127 & n18764 ;
  assign n53238 = ~n18028 & ~n53237 ;
  assign n53239 = ~n27365 & ~n53237 ;
  assign n53240 = ~n53238 & ~n53239 ;
  assign n53241 = ~x53 & ~n53240 ;
  assign n53242 = x53 & n53240 ;
  assign n53243 = ~n53241 & ~n53242 ;
  assign n53244 = ~n53236 & ~n53243 ;
  assign n53245 = n53236 & n53243 ;
  assign n53246 = ~n53244 & ~n53245 ;
  assign n53247 = ~n53235 & n53246 ;
  assign n53248 = ~n53235 & ~n53247 ;
  assign n53249 = n53246 & ~n53247 ;
  assign n53250 = ~n53248 & ~n53249 ;
  assign n53251 = ~n53067 & ~n53079 ;
  assign n53252 = n53250 & n53251 ;
  assign n53253 = ~n53250 & ~n53251 ;
  assign n53254 = ~n53252 & ~n53253 ;
  assign n53255 = ~n53085 & ~n53088 ;
  assign n53256 = n53254 & ~n53255 ;
  assign n53257 = ~n53254 & n53255 ;
  assign n53258 = ~n53256 & ~n53257 ;
  assign n53261 = ~n53258 & ~x244 ;
  assign n53262 = ~n53260 & ~n53261 ;
  assign n53263 = ~n53171 & ~n53174 ;
  assign n53264 = ~n53162 & ~n53165 ;
  assign n53265 = ~n53137 & ~n53150 ;
  assign n53266 = x127 & n20143 ;
  assign n53267 = x125 & n20854 ;
  assign n53268 = x126 & n20138 ;
  assign n53269 = ~n53267 & ~n53268 ;
  assign n53270 = ~n53266 & n53269 ;
  assign n53271 = n20146 & n26533 ;
  assign n53272 = n53270 & ~n53271 ;
  assign n53273 = x56 & ~n53272 ;
  assign n53274 = x56 & ~n53273 ;
  assign n53275 = ~n53272 & ~n53273 ;
  assign n53276 = ~n53274 & ~n53275 ;
  assign n53277 = ~n53265 & ~n53276 ;
  assign n53278 = ~n53265 & ~n53277 ;
  assign n53279 = ~n53276 & ~n53277 ;
  assign n53280 = ~n53278 & ~n53279 ;
  assign n53281 = ~n53107 & ~n53118 ;
  assign n53282 = ~n53133 & ~n53281 ;
  assign n53283 = x124 & n22325 ;
  assign n53284 = x122 & n23066 ;
  assign n53285 = x123 & n22320 ;
  assign n53286 = ~n53284 & ~n53285 ;
  assign n53287 = ~n53283 & n53286 ;
  assign n53288 = n22328 & n23796 ;
  assign n53289 = n53287 & ~n53288 ;
  assign n53290 = x59 & ~n53289 ;
  assign n53291 = x59 & ~n53290 ;
  assign n53292 = ~n53289 & ~n53290 ;
  assign n53293 = ~n53291 & ~n53292 ;
  assign n53294 = x53 & ~n53099 ;
  assign n53295 = ~x53 & n53099 ;
  assign n53296 = ~n53294 & ~n53295 ;
  assign n53297 = x117 & n27024 ;
  assign n53298 = x118 & ~n26217 ;
  assign n53299 = ~n53297 & ~n53298 ;
  assign n53300 = n53296 & n53299 ;
  assign n53301 = ~n53296 & ~n53299 ;
  assign n53302 = ~n53300 & ~n53301 ;
  assign n53303 = x121 & n24612 ;
  assign n53304 = x119 & n25390 ;
  assign n53305 = x120 & n24607 ;
  assign n53306 = ~n53304 & ~n53305 ;
  assign n53307 = ~n53303 & n53306 ;
  assign n53308 = n21870 & n24615 ;
  assign n53309 = n53307 & ~n53308 ;
  assign n53310 = x62 & ~n53309 ;
  assign n53311 = x62 & ~n53310 ;
  assign n53312 = ~n53309 & ~n53310 ;
  assign n53313 = ~n53311 & ~n53312 ;
  assign n53314 = n53302 & ~n53313 ;
  assign n53315 = n53302 & ~n53314 ;
  assign n53316 = ~n53313 & ~n53314 ;
  assign n53317 = ~n53315 & ~n53316 ;
  assign n53318 = ~n53105 & ~n53317 ;
  assign n53319 = n53105 & n53317 ;
  assign n53320 = ~n53318 & ~n53319 ;
  assign n53321 = ~n53293 & n53320 ;
  assign n53322 = ~n53293 & ~n53321 ;
  assign n53323 = n53320 & ~n53321 ;
  assign n53324 = ~n53322 & ~n53323 ;
  assign n53325 = ~n53282 & ~n53324 ;
  assign n53326 = ~n53282 & ~n53325 ;
  assign n53327 = ~n53324 & ~n53325 ;
  assign n53328 = ~n53326 & ~n53327 ;
  assign n53329 = ~n53280 & n53328 ;
  assign n53330 = n53280 & ~n53328 ;
  assign n53331 = ~n53329 & ~n53330 ;
  assign n53332 = ~n53264 & ~n53331 ;
  assign n53333 = n53264 & n53331 ;
  assign n53334 = ~n53332 & ~n53333 ;
  assign n53335 = ~n53263 & n53334 ;
  assign n53336 = n53263 & ~n53334 ;
  assign n53337 = ~n53335 & ~n53336 ;
  assign n53414 = n53337 & x245 ;
  assign n53338 = ~n53253 & ~n53256 ;
  assign n53339 = ~n53244 & ~n53247 ;
  assign n53340 = ~n53219 & ~n53232 ;
  assign n53341 = ~x127 & n20143 ;
  assign n53342 = ~x125 & n20854 ;
  assign n53343 = ~x126 & n20138 ;
  assign n53344 = ~n53342 & ~n53343 ;
  assign n53345 = ~n53341 & n53344 ;
  assign n53346 = n20146 & n26932 ;
  assign n53347 = n53345 & ~n53346 ;
  assign n53348 = ~x56 & ~n53347 ;
  assign n53349 = ~x56 & ~n53348 ;
  assign n53350 = ~n53347 & ~n53348 ;
  assign n53351 = ~n53349 & ~n53350 ;
  assign n53352 = ~n53340 & ~n53351 ;
  assign n53353 = ~n53340 & ~n53352 ;
  assign n53354 = ~n53351 & ~n53352 ;
  assign n53355 = ~n53353 & ~n53354 ;
  assign n53356 = ~n53189 & ~n53200 ;
  assign n53357 = ~n53215 & ~n53356 ;
  assign n53358 = ~x124 & n22325 ;
  assign n53359 = ~x122 & n23066 ;
  assign n53360 = ~x123 & n22320 ;
  assign n53361 = ~n53359 & ~n53360 ;
  assign n53362 = ~n53358 & n53361 ;
  assign n53363 = n22328 & n24176 ;
  assign n53364 = n53362 & ~n53363 ;
  assign n53365 = ~x59 & ~n53364 ;
  assign n53366 = ~x59 & ~n53365 ;
  assign n53367 = ~n53364 & ~n53365 ;
  assign n53368 = ~n53366 & ~n53367 ;
  assign n53369 = ~x53 & ~n53181 ;
  assign n53370 = x53 & n53181 ;
  assign n53371 = ~n53369 & ~n53370 ;
  assign n53372 = ~x117 & n27427 ;
  assign n53373 = ~x118 & ~n26217 ;
  assign n53374 = ~n53372 & ~n53373 ;
  assign n53375 = n53371 & n53374 ;
  assign n53376 = ~n53371 & ~n53374 ;
  assign n53377 = ~n53375 & ~n53376 ;
  assign n53378 = ~x121 & n24612 ;
  assign n53379 = ~x119 & n25390 ;
  assign n53380 = ~x120 & n24607 ;
  assign n53381 = ~n53379 & ~n53380 ;
  assign n53382 = ~n53378 & n53381 ;
  assign n53383 = n22229 & n24615 ;
  assign n53384 = n53382 & ~n53383 ;
  assign n53385 = ~x62 & ~n53384 ;
  assign n53386 = ~x62 & ~n53385 ;
  assign n53387 = ~n53384 & ~n53385 ;
  assign n53388 = ~n53386 & ~n53387 ;
  assign n53389 = n53377 & ~n53388 ;
  assign n53390 = n53377 & ~n53389 ;
  assign n53391 = ~n53388 & ~n53389 ;
  assign n53392 = ~n53390 & ~n53391 ;
  assign n53393 = ~n53187 & ~n53392 ;
  assign n53394 = n53187 & n53392 ;
  assign n53395 = ~n53393 & ~n53394 ;
  assign n53396 = ~n53368 & n53395 ;
  assign n53397 = ~n53368 & ~n53396 ;
  assign n53398 = n53395 & ~n53396 ;
  assign n53399 = ~n53397 & ~n53398 ;
  assign n53400 = ~n53357 & ~n53399 ;
  assign n53401 = ~n53357 & ~n53400 ;
  assign n53402 = ~n53399 & ~n53400 ;
  assign n53403 = ~n53401 & ~n53402 ;
  assign n53404 = ~n53355 & n53403 ;
  assign n53405 = n53355 & ~n53403 ;
  assign n53406 = ~n53404 & ~n53405 ;
  assign n53407 = ~n53339 & ~n53406 ;
  assign n53408 = n53339 & n53406 ;
  assign n53409 = ~n53407 & ~n53408 ;
  assign n53410 = ~n53338 & n53409 ;
  assign n53411 = n53338 & ~n53409 ;
  assign n53412 = ~n53410 & ~n53411 ;
  assign n53415 = ~n53412 & ~x245 ;
  assign n53416 = ~n53414 & ~n53415 ;
  assign n53417 = ~n53321 & ~n53325 ;
  assign n53418 = x125 & n22325 ;
  assign n53419 = x123 & n23066 ;
  assign n53420 = x124 & n22320 ;
  assign n53421 = ~n53419 & ~n53420 ;
  assign n53422 = ~n53418 & n53421 ;
  assign n53423 = n22328 & n24935 ;
  assign n53424 = n53422 & ~n53423 ;
  assign n53425 = x59 & ~n53424 ;
  assign n53426 = x59 & ~n53425 ;
  assign n53427 = ~n53424 & ~n53425 ;
  assign n53428 = ~n53426 & ~n53427 ;
  assign n53429 = ~n53314 & ~n53318 ;
  assign n53430 = x118 & n27024 ;
  assign n53431 = x119 & ~n26217 ;
  assign n53432 = ~n53430 & ~n53431 ;
  assign n53433 = ~x53 & ~n53099 ;
  assign n53434 = ~n53301 & ~n53433 ;
  assign n53435 = n53432 & ~n53434 ;
  assign n53436 = ~n53432 & n53434 ;
  assign n53437 = ~n53435 & ~n53436 ;
  assign n53438 = x122 & n24612 ;
  assign n53439 = x120 & n25390 ;
  assign n53440 = x121 & n24607 ;
  assign n53441 = ~n53439 & ~n53440 ;
  assign n53442 = ~n53438 & n53441 ;
  assign n53443 = ~n24615 & n53442 ;
  assign n53444 = ~n22622 & n53442 ;
  assign n53445 = ~n53443 & ~n53444 ;
  assign n53446 = x62 & ~n53445 ;
  assign n53447 = ~x62 & n53445 ;
  assign n53448 = ~n53446 & ~n53447 ;
  assign n53449 = n53437 & ~n53448 ;
  assign n53450 = ~n53437 & n53448 ;
  assign n53451 = ~n53449 & ~n53450 ;
  assign n53452 = ~n53429 & n53451 ;
  assign n53453 = ~n53429 & ~n53452 ;
  assign n53454 = n53451 & ~n53452 ;
  assign n53455 = ~n53453 & ~n53454 ;
  assign n53456 = ~n53428 & ~n53455 ;
  assign n53457 = n53428 & ~n53454 ;
  assign n53458 = ~n53453 & n53457 ;
  assign n53459 = ~n53456 & ~n53458 ;
  assign n53460 = ~n53417 & n53459 ;
  assign n53461 = n53417 & ~n53459 ;
  assign n53462 = ~n53460 & ~n53461 ;
  assign n53463 = x126 & n20854 ;
  assign n53464 = x127 & n20138 ;
  assign n53465 = ~n53463 & ~n53464 ;
  assign n53466 = n20146 & ~n26965 ;
  assign n53467 = n53465 & ~n53466 ;
  assign n53468 = x56 & ~n53467 ;
  assign n53469 = x56 & ~n53468 ;
  assign n53470 = ~n53467 & ~n53468 ;
  assign n53471 = ~n53469 & ~n53470 ;
  assign n53472 = n53462 & ~n53471 ;
  assign n53473 = n53462 & ~n53472 ;
  assign n53474 = ~n53471 & ~n53472 ;
  assign n53475 = ~n53473 & ~n53474 ;
  assign n53476 = ~n53280 & ~n53328 ;
  assign n53477 = ~n53277 & ~n53476 ;
  assign n53478 = ~n53475 & ~n53477 ;
  assign n53479 = ~n53475 & ~n53478 ;
  assign n53480 = ~n53477 & ~n53478 ;
  assign n53481 = ~n53479 & ~n53480 ;
  assign n53482 = ~n53332 & ~n53335 ;
  assign n53483 = ~n53481 & ~n53482 ;
  assign n53484 = n53481 & n53482 ;
  assign n53485 = ~n53483 & ~n53484 ;
  assign n53556 = n53485 & x246 ;
  assign n53486 = ~n53396 & ~n53400 ;
  assign n53487 = ~x125 & n22325 ;
  assign n53488 = ~x123 & n23066 ;
  assign n53489 = ~x124 & n22320 ;
  assign n53490 = ~n53488 & ~n53489 ;
  assign n53491 = ~n53487 & n53490 ;
  assign n53492 = n22328 & n25330 ;
  assign n53493 = n53491 & ~n53492 ;
  assign n53494 = ~x59 & ~n53493 ;
  assign n53495 = ~x59 & ~n53494 ;
  assign n53496 = ~n53493 & ~n53494 ;
  assign n53497 = ~n53495 & ~n53496 ;
  assign n53498 = ~n53389 & ~n53393 ;
  assign n53499 = ~x118 & n27427 ;
  assign n53500 = ~x119 & ~n26217 ;
  assign n53501 = ~n53499 & ~n53500 ;
  assign n53502 = x53 & ~n53181 ;
  assign n53503 = ~n53376 & ~n53502 ;
  assign n53504 = n53501 & ~n53503 ;
  assign n53505 = ~n53501 & n53503 ;
  assign n53506 = ~n53504 & ~n53505 ;
  assign n53507 = ~x122 & n24612 ;
  assign n53508 = ~x120 & n25390 ;
  assign n53509 = ~x121 & n24607 ;
  assign n53510 = ~n53508 & ~n53509 ;
  assign n53511 = ~n53507 & n53510 ;
  assign n53512 = ~n24615 & n53511 ;
  assign n53513 = ~n22998 & n53511 ;
  assign n53514 = ~n53512 & ~n53513 ;
  assign n53515 = ~x62 & ~n53514 ;
  assign n53516 = x62 & n53514 ;
  assign n53517 = ~n53515 & ~n53516 ;
  assign n53518 = n53506 & ~n53517 ;
  assign n53519 = ~n53506 & n53517 ;
  assign n53520 = ~n53518 & ~n53519 ;
  assign n53521 = ~n53498 & n53520 ;
  assign n53522 = ~n53498 & ~n53521 ;
  assign n53523 = n53520 & ~n53521 ;
  assign n53524 = ~n53522 & ~n53523 ;
  assign n53525 = ~n53497 & ~n53524 ;
  assign n53526 = n53497 & ~n53523 ;
  assign n53527 = ~n53522 & n53526 ;
  assign n53528 = ~n53525 & ~n53527 ;
  assign n53529 = ~n53486 & n53528 ;
  assign n53530 = n53486 & ~n53528 ;
  assign n53531 = ~n53529 & ~n53530 ;
  assign n53532 = ~x126 & n20854 ;
  assign n53533 = ~x127 & n20138 ;
  assign n53534 = ~n53532 & ~n53533 ;
  assign n53535 = n20146 & ~n27368 ;
  assign n53536 = n53534 & ~n53535 ;
  assign n53537 = ~x56 & ~n53536 ;
  assign n53538 = ~x56 & ~n53537 ;
  assign n53539 = ~n53536 & ~n53537 ;
  assign n53540 = ~n53538 & ~n53539 ;
  assign n53541 = n53531 & ~n53540 ;
  assign n53542 = n53531 & ~n53541 ;
  assign n53543 = ~n53540 & ~n53541 ;
  assign n53544 = ~n53542 & ~n53543 ;
  assign n53545 = ~n53355 & ~n53403 ;
  assign n53546 = ~n53352 & ~n53545 ;
  assign n53547 = ~n53544 & ~n53546 ;
  assign n53548 = ~n53544 & ~n53547 ;
  assign n53549 = ~n53546 & ~n53547 ;
  assign n53550 = ~n53548 & ~n53549 ;
  assign n53551 = ~n53407 & ~n53410 ;
  assign n53552 = ~n53550 & ~n53551 ;
  assign n53553 = n53550 & n53551 ;
  assign n53554 = ~n53552 & ~n53553 ;
  assign n53557 = ~n53554 & ~x246 ;
  assign n53558 = ~n53556 & ~n53557 ;
  assign n53559 = x123 & n24612 ;
  assign n53560 = x121 & n25390 ;
  assign n53561 = x122 & n24607 ;
  assign n53562 = ~n53560 & ~n53561 ;
  assign n53563 = ~n53559 & n53562 ;
  assign n53564 = n23382 & n24615 ;
  assign n53565 = n53563 & ~n53564 ;
  assign n53566 = x62 & ~n53565 ;
  assign n53567 = x62 & ~n53566 ;
  assign n53568 = ~n53565 & ~n53566 ;
  assign n53569 = ~n53567 & ~n53568 ;
  assign n53570 = x119 & n27024 ;
  assign n53571 = x120 & ~n26217 ;
  assign n53572 = ~n53570 & ~n53571 ;
  assign n53573 = n53432 & ~n53572 ;
  assign n53574 = n53432 & ~n53573 ;
  assign n53575 = ~n53572 & ~n53573 ;
  assign n53576 = ~n53574 & ~n53575 ;
  assign n53577 = ~n53569 & ~n53576 ;
  assign n53578 = ~n53569 & ~n53577 ;
  assign n53579 = ~n53576 & ~n53577 ;
  assign n53580 = ~n53578 & ~n53579 ;
  assign n53581 = ~n53435 & ~n53449 ;
  assign n53582 = n53580 & n53581 ;
  assign n53583 = ~n53580 & ~n53581 ;
  assign n53584 = ~n53582 & ~n53583 ;
  assign n53585 = x126 & n22325 ;
  assign n53586 = x124 & n23066 ;
  assign n53587 = x125 & n22320 ;
  assign n53588 = ~n53586 & ~n53587 ;
  assign n53589 = ~n53585 & n53588 ;
  assign n53590 = n22328 & n25735 ;
  assign n53591 = n53589 & ~n53590 ;
  assign n53592 = x59 & ~n53591 ;
  assign n53593 = x59 & ~n53592 ;
  assign n53594 = ~n53591 & ~n53592 ;
  assign n53595 = ~n53593 & ~n53594 ;
  assign n53596 = n53584 & ~n53595 ;
  assign n53597 = n53584 & ~n53596 ;
  assign n53598 = ~n53595 & ~n53596 ;
  assign n53599 = ~n53597 & ~n53598 ;
  assign n53600 = ~n53452 & ~n53456 ;
  assign n53601 = x127 & n20854 ;
  assign n53602 = ~n20146 & ~n53601 ;
  assign n53603 = ~n26962 & ~n53601 ;
  assign n53604 = ~n53602 & ~n53603 ;
  assign n53605 = x56 & ~n53604 ;
  assign n53606 = ~x56 & n53604 ;
  assign n53607 = ~n53605 & ~n53606 ;
  assign n53608 = ~n53600 & ~n53607 ;
  assign n53609 = n53600 & n53607 ;
  assign n53610 = ~n53608 & ~n53609 ;
  assign n53611 = ~n53599 & n53610 ;
  assign n53612 = ~n53599 & ~n53611 ;
  assign n53613 = n53610 & ~n53611 ;
  assign n53614 = ~n53612 & ~n53613 ;
  assign n53615 = ~n53460 & ~n53472 ;
  assign n53616 = n53614 & n53615 ;
  assign n53617 = ~n53614 & ~n53615 ;
  assign n53618 = ~n53616 & ~n53617 ;
  assign n53619 = ~n53478 & ~n53483 ;
  assign n53620 = n53618 & ~n53619 ;
  assign n53621 = ~n53618 & n53619 ;
  assign n53622 = ~n53620 & ~n53621 ;
  assign n53688 = n53622 & x247 ;
  assign n53623 = ~x123 & n24612 ;
  assign n53624 = ~x121 & n25390 ;
  assign n53625 = ~x122 & n24607 ;
  assign n53626 = ~n53624 & ~n53625 ;
  assign n53627 = ~n53623 & n53626 ;
  assign n53628 = n23760 & n24615 ;
  assign n53629 = n53627 & ~n53628 ;
  assign n53630 = ~x62 & ~n53629 ;
  assign n53631 = ~x62 & ~n53630 ;
  assign n53632 = ~n53629 & ~n53630 ;
  assign n53633 = ~n53631 & ~n53632 ;
  assign n53634 = ~x119 & n27427 ;
  assign n53635 = ~x120 & ~n26217 ;
  assign n53636 = ~n53634 & ~n53635 ;
  assign n53637 = n53501 & ~n53636 ;
  assign n53638 = n53501 & ~n53637 ;
  assign n53639 = ~n53636 & ~n53637 ;
  assign n53640 = ~n53638 & ~n53639 ;
  assign n53641 = ~n53633 & ~n53640 ;
  assign n53642 = ~n53633 & ~n53641 ;
  assign n53643 = ~n53640 & ~n53641 ;
  assign n53644 = ~n53642 & ~n53643 ;
  assign n53645 = ~n53504 & ~n53518 ;
  assign n53646 = n53644 & n53645 ;
  assign n53647 = ~n53644 & ~n53645 ;
  assign n53648 = ~n53646 & ~n53647 ;
  assign n53649 = ~x126 & n22325 ;
  assign n53650 = ~x124 & n23066 ;
  assign n53651 = ~x125 & n22320 ;
  assign n53652 = ~n53650 & ~n53651 ;
  assign n53653 = ~n53649 & n53652 ;
  assign n53654 = n22328 & n26128 ;
  assign n53655 = n53653 & ~n53654 ;
  assign n53656 = ~x59 & ~n53655 ;
  assign n53657 = ~x59 & ~n53656 ;
  assign n53658 = ~n53655 & ~n53656 ;
  assign n53659 = ~n53657 & ~n53658 ;
  assign n53660 = n53648 & ~n53659 ;
  assign n53661 = n53648 & ~n53660 ;
  assign n53662 = ~n53659 & ~n53660 ;
  assign n53663 = ~n53661 & ~n53662 ;
  assign n53664 = ~n53521 & ~n53525 ;
  assign n53665 = ~x127 & n20854 ;
  assign n53666 = ~n20146 & ~n53665 ;
  assign n53667 = ~n27365 & ~n53665 ;
  assign n53668 = ~n53666 & ~n53667 ;
  assign n53669 = ~x56 & ~n53668 ;
  assign n53670 = x56 & n53668 ;
  assign n53671 = ~n53669 & ~n53670 ;
  assign n53672 = ~n53664 & ~n53671 ;
  assign n53673 = n53664 & n53671 ;
  assign n53674 = ~n53672 & ~n53673 ;
  assign n53675 = ~n53663 & n53674 ;
  assign n53676 = ~n53663 & ~n53675 ;
  assign n53677 = n53674 & ~n53675 ;
  assign n53678 = ~n53676 & ~n53677 ;
  assign n53679 = ~n53529 & ~n53541 ;
  assign n53680 = n53678 & n53679 ;
  assign n53681 = ~n53678 & ~n53679 ;
  assign n53682 = ~n53680 & ~n53681 ;
  assign n53683 = ~n53547 & ~n53552 ;
  assign n53684 = n53682 & ~n53683 ;
  assign n53685 = ~n53682 & n53683 ;
  assign n53686 = ~n53684 & ~n53685 ;
  assign n53689 = ~n53686 & ~x247 ;
  assign n53690 = ~n53688 & ~n53689 ;
  assign n53691 = ~n53583 & ~n53596 ;
  assign n53692 = x127 & n22325 ;
  assign n53693 = x125 & n23066 ;
  assign n53694 = x126 & n22320 ;
  assign n53695 = ~n53693 & ~n53694 ;
  assign n53696 = ~n53692 & n53695 ;
  assign n53697 = n22328 & n26533 ;
  assign n53698 = n53696 & ~n53697 ;
  assign n53699 = x59 & ~n53698 ;
  assign n53700 = x59 & ~n53699 ;
  assign n53701 = ~n53698 & ~n53699 ;
  assign n53702 = ~n53700 & ~n53701 ;
  assign n53703 = ~n53691 & ~n53702 ;
  assign n53704 = ~n53691 & ~n53703 ;
  assign n53705 = ~n53702 & ~n53703 ;
  assign n53706 = ~n53704 & ~n53705 ;
  assign n53707 = x120 & n27024 ;
  assign n53708 = x121 & ~n26217 ;
  assign n53709 = ~n53707 & ~n53708 ;
  assign n53710 = ~x56 & ~n53709 ;
  assign n53711 = ~x56 & ~n53710 ;
  assign n53712 = ~n53709 & ~n53710 ;
  assign n53713 = ~n53711 & ~n53712 ;
  assign n53714 = ~n53432 & ~n53713 ;
  assign n53715 = ~n53432 & ~n53714 ;
  assign n53716 = ~n53713 & ~n53714 ;
  assign n53717 = ~n53715 & ~n53716 ;
  assign n53718 = ~n53573 & ~n53577 ;
  assign n53719 = n53717 & n53718 ;
  assign n53720 = ~n53717 & ~n53718 ;
  assign n53721 = ~n53719 & ~n53720 ;
  assign n53722 = x124 & n24612 ;
  assign n53723 = x122 & n25390 ;
  assign n53724 = x123 & n24607 ;
  assign n53725 = ~n53723 & ~n53724 ;
  assign n53726 = ~n53722 & n53725 ;
  assign n53727 = n23796 & n24615 ;
  assign n53728 = n53726 & ~n53727 ;
  assign n53729 = x62 & ~n53728 ;
  assign n53730 = x62 & ~n53729 ;
  assign n53731 = ~n53728 & ~n53729 ;
  assign n53732 = ~n53730 & ~n53731 ;
  assign n53733 = n53721 & ~n53732 ;
  assign n53734 = ~n53721 & n53732 ;
  assign n53735 = ~n53706 & ~n53734 ;
  assign n53736 = ~n53733 & n53735 ;
  assign n53737 = ~n53706 & ~n53736 ;
  assign n53738 = ~n53734 & ~n53736 ;
  assign n53739 = ~n53733 & n53738 ;
  assign n53740 = ~n53737 & ~n53739 ;
  assign n53741 = ~n53608 & ~n53611 ;
  assign n53742 = n53740 & n53741 ;
  assign n53743 = ~n53740 & ~n53741 ;
  assign n53744 = ~n53742 & ~n53743 ;
  assign n53745 = ~n53617 & ~n53620 ;
  assign n53746 = n53744 & ~n53745 ;
  assign n53747 = ~n53744 & n53745 ;
  assign n53748 = ~n53746 & ~n53747 ;
  assign n53808 = n53748 & x248 ;
  assign n53749 = ~n53647 & ~n53660 ;
  assign n53750 = ~x127 & n22325 ;
  assign n53751 = ~x125 & n23066 ;
  assign n53752 = ~x126 & n22320 ;
  assign n53753 = ~n53751 & ~n53752 ;
  assign n53754 = ~n53750 & n53753 ;
  assign n53755 = n22328 & n26932 ;
  assign n53756 = n53754 & ~n53755 ;
  assign n53757 = ~x59 & ~n53756 ;
  assign n53758 = ~x59 & ~n53757 ;
  assign n53759 = ~n53756 & ~n53757 ;
  assign n53760 = ~n53758 & ~n53759 ;
  assign n53761 = ~n53749 & ~n53760 ;
  assign n53762 = ~n53749 & ~n53761 ;
  assign n53763 = ~n53760 & ~n53761 ;
  assign n53764 = ~n53762 & ~n53763 ;
  assign n53765 = ~x120 & n27427 ;
  assign n53766 = ~x121 & ~n26217 ;
  assign n53767 = ~n53765 & ~n53766 ;
  assign n53768 = x56 & ~n53767 ;
  assign n53769 = x56 & ~n53768 ;
  assign n53770 = ~n53767 & ~n53768 ;
  assign n53771 = ~n53769 & ~n53770 ;
  assign n53772 = ~n53501 & ~n53771 ;
  assign n53773 = ~n53501 & ~n53772 ;
  assign n53774 = ~n53771 & ~n53772 ;
  assign n53775 = ~n53773 & ~n53774 ;
  assign n53776 = ~n53637 & ~n53641 ;
  assign n53777 = n53775 & n53776 ;
  assign n53778 = ~n53775 & ~n53776 ;
  assign n53779 = ~n53777 & ~n53778 ;
  assign n53780 = ~x124 & n24612 ;
  assign n53781 = ~x122 & n25390 ;
  assign n53782 = ~x123 & n24607 ;
  assign n53783 = ~n53781 & ~n53782 ;
  assign n53784 = ~n53780 & n53783 ;
  assign n53785 = n24176 & n24615 ;
  assign n53786 = n53784 & ~n53785 ;
  assign n53787 = ~x62 & ~n53786 ;
  assign n53788 = ~x62 & ~n53787 ;
  assign n53789 = ~n53786 & ~n53787 ;
  assign n53790 = ~n53788 & ~n53789 ;
  assign n53791 = n53779 & ~n53790 ;
  assign n53792 = ~n53779 & n53790 ;
  assign n53793 = ~n53764 & ~n53792 ;
  assign n53794 = ~n53791 & n53793 ;
  assign n53795 = ~n53764 & ~n53794 ;
  assign n53796 = ~n53792 & ~n53794 ;
  assign n53797 = ~n53791 & n53796 ;
  assign n53798 = ~n53795 & ~n53797 ;
  assign n53799 = ~n53672 & ~n53675 ;
  assign n53800 = n53798 & n53799 ;
  assign n53801 = ~n53798 & ~n53799 ;
  assign n53802 = ~n53800 & ~n53801 ;
  assign n53803 = ~n53681 & ~n53684 ;
  assign n53804 = n53802 & ~n53803 ;
  assign n53805 = ~n53802 & n53803 ;
  assign n53806 = ~n53804 & ~n53805 ;
  assign n53809 = ~n53806 & ~x248 ;
  assign n53810 = ~n53808 & ~n53809 ;
  assign n53811 = ~n53720 & ~n53733 ;
  assign n53812 = x121 & n27024 ;
  assign n53813 = x122 & ~n26217 ;
  assign n53814 = ~n53812 & ~n53813 ;
  assign n53815 = ~n53710 & ~n53714 ;
  assign n53816 = ~n53814 & n53815 ;
  assign n53817 = n53814 & ~n53815 ;
  assign n53818 = ~n53816 & ~n53817 ;
  assign n53819 = x125 & n24612 ;
  assign n53820 = x123 & n25390 ;
  assign n53821 = x124 & n24607 ;
  assign n53822 = ~n53820 & ~n53821 ;
  assign n53823 = ~n53819 & n53822 ;
  assign n53824 = ~n24615 & n53823 ;
  assign n53825 = ~n24935 & n53823 ;
  assign n53826 = ~n53824 & ~n53825 ;
  assign n53827 = x62 & ~n53826 ;
  assign n53828 = ~x62 & n53826 ;
  assign n53829 = ~n53827 & ~n53828 ;
  assign n53830 = n53818 & ~n53829 ;
  assign n53831 = ~n53818 & n53829 ;
  assign n53832 = ~n53830 & ~n53831 ;
  assign n53833 = ~n53811 & n53832 ;
  assign n53834 = n53811 & ~n53832 ;
  assign n53835 = ~n53833 & ~n53834 ;
  assign n53836 = x126 & n23066 ;
  assign n53837 = x127 & n22320 ;
  assign n53838 = ~n53836 & ~n53837 ;
  assign n53839 = n22328 & ~n26965 ;
  assign n53840 = n53838 & ~n53839 ;
  assign n53841 = x59 & ~n53840 ;
  assign n53842 = x59 & ~n53841 ;
  assign n53843 = ~n53840 & ~n53841 ;
  assign n53844 = ~n53842 & ~n53843 ;
  assign n53845 = n53835 & ~n53844 ;
  assign n53846 = n53835 & ~n53845 ;
  assign n53847 = ~n53844 & ~n53845 ;
  assign n53848 = ~n53846 & ~n53847 ;
  assign n53849 = ~n53703 & ~n53736 ;
  assign n53850 = n53848 & n53849 ;
  assign n53851 = ~n53848 & ~n53849 ;
  assign n53852 = ~n53850 & ~n53851 ;
  assign n53853 = ~n53743 & ~n53746 ;
  assign n53854 = n53852 & ~n53853 ;
  assign n53855 = ~n53852 & n53853 ;
  assign n53856 = ~n53854 & ~n53855 ;
  assign n53904 = n53856 & x249 ;
  assign n53857 = ~n53778 & ~n53791 ;
  assign n53858 = ~x121 & n27427 ;
  assign n53859 = ~x122 & ~n26217 ;
  assign n53860 = ~n53858 & ~n53859 ;
  assign n53861 = ~n53768 & ~n53772 ;
  assign n53862 = ~n53860 & n53861 ;
  assign n53863 = n53860 & ~n53861 ;
  assign n53864 = ~n53862 & ~n53863 ;
  assign n53865 = ~x125 & n24612 ;
  assign n53866 = ~x123 & n25390 ;
  assign n53867 = ~x124 & n24607 ;
  assign n53868 = ~n53866 & ~n53867 ;
  assign n53869 = ~n53865 & n53868 ;
  assign n53870 = ~n24615 & n53869 ;
  assign n53871 = ~n25330 & n53869 ;
  assign n53872 = ~n53870 & ~n53871 ;
  assign n53873 = ~x62 & ~n53872 ;
  assign n53874 = x62 & n53872 ;
  assign n53875 = ~n53873 & ~n53874 ;
  assign n53876 = n53864 & ~n53875 ;
  assign n53877 = ~n53864 & n53875 ;
  assign n53878 = ~n53876 & ~n53877 ;
  assign n53879 = ~n53857 & n53878 ;
  assign n53880 = n53857 & ~n53878 ;
  assign n53881 = ~n53879 & ~n53880 ;
  assign n53882 = ~x126 & n23066 ;
  assign n53883 = ~x127 & n22320 ;
  assign n53884 = ~n53882 & ~n53883 ;
  assign n53885 = n22328 & ~n27368 ;
  assign n53886 = n53884 & ~n53885 ;
  assign n53887 = ~x59 & ~n53886 ;
  assign n53888 = ~x59 & ~n53887 ;
  assign n53889 = ~n53886 & ~n53887 ;
  assign n53890 = ~n53888 & ~n53889 ;
  assign n53891 = n53881 & ~n53890 ;
  assign n53892 = n53881 & ~n53891 ;
  assign n53893 = ~n53890 & ~n53891 ;
  assign n53894 = ~n53892 & ~n53893 ;
  assign n53895 = ~n53761 & ~n53794 ;
  assign n53896 = n53894 & n53895 ;
  assign n53897 = ~n53894 & ~n53895 ;
  assign n53898 = ~n53896 & ~n53897 ;
  assign n53899 = ~n53801 & ~n53804 ;
  assign n53900 = n53898 & ~n53899 ;
  assign n53901 = ~n53898 & n53899 ;
  assign n53902 = ~n53900 & ~n53901 ;
  assign n53905 = ~n53902 & ~x249 ;
  assign n53906 = ~n53904 & ~n53905 ;
  assign n53907 = ~n53851 & ~n53854 ;
  assign n53908 = ~n53833 & ~n53845 ;
  assign n53909 = ~n53817 & ~n53830 ;
  assign n53910 = x122 & n27024 ;
  assign n53911 = x123 & ~n26217 ;
  assign n53912 = ~n53910 & ~n53911 ;
  assign n53913 = n53814 & ~n53912 ;
  assign n53914 = ~n53814 & n53912 ;
  assign n53915 = ~n53909 & ~n53914 ;
  assign n53916 = ~n53913 & n53915 ;
  assign n53917 = ~n53909 & ~n53916 ;
  assign n53918 = ~n53914 & ~n53916 ;
  assign n53919 = ~n53913 & n53918 ;
  assign n53920 = ~n53917 & ~n53919 ;
  assign n53921 = x126 & n24612 ;
  assign n53922 = x124 & n25390 ;
  assign n53923 = x125 & n24607 ;
  assign n53924 = ~n53922 & ~n53923 ;
  assign n53925 = ~n53921 & n53924 ;
  assign n53926 = n24615 & n25735 ;
  assign n53927 = n53925 & ~n53926 ;
  assign n53928 = x62 & ~n53927 ;
  assign n53929 = x62 & ~n53928 ;
  assign n53930 = ~n53927 & ~n53928 ;
  assign n53931 = ~n53929 & ~n53930 ;
  assign n53932 = x127 & n23066 ;
  assign n53933 = n22328 & n26962 ;
  assign n53934 = ~n53932 & ~n53933 ;
  assign n53935 = x59 & ~n53934 ;
  assign n53936 = x59 & ~n53935 ;
  assign n53937 = ~n53934 & ~n53935 ;
  assign n53938 = ~n53936 & ~n53937 ;
  assign n53939 = ~n53931 & ~n53938 ;
  assign n53940 = ~n53931 & ~n53939 ;
  assign n53941 = ~n53938 & ~n53939 ;
  assign n53942 = ~n53940 & ~n53941 ;
  assign n53943 = ~n53920 & n53942 ;
  assign n53944 = n53920 & ~n53942 ;
  assign n53945 = ~n53943 & ~n53944 ;
  assign n53946 = ~n53908 & ~n53945 ;
  assign n53947 = ~n53908 & ~n53946 ;
  assign n53948 = ~n53945 & ~n53946 ;
  assign n53949 = ~n53947 & ~n53948 ;
  assign n53950 = ~n53907 & ~n53949 ;
  assign n53951 = n53907 & ~n53948 ;
  assign n53952 = ~n53947 & n53951 ;
  assign n53953 = ~n53950 & ~n53952 ;
  assign n54002 = n53953 & x250 ;
  assign n53954 = ~n53897 & ~n53900 ;
  assign n53955 = ~n53879 & ~n53891 ;
  assign n53956 = ~n53863 & ~n53876 ;
  assign n53957 = ~x122 & n27427 ;
  assign n53958 = ~x123 & ~n26217 ;
  assign n53959 = ~n53957 & ~n53958 ;
  assign n53960 = n53860 & ~n53959 ;
  assign n53961 = ~n53860 & n53959 ;
  assign n53962 = ~n53956 & ~n53961 ;
  assign n53963 = ~n53960 & n53962 ;
  assign n53964 = ~n53956 & ~n53963 ;
  assign n53965 = ~n53961 & ~n53963 ;
  assign n53966 = ~n53960 & n53965 ;
  assign n53967 = ~n53964 & ~n53966 ;
  assign n53968 = ~x126 & n24612 ;
  assign n53969 = ~x124 & n25390 ;
  assign n53970 = ~x125 & n24607 ;
  assign n53971 = ~n53969 & ~n53970 ;
  assign n53972 = ~n53968 & n53971 ;
  assign n53973 = n24615 & n26128 ;
  assign n53974 = n53972 & ~n53973 ;
  assign n53975 = ~x62 & ~n53974 ;
  assign n53976 = ~x62 & ~n53975 ;
  assign n53977 = ~n53974 & ~n53975 ;
  assign n53978 = ~n53976 & ~n53977 ;
  assign n53979 = ~x127 & n23066 ;
  assign n53980 = n22328 & n27365 ;
  assign n53981 = ~n53979 & ~n53980 ;
  assign n53982 = ~x59 & ~n53981 ;
  assign n53983 = ~x59 & ~n53982 ;
  assign n53984 = ~n53981 & ~n53982 ;
  assign n53985 = ~n53983 & ~n53984 ;
  assign n53986 = ~n53978 & ~n53985 ;
  assign n53987 = ~n53978 & ~n53986 ;
  assign n53988 = ~n53985 & ~n53986 ;
  assign n53989 = ~n53987 & ~n53988 ;
  assign n53990 = ~n53967 & n53989 ;
  assign n53991 = n53967 & ~n53989 ;
  assign n53992 = ~n53990 & ~n53991 ;
  assign n53993 = ~n53955 & ~n53992 ;
  assign n53994 = ~n53955 & ~n53993 ;
  assign n53995 = ~n53992 & ~n53993 ;
  assign n53996 = ~n53994 & ~n53995 ;
  assign n53997 = ~n53954 & ~n53996 ;
  assign n53998 = n53954 & ~n53995 ;
  assign n53999 = ~n53994 & n53998 ;
  assign n54000 = ~n53997 & ~n53999 ;
  assign n54003 = ~n54000 & ~x250 ;
  assign n54004 = ~n54002 & ~n54003 ;
  assign n54005 = ~n53946 & ~n53950 ;
  assign n54006 = ~n53920 & ~n53942 ;
  assign n54007 = ~n53939 & ~n54006 ;
  assign n54008 = x59 & ~n53912 ;
  assign n54009 = ~x59 & n53912 ;
  assign n54010 = ~n54008 & ~n54009 ;
  assign n54011 = x123 & n27024 ;
  assign n54012 = x124 & ~n26217 ;
  assign n54013 = ~n54011 & ~n54012 ;
  assign n54014 = n54010 & n54013 ;
  assign n54015 = ~n54010 & ~n54013 ;
  assign n54016 = ~n54014 & ~n54015 ;
  assign n54017 = x127 & n24612 ;
  assign n54018 = x125 & n25390 ;
  assign n54019 = x126 & n24607 ;
  assign n54020 = ~n54018 & ~n54019 ;
  assign n54021 = ~n54017 & n54020 ;
  assign n54022 = n24615 & n26533 ;
  assign n54023 = n54021 & ~n54022 ;
  assign n54024 = x62 & ~n54023 ;
  assign n54025 = x62 & ~n54024 ;
  assign n54026 = ~n54023 & ~n54024 ;
  assign n54027 = ~n54025 & ~n54026 ;
  assign n54028 = n54016 & ~n54027 ;
  assign n54029 = n54016 & ~n54028 ;
  assign n54030 = ~n54027 & ~n54028 ;
  assign n54031 = ~n54029 & ~n54030 ;
  assign n54032 = ~n53918 & ~n54031 ;
  assign n54033 = n53918 & n54031 ;
  assign n54034 = ~n54032 & ~n54033 ;
  assign n54035 = ~n54007 & n54034 ;
  assign n54036 = ~n54007 & ~n54035 ;
  assign n54037 = n54034 & ~n54035 ;
  assign n54038 = ~n54036 & ~n54037 ;
  assign n54039 = ~n54005 & ~n54038 ;
  assign n54040 = n54005 & ~n54037 ;
  assign n54041 = ~n54036 & n54040 ;
  assign n54042 = ~n54039 & ~n54041 ;
  assign n54082 = n54042 & x251 ;
  assign n54043 = ~n53993 & ~n53997 ;
  assign n54044 = ~n53967 & ~n53989 ;
  assign n54045 = ~n53986 & ~n54044 ;
  assign n54046 = ~x59 & ~n53959 ;
  assign n54047 = x59 & n53959 ;
  assign n54048 = ~n54046 & ~n54047 ;
  assign n54049 = ~x123 & n27427 ;
  assign n54050 = ~x124 & ~n26217 ;
  assign n54051 = ~n54049 & ~n54050 ;
  assign n54052 = n54048 & n54051 ;
  assign n54053 = ~n54048 & ~n54051 ;
  assign n54054 = ~n54052 & ~n54053 ;
  assign n54055 = ~x127 & n24612 ;
  assign n54056 = ~x125 & n25390 ;
  assign n54057 = ~x126 & n24607 ;
  assign n54058 = ~n54056 & ~n54057 ;
  assign n54059 = ~n54055 & n54058 ;
  assign n54060 = n24615 & n26932 ;
  assign n54061 = n54059 & ~n54060 ;
  assign n54062 = ~x62 & ~n54061 ;
  assign n54063 = ~x62 & ~n54062 ;
  assign n54064 = ~n54061 & ~n54062 ;
  assign n54065 = ~n54063 & ~n54064 ;
  assign n54066 = n54054 & ~n54065 ;
  assign n54067 = n54054 & ~n54066 ;
  assign n54068 = ~n54065 & ~n54066 ;
  assign n54069 = ~n54067 & ~n54068 ;
  assign n54070 = ~n53965 & ~n54069 ;
  assign n54071 = n53965 & n54069 ;
  assign n54072 = ~n54070 & ~n54071 ;
  assign n54073 = ~n54045 & n54072 ;
  assign n54074 = ~n54045 & ~n54073 ;
  assign n54075 = n54072 & ~n54073 ;
  assign n54076 = ~n54074 & ~n54075 ;
  assign n54077 = ~n54043 & ~n54076 ;
  assign n54078 = n54043 & ~n54075 ;
  assign n54079 = ~n54074 & n54078 ;
  assign n54080 = ~n54077 & ~n54079 ;
  assign n54083 = ~n54080 & ~x251 ;
  assign n54084 = ~n54082 & ~n54083 ;
  assign n54085 = ~n54035 & ~n54039 ;
  assign n54086 = ~n54028 & ~n54032 ;
  assign n54087 = x124 & n27024 ;
  assign n54088 = x125 & ~n26217 ;
  assign n54089 = ~n54087 & ~n54088 ;
  assign n54090 = ~x59 & ~n53912 ;
  assign n54091 = ~n54015 & ~n54090 ;
  assign n54092 = n54089 & ~n54091 ;
  assign n54093 = ~n54089 & n54091 ;
  assign n54094 = ~n54092 & ~n54093 ;
  assign n54095 = x126 & n25390 ;
  assign n54096 = x127 & n24607 ;
  assign n54097 = ~n54095 & ~n54096 ;
  assign n54098 = ~n24615 & n54097 ;
  assign n54099 = n26965 & n54097 ;
  assign n54100 = ~n54098 & ~n54099 ;
  assign n54101 = x62 & ~n54100 ;
  assign n54102 = ~x62 & n54100 ;
  assign n54103 = ~n54101 & ~n54102 ;
  assign n54104 = n54094 & ~n54103 ;
  assign n54105 = ~n54094 & n54103 ;
  assign n54106 = ~n54104 & ~n54105 ;
  assign n54107 = ~n54086 & n54106 ;
  assign n54108 = ~n54086 & ~n54107 ;
  assign n54109 = n54106 & ~n54107 ;
  assign n54110 = ~n54108 & ~n54109 ;
  assign n54111 = ~n54085 & ~n54110 ;
  assign n54112 = n54085 & ~n54109 ;
  assign n54113 = ~n54108 & n54112 ;
  assign n54114 = ~n54111 & ~n54113 ;
  assign n54146 = n54114 & x252 ;
  assign n54115 = ~n54073 & ~n54077 ;
  assign n54116 = ~n54066 & ~n54070 ;
  assign n54117 = ~x124 & n27427 ;
  assign n54118 = ~x125 & ~n26217 ;
  assign n54119 = ~n54117 & ~n54118 ;
  assign n54120 = x59 & ~n53959 ;
  assign n54121 = ~n54053 & ~n54120 ;
  assign n54122 = n54119 & ~n54121 ;
  assign n54123 = ~n54119 & n54121 ;
  assign n54124 = ~n54122 & ~n54123 ;
  assign n54125 = ~x126 & n25390 ;
  assign n54126 = ~x127 & n24607 ;
  assign n54127 = ~n54125 & ~n54126 ;
  assign n54128 = ~n24615 & n54127 ;
  assign n54129 = n27368 & n54127 ;
  assign n54130 = ~n54128 & ~n54129 ;
  assign n54131 = ~x62 & ~n54130 ;
  assign n54132 = x62 & n54130 ;
  assign n54133 = ~n54131 & ~n54132 ;
  assign n54134 = n54124 & ~n54133 ;
  assign n54135 = ~n54124 & n54133 ;
  assign n54136 = ~n54134 & ~n54135 ;
  assign n54137 = ~n54116 & n54136 ;
  assign n54138 = ~n54116 & ~n54137 ;
  assign n54139 = n54136 & ~n54137 ;
  assign n54140 = ~n54138 & ~n54139 ;
  assign n54141 = ~n54115 & ~n54140 ;
  assign n54142 = n54115 & ~n54139 ;
  assign n54143 = ~n54138 & n54142 ;
  assign n54144 = ~n54141 & ~n54143 ;
  assign n54147 = ~n54144 & ~x252 ;
  assign n54148 = ~n54146 & ~n54147 ;
  assign n54149 = ~n54107 & ~n54111 ;
  assign n54150 = ~n54092 & ~n54104 ;
  assign n54151 = x125 & n27024 ;
  assign n54152 = x126 & ~n26217 ;
  assign n54153 = ~n54151 & ~n54152 ;
  assign n54154 = n54089 & ~n54153 ;
  assign n54155 = ~n54089 & n54153 ;
  assign n54156 = ~n54154 & ~n54155 ;
  assign n54157 = x127 & n25390 ;
  assign n54158 = ~n24615 & ~n54157 ;
  assign n54159 = ~n26962 & ~n54157 ;
  assign n54160 = ~n54158 & ~n54159 ;
  assign n54161 = x62 & ~n54160 ;
  assign n54162 = ~x62 & n54160 ;
  assign n54163 = ~n54161 & ~n54162 ;
  assign n54164 = n54156 & ~n54163 ;
  assign n54165 = ~n54156 & n54163 ;
  assign n54166 = ~n54164 & ~n54165 ;
  assign n54167 = ~n54150 & n54166 ;
  assign n54168 = ~n54150 & ~n54167 ;
  assign n54169 = n54166 & ~n54167 ;
  assign n54170 = ~n54168 & ~n54169 ;
  assign n54171 = ~n54149 & ~n54170 ;
  assign n54172 = n54149 & ~n54169 ;
  assign n54173 = ~n54168 & n54172 ;
  assign n54174 = ~n54171 & ~n54173 ;
  assign n54202 = n54174 & x253 ;
  assign n54175 = ~n54137 & ~n54141 ;
  assign n54176 = ~n54122 & ~n54134 ;
  assign n54177 = ~x125 & n27427 ;
  assign n54178 = ~x126 & ~n26217 ;
  assign n54179 = ~n54177 & ~n54178 ;
  assign n54180 = n54119 & ~n54179 ;
  assign n54181 = ~n54119 & n54179 ;
  assign n54182 = ~n54180 & ~n54181 ;
  assign n54183 = ~x127 & n25390 ;
  assign n54184 = ~n24615 & ~n54183 ;
  assign n54185 = ~n27365 & ~n54183 ;
  assign n54186 = ~n54184 & ~n54185 ;
  assign n54187 = ~x62 & ~n54186 ;
  assign n54188 = x62 & n54186 ;
  assign n54189 = ~n54187 & ~n54188 ;
  assign n54190 = n54182 & ~n54189 ;
  assign n54191 = ~n54182 & n54189 ;
  assign n54192 = ~n54190 & ~n54191 ;
  assign n54193 = ~n54176 & n54192 ;
  assign n54194 = ~n54176 & ~n54193 ;
  assign n54195 = n54192 & ~n54193 ;
  assign n54196 = ~n54194 & ~n54195 ;
  assign n54197 = ~n54175 & ~n54196 ;
  assign n54198 = n54175 & ~n54195 ;
  assign n54199 = ~n54194 & n54198 ;
  assign n54200 = ~n54197 & ~n54199 ;
  assign n54203 = ~n54200 & ~x253 ;
  assign n54204 = ~n54202 & ~n54203 ;
  assign n54205 = ~n54167 & ~n54171 ;
  assign n54206 = ~n54154 & ~n54164 ;
  assign n54207 = x126 & n27024 ;
  assign n54208 = x127 & ~n26217 ;
  assign n54209 = ~n54207 & ~n54208 ;
  assign n54210 = ~x62 & ~n54209 ;
  assign n54211 = x62 & n54209 ;
  assign n54212 = ~n54210 & ~n54211 ;
  assign n54213 = ~n54089 & n54212 ;
  assign n54214 = n54089 & ~n54212 ;
  assign n54215 = ~n54213 & ~n54214 ;
  assign n54216 = ~n54206 & n54215 ;
  assign n54217 = n54206 & ~n54215 ;
  assign n54218 = ~n54216 & ~n54217 ;
  assign n54219 = ~n54205 & n54218 ;
  assign n54220 = n54205 & ~n54218 ;
  assign n54221 = ~n54219 & ~n54220 ;
  assign n54240 = n54221 & x254 ;
  assign n54222 = ~n54193 & ~n54197 ;
  assign n54223 = ~n54180 & ~n54190 ;
  assign n54224 = ~x126 & n27427 ;
  assign n54225 = ~x127 & ~n26217 ;
  assign n54226 = ~n54224 & ~n54225 ;
  assign n54227 = x62 & ~n54226 ;
  assign n54228 = ~x62 & n54226 ;
  assign n54229 = ~n54227 & ~n54228 ;
  assign n54230 = ~n54119 & n54229 ;
  assign n54231 = n54119 & ~n54229 ;
  assign n54232 = ~n54230 & ~n54231 ;
  assign n54233 = ~n54223 & n54232 ;
  assign n54234 = n54223 & ~n54232 ;
  assign n54235 = ~n54233 & ~n54234 ;
  assign n54236 = ~n54222 & n54235 ;
  assign n54237 = n54222 & ~n54235 ;
  assign n54238 = ~n54236 & ~n54237 ;
  assign n54241 = ~n54238 & ~x254 ;
  assign n54242 = ~n54240 & ~n54241 ;
  assign n54243 = ~n54210 & ~n54213 ;
  assign n54244 = x127 & n27024 ;
  assign n54245 = ~n54243 & n54244 ;
  assign n54246 = n54243 & ~n54244 ;
  assign n54247 = ~n54245 & ~n54246 ;
  assign n54248 = ~n54216 & ~n54219 ;
  assign n54249 = n54247 & n54248 ;
  assign n54250 = ~n54247 & ~n54248 ;
  assign n54251 = ~n54249 & ~n54250 ;
  assign n54262 = n54251 & x255 ;
  assign n54252 = ~n54227 & ~n54230 ;
  assign n54253 = ~x127 & n27427 ;
  assign n54254 = ~n54252 & n54253 ;
  assign n54255 = n54252 & ~n54253 ;
  assign n54256 = ~n54254 & ~n54255 ;
  assign n54257 = ~n54233 & ~n54236 ;
  assign n54258 = n54256 & n54257 ;
  assign n54259 = ~n54256 & ~n54257 ;
  assign n54260 = ~n54258 & ~n54259 ;
  assign n54263 = ~n54260 & ~x255 ;
  assign n54264 = ~n54262 & ~n54263 ;
  assign y0 = ~n140 ;
  assign y1 = ~n180 ;
  assign y2 = ~n227 ;
  assign y3 = ~n283 ;
  assign y4 = ~n370 ;
  assign y5 = ~n453 ;
  assign y6 = ~n545 ;
  assign y7 = ~n670 ;
  assign y8 = ~n791 ;
  assign y9 = ~n921 ;
  assign y10 = ~n1082 ;
  assign y11 = ~n1241 ;
  assign y12 = ~n1409 ;
  assign y13 = ~n1610 ;
  assign y14 = ~n1803 ;
  assign y15 = ~n2015 ;
  assign y16 = ~n2246 ;
  assign y17 = ~n2479 ;
  assign y18 = ~n2715 ;
  assign y19 = ~n2990 ;
  assign y20 = ~n3265 ;
  assign y21 = ~n3539 ;
  assign y22 = ~n3848 ;
  assign y23 = ~n4161 ;
  assign y24 = ~n4475 ;
  assign y25 = ~n4824 ;
  assign y26 = ~n5171 ;
  assign y27 = ~n5523 ;
  assign y28 = ~n5912 ;
  assign y29 = ~n6303 ;
  assign y30 = ~n6689 ;
  assign y31 = ~n7118 ;
  assign y32 = ~n7547 ;
  assign y33 = ~n7965 ;
  assign y34 = ~n8442 ;
  assign y35 = ~n8901 ;
  assign y36 = ~n9357 ;
  assign y37 = ~n9860 ;
  assign y38 = ~n10351 ;
  assign y39 = ~n10851 ;
  assign y40 = ~n11396 ;
  assign y41 = ~n11923 ;
  assign y42 = ~n12465 ;
  assign y43 = ~n13052 ;
  assign y44 = ~n13617 ;
  assign y45 = ~n14193 ;
  assign y46 = ~n14820 ;
  assign y47 = ~n15429 ;
  assign y48 = ~n16037 ;
  assign y49 = ~n16700 ;
  assign y50 = ~n17351 ;
  assign y51 = ~n17993 ;
  assign y52 = ~n18694 ;
  assign y53 = ~n19381 ;
  assign y54 = ~n20067 ;
  assign y55 = ~n20794 ;
  assign y56 = ~n21519 ;
  assign y57 = ~n22247 ;
  assign y58 = ~n23016 ;
  assign y59 = ~n23781 ;
  assign y60 = ~n24545 ;
  assign y61 = ~n25352 ;
  assign y62 = ~n26147 ;
  assign y63 = ~n26955 ;
  assign y64 = ~n27765 ;
  assign y65 = ~n28565 ;
  assign y66 = ~n29347 ;
  assign y67 = ~n30143 ;
  assign y68 = ~n30929 ;
  assign y69 = ~n31686 ;
  assign y70 = ~n32434 ;
  assign y71 = ~n33184 ;
  assign y72 = ~n33916 ;
  assign y73 = ~n34650 ;
  assign y74 = ~n35356 ;
  assign y75 = ~n36052 ;
  assign y76 = ~n36748 ;
  assign y77 = ~n37404 ;
  assign y78 = ~n38058 ;
  assign y79 = ~n38692 ;
  assign y80 = ~n39318 ;
  assign y81 = ~n39926 ;
  assign y82 = ~n40526 ;
  assign y83 = ~n41102 ;
  assign y84 = ~n41680 ;
  assign y85 = ~n42232 ;
  assign y86 = ~n42778 ;
  assign y87 = ~n43314 ;
  assign y88 = ~n43838 ;
  assign y89 = ~n44340 ;
  assign y90 = ~n44830 ;
  assign y91 = ~n45308 ;
  assign y92 = ~n45782 ;
  assign y93 = ~n46238 ;
  assign y94 = ~n46682 ;
  assign y95 = ~n47118 ;
  assign y96 = ~n47538 ;
  assign y97 = ~n47940 ;
  assign y98 = ~n48336 ;
  assign y99 = ~n48714 ;
  assign y100 = ~n49084 ;
  assign y101 = ~n49442 ;
  assign y102 = ~n49786 ;
  assign y103 = ~n50114 ;
  assign y104 = ~n50436 ;
  assign y105 = ~n50742 ;
  assign y106 = ~n51032 ;
  assign y107 = ~n51322 ;
  assign y108 = ~n51586 ;
  assign y109 = ~n51836 ;
  assign y110 = ~n52086 ;
  assign y111 = ~n52310 ;
  assign y112 = ~n52524 ;
  assign y113 = ~n52730 ;
  assign y114 = ~n52922 ;
  assign y115 = ~n53094 ;
  assign y116 = ~n53262 ;
  assign y117 = ~n53416 ;
  assign y118 = ~n53558 ;
  assign y119 = ~n53690 ;
  assign y120 = ~n53810 ;
  assign y121 = ~n53906 ;
  assign y122 = ~n54004 ;
  assign y123 = ~n54084 ;
  assign y124 = ~n54148 ;
  assign y125 = ~n54204 ;
  assign y126 = ~n54242 ;
  assign y127 = ~n54264 ;
endmodule
