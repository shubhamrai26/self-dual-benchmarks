module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 , y15409 , y15410 , y15411 , y15412 , y15413 , y15414 , y15415 , y15416 , y15417 , y15418 , y15419 , y15420 , y15421 , y15422 , y15423 , y15424 , y15425 , y15426 , y15427 , y15428 , y15429 , y15430 , y15431 , y15432 , y15433 , y15434 , y15435 , y15436 , y15437 , y15438 , y15439 , y15440 , y15441 , y15442 , y15443 , y15444 , y15445 , y15446 , y15447 , y15448 , y15449 , y15450 , y15451 , y15452 , y15453 , y15454 , y15455 , y15456 , y15457 , y15458 , y15459 , y15460 , y15461 , y15462 , y15463 , y15464 , y15465 , y15466 , y15467 , y15468 , y15469 , y15470 , y15471 , y15472 , y15473 , y15474 , y15475 , y15476 , y15477 , y15478 , y15479 , y15480 , y15481 , y15482 , y15483 , y15484 , y15485 , y15486 , y15487 , y15488 , y15489 , y15490 , y15491 , y15492 , y15493 , y15494 , y15495 , y15496 , y15497 , y15498 , y15499 , y15500 , y15501 , y15502 , y15503 , y15504 , y15505 , y15506 , y15507 , y15508 , y15509 , y15510 , y15511 , y15512 , y15513 , y15514 , y15515 , y15516 , y15517 , y15518 , y15519 , y15520 , y15521 , y15522 , y15523 , y15524 , y15525 , y15526 , y15527 , y15528 , y15529 , y15530 , y15531 , y15532 , y15533 , y15534 , y15535 , y15536 , y15537 , y15538 , y15539 , y15540 , y15541 , y15542 , y15543 , y15544 , y15545 , y15546 , y15547 , y15548 , y15549 , y15550 , y15551 , y15552 , y15553 , y15554 , y15555 , y15556 , y15557 , y15558 , y15559 , y15560 , y15561 , y15562 , y15563 , y15564 , y15565 , y15566 , y15567 , y15568 , y15569 , y15570 , y15571 , y15572 , y15573 , y15574 , y15575 , y15576 , y15577 , y15578 , y15579 , y15580 , y15581 , y15582 , y15583 , y15584 , y15585 , y15586 , y15587 , y15588 , y15589 , y15590 , y15591 , y15592 , y15593 , y15594 , y15595 , y15596 , y15597 , y15598 , y15599 , y15600 , y15601 , y15602 , y15603 , y15604 , y15605 , y15606 , y15607 , y15608 , y15609 , y15610 , y15611 , y15612 , y15613 , y15614 , y15615 , y15616 , y15617 , y15618 , y15619 , y15620 , y15621 , y15622 , y15623 , y15624 , y15625 , y15626 , y15627 , y15628 , y15629 , y15630 , y15631 , y15632 , y15633 , y15634 , y15635 , y15636 , y15637 , y15638 , y15639 , y15640 , y15641 , y15642 , y15643 , y15644 , y15645 , y15646 , y15647 , y15648 , y15649 , y15650 , y15651 , y15652 , y15653 , y15654 , y15655 , y15656 , y15657 , y15658 , y15659 , y15660 , y15661 , y15662 , y15663 , y15664 , y15665 , y15666 , y15667 , y15668 , y15669 , y15670 , y15671 , y15672 , y15673 , y15674 , y15675 , y15676 , y15677 , y15678 , y15679 , y15680 , y15681 , y15682 , y15683 , y15684 , y15685 , y15686 , y15687 , y15688 , y15689 , y15690 , y15691 , y15692 , y15693 , y15694 , y15695 , y15696 , y15697 , y15698 , y15699 , y15700 , y15701 , y15702 , y15703 , y15704 , y15705 , y15706 , y15707 , y15708 , y15709 , y15710 , y15711 , y15712 , y15713 , y15714 , y15715 , y15716 , y15717 , y15718 , y15719 , y15720 , y15721 , y15722 , y15723 , y15724 , y15725 , y15726 , y15727 , y15728 , y15729 , y15730 , y15731 , y15732 , y15733 , y15734 , y15735 , y15736 , y15737 , y15738 , y15739 , y15740 , y15741 , y15742 , y15743 , y15744 , y15745 , y15746 , y15747 , y15748 , y15749 , y15750 , y15751 , y15752 , y15753 , y15754 , y15755 , y15756 , y15757 , y15758 , y15759 , y15760 , y15761 , y15762 , y15763 , y15764 , y15765 , y15766 , y15767 , y15768 , y15769 , y15770 , y15771 , y15772 , y15773 , y15774 , y15775 , y15776 , y15777 , y15778 , y15779 , y15780 , y15781 , y15782 , y15783 , y15784 , y15785 , y15786 , y15787 , y15788 , y15789 , y15790 , y15791 , y15792 , y15793 , y15794 , y15795 , y15796 , y15797 , y15798 , y15799 , y15800 , y15801 , y15802 , y15803 , y15804 , y15805 , y15806 , y15807 , y15808 , y15809 , y15810 , y15811 , y15812 , y15813 , y15814 , y15815 , y15816 , y15817 , y15818 , y15819 , y15820 , y15821 , y15822 , y15823 , y15824 , y15825 , y15826 , y15827 , y15828 , y15829 , y15830 , y15831 , y15832 , y15833 , y15834 , y15835 , y15836 , y15837 , y15838 , y15839 , y15840 , y15841 , y15842 , y15843 , y15844 , y15845 , y15846 , y15847 , y15848 , y15849 , y15850 , y15851 , y15852 , y15853 , y15854 , y15855 , y15856 , y15857 , y15858 , y15859 , y15860 , y15861 , y15862 , y15863 , y15864 , y15865 , y15866 , y15867 , y15868 , y15869 , y15870 , y15871 , y15872 , y15873 , y15874 , y15875 , y15876 , y15877 , y15878 , y15879 , y15880 , y15881 , y15882 , y15883 , y15884 , y15885 , y15886 , y15887 , y15888 , y15889 , y15890 , y15891 , y15892 , y15893 , y15894 , y15895 , y15896 , y15897 , y15898 , y15899 , y15900 , y15901 , y15902 , y15903 , y15904 , y15905 , y15906 , y15907 , y15908 , y15909 , y15910 , y15911 , y15912 , y15913 , y15914 , y15915 , y15916 , y15917 , y15918 , y15919 , y15920 , y15921 , y15922 , y15923 , y15924 , y15925 , y15926 , y15927 , y15928 , y15929 , y15930 , y15931 , y15932 , y15933 , y15934 , y15935 , y15936 , y15937 , y15938 , y15939 , y15940 , y15941 , y15942 , y15943 , y15944 , y15945 , y15946 , y15947 , y15948 , y15949 , y15950 , y15951 , y15952 , y15953 , y15954 , y15955 , y15956 , y15957 , y15958 , y15959 , y15960 , y15961 , y15962 , y15963 , y15964 , y15965 , y15966 , y15967 , y15968 , y15969 , y15970 , y15971 , y15972 , y15973 , y15974 , y15975 , y15976 , y15977 , y15978 , y15979 , y15980 , y15981 , y15982 , y15983 , y15984 , y15985 , y15986 , y15987 , y15988 , y15989 , y15990 , y15991 , y15992 , y15993 , y15994 , y15995 , y15996 , y15997 , y15998 , y15999 , y16000 , y16001 , y16002 , y16003 , y16004 , y16005 , y16006 , y16007 , y16008 , y16009 , y16010 , y16011 , y16012 , y16013 , y16014 , y16015 , y16016 , y16017 , y16018 , y16019 , y16020 , y16021 , y16022 , y16023 , y16024 , y16025 , y16026 , y16027 , y16028 , y16029 , y16030 , y16031 , y16032 , y16033 , y16034 , y16035 , y16036 , y16037 , y16038 , y16039 , y16040 , y16041 , y16042 , y16043 , y16044 , y16045 , y16046 , y16047 , y16048 , y16049 , y16050 , y16051 , y16052 , y16053 , y16054 , y16055 , y16056 , y16057 , y16058 , y16059 , y16060 , y16061 , y16062 , y16063 , y16064 , y16065 , y16066 , y16067 , y16068 , y16069 , y16070 , y16071 , y16072 , y16073 , y16074 , y16075 , y16076 , y16077 , y16078 , y16079 , y16080 , y16081 , y16082 , y16083 , y16084 , y16085 , y16086 , y16087 , y16088 , y16089 , y16090 , y16091 , y16092 , y16093 , y16094 , y16095 , y16096 , y16097 , y16098 , y16099 , y16100 , y16101 , y16102 , y16103 , y16104 , y16105 , y16106 , y16107 , y16108 , y16109 , y16110 , y16111 , y16112 , y16113 , y16114 , y16115 , y16116 , y16117 , y16118 , y16119 , y16120 , y16121 , y16122 , y16123 , y16124 , y16125 , y16126 , y16127 , y16128 , y16129 , y16130 , y16131 , y16132 , y16133 , y16134 , y16135 , y16136 , y16137 , y16138 , y16139 , y16140 , y16141 , y16142 , y16143 , y16144 , y16145 , y16146 , y16147 , y16148 , y16149 , y16150 , y16151 , y16152 , y16153 , y16154 , y16155 , y16156 , y16157 , y16158 , y16159 , y16160 , y16161 , y16162 , y16163 , y16164 , y16165 , y16166 , y16167 , y16168 , y16169 , y16170 , y16171 , y16172 , y16173 , y16174 , y16175 , y16176 , y16177 , y16178 , y16179 , y16180 , y16181 , y16182 , y16183 , y16184 , y16185 , y16186 , y16187 , y16188 , y16189 , y16190 , y16191 , y16192 , y16193 , y16194 , y16195 , y16196 , y16197 , y16198 , y16199 , y16200 , y16201 , y16202 , y16203 , y16204 , y16205 , y16206 , y16207 , y16208 , y16209 , y16210 , y16211 , y16212 , y16213 , y16214 , y16215 , y16216 , y16217 , y16218 , y16219 , y16220 , y16221 , y16222 , y16223 , y16224 , y16225 , y16226 , y16227 , y16228 , y16229 , y16230 , y16231 , y16232 , y16233 , y16234 , y16235 , y16236 , y16237 , y16238 , y16239 , y16240 , y16241 , y16242 , y16243 , y16244 , y16245 , y16246 , y16247 , y16248 , y16249 , y16250 , y16251 , y16252 , y16253 , y16254 , y16255 , y16256 , y16257 , y16258 , y16259 , y16260 , y16261 , y16262 , y16263 , y16264 , y16265 , y16266 , y16267 , y16268 , y16269 , y16270 , y16271 , y16272 , y16273 , y16274 , y16275 , y16276 , y16277 , y16278 , y16279 , y16280 , y16281 , y16282 , y16283 , y16284 , y16285 , y16286 , y16287 , y16288 , y16289 , y16290 , y16291 , y16292 , y16293 , y16294 , y16295 , y16296 , y16297 , y16298 , y16299 , y16300 , y16301 , y16302 , y16303 , y16304 , y16305 , y16306 , y16307 , y16308 , y16309 , y16310 , y16311 , y16312 , y16313 , y16314 , y16315 , y16316 , y16317 , y16318 , y16319 , y16320 , y16321 , y16322 , y16323 , y16324 , y16325 , y16326 , y16327 , y16328 , y16329 , y16330 , y16331 , y16332 , y16333 , y16334 , y16335 , y16336 , y16337 , y16338 , y16339 , y16340 , y16341 , y16342 , y16343 , y16344 , y16345 , y16346 , y16347 , y16348 , y16349 , y16350 , y16351 , y16352 , y16353 , y16354 , y16355 , y16356 , y16357 , y16358 , y16359 , y16360 , y16361 , y16362 , y16363 , y16364 , y16365 , y16366 , y16367 , y16368 , y16369 , y16370 , y16371 , y16372 , y16373 , y16374 , y16375 , y16376 , y16377 , y16378 , y16379 , y16380 , y16381 , y16382 , y16383 , y16384 , y16385 , y16386 , y16387 , y16388 , y16389 , y16390 , y16391 , y16392 , y16393 , y16394 , y16395 , y16396 , y16397 , y16398 , y16399 , y16400 , y16401 , y16402 , y16403 , y16404 , y16405 , y16406 , y16407 , y16408 , y16409 , y16410 , y16411 , y16412 , y16413 , y16414 , y16415 , y16416 , y16417 , y16418 , y16419 , y16420 , y16421 , y16422 , y16423 , y16424 , y16425 , y16426 , y16427 , y16428 , y16429 , y16430 , y16431 , y16432 , y16433 , y16434 , y16435 , y16436 , y16437 , y16438 , y16439 , y16440 , y16441 , y16442 , y16443 , y16444 , y16445 , y16446 , y16447 , y16448 , y16449 , y16450 , y16451 , y16452 , y16453 , y16454 , y16455 , y16456 , y16457 , y16458 , y16459 , y16460 , y16461 , y16462 , y16463 , y16464 , y16465 , y16466 , y16467 , y16468 , y16469 , y16470 , y16471 , y16472 , y16473 , y16474 , y16475 , y16476 , y16477 , y16478 , y16479 , y16480 , y16481 , y16482 , y16483 , y16484 , y16485 , y16486 , y16487 , y16488 , y16489 , y16490 , y16491 , y16492 , y16493 , y16494 , y16495 , y16496 , y16497 , y16498 , y16499 , y16500 , y16501 , y16502 , y16503 , y16504 , y16505 , y16506 , y16507 , y16508 , y16509 , y16510 , y16511 , y16512 , y16513 , y16514 , y16515 , y16516 , y16517 , y16518 , y16519 , y16520 , y16521 , y16522 , y16523 , y16524 , y16525 , y16526 , y16527 , y16528 , y16529 , y16530 , y16531 , y16532 , y16533 , y16534 , y16535 , y16536 , y16537 , y16538 , y16539 , y16540 , y16541 , y16542 , y16543 , y16544 , y16545 , y16546 , y16547 , y16548 , y16549 , y16550 , y16551 , y16552 , y16553 , y16554 , y16555 , y16556 , y16557 , y16558 , y16559 , y16560 , y16561 , y16562 , y16563 , y16564 , y16565 , y16566 , y16567 , y16568 , y16569 , y16570 , y16571 , y16572 , y16573 , y16574 , y16575 , y16576 , y16577 , y16578 , y16579 , y16580 , y16581 , y16582 , y16583 , y16584 , y16585 , y16586 , y16587 , y16588 , y16589 , y16590 , y16591 , y16592 , y16593 , y16594 , y16595 , y16596 , y16597 , y16598 , y16599 , y16600 , y16601 , y16602 , y16603 , y16604 , y16605 , y16606 , y16607 , y16608 , y16609 , y16610 , y16611 , y16612 , y16613 , y16614 , y16615 , y16616 , y16617 , y16618 , y16619 , y16620 , y16621 , y16622 , y16623 , y16624 , y16625 , y16626 , y16627 , y16628 , y16629 , y16630 , y16631 , y16632 , y16633 , y16634 , y16635 , y16636 , y16637 , y16638 , y16639 , y16640 , y16641 , y16642 , y16643 , y16644 , y16645 , y16646 , y16647 , y16648 , y16649 , y16650 , y16651 , y16652 , y16653 , y16654 , y16655 , y16656 , y16657 , y16658 , y16659 , y16660 , y16661 , y16662 , y16663 , y16664 , y16665 , y16666 , y16667 , y16668 , y16669 , y16670 , y16671 , y16672 , y16673 , y16674 , y16675 , y16676 , y16677 , y16678 , y16679 , y16680 , y16681 , y16682 , y16683 , y16684 , y16685 , y16686 , y16687 , y16688 , y16689 , y16690 , y16691 , y16692 , y16693 , y16694 , y16695 , y16696 , y16697 , y16698 , y16699 , y16700 , y16701 , y16702 , y16703 , y16704 , y16705 , y16706 , y16707 , y16708 , y16709 , y16710 , y16711 , y16712 , y16713 , y16714 , y16715 , y16716 , y16717 , y16718 , y16719 , y16720 , y16721 , y16722 , y16723 , y16724 , y16725 , y16726 , y16727 , y16728 , y16729 , y16730 , y16731 , y16732 , y16733 , y16734 , y16735 , y16736 , y16737 , y16738 , y16739 , y16740 , y16741 , y16742 , y16743 , y16744 , y16745 , y16746 , y16747 , y16748 , y16749 , y16750 , y16751 , y16752 , y16753 , y16754 , y16755 , y16756 , y16757 , y16758 , y16759 , y16760 , y16761 , y16762 , y16763 , y16764 , y16765 , y16766 , y16767 , y16768 , y16769 , y16770 , y16771 , y16772 , y16773 , y16774 , y16775 , y16776 , y16777 , y16778 , y16779 , y16780 , y16781 , y16782 , y16783 , y16784 , y16785 , y16786 , y16787 , y16788 , y16789 , y16790 , y16791 , y16792 , y16793 , y16794 , y16795 , y16796 , y16797 , y16798 , y16799 , y16800 , y16801 , y16802 , y16803 , y16804 , y16805 , y16806 , y16807 , y16808 , y16809 , y16810 , y16811 , y16812 , y16813 , y16814 , y16815 , y16816 , y16817 , y16818 , y16819 , y16820 , y16821 , y16822 , y16823 , y16824 , y16825 , y16826 , y16827 , y16828 , y16829 , y16830 , y16831 , y16832 , y16833 , y16834 , y16835 , y16836 , y16837 , y16838 , y16839 , y16840 , y16841 , y16842 , y16843 , y16844 , y16845 , y16846 , y16847 , y16848 , y16849 , y16850 , y16851 , y16852 , y16853 , y16854 , y16855 , y16856 , y16857 , y16858 , y16859 , y16860 , y16861 , y16862 , y16863 , y16864 , y16865 , y16866 , y16867 , y16868 , y16869 , y16870 , y16871 , y16872 , y16873 , y16874 , y16875 , y16876 , y16877 , y16878 , y16879 , y16880 , y16881 , y16882 , y16883 , y16884 , y16885 , y16886 , y16887 , y16888 , y16889 , y16890 , y16891 , y16892 , y16893 , y16894 , y16895 , y16896 , y16897 , y16898 , y16899 , y16900 , y16901 , y16902 , y16903 , y16904 , y16905 , y16906 , y16907 , y16908 , y16909 , y16910 , y16911 , y16912 , y16913 , y16914 , y16915 , y16916 , y16917 , y16918 , y16919 , y16920 , y16921 , y16922 , y16923 , y16924 , y16925 , y16926 , y16927 , y16928 , y16929 , y16930 , y16931 , y16932 , y16933 , y16934 , y16935 , y16936 , y16937 , y16938 , y16939 , y16940 , y16941 , y16942 , y16943 , y16944 , y16945 , y16946 , y16947 , y16948 , y16949 , y16950 , y16951 , y16952 , y16953 , y16954 , y16955 , y16956 , y16957 , y16958 , y16959 , y16960 , y16961 , y16962 , y16963 , y16964 , y16965 , y16966 , y16967 , y16968 , y16969 , y16970 , y16971 , y16972 , y16973 , y16974 , y16975 , y16976 , y16977 , y16978 , y16979 , y16980 , y16981 , y16982 , y16983 , y16984 , y16985 , y16986 , y16987 , y16988 , y16989 , y16990 , y16991 , y16992 , y16993 , y16994 , y16995 , y16996 , y16997 , y16998 , y16999 , y17000 , y17001 , y17002 , y17003 , y17004 , y17005 , y17006 , y17007 , y17008 , y17009 , y17010 , y17011 , y17012 , y17013 , y17014 , y17015 , y17016 , y17017 , y17018 , y17019 , y17020 , y17021 , y17022 , y17023 , y17024 , y17025 , y17026 , y17027 , y17028 , y17029 , y17030 , y17031 , y17032 , y17033 , y17034 , y17035 , y17036 , y17037 , y17038 , y17039 , y17040 , y17041 , y17042 , y17043 , y17044 , y17045 , y17046 , y17047 , y17048 , y17049 , y17050 , y17051 , y17052 , y17053 , y17054 , y17055 , y17056 , y17057 , y17058 , y17059 , y17060 , y17061 , y17062 , y17063 , y17064 , y17065 , y17066 , y17067 , y17068 , y17069 , y17070 , y17071 , y17072 , y17073 , y17074 , y17075 , y17076 , y17077 , y17078 , y17079 , y17080 , y17081 , y17082 , y17083 , y17084 , y17085 , y17086 , y17087 , y17088 , y17089 , y17090 , y17091 , y17092 , y17093 , y17094 , y17095 , y17096 , y17097 , y17098 , y17099 , y17100 , y17101 , y17102 , y17103 , y17104 , y17105 , y17106 , y17107 , y17108 , y17109 , y17110 , y17111 , y17112 , y17113 , y17114 , y17115 , y17116 , y17117 , y17118 , y17119 , y17120 , y17121 , y17122 , y17123 , y17124 , y17125 , y17126 , y17127 , y17128 , y17129 , y17130 , y17131 , y17132 , y17133 , y17134 , y17135 , y17136 , y17137 , y17138 , y17139 , y17140 , y17141 , y17142 , y17143 , y17144 , y17145 , y17146 , y17147 , y17148 , y17149 , y17150 , y17151 , y17152 , y17153 , y17154 , y17155 , y17156 , y17157 , y17158 , y17159 , y17160 , y17161 , y17162 , y17163 , y17164 , y17165 , y17166 , y17167 , y17168 , y17169 , y17170 , y17171 , y17172 , y17173 , y17174 , y17175 , y17176 , y17177 , y17178 , y17179 , y17180 , y17181 , y17182 , y17183 , y17184 , y17185 , y17186 , y17187 , y17188 , y17189 , y17190 , y17191 , y17192 , y17193 , y17194 , y17195 , y17196 , y17197 , y17198 , y17199 , y17200 , y17201 , y17202 , y17203 , y17204 , y17205 , y17206 , y17207 , y17208 , y17209 , y17210 , y17211 , y17212 , y17213 , y17214 , y17215 , y17216 , y17217 , y17218 , y17219 , y17220 , y17221 , y17222 , y17223 , y17224 , y17225 , y17226 , y17227 , y17228 , y17229 , y17230 , y17231 , y17232 , y17233 , y17234 , y17235 , y17236 , y17237 , y17238 , y17239 , y17240 , y17241 , y17242 , y17243 , y17244 , y17245 , y17246 , y17247 , y17248 , y17249 , y17250 , y17251 , y17252 , y17253 , y17254 , y17255 , y17256 , y17257 , y17258 , y17259 , y17260 , y17261 , y17262 , y17263 , y17264 , y17265 , y17266 , y17267 , y17268 , y17269 , y17270 , y17271 , y17272 , y17273 , y17274 , y17275 , y17276 , y17277 , y17278 , y17279 , y17280 , y17281 , y17282 , y17283 , y17284 , y17285 , y17286 , y17287 , y17288 , y17289 , y17290 , y17291 , y17292 , y17293 , y17294 , y17295 , y17296 , y17297 , y17298 , y17299 , y17300 , y17301 , y17302 , y17303 , y17304 , y17305 , y17306 , y17307 , y17308 , y17309 , y17310 , y17311 , y17312 , y17313 , y17314 , y17315 , y17316 , y17317 , y17318 , y17319 , y17320 , y17321 , y17322 , y17323 , y17324 , y17325 , y17326 , y17327 , y17328 , y17329 , y17330 , y17331 , y17332 , y17333 , y17334 , y17335 , y17336 , y17337 , y17338 , y17339 , y17340 , y17341 , y17342 , y17343 , y17344 , y17345 , y17346 , y17347 , y17348 , y17349 , y17350 , y17351 , y17352 , y17353 , y17354 , y17355 , y17356 , y17357 , y17358 , y17359 , y17360 , y17361 , y17362 , y17363 , y17364 , y17365 , y17366 , y17367 , y17368 , y17369 , y17370 , y17371 , y17372 , y17373 , y17374 , y17375 , y17376 , y17377 , y17378 , y17379 , y17380 , y17381 , y17382 , y17383 , y17384 , y17385 , y17386 , y17387 , y17388 , y17389 , y17390 , y17391 , y17392 , y17393 , y17394 , y17395 , y17396 , y17397 , y17398 , y17399 , y17400 , y17401 , y17402 , y17403 , y17404 , y17405 , y17406 , y17407 , y17408 , y17409 , y17410 , y17411 , y17412 , y17413 , y17414 , y17415 , y17416 , y17417 , y17418 , y17419 , y17420 , y17421 , y17422 , y17423 , y17424 , y17425 , y17426 , y17427 , y17428 , y17429 , y17430 , y17431 , y17432 , y17433 , y17434 , y17435 , y17436 , y17437 , y17438 , y17439 , y17440 , y17441 , y17442 , y17443 , y17444 , y17445 , y17446 , y17447 , y17448 , y17449 , y17450 , y17451 , y17452 , y17453 , y17454 , y17455 , y17456 , y17457 , y17458 , y17459 , y17460 , y17461 , y17462 , y17463 , y17464 , y17465 , y17466 , y17467 , y17468 , y17469 , y17470 , y17471 , y17472 , y17473 , y17474 , y17475 , y17476 , y17477 , y17478 , y17479 , y17480 , y17481 , y17482 , y17483 , y17484 , y17485 , y17486 , y17487 , y17488 , y17489 , y17490 , y17491 , y17492 , y17493 , y17494 , y17495 , y17496 , y17497 , y17498 , y17499 , y17500 , y17501 , y17502 , y17503 , y17504 , y17505 , y17506 , y17507 , y17508 , y17509 , y17510 , y17511 , y17512 , y17513 , y17514 , y17515 , y17516 , y17517 , y17518 , y17519 , y17520 , y17521 , y17522 , y17523 , y17524 , y17525 , y17526 , y17527 , y17528 , y17529 , y17530 , y17531 , y17532 , y17533 , y17534 , y17535 , y17536 , y17537 , y17538 , y17539 , y17540 , y17541 , y17542 , y17543 , y17544 , y17545 , y17546 , y17547 , y17548 , y17549 , y17550 , y17551 , y17552 , y17553 , y17554 , y17555 , y17556 , y17557 , y17558 , y17559 , y17560 , y17561 , y17562 , y17563 , y17564 , y17565 , y17566 , y17567 , y17568 , y17569 , y17570 , y17571 , y17572 , y17573 , y17574 , y17575 , y17576 , y17577 , y17578 , y17579 , y17580 , y17581 , y17582 , y17583 , y17584 , y17585 , y17586 , y17587 , y17588 , y17589 , y17590 , y17591 , y17592 , y17593 , y17594 , y17595 , y17596 , y17597 , y17598 , y17599 , y17600 , y17601 , y17602 , y17603 , y17604 , y17605 , y17606 , y17607 , y17608 , y17609 , y17610 , y17611 , y17612 , y17613 , y17614 , y17615 , y17616 , y17617 , y17618 , y17619 , y17620 , y17621 , y17622 , y17623 , y17624 , y17625 , y17626 , y17627 , y17628 , y17629 , y17630 , y17631 , y17632 , y17633 , y17634 , y17635 , y17636 , y17637 , y17638 , y17639 , y17640 , y17641 , y17642 , y17643 , y17644 , y17645 , y17646 , y17647 , y17648 , y17649 , y17650 , y17651 , y17652 , y17653 , y17654 , y17655 , y17656 , y17657 , y17658 , y17659 , y17660 , y17661 , y17662 , y17663 , y17664 , y17665 , y17666 , y17667 , y17668 , y17669 , y17670 , y17671 , y17672 , y17673 , y17674 , y17675 , y17676 , y17677 , y17678 , y17679 , y17680 , y17681 , y17682 , y17683 , y17684 , y17685 , y17686 , y17687 , y17688 , y17689 , y17690 , y17691 , y17692 , y17693 , y17694 , y17695 , y17696 , y17697 , y17698 , y17699 , y17700 , y17701 , y17702 , y17703 , y17704 , y17705 , y17706 , y17707 , y17708 , y17709 , y17710 , y17711 , y17712 , y17713 , y17714 , y17715 , y17716 , y17717 , y17718 , y17719 , y17720 , y17721 , y17722 , y17723 , y17724 , y17725 , y17726 , y17727 , y17728 , y17729 , y17730 , y17731 , y17732 , y17733 , y17734 , y17735 , y17736 , y17737 , y17738 , y17739 , y17740 , y17741 , y17742 , y17743 , y17744 , y17745 , y17746 , y17747 , y17748 , y17749 , y17750 , y17751 , y17752 , y17753 , y17754 , y17755 , y17756 , y17757 , y17758 , y17759 , y17760 , y17761 , y17762 , y17763 , y17764 , y17765 , y17766 , y17767 , y17768 , y17769 , y17770 , y17771 , y17772 , y17773 , y17774 , y17775 , y17776 , y17777 , y17778 , y17779 , y17780 , y17781 , y17782 , y17783 , y17784 , y17785 , y17786 , y17787 , y17788 , y17789 , y17790 , y17791 , y17792 , y17793 , y17794 , y17795 , y17796 , y17797 , y17798 , y17799 , y17800 , y17801 , y17802 , y17803 , y17804 , y17805 , y17806 , y17807 , y17808 , y17809 , y17810 , y17811 , y17812 , y17813 , y17814 , y17815 , y17816 , y17817 , y17818 , y17819 , y17820 , y17821 , y17822 , y17823 , y17824 , y17825 , y17826 , y17827 , y17828 , y17829 , y17830 , y17831 , y17832 , y17833 , y17834 , y17835 , y17836 , y17837 , y17838 , y17839 , y17840 , y17841 , y17842 , y17843 , y17844 , y17845 , y17846 , y17847 , y17848 , y17849 , y17850 , y17851 , y17852 , y17853 , y17854 , y17855 , y17856 , y17857 , y17858 , y17859 , y17860 , y17861 , y17862 , y17863 , y17864 , y17865 , y17866 , y17867 , y17868 , y17869 , y17870 , y17871 , y17872 , y17873 , y17874 , y17875 , y17876 , y17877 , y17878 , y17879 , y17880 , y17881 , y17882 , y17883 , y17884 , y17885 , y17886 , y17887 , y17888 , y17889 , y17890 , y17891 , y17892 , y17893 , y17894 , y17895 , y17896 , y17897 , y17898 , y17899 , y17900 , y17901 , y17902 , y17903 , y17904 , y17905 , y17906 , y17907 , y17908 , y17909 , y17910 , y17911 , y17912 , y17913 , y17914 , y17915 , y17916 , y17917 , y17918 , y17919 , y17920 , y17921 , y17922 , y17923 , y17924 , y17925 , y17926 , y17927 , y17928 , y17929 , y17930 , y17931 , y17932 , y17933 , y17934 , y17935 , y17936 , y17937 , y17938 , y17939 , y17940 , y17941 , y17942 , y17943 , y17944 , y17945 , y17946 , y17947 , y17948 , y17949 , y17950 , y17951 , y17952 , y17953 , y17954 , y17955 , y17956 , y17957 , y17958 , y17959 , y17960 , y17961 , y17962 , y17963 , y17964 , y17965 , y17966 , y17967 , y17968 , y17969 , y17970 , y17971 , y17972 , y17973 , y17974 , y17975 , y17976 , y17977 , y17978 , y17979 , y17980 , y17981 , y17982 , y17983 , y17984 , y17985 , y17986 , y17987 , y17988 , y17989 , y17990 , y17991 , y17992 , y17993 , y17994 , y17995 , y17996 , y17997 , y17998 , y17999 , y18000 , y18001 , y18002 , y18003 , y18004 , y18005 , y18006 , y18007 , y18008 , y18009 , y18010 , y18011 , y18012 , y18013 , y18014 , y18015 , y18016 , y18017 , y18018 , y18019 , y18020 , y18021 , y18022 , y18023 , y18024 , y18025 , y18026 , y18027 , y18028 , y18029 , y18030 , y18031 , y18032 , y18033 , y18034 , y18035 , y18036 , y18037 , y18038 , y18039 , y18040 , y18041 , y18042 , y18043 , y18044 , y18045 , y18046 , y18047 , y18048 , y18049 , y18050 , y18051 , y18052 , y18053 , y18054 , y18055 , y18056 , y18057 , y18058 , y18059 , y18060 , y18061 , y18062 , y18063 , y18064 , y18065 , y18066 , y18067 , y18068 , y18069 , y18070 , y18071 , y18072 , y18073 , y18074 , y18075 , y18076 , y18077 , y18078 , y18079 , y18080 , y18081 , y18082 , y18083 , y18084 , y18085 , y18086 , y18087 , y18088 , y18089 , y18090 , y18091 , y18092 , y18093 , y18094 , y18095 , y18096 , y18097 , y18098 , y18099 , y18100 , y18101 , y18102 , y18103 , y18104 , y18105 , y18106 , y18107 , y18108 , y18109 , y18110 , y18111 , y18112 , y18113 , y18114 , y18115 , y18116 , y18117 , y18118 , y18119 , y18120 , y18121 , y18122 , y18123 , y18124 , y18125 , y18126 , y18127 , y18128 , y18129 , y18130 , y18131 , y18132 , y18133 , y18134 , y18135 , y18136 , y18137 , y18138 , y18139 , y18140 , y18141 , y18142 , y18143 , y18144 , y18145 , y18146 , y18147 , y18148 , y18149 , y18150 , y18151 , y18152 , y18153 , y18154 , y18155 , y18156 , y18157 , y18158 , y18159 , y18160 , y18161 , y18162 , y18163 , y18164 , y18165 , y18166 , y18167 , y18168 , y18169 , y18170 , y18171 , y18172 , y18173 , y18174 , y18175 , y18176 , y18177 , y18178 , y18179 , y18180 , y18181 , y18182 , y18183 , y18184 , y18185 , y18186 , y18187 , y18188 , y18189 , y18190 , y18191 , y18192 , y18193 , y18194 , y18195 , y18196 , y18197 , y18198 , y18199 , y18200 , y18201 , y18202 , y18203 , y18204 , y18205 , y18206 , y18207 , y18208 , y18209 , y18210 , y18211 , y18212 , y18213 , y18214 , y18215 , y18216 , y18217 , y18218 , y18219 , y18220 , y18221 , y18222 , y18223 , y18224 , y18225 , y18226 , y18227 , y18228 , y18229 , y18230 , y18231 , y18232 , y18233 , y18234 , y18235 , y18236 , y18237 , y18238 , y18239 , y18240 , y18241 , y18242 , y18243 , y18244 , y18245 , y18246 , y18247 , y18248 , y18249 , y18250 , y18251 , y18252 , y18253 , y18254 , y18255 , y18256 , y18257 , y18258 , y18259 , y18260 , y18261 , y18262 , y18263 , y18264 , y18265 , y18266 , y18267 , y18268 , y18269 , y18270 , y18271 , y18272 , y18273 , y18274 , y18275 , y18276 , y18277 , y18278 , y18279 , y18280 , y18281 , y18282 , y18283 , y18284 , y18285 , y18286 , y18287 , y18288 , y18289 , y18290 , y18291 , y18292 , y18293 , y18294 , y18295 , y18296 , y18297 , y18298 , y18299 , y18300 , y18301 , y18302 , y18303 , y18304 , y18305 , y18306 , y18307 , y18308 , y18309 , y18310 , y18311 , y18312 , y18313 , y18314 , y18315 , y18316 , y18317 , y18318 , y18319 , y18320 , y18321 , y18322 , y18323 , y18324 , y18325 , y18326 , y18327 , y18328 , y18329 , y18330 , y18331 , y18332 , y18333 , y18334 , y18335 , y18336 , y18337 , y18338 , y18339 , y18340 , y18341 , y18342 , y18343 , y18344 , y18345 , y18346 , y18347 , y18348 , y18349 , y18350 , y18351 , y18352 , y18353 , y18354 , y18355 , y18356 , y18357 , y18358 , y18359 , y18360 , y18361 , y18362 , y18363 , y18364 , y18365 , y18366 , y18367 , y18368 , y18369 , y18370 , y18371 , y18372 , y18373 , y18374 , y18375 , y18376 , y18377 , y18378 , y18379 , y18380 , y18381 , y18382 , y18383 , y18384 , y18385 , y18386 , y18387 , y18388 , y18389 , y18390 , y18391 , y18392 , y18393 , y18394 , y18395 , y18396 , y18397 , y18398 , y18399 , y18400 , y18401 , y18402 , y18403 , y18404 , y18405 , y18406 , y18407 , y18408 , y18409 , y18410 , y18411 , y18412 , y18413 , y18414 , y18415 , y18416 , y18417 , y18418 , y18419 , y18420 , y18421 , y18422 , y18423 , y18424 , y18425 , y18426 , y18427 , y18428 , y18429 , y18430 , y18431 , y18432 , y18433 , y18434 , y18435 , y18436 , y18437 , y18438 , y18439 , y18440 , y18441 , y18442 , y18443 , y18444 , y18445 , y18446 , y18447 , y18448 , y18449 , y18450 , y18451 , y18452 , y18453 , y18454 , y18455 , y18456 , y18457 , y18458 , y18459 , y18460 , y18461 , y18462 , y18463 , y18464 , y18465 , y18466 , y18467 , y18468 , y18469 , y18470 , y18471 , y18472 , y18473 , y18474 , y18475 , y18476 , y18477 , y18478 , y18479 , y18480 , y18481 , y18482 , y18483 , y18484 , y18485 , y18486 , y18487 , y18488 , y18489 , y18490 , y18491 , y18492 , y18493 , y18494 , y18495 , y18496 , y18497 , y18498 , y18499 , y18500 , y18501 , y18502 , y18503 , y18504 , y18505 , y18506 , y18507 , y18508 , y18509 , y18510 , y18511 , y18512 , y18513 , y18514 , y18515 , y18516 , y18517 , y18518 , y18519 , y18520 , y18521 , y18522 , y18523 , y18524 , y18525 , y18526 , y18527 , y18528 , y18529 , y18530 , y18531 , y18532 , y18533 , y18534 , y18535 , y18536 , y18537 , y18538 , y18539 , y18540 , y18541 , y18542 , y18543 , y18544 , y18545 , y18546 , y18547 , y18548 , y18549 , y18550 , y18551 , y18552 , y18553 , y18554 , y18555 , y18556 , y18557 , y18558 , y18559 , y18560 , y18561 , y18562 , y18563 , y18564 , y18565 , y18566 , y18567 , y18568 , y18569 , y18570 , y18571 , y18572 , y18573 , y18574 , y18575 , y18576 , y18577 , y18578 , y18579 , y18580 , y18581 , y18582 , y18583 , y18584 , y18585 , y18586 , y18587 , y18588 , y18589 , y18590 , y18591 , y18592 , y18593 , y18594 , y18595 , y18596 , y18597 , y18598 , y18599 , y18600 , y18601 , y18602 , y18603 , y18604 , y18605 , y18606 , y18607 , y18608 , y18609 , y18610 , y18611 , y18612 , y18613 , y18614 , y18615 , y18616 , y18617 , y18618 , y18619 , y18620 , y18621 , y18622 , y18623 , y18624 , y18625 , y18626 , y18627 , y18628 , y18629 , y18630 , y18631 , y18632 , y18633 , y18634 , y18635 , y18636 , y18637 , y18638 , y18639 , y18640 , y18641 , y18642 , y18643 , y18644 , y18645 , y18646 , y18647 , y18648 , y18649 , y18650 , y18651 , y18652 , y18653 , y18654 , y18655 , y18656 , y18657 , y18658 , y18659 , y18660 , y18661 , y18662 , y18663 , y18664 , y18665 , y18666 , y18667 , y18668 , y18669 , y18670 , y18671 , y18672 , y18673 , y18674 , y18675 , y18676 , y18677 , y18678 , y18679 , y18680 , y18681 , y18682 , y18683 , y18684 , y18685 , y18686 , y18687 , y18688 , y18689 , y18690 , y18691 , y18692 , y18693 , y18694 , y18695 , y18696 , y18697 , y18698 , y18699 , y18700 , y18701 , y18702 , y18703 , y18704 , y18705 , y18706 , y18707 , y18708 , y18709 , y18710 , y18711 , y18712 , y18713 , y18714 , y18715 , y18716 , y18717 , y18718 , y18719 , y18720 , y18721 , y18722 , y18723 , y18724 , y18725 , y18726 , y18727 , y18728 , y18729 , y18730 , y18731 , y18732 , y18733 , y18734 , y18735 , y18736 , y18737 , y18738 , y18739 , y18740 , y18741 , y18742 , y18743 , y18744 , y18745 , y18746 , y18747 , y18748 , y18749 , y18750 , y18751 , y18752 , y18753 , y18754 , y18755 , y18756 , y18757 , y18758 , y18759 , y18760 , y18761 , y18762 , y18763 , y18764 , y18765 , y18766 , y18767 , y18768 , y18769 , y18770 , y18771 , y18772 , y18773 , y18774 , y18775 , y18776 , y18777 , y18778 , y18779 , y18780 , y18781 , y18782 , y18783 , y18784 , y18785 , y18786 , y18787 , y18788 , y18789 , y18790 , y18791 , y18792 , y18793 , y18794 , y18795 , y18796 , y18797 , y18798 , y18799 , y18800 , y18801 , y18802 , y18803 , y18804 , y18805 , y18806 , y18807 , y18808 , y18809 , y18810 , y18811 , y18812 , y18813 , y18814 , y18815 , y18816 , y18817 , y18818 , y18819 , y18820 , y18821 , y18822 , y18823 , y18824 , y18825 , y18826 , y18827 , y18828 , y18829 , y18830 , y18831 , y18832 , y18833 , y18834 , y18835 , y18836 , y18837 , y18838 , y18839 , y18840 , y18841 , y18842 , y18843 , y18844 , y18845 , y18846 , y18847 , y18848 , y18849 , y18850 , y18851 , y18852 , y18853 , y18854 , y18855 , y18856 , y18857 , y18858 , y18859 , y18860 , y18861 , y18862 , y18863 , y18864 , y18865 , y18866 , y18867 , y18868 , y18869 , y18870 , y18871 , y18872 , y18873 , y18874 , y18875 , y18876 , y18877 , y18878 , y18879 , y18880 , y18881 , y18882 , y18883 , y18884 , y18885 , y18886 , y18887 , y18888 , y18889 , y18890 , y18891 , y18892 , y18893 , y18894 , y18895 , y18896 , y18897 , y18898 , y18899 , y18900 , y18901 , y18902 , y18903 , y18904 , y18905 , y18906 , y18907 , y18908 , y18909 , y18910 , y18911 , y18912 , y18913 , y18914 , y18915 , y18916 , y18917 , y18918 , y18919 , y18920 , y18921 , y18922 , y18923 , y18924 , y18925 , y18926 , y18927 , y18928 , y18929 , y18930 , y18931 , y18932 , y18933 , y18934 , y18935 , y18936 , y18937 , y18938 , y18939 , y18940 , y18941 , y18942 , y18943 , y18944 , y18945 , y18946 , y18947 , y18948 , y18949 , y18950 , y18951 , y18952 , y18953 , y18954 , y18955 , y18956 , y18957 , y18958 , y18959 , y18960 , y18961 , y18962 , y18963 , y18964 , y18965 , y18966 , y18967 , y18968 , y18969 , y18970 , y18971 , y18972 , y18973 , y18974 , y18975 , y18976 , y18977 , y18978 , y18979 , y18980 , y18981 , y18982 , y18983 , y18984 , y18985 , y18986 , y18987 , y18988 , y18989 , y18990 , y18991 , y18992 , y18993 , y18994 , y18995 , y18996 , y18997 , y18998 , y18999 , y19000 , y19001 , y19002 , y19003 , y19004 , y19005 , y19006 , y19007 , y19008 , y19009 , y19010 , y19011 , y19012 , y19013 , y19014 , y19015 , y19016 , y19017 , y19018 , y19019 , y19020 , y19021 , y19022 , y19023 , y19024 , y19025 , y19026 , y19027 , y19028 , y19029 , y19030 , y19031 , y19032 , y19033 , y19034 , y19035 , y19036 , y19037 , y19038 , y19039 , y19040 , y19041 , y19042 , y19043 , y19044 , y19045 , y19046 , y19047 , y19048 , y19049 , y19050 , y19051 , y19052 , y19053 , y19054 , y19055 , y19056 , y19057 , y19058 , y19059 , y19060 , y19061 , y19062 , y19063 , y19064 , y19065 , y19066 , y19067 , y19068 , y19069 , y19070 , y19071 , y19072 , y19073 , y19074 , y19075 , y19076 , y19077 , y19078 , y19079 , y19080 , y19081 , y19082 , y19083 , y19084 , y19085 , y19086 , y19087 , y19088 , y19089 , y19090 , y19091 , y19092 , y19093 , y19094 , y19095 , y19096 , y19097 , y19098 , y19099 , y19100 , y19101 , y19102 , y19103 , y19104 , y19105 , y19106 , y19107 , y19108 , y19109 , y19110 , y19111 , y19112 , y19113 , y19114 , y19115 , y19116 , y19117 , y19118 , y19119 , y19120 , y19121 , y19122 , y19123 , y19124 , y19125 , y19126 , y19127 , y19128 , y19129 , y19130 , y19131 , y19132 , y19133 , y19134 , y19135 , y19136 , y19137 , y19138 , y19139 , y19140 , y19141 , y19142 , y19143 , y19144 , y19145 , y19146 , y19147 , y19148 , y19149 , y19150 , y19151 , y19152 , y19153 , y19154 , y19155 , y19156 , y19157 , y19158 , y19159 , y19160 , y19161 , y19162 , y19163 , y19164 , y19165 , y19166 , y19167 , y19168 , y19169 , y19170 , y19171 , y19172 , y19173 , y19174 , y19175 , y19176 , y19177 , y19178 , y19179 , y19180 , y19181 , y19182 , y19183 , y19184 , y19185 , y19186 , y19187 , y19188 , y19189 , y19190 , y19191 , y19192 , y19193 , y19194 , y19195 , y19196 , y19197 , y19198 , y19199 , y19200 , y19201 , y19202 , y19203 , y19204 , y19205 , y19206 , y19207 , y19208 , y19209 , y19210 , y19211 , y19212 , y19213 , y19214 , y19215 , y19216 , y19217 , y19218 , y19219 , y19220 , y19221 , y19222 , y19223 , y19224 , y19225 , y19226 , y19227 , y19228 , y19229 , y19230 , y19231 , y19232 , y19233 , y19234 , y19235 , y19236 , y19237 , y19238 , y19239 , y19240 , y19241 , y19242 , y19243 , y19244 , y19245 , y19246 , y19247 , y19248 , y19249 , y19250 , y19251 , y19252 , y19253 , y19254 , y19255 , y19256 , y19257 , y19258 , y19259 , y19260 , y19261 , y19262 , y19263 , y19264 , y19265 , y19266 , y19267 , y19268 , y19269 , y19270 , y19271 , y19272 , y19273 , y19274 , y19275 , y19276 , y19277 , y19278 , y19279 , y19280 , y19281 , y19282 , y19283 , y19284 , y19285 , y19286 , y19287 , y19288 , y19289 , y19290 , y19291 , y19292 , y19293 , y19294 , y19295 , y19296 , y19297 , y19298 , y19299 , y19300 , y19301 , y19302 , y19303 , y19304 , y19305 , y19306 , y19307 , y19308 , y19309 , y19310 , y19311 , y19312 , y19313 , y19314 , y19315 , y19316 , y19317 , y19318 , y19319 , y19320 , y19321 , y19322 , y19323 , y19324 , y19325 , y19326 , y19327 , y19328 , y19329 , y19330 , y19331 , y19332 , y19333 , y19334 , y19335 , y19336 , y19337 , y19338 , y19339 , y19340 , y19341 , y19342 , y19343 , y19344 , y19345 , y19346 , y19347 , y19348 , y19349 , y19350 , y19351 , y19352 , y19353 , y19354 , y19355 , y19356 , y19357 , y19358 , y19359 , y19360 , y19361 , y19362 , y19363 , y19364 , y19365 , y19366 , y19367 , y19368 , y19369 , y19370 , y19371 , y19372 , y19373 , y19374 , y19375 , y19376 , y19377 , y19378 , y19379 , y19380 , y19381 , y19382 , y19383 , y19384 , y19385 , y19386 , y19387 , y19388 , y19389 , y19390 , y19391 , y19392 , y19393 , y19394 , y19395 , y19396 , y19397 , y19398 , y19399 , y19400 , y19401 , y19402 , y19403 , y19404 , y19405 , y19406 , y19407 , y19408 , y19409 , y19410 , y19411 , y19412 , y19413 , y19414 , y19415 , y19416 , y19417 , y19418 , y19419 , y19420 , y19421 , y19422 , y19423 , y19424 , y19425 , y19426 , y19427 , y19428 , y19429 , y19430 , y19431 , y19432 , y19433 , y19434 , y19435 , y19436 , y19437 , y19438 , y19439 , y19440 , y19441 , y19442 , y19443 , y19444 , y19445 , y19446 , y19447 , y19448 , y19449 , y19450 , y19451 , y19452 , y19453 , y19454 , y19455 , y19456 , y19457 , y19458 , y19459 , y19460 , y19461 , y19462 , y19463 , y19464 , y19465 , y19466 , y19467 , y19468 , y19469 , y19470 , y19471 , y19472 , y19473 , y19474 , y19475 , y19476 , y19477 , y19478 , y19479 , y19480 , y19481 , y19482 , y19483 , y19484 , y19485 , y19486 , y19487 , y19488 , y19489 , y19490 , y19491 , y19492 , y19493 , y19494 , y19495 , y19496 , y19497 , y19498 , y19499 , y19500 , y19501 , y19502 , y19503 , y19504 , y19505 , y19506 , y19507 , y19508 , y19509 , y19510 , y19511 , y19512 , y19513 , y19514 , y19515 , y19516 , y19517 , y19518 , y19519 , y19520 , y19521 , y19522 , y19523 , y19524 , y19525 , y19526 , y19527 , y19528 , y19529 , y19530 , y19531 , y19532 , y19533 , y19534 , y19535 , y19536 , y19537 , y19538 , y19539 , y19540 , y19541 , y19542 , y19543 , y19544 , y19545 , y19546 , y19547 , y19548 , y19549 , y19550 , y19551 , y19552 , y19553 , y19554 , y19555 , y19556 , y19557 , y19558 , y19559 , y19560 , y19561 , y19562 , y19563 , y19564 , y19565 , y19566 , y19567 , y19568 , y19569 , y19570 , y19571 , y19572 , y19573 , y19574 , y19575 , y19576 , y19577 , y19578 , y19579 , y19580 , y19581 , y19582 , y19583 , y19584 , y19585 , y19586 , y19587 , y19588 , y19589 , y19590 , y19591 , y19592 , y19593 , y19594 , y19595 , y19596 , y19597 , y19598 , y19599 , y19600 , y19601 , y19602 , y19603 , y19604 , y19605 , y19606 , y19607 , y19608 , y19609 , y19610 , y19611 , y19612 , y19613 , y19614 , y19615 , y19616 , y19617 , y19618 , y19619 , y19620 , y19621 , y19622 , y19623 , y19624 , y19625 , y19626 , y19627 , y19628 , y19629 , y19630 , y19631 , y19632 , y19633 , y19634 , y19635 , y19636 , y19637 , y19638 , y19639 , y19640 , y19641 , y19642 , y19643 , y19644 , y19645 , y19646 , y19647 , y19648 , y19649 , y19650 , y19651 , y19652 , y19653 , y19654 , y19655 , y19656 , y19657 , y19658 , y19659 , y19660 , y19661 , y19662 , y19663 , y19664 , y19665 , y19666 , y19667 , y19668 , y19669 , y19670 , y19671 , y19672 , y19673 , y19674 , y19675 , y19676 , y19677 , y19678 , y19679 , y19680 , y19681 , y19682 , y19683 , y19684 , y19685 , y19686 , y19687 , y19688 , y19689 , y19690 , y19691 , y19692 , y19693 , y19694 , y19695 , y19696 , y19697 , y19698 , y19699 , y19700 , y19701 , y19702 , y19703 , y19704 , y19705 , y19706 , y19707 , y19708 , y19709 , y19710 , y19711 , y19712 , y19713 , y19714 , y19715 , y19716 , y19717 , y19718 , y19719 , y19720 , y19721 , y19722 , y19723 , y19724 , y19725 , y19726 , y19727 , y19728 , y19729 , y19730 , y19731 , y19732 , y19733 , y19734 , y19735 , y19736 , y19737 , y19738 , y19739 , y19740 , y19741 , y19742 , y19743 , y19744 , y19745 , y19746 , y19747 , y19748 , y19749 , y19750 , y19751 , y19752 , y19753 , y19754 , y19755 , y19756 , y19757 , y19758 , y19759 , y19760 , y19761 , y19762 , y19763 , y19764 , y19765 , y19766 , y19767 , y19768 , y19769 , y19770 , y19771 , y19772 , y19773 , y19774 , y19775 , y19776 , y19777 , y19778 , y19779 , y19780 , y19781 , y19782 , y19783 , y19784 , y19785 , y19786 , y19787 , y19788 , y19789 , y19790 , y19791 , y19792 , y19793 , y19794 , y19795 , y19796 , y19797 , y19798 , y19799 , y19800 , y19801 , y19802 , y19803 , y19804 , y19805 , y19806 , y19807 , y19808 , y19809 , y19810 , y19811 , y19812 , y19813 , y19814 , y19815 , y19816 , y19817 , y19818 , y19819 , y19820 , y19821 , y19822 , y19823 , y19824 , y19825 , y19826 , y19827 , y19828 , y19829 , y19830 , y19831 , y19832 , y19833 , y19834 , y19835 , y19836 , y19837 , y19838 , y19839 , y19840 , y19841 , y19842 , y19843 , y19844 , y19845 , y19846 , y19847 , y19848 , y19849 , y19850 , y19851 , y19852 , y19853 , y19854 , y19855 , y19856 , y19857 , y19858 , y19859 , y19860 , y19861 , y19862 , y19863 , y19864 , y19865 , y19866 , y19867 , y19868 , y19869 , y19870 , y19871 , y19872 , y19873 , y19874 , y19875 , y19876 , y19877 , y19878 , y19879 , y19880 , y19881 , y19882 , y19883 , y19884 , y19885 , y19886 , y19887 , y19888 , y19889 , y19890 , y19891 , y19892 , y19893 , y19894 , y19895 , y19896 , y19897 , y19898 , y19899 , y19900 , y19901 , y19902 , y19903 , y19904 , y19905 , y19906 , y19907 , y19908 , y19909 , y19910 , y19911 , y19912 , y19913 , y19914 , y19915 , y19916 , y19917 , y19918 , y19919 , y19920 , y19921 , y19922 , y19923 , y19924 , y19925 , y19926 , y19927 , y19928 , y19929 , y19930 , y19931 , y19932 , y19933 , y19934 , y19935 , y19936 , y19937 , y19938 , y19939 , y19940 , y19941 , y19942 , y19943 , y19944 , y19945 , y19946 , y19947 , y19948 , y19949 , y19950 , y19951 , y19952 , y19953 , y19954 , y19955 , y19956 , y19957 , y19958 , y19959 , y19960 , y19961 , y19962 , y19963 , y19964 , y19965 , y19966 , y19967 , y19968 , y19969 , y19970 , y19971 , y19972 , y19973 , y19974 , y19975 , y19976 , y19977 , y19978 , y19979 , y19980 , y19981 , y19982 , y19983 , y19984 , y19985 , y19986 , y19987 , y19988 , y19989 , y19990 , y19991 , y19992 , y19993 , y19994 , y19995 , y19996 , y19997 , y19998 , y19999 , y20000 , y20001 , y20002 , y20003 , y20004 , y20005 , y20006 , y20007 , y20008 , y20009 , y20010 , y20011 , y20012 , y20013 , y20014 , y20015 , y20016 , y20017 , y20018 , y20019 , y20020 , y20021 , y20022 , y20023 , y20024 , y20025 , y20026 , y20027 , y20028 , y20029 , y20030 , y20031 , y20032 , y20033 , y20034 , y20035 , y20036 , y20037 , y20038 , y20039 , y20040 , y20041 , y20042 , y20043 , y20044 , y20045 , y20046 , y20047 , y20048 , y20049 , y20050 , y20051 , y20052 , y20053 , y20054 , y20055 , y20056 , y20057 , y20058 , y20059 , y20060 , y20061 , y20062 , y20063 , y20064 , y20065 , y20066 , y20067 , y20068 , y20069 , y20070 , y20071 , y20072 , y20073 , y20074 , y20075 , y20076 , y20077 , y20078 , y20079 , y20080 , y20081 , y20082 , y20083 , y20084 , y20085 , y20086 , y20087 , y20088 , y20089 , y20090 , y20091 , y20092 , y20093 , y20094 , y20095 , y20096 , y20097 , y20098 , y20099 , y20100 , y20101 , y20102 , y20103 , y20104 , y20105 , y20106 , y20107 , y20108 , y20109 , y20110 , y20111 , y20112 , y20113 , y20114 , y20115 , y20116 , y20117 , y20118 , y20119 , y20120 , y20121 , y20122 , y20123 , y20124 , y20125 , y20126 , y20127 , y20128 , y20129 , y20130 , y20131 , y20132 , y20133 , y20134 , y20135 , y20136 , y20137 , y20138 , y20139 , y20140 , y20141 , y20142 , y20143 , y20144 , y20145 , y20146 , y20147 , y20148 , y20149 , y20150 , y20151 , y20152 , y20153 , y20154 , y20155 , y20156 , y20157 , y20158 , y20159 , y20160 , y20161 , y20162 , y20163 , y20164 , y20165 , y20166 , y20167 , y20168 , y20169 , y20170 , y20171 , y20172 , y20173 , y20174 , y20175 , y20176 , y20177 , y20178 , y20179 , y20180 , y20181 , y20182 , y20183 , y20184 , y20185 , y20186 , y20187 , y20188 , y20189 , y20190 , y20191 , y20192 , y20193 , y20194 , y20195 , y20196 , y20197 , y20198 , y20199 , y20200 , y20201 , y20202 , y20203 , y20204 , y20205 , y20206 , y20207 , y20208 , y20209 , y20210 , y20211 , y20212 , y20213 , y20214 , y20215 , y20216 , y20217 , y20218 , y20219 , y20220 , y20221 , y20222 , y20223 , y20224 , y20225 , y20226 , y20227 , y20228 , y20229 , y20230 , y20231 , y20232 , y20233 , y20234 , y20235 , y20236 , y20237 , y20238 , y20239 , y20240 , y20241 , y20242 , y20243 , y20244 , y20245 , y20246 , y20247 , y20248 , y20249 , y20250 , y20251 , y20252 , y20253 , y20254 , y20255 , y20256 , y20257 , y20258 , y20259 , y20260 , y20261 , y20262 , y20263 , y20264 , y20265 , y20266 , y20267 , y20268 , y20269 , y20270 , y20271 , y20272 , y20273 , y20274 , y20275 , y20276 , y20277 , y20278 , y20279 , y20280 , y20281 , y20282 , y20283 , y20284 , y20285 , y20286 , y20287 , y20288 , y20289 , y20290 , y20291 , y20292 , y20293 , y20294 , y20295 , y20296 , y20297 , y20298 , y20299 , y20300 , y20301 , y20302 , y20303 , y20304 , y20305 , y20306 , y20307 , y20308 , y20309 , y20310 , y20311 , y20312 , y20313 , y20314 , y20315 , y20316 , y20317 , y20318 , y20319 , y20320 , y20321 , y20322 , y20323 , y20324 , y20325 , y20326 , y20327 , y20328 , y20329 , y20330 , y20331 , y20332 , y20333 , y20334 , y20335 , y20336 , y20337 , y20338 , y20339 , y20340 , y20341 , y20342 , y20343 , y20344 , y20345 , y20346 , y20347 , y20348 , y20349 , y20350 , y20351 , y20352 , y20353 , y20354 , y20355 , y20356 , y20357 , y20358 , y20359 , y20360 , y20361 , y20362 , y20363 , y20364 , y20365 , y20366 , y20367 , y20368 , y20369 , y20370 , y20371 , y20372 , y20373 , y20374 , y20375 , y20376 , y20377 , y20378 , y20379 , y20380 , y20381 , y20382 , y20383 , y20384 , y20385 , y20386 , y20387 , y20388 , y20389 , y20390 , y20391 , y20392 , y20393 , y20394 , y20395 , y20396 , y20397 , y20398 , y20399 , y20400 , y20401 , y20402 , y20403 , y20404 , y20405 , y20406 , y20407 , y20408 , y20409 , y20410 , y20411 , y20412 , y20413 , y20414 , y20415 , y20416 , y20417 , y20418 , y20419 , y20420 , y20421 , y20422 , y20423 , y20424 , y20425 , y20426 , y20427 , y20428 , y20429 , y20430 , y20431 , y20432 , y20433 , y20434 , y20435 , y20436 , y20437 , y20438 , y20439 , y20440 , y20441 , y20442 , y20443 , y20444 , y20445 , y20446 , y20447 , y20448 , y20449 , y20450 , y20451 , y20452 , y20453 , y20454 , y20455 , y20456 , y20457 , y20458 , y20459 , y20460 , y20461 , y20462 , y20463 , y20464 , y20465 , y20466 , y20467 , y20468 , y20469 , y20470 , y20471 , y20472 , y20473 , y20474 , y20475 , y20476 , y20477 , y20478 , y20479 , y20480 , y20481 , y20482 , y20483 , y20484 , y20485 , y20486 , y20487 , y20488 , y20489 , y20490 , y20491 , y20492 , y20493 , y20494 , y20495 , y20496 , y20497 , y20498 , y20499 , y20500 , y20501 , y20502 , y20503 , y20504 , y20505 , y20506 , y20507 , y20508 , y20509 , y20510 , y20511 , y20512 , y20513 , y20514 , y20515 , y20516 , y20517 , y20518 , y20519 , y20520 , y20521 , y20522 , y20523 , y20524 , y20525 , y20526 , y20527 , y20528 , y20529 , y20530 , y20531 , y20532 , y20533 , y20534 , y20535 , y20536 , y20537 , y20538 , y20539 , y20540 , y20541 , y20542 , y20543 , y20544 , y20545 , y20546 , y20547 , y20548 , y20549 , y20550 , y20551 , y20552 , y20553 , y20554 , y20555 , y20556 , y20557 , y20558 , y20559 , y20560 , y20561 , y20562 , y20563 , y20564 , y20565 , y20566 , y20567 , y20568 , y20569 , y20570 , y20571 , y20572 , y20573 , y20574 , y20575 , y20576 , y20577 , y20578 , y20579 , y20580 , y20581 , y20582 , y20583 , y20584 , y20585 , y20586 , y20587 , y20588 , y20589 , y20590 , y20591 , y20592 , y20593 , y20594 , y20595 , y20596 , y20597 , y20598 , y20599 , y20600 , y20601 , y20602 , y20603 , y20604 , y20605 , y20606 , y20607 , y20608 , y20609 , y20610 , y20611 , y20612 , y20613 , y20614 , y20615 , y20616 , y20617 , y20618 , y20619 , y20620 , y20621 , y20622 , y20623 , y20624 , y20625 , y20626 , y20627 , y20628 , y20629 , y20630 , y20631 , y20632 , y20633 , y20634 , y20635 , y20636 , y20637 , y20638 , y20639 , y20640 , y20641 , y20642 , y20643 , y20644 , y20645 , y20646 , y20647 , y20648 , y20649 , y20650 , y20651 , y20652 , y20653 , y20654 , y20655 , y20656 , y20657 , y20658 , y20659 , y20660 , y20661 , y20662 , y20663 , y20664 , y20665 , y20666 , y20667 , y20668 , y20669 , y20670 , y20671 , y20672 , y20673 , y20674 , y20675 , y20676 , y20677 , y20678 , y20679 , y20680 , y20681 , y20682 , y20683 , y20684 , y20685 , y20686 , y20687 , y20688 , y20689 , y20690 , y20691 , y20692 , y20693 , y20694 , y20695 , y20696 , y20697 , y20698 , y20699 , y20700 , y20701 , y20702 , y20703 , y20704 , y20705 , y20706 , y20707 , y20708 , y20709 , y20710 , y20711 , y20712 , y20713 , y20714 , y20715 , y20716 , y20717 , y20718 , y20719 , y20720 , y20721 , y20722 , y20723 , y20724 , y20725 , y20726 , y20727 , y20728 , y20729 , y20730 , y20731 , y20732 , y20733 , y20734 , y20735 , y20736 , y20737 , y20738 , y20739 , y20740 , y20741 , y20742 , y20743 , y20744 , y20745 , y20746 , y20747 , y20748 , y20749 , y20750 , y20751 , y20752 , y20753 , y20754 , y20755 , y20756 , y20757 , y20758 , y20759 , y20760 , y20761 , y20762 , y20763 , y20764 , y20765 , y20766 , y20767 , y20768 , y20769 , y20770 , y20771 , y20772 , y20773 , y20774 , y20775 , y20776 , y20777 , y20778 , y20779 , y20780 , y20781 , y20782 , y20783 , y20784 , y20785 , y20786 , y20787 , y20788 , y20789 , y20790 , y20791 , y20792 , y20793 , y20794 , y20795 , y20796 , y20797 , y20798 , y20799 , y20800 , y20801 , y20802 , y20803 , y20804 , y20805 , y20806 , y20807 , y20808 , y20809 , y20810 , y20811 , y20812 , y20813 , y20814 , y20815 , y20816 , y20817 , y20818 , y20819 , y20820 , y20821 , y20822 , y20823 , y20824 , y20825 , y20826 , y20827 , y20828 , y20829 , y20830 , y20831 , y20832 , y20833 , y20834 , y20835 , y20836 , y20837 , y20838 , y20839 , y20840 , y20841 , y20842 , y20843 , y20844 , y20845 , y20846 , y20847 , y20848 , y20849 , y20850 , y20851 , y20852 , y20853 , y20854 , y20855 , y20856 , y20857 , y20858 , y20859 , y20860 , y20861 , y20862 , y20863 , y20864 , y20865 , y20866 , y20867 , y20868 , y20869 , y20870 , y20871 , y20872 , y20873 , y20874 , y20875 , y20876 , y20877 , y20878 , y20879 , y20880 , y20881 , y20882 , y20883 , y20884 , y20885 , y20886 , y20887 , y20888 , y20889 , y20890 , y20891 , y20892 , y20893 , y20894 , y20895 , y20896 , y20897 , y20898 , y20899 , y20900 , y20901 , y20902 , y20903 , y20904 , y20905 , y20906 , y20907 , y20908 , y20909 , y20910 , y20911 , y20912 , y20913 , y20914 , y20915 , y20916 , y20917 , y20918 , y20919 , y20920 , y20921 , y20922 , y20923 , y20924 , y20925 , y20926 , y20927 , y20928 , y20929 , y20930 , y20931 , y20932 , y20933 , y20934 , y20935 , y20936 , y20937 , y20938 , y20939 , y20940 , y20941 , y20942 , y20943 , y20944 , y20945 , y20946 , y20947 , y20948 , y20949 , y20950 , y20951 , y20952 , y20953 , y20954 , y20955 , y20956 , y20957 , y20958 , y20959 , y20960 , y20961 , y20962 , y20963 , y20964 , y20965 , y20966 , y20967 , y20968 , y20969 , y20970 , y20971 , y20972 , y20973 , y20974 , y20975 , y20976 , y20977 , y20978 , y20979 , y20980 , y20981 , y20982 , y20983 , y20984 , y20985 , y20986 , y20987 , y20988 , y20989 , y20990 , y20991 , y20992 , y20993 , y20994 , y20995 , y20996 , y20997 , y20998 , y20999 , y21000 , y21001 , y21002 , y21003 , y21004 , y21005 , y21006 , y21007 , y21008 , y21009 , y21010 , y21011 , y21012 , y21013 , y21014 , y21015 , y21016 , y21017 , y21018 , y21019 , y21020 , y21021 , y21022 , y21023 , y21024 , y21025 , y21026 , y21027 , y21028 , y21029 , y21030 , y21031 , y21032 , y21033 , y21034 , y21035 , y21036 , y21037 , y21038 , y21039 , y21040 , y21041 , y21042 , y21043 , y21044 , y21045 , y21046 , y21047 , y21048 , y21049 , y21050 , y21051 , y21052 , y21053 , y21054 , y21055 , y21056 , y21057 , y21058 , y21059 , y21060 , y21061 , y21062 , y21063 , y21064 , y21065 , y21066 , y21067 , y21068 , y21069 , y21070 , y21071 , y21072 , y21073 , y21074 , y21075 , y21076 , y21077 , y21078 , y21079 , y21080 , y21081 , y21082 , y21083 , y21084 , y21085 , y21086 , y21087 , y21088 , y21089 , y21090 , y21091 , y21092 , y21093 , y21094 , y21095 , y21096 , y21097 , y21098 , y21099 , y21100 , y21101 , y21102 , y21103 , y21104 , y21105 , y21106 , y21107 , y21108 , y21109 , y21110 , y21111 , y21112 , y21113 , y21114 , y21115 , y21116 , y21117 , y21118 , y21119 , y21120 , y21121 , y21122 , y21123 , y21124 , y21125 , y21126 , y21127 , y21128 , y21129 , y21130 , y21131 , y21132 , y21133 , y21134 , y21135 , y21136 , y21137 , y21138 , y21139 , y21140 , y21141 , y21142 , y21143 , y21144 , y21145 , y21146 , y21147 , y21148 , y21149 , y21150 , y21151 , y21152 , y21153 , y21154 , y21155 , y21156 , y21157 , y21158 , y21159 , y21160 , y21161 , y21162 , y21163 , y21164 , y21165 , y21166 , y21167 , y21168 , y21169 , y21170 , y21171 , y21172 , y21173 , y21174 , y21175 , y21176 , y21177 , y21178 , y21179 , y21180 , y21181 , y21182 , y21183 , y21184 , y21185 , y21186 , y21187 , y21188 , y21189 , y21190 , y21191 , y21192 , y21193 , y21194 , y21195 , y21196 , y21197 , y21198 , y21199 , y21200 , y21201 , y21202 , y21203 , y21204 , y21205 , y21206 , y21207 , y21208 , y21209 , y21210 , y21211 , y21212 , y21213 , y21214 , y21215 , y21216 , y21217 , y21218 , y21219 , y21220 , y21221 , y21222 , y21223 , y21224 , y21225 , y21226 , y21227 , y21228 , y21229 , y21230 , y21231 , y21232 , y21233 , y21234 , y21235 , y21236 , y21237 , y21238 , y21239 , y21240 , y21241 , y21242 , y21243 , y21244 , y21245 , y21246 , y21247 , y21248 , y21249 , y21250 , y21251 , y21252 , y21253 , y21254 , y21255 , y21256 , y21257 , y21258 , y21259 , y21260 , y21261 , y21262 , y21263 , y21264 , y21265 , y21266 , y21267 , y21268 , y21269 , y21270 , y21271 , y21272 , y21273 , y21274 , y21275 , y21276 , y21277 , y21278 , y21279 , y21280 , y21281 , y21282 , y21283 , y21284 , y21285 , y21286 , y21287 , y21288 , y21289 , y21290 , y21291 , y21292 , y21293 , y21294 , y21295 , y21296 , y21297 , y21298 , y21299 , y21300 , y21301 , y21302 , y21303 , y21304 , y21305 , y21306 , y21307 , y21308 , y21309 , y21310 , y21311 , y21312 , y21313 , y21314 , y21315 , y21316 , y21317 , y21318 , y21319 , y21320 , y21321 , y21322 , y21323 , y21324 , y21325 , y21326 , y21327 , y21328 , y21329 , y21330 , y21331 , y21332 , y21333 , y21334 , y21335 , y21336 , y21337 , y21338 , y21339 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 , y15409 , y15410 , y15411 , y15412 , y15413 , y15414 , y15415 , y15416 , y15417 , y15418 , y15419 , y15420 , y15421 , y15422 , y15423 , y15424 , y15425 , y15426 , y15427 , y15428 , y15429 , y15430 , y15431 , y15432 , y15433 , y15434 , y15435 , y15436 , y15437 , y15438 , y15439 , y15440 , y15441 , y15442 , y15443 , y15444 , y15445 , y15446 , y15447 , y15448 , y15449 , y15450 , y15451 , y15452 , y15453 , y15454 , y15455 , y15456 , y15457 , y15458 , y15459 , y15460 , y15461 , y15462 , y15463 , y15464 , y15465 , y15466 , y15467 , y15468 , y15469 , y15470 , y15471 , y15472 , y15473 , y15474 , y15475 , y15476 , y15477 , y15478 , y15479 , y15480 , y15481 , y15482 , y15483 , y15484 , y15485 , y15486 , y15487 , y15488 , y15489 , y15490 , y15491 , y15492 , y15493 , y15494 , y15495 , y15496 , y15497 , y15498 , y15499 , y15500 , y15501 , y15502 , y15503 , y15504 , y15505 , y15506 , y15507 , y15508 , y15509 , y15510 , y15511 , y15512 , y15513 , y15514 , y15515 , y15516 , y15517 , y15518 , y15519 , y15520 , y15521 , y15522 , y15523 , y15524 , y15525 , y15526 , y15527 , y15528 , y15529 , y15530 , y15531 , y15532 , y15533 , y15534 , y15535 , y15536 , y15537 , y15538 , y15539 , y15540 , y15541 , y15542 , y15543 , y15544 , y15545 , y15546 , y15547 , y15548 , y15549 , y15550 , y15551 , y15552 , y15553 , y15554 , y15555 , y15556 , y15557 , y15558 , y15559 , y15560 , y15561 , y15562 , y15563 , y15564 , y15565 , y15566 , y15567 , y15568 , y15569 , y15570 , y15571 , y15572 , y15573 , y15574 , y15575 , y15576 , y15577 , y15578 , y15579 , y15580 , y15581 , y15582 , y15583 , y15584 , y15585 , y15586 , y15587 , y15588 , y15589 , y15590 , y15591 , y15592 , y15593 , y15594 , y15595 , y15596 , y15597 , y15598 , y15599 , y15600 , y15601 , y15602 , y15603 , y15604 , y15605 , y15606 , y15607 , y15608 , y15609 , y15610 , y15611 , y15612 , y15613 , y15614 , y15615 , y15616 , y15617 , y15618 , y15619 , y15620 , y15621 , y15622 , y15623 , y15624 , y15625 , y15626 , y15627 , y15628 , y15629 , y15630 , y15631 , y15632 , y15633 , y15634 , y15635 , y15636 , y15637 , y15638 , y15639 , y15640 , y15641 , y15642 , y15643 , y15644 , y15645 , y15646 , y15647 , y15648 , y15649 , y15650 , y15651 , y15652 , y15653 , y15654 , y15655 , y15656 , y15657 , y15658 , y15659 , y15660 , y15661 , y15662 , y15663 , y15664 , y15665 , y15666 , y15667 , y15668 , y15669 , y15670 , y15671 , y15672 , y15673 , y15674 , y15675 , y15676 , y15677 , y15678 , y15679 , y15680 , y15681 , y15682 , y15683 , y15684 , y15685 , y15686 , y15687 , y15688 , y15689 , y15690 , y15691 , y15692 , y15693 , y15694 , y15695 , y15696 , y15697 , y15698 , y15699 , y15700 , y15701 , y15702 , y15703 , y15704 , y15705 , y15706 , y15707 , y15708 , y15709 , y15710 , y15711 , y15712 , y15713 , y15714 , y15715 , y15716 , y15717 , y15718 , y15719 , y15720 , y15721 , y15722 , y15723 , y15724 , y15725 , y15726 , y15727 , y15728 , y15729 , y15730 , y15731 , y15732 , y15733 , y15734 , y15735 , y15736 , y15737 , y15738 , y15739 , y15740 , y15741 , y15742 , y15743 , y15744 , y15745 , y15746 , y15747 , y15748 , y15749 , y15750 , y15751 , y15752 , y15753 , y15754 , y15755 , y15756 , y15757 , y15758 , y15759 , y15760 , y15761 , y15762 , y15763 , y15764 , y15765 , y15766 , y15767 , y15768 , y15769 , y15770 , y15771 , y15772 , y15773 , y15774 , y15775 , y15776 , y15777 , y15778 , y15779 , y15780 , y15781 , y15782 , y15783 , y15784 , y15785 , y15786 , y15787 , y15788 , y15789 , y15790 , y15791 , y15792 , y15793 , y15794 , y15795 , y15796 , y15797 , y15798 , y15799 , y15800 , y15801 , y15802 , y15803 , y15804 , y15805 , y15806 , y15807 , y15808 , y15809 , y15810 , y15811 , y15812 , y15813 , y15814 , y15815 , y15816 , y15817 , y15818 , y15819 , y15820 , y15821 , y15822 , y15823 , y15824 , y15825 , y15826 , y15827 , y15828 , y15829 , y15830 , y15831 , y15832 , y15833 , y15834 , y15835 , y15836 , y15837 , y15838 , y15839 , y15840 , y15841 , y15842 , y15843 , y15844 , y15845 , y15846 , y15847 , y15848 , y15849 , y15850 , y15851 , y15852 , y15853 , y15854 , y15855 , y15856 , y15857 , y15858 , y15859 , y15860 , y15861 , y15862 , y15863 , y15864 , y15865 , y15866 , y15867 , y15868 , y15869 , y15870 , y15871 , y15872 , y15873 , y15874 , y15875 , y15876 , y15877 , y15878 , y15879 , y15880 , y15881 , y15882 , y15883 , y15884 , y15885 , y15886 , y15887 , y15888 , y15889 , y15890 , y15891 , y15892 , y15893 , y15894 , y15895 , y15896 , y15897 , y15898 , y15899 , y15900 , y15901 , y15902 , y15903 , y15904 , y15905 , y15906 , y15907 , y15908 , y15909 , y15910 , y15911 , y15912 , y15913 , y15914 , y15915 , y15916 , y15917 , y15918 , y15919 , y15920 , y15921 , y15922 , y15923 , y15924 , y15925 , y15926 , y15927 , y15928 , y15929 , y15930 , y15931 , y15932 , y15933 , y15934 , y15935 , y15936 , y15937 , y15938 , y15939 , y15940 , y15941 , y15942 , y15943 , y15944 , y15945 , y15946 , y15947 , y15948 , y15949 , y15950 , y15951 , y15952 , y15953 , y15954 , y15955 , y15956 , y15957 , y15958 , y15959 , y15960 , y15961 , y15962 , y15963 , y15964 , y15965 , y15966 , y15967 , y15968 , y15969 , y15970 , y15971 , y15972 , y15973 , y15974 , y15975 , y15976 , y15977 , y15978 , y15979 , y15980 , y15981 , y15982 , y15983 , y15984 , y15985 , y15986 , y15987 , y15988 , y15989 , y15990 , y15991 , y15992 , y15993 , y15994 , y15995 , y15996 , y15997 , y15998 , y15999 , y16000 , y16001 , y16002 , y16003 , y16004 , y16005 , y16006 , y16007 , y16008 , y16009 , y16010 , y16011 , y16012 , y16013 , y16014 , y16015 , y16016 , y16017 , y16018 , y16019 , y16020 , y16021 , y16022 , y16023 , y16024 , y16025 , y16026 , y16027 , y16028 , y16029 , y16030 , y16031 , y16032 , y16033 , y16034 , y16035 , y16036 , y16037 , y16038 , y16039 , y16040 , y16041 , y16042 , y16043 , y16044 , y16045 , y16046 , y16047 , y16048 , y16049 , y16050 , y16051 , y16052 , y16053 , y16054 , y16055 , y16056 , y16057 , y16058 , y16059 , y16060 , y16061 , y16062 , y16063 , y16064 , y16065 , y16066 , y16067 , y16068 , y16069 , y16070 , y16071 , y16072 , y16073 , y16074 , y16075 , y16076 , y16077 , y16078 , y16079 , y16080 , y16081 , y16082 , y16083 , y16084 , y16085 , y16086 , y16087 , y16088 , y16089 , y16090 , y16091 , y16092 , y16093 , y16094 , y16095 , y16096 , y16097 , y16098 , y16099 , y16100 , y16101 , y16102 , y16103 , y16104 , y16105 , y16106 , y16107 , y16108 , y16109 , y16110 , y16111 , y16112 , y16113 , y16114 , y16115 , y16116 , y16117 , y16118 , y16119 , y16120 , y16121 , y16122 , y16123 , y16124 , y16125 , y16126 , y16127 , y16128 , y16129 , y16130 , y16131 , y16132 , y16133 , y16134 , y16135 , y16136 , y16137 , y16138 , y16139 , y16140 , y16141 , y16142 , y16143 , y16144 , y16145 , y16146 , y16147 , y16148 , y16149 , y16150 , y16151 , y16152 , y16153 , y16154 , y16155 , y16156 , y16157 , y16158 , y16159 , y16160 , y16161 , y16162 , y16163 , y16164 , y16165 , y16166 , y16167 , y16168 , y16169 , y16170 , y16171 , y16172 , y16173 , y16174 , y16175 , y16176 , y16177 , y16178 , y16179 , y16180 , y16181 , y16182 , y16183 , y16184 , y16185 , y16186 , y16187 , y16188 , y16189 , y16190 , y16191 , y16192 , y16193 , y16194 , y16195 , y16196 , y16197 , y16198 , y16199 , y16200 , y16201 , y16202 , y16203 , y16204 , y16205 , y16206 , y16207 , y16208 , y16209 , y16210 , y16211 , y16212 , y16213 , y16214 , y16215 , y16216 , y16217 , y16218 , y16219 , y16220 , y16221 , y16222 , y16223 , y16224 , y16225 , y16226 , y16227 , y16228 , y16229 , y16230 , y16231 , y16232 , y16233 , y16234 , y16235 , y16236 , y16237 , y16238 , y16239 , y16240 , y16241 , y16242 , y16243 , y16244 , y16245 , y16246 , y16247 , y16248 , y16249 , y16250 , y16251 , y16252 , y16253 , y16254 , y16255 , y16256 , y16257 , y16258 , y16259 , y16260 , y16261 , y16262 , y16263 , y16264 , y16265 , y16266 , y16267 , y16268 , y16269 , y16270 , y16271 , y16272 , y16273 , y16274 , y16275 , y16276 , y16277 , y16278 , y16279 , y16280 , y16281 , y16282 , y16283 , y16284 , y16285 , y16286 , y16287 , y16288 , y16289 , y16290 , y16291 , y16292 , y16293 , y16294 , y16295 , y16296 , y16297 , y16298 , y16299 , y16300 , y16301 , y16302 , y16303 , y16304 , y16305 , y16306 , y16307 , y16308 , y16309 , y16310 , y16311 , y16312 , y16313 , y16314 , y16315 , y16316 , y16317 , y16318 , y16319 , y16320 , y16321 , y16322 , y16323 , y16324 , y16325 , y16326 , y16327 , y16328 , y16329 , y16330 , y16331 , y16332 , y16333 , y16334 , y16335 , y16336 , y16337 , y16338 , y16339 , y16340 , y16341 , y16342 , y16343 , y16344 , y16345 , y16346 , y16347 , y16348 , y16349 , y16350 , y16351 , y16352 , y16353 , y16354 , y16355 , y16356 , y16357 , y16358 , y16359 , y16360 , y16361 , y16362 , y16363 , y16364 , y16365 , y16366 , y16367 , y16368 , y16369 , y16370 , y16371 , y16372 , y16373 , y16374 , y16375 , y16376 , y16377 , y16378 , y16379 , y16380 , y16381 , y16382 , y16383 , y16384 , y16385 , y16386 , y16387 , y16388 , y16389 , y16390 , y16391 , y16392 , y16393 , y16394 , y16395 , y16396 , y16397 , y16398 , y16399 , y16400 , y16401 , y16402 , y16403 , y16404 , y16405 , y16406 , y16407 , y16408 , y16409 , y16410 , y16411 , y16412 , y16413 , y16414 , y16415 , y16416 , y16417 , y16418 , y16419 , y16420 , y16421 , y16422 , y16423 , y16424 , y16425 , y16426 , y16427 , y16428 , y16429 , y16430 , y16431 , y16432 , y16433 , y16434 , y16435 , y16436 , y16437 , y16438 , y16439 , y16440 , y16441 , y16442 , y16443 , y16444 , y16445 , y16446 , y16447 , y16448 , y16449 , y16450 , y16451 , y16452 , y16453 , y16454 , y16455 , y16456 , y16457 , y16458 , y16459 , y16460 , y16461 , y16462 , y16463 , y16464 , y16465 , y16466 , y16467 , y16468 , y16469 , y16470 , y16471 , y16472 , y16473 , y16474 , y16475 , y16476 , y16477 , y16478 , y16479 , y16480 , y16481 , y16482 , y16483 , y16484 , y16485 , y16486 , y16487 , y16488 , y16489 , y16490 , y16491 , y16492 , y16493 , y16494 , y16495 , y16496 , y16497 , y16498 , y16499 , y16500 , y16501 , y16502 , y16503 , y16504 , y16505 , y16506 , y16507 , y16508 , y16509 , y16510 , y16511 , y16512 , y16513 , y16514 , y16515 , y16516 , y16517 , y16518 , y16519 , y16520 , y16521 , y16522 , y16523 , y16524 , y16525 , y16526 , y16527 , y16528 , y16529 , y16530 , y16531 , y16532 , y16533 , y16534 , y16535 , y16536 , y16537 , y16538 , y16539 , y16540 , y16541 , y16542 , y16543 , y16544 , y16545 , y16546 , y16547 , y16548 , y16549 , y16550 , y16551 , y16552 , y16553 , y16554 , y16555 , y16556 , y16557 , y16558 , y16559 , y16560 , y16561 , y16562 , y16563 , y16564 , y16565 , y16566 , y16567 , y16568 , y16569 , y16570 , y16571 , y16572 , y16573 , y16574 , y16575 , y16576 , y16577 , y16578 , y16579 , y16580 , y16581 , y16582 , y16583 , y16584 , y16585 , y16586 , y16587 , y16588 , y16589 , y16590 , y16591 , y16592 , y16593 , y16594 , y16595 , y16596 , y16597 , y16598 , y16599 , y16600 , y16601 , y16602 , y16603 , y16604 , y16605 , y16606 , y16607 , y16608 , y16609 , y16610 , y16611 , y16612 , y16613 , y16614 , y16615 , y16616 , y16617 , y16618 , y16619 , y16620 , y16621 , y16622 , y16623 , y16624 , y16625 , y16626 , y16627 , y16628 , y16629 , y16630 , y16631 , y16632 , y16633 , y16634 , y16635 , y16636 , y16637 , y16638 , y16639 , y16640 , y16641 , y16642 , y16643 , y16644 , y16645 , y16646 , y16647 , y16648 , y16649 , y16650 , y16651 , y16652 , y16653 , y16654 , y16655 , y16656 , y16657 , y16658 , y16659 , y16660 , y16661 , y16662 , y16663 , y16664 , y16665 , y16666 , y16667 , y16668 , y16669 , y16670 , y16671 , y16672 , y16673 , y16674 , y16675 , y16676 , y16677 , y16678 , y16679 , y16680 , y16681 , y16682 , y16683 , y16684 , y16685 , y16686 , y16687 , y16688 , y16689 , y16690 , y16691 , y16692 , y16693 , y16694 , y16695 , y16696 , y16697 , y16698 , y16699 , y16700 , y16701 , y16702 , y16703 , y16704 , y16705 , y16706 , y16707 , y16708 , y16709 , y16710 , y16711 , y16712 , y16713 , y16714 , y16715 , y16716 , y16717 , y16718 , y16719 , y16720 , y16721 , y16722 , y16723 , y16724 , y16725 , y16726 , y16727 , y16728 , y16729 , y16730 , y16731 , y16732 , y16733 , y16734 , y16735 , y16736 , y16737 , y16738 , y16739 , y16740 , y16741 , y16742 , y16743 , y16744 , y16745 , y16746 , y16747 , y16748 , y16749 , y16750 , y16751 , y16752 , y16753 , y16754 , y16755 , y16756 , y16757 , y16758 , y16759 , y16760 , y16761 , y16762 , y16763 , y16764 , y16765 , y16766 , y16767 , y16768 , y16769 , y16770 , y16771 , y16772 , y16773 , y16774 , y16775 , y16776 , y16777 , y16778 , y16779 , y16780 , y16781 , y16782 , y16783 , y16784 , y16785 , y16786 , y16787 , y16788 , y16789 , y16790 , y16791 , y16792 , y16793 , y16794 , y16795 , y16796 , y16797 , y16798 , y16799 , y16800 , y16801 , y16802 , y16803 , y16804 , y16805 , y16806 , y16807 , y16808 , y16809 , y16810 , y16811 , y16812 , y16813 , y16814 , y16815 , y16816 , y16817 , y16818 , y16819 , y16820 , y16821 , y16822 , y16823 , y16824 , y16825 , y16826 , y16827 , y16828 , y16829 , y16830 , y16831 , y16832 , y16833 , y16834 , y16835 , y16836 , y16837 , y16838 , y16839 , y16840 , y16841 , y16842 , y16843 , y16844 , y16845 , y16846 , y16847 , y16848 , y16849 , y16850 , y16851 , y16852 , y16853 , y16854 , y16855 , y16856 , y16857 , y16858 , y16859 , y16860 , y16861 , y16862 , y16863 , y16864 , y16865 , y16866 , y16867 , y16868 , y16869 , y16870 , y16871 , y16872 , y16873 , y16874 , y16875 , y16876 , y16877 , y16878 , y16879 , y16880 , y16881 , y16882 , y16883 , y16884 , y16885 , y16886 , y16887 , y16888 , y16889 , y16890 , y16891 , y16892 , y16893 , y16894 , y16895 , y16896 , y16897 , y16898 , y16899 , y16900 , y16901 , y16902 , y16903 , y16904 , y16905 , y16906 , y16907 , y16908 , y16909 , y16910 , y16911 , y16912 , y16913 , y16914 , y16915 , y16916 , y16917 , y16918 , y16919 , y16920 , y16921 , y16922 , y16923 , y16924 , y16925 , y16926 , y16927 , y16928 , y16929 , y16930 , y16931 , y16932 , y16933 , y16934 , y16935 , y16936 , y16937 , y16938 , y16939 , y16940 , y16941 , y16942 , y16943 , y16944 , y16945 , y16946 , y16947 , y16948 , y16949 , y16950 , y16951 , y16952 , y16953 , y16954 , y16955 , y16956 , y16957 , y16958 , y16959 , y16960 , y16961 , y16962 , y16963 , y16964 , y16965 , y16966 , y16967 , y16968 , y16969 , y16970 , y16971 , y16972 , y16973 , y16974 , y16975 , y16976 , y16977 , y16978 , y16979 , y16980 , y16981 , y16982 , y16983 , y16984 , y16985 , y16986 , y16987 , y16988 , y16989 , y16990 , y16991 , y16992 , y16993 , y16994 , y16995 , y16996 , y16997 , y16998 , y16999 , y17000 , y17001 , y17002 , y17003 , y17004 , y17005 , y17006 , y17007 , y17008 , y17009 , y17010 , y17011 , y17012 , y17013 , y17014 , y17015 , y17016 , y17017 , y17018 , y17019 , y17020 , y17021 , y17022 , y17023 , y17024 , y17025 , y17026 , y17027 , y17028 , y17029 , y17030 , y17031 , y17032 , y17033 , y17034 , y17035 , y17036 , y17037 , y17038 , y17039 , y17040 , y17041 , y17042 , y17043 , y17044 , y17045 , y17046 , y17047 , y17048 , y17049 , y17050 , y17051 , y17052 , y17053 , y17054 , y17055 , y17056 , y17057 , y17058 , y17059 , y17060 , y17061 , y17062 , y17063 , y17064 , y17065 , y17066 , y17067 , y17068 , y17069 , y17070 , y17071 , y17072 , y17073 , y17074 , y17075 , y17076 , y17077 , y17078 , y17079 , y17080 , y17081 , y17082 , y17083 , y17084 , y17085 , y17086 , y17087 , y17088 , y17089 , y17090 , y17091 , y17092 , y17093 , y17094 , y17095 , y17096 , y17097 , y17098 , y17099 , y17100 , y17101 , y17102 , y17103 , y17104 , y17105 , y17106 , y17107 , y17108 , y17109 , y17110 , y17111 , y17112 , y17113 , y17114 , y17115 , y17116 , y17117 , y17118 , y17119 , y17120 , y17121 , y17122 , y17123 , y17124 , y17125 , y17126 , y17127 , y17128 , y17129 , y17130 , y17131 , y17132 , y17133 , y17134 , y17135 , y17136 , y17137 , y17138 , y17139 , y17140 , y17141 , y17142 , y17143 , y17144 , y17145 , y17146 , y17147 , y17148 , y17149 , y17150 , y17151 , y17152 , y17153 , y17154 , y17155 , y17156 , y17157 , y17158 , y17159 , y17160 , y17161 , y17162 , y17163 , y17164 , y17165 , y17166 , y17167 , y17168 , y17169 , y17170 , y17171 , y17172 , y17173 , y17174 , y17175 , y17176 , y17177 , y17178 , y17179 , y17180 , y17181 , y17182 , y17183 , y17184 , y17185 , y17186 , y17187 , y17188 , y17189 , y17190 , y17191 , y17192 , y17193 , y17194 , y17195 , y17196 , y17197 , y17198 , y17199 , y17200 , y17201 , y17202 , y17203 , y17204 , y17205 , y17206 , y17207 , y17208 , y17209 , y17210 , y17211 , y17212 , y17213 , y17214 , y17215 , y17216 , y17217 , y17218 , y17219 , y17220 , y17221 , y17222 , y17223 , y17224 , y17225 , y17226 , y17227 , y17228 , y17229 , y17230 , y17231 , y17232 , y17233 , y17234 , y17235 , y17236 , y17237 , y17238 , y17239 , y17240 , y17241 , y17242 , y17243 , y17244 , y17245 , y17246 , y17247 , y17248 , y17249 , y17250 , y17251 , y17252 , y17253 , y17254 , y17255 , y17256 , y17257 , y17258 , y17259 , y17260 , y17261 , y17262 , y17263 , y17264 , y17265 , y17266 , y17267 , y17268 , y17269 , y17270 , y17271 , y17272 , y17273 , y17274 , y17275 , y17276 , y17277 , y17278 , y17279 , y17280 , y17281 , y17282 , y17283 , y17284 , y17285 , y17286 , y17287 , y17288 , y17289 , y17290 , y17291 , y17292 , y17293 , y17294 , y17295 , y17296 , y17297 , y17298 , y17299 , y17300 , y17301 , y17302 , y17303 , y17304 , y17305 , y17306 , y17307 , y17308 , y17309 , y17310 , y17311 , y17312 , y17313 , y17314 , y17315 , y17316 , y17317 , y17318 , y17319 , y17320 , y17321 , y17322 , y17323 , y17324 , y17325 , y17326 , y17327 , y17328 , y17329 , y17330 , y17331 , y17332 , y17333 , y17334 , y17335 , y17336 , y17337 , y17338 , y17339 , y17340 , y17341 , y17342 , y17343 , y17344 , y17345 , y17346 , y17347 , y17348 , y17349 , y17350 , y17351 , y17352 , y17353 , y17354 , y17355 , y17356 , y17357 , y17358 , y17359 , y17360 , y17361 , y17362 , y17363 , y17364 , y17365 , y17366 , y17367 , y17368 , y17369 , y17370 , y17371 , y17372 , y17373 , y17374 , y17375 , y17376 , y17377 , y17378 , y17379 , y17380 , y17381 , y17382 , y17383 , y17384 , y17385 , y17386 , y17387 , y17388 , y17389 , y17390 , y17391 , y17392 , y17393 , y17394 , y17395 , y17396 , y17397 , y17398 , y17399 , y17400 , y17401 , y17402 , y17403 , y17404 , y17405 , y17406 , y17407 , y17408 , y17409 , y17410 , y17411 , y17412 , y17413 , y17414 , y17415 , y17416 , y17417 , y17418 , y17419 , y17420 , y17421 , y17422 , y17423 , y17424 , y17425 , y17426 , y17427 , y17428 , y17429 , y17430 , y17431 , y17432 , y17433 , y17434 , y17435 , y17436 , y17437 , y17438 , y17439 , y17440 , y17441 , y17442 , y17443 , y17444 , y17445 , y17446 , y17447 , y17448 , y17449 , y17450 , y17451 , y17452 , y17453 , y17454 , y17455 , y17456 , y17457 , y17458 , y17459 , y17460 , y17461 , y17462 , y17463 , y17464 , y17465 , y17466 , y17467 , y17468 , y17469 , y17470 , y17471 , y17472 , y17473 , y17474 , y17475 , y17476 , y17477 , y17478 , y17479 , y17480 , y17481 , y17482 , y17483 , y17484 , y17485 , y17486 , y17487 , y17488 , y17489 , y17490 , y17491 , y17492 , y17493 , y17494 , y17495 , y17496 , y17497 , y17498 , y17499 , y17500 , y17501 , y17502 , y17503 , y17504 , y17505 , y17506 , y17507 , y17508 , y17509 , y17510 , y17511 , y17512 , y17513 , y17514 , y17515 , y17516 , y17517 , y17518 , y17519 , y17520 , y17521 , y17522 , y17523 , y17524 , y17525 , y17526 , y17527 , y17528 , y17529 , y17530 , y17531 , y17532 , y17533 , y17534 , y17535 , y17536 , y17537 , y17538 , y17539 , y17540 , y17541 , y17542 , y17543 , y17544 , y17545 , y17546 , y17547 , y17548 , y17549 , y17550 , y17551 , y17552 , y17553 , y17554 , y17555 , y17556 , y17557 , y17558 , y17559 , y17560 , y17561 , y17562 , y17563 , y17564 , y17565 , y17566 , y17567 , y17568 , y17569 , y17570 , y17571 , y17572 , y17573 , y17574 , y17575 , y17576 , y17577 , y17578 , y17579 , y17580 , y17581 , y17582 , y17583 , y17584 , y17585 , y17586 , y17587 , y17588 , y17589 , y17590 , y17591 , y17592 , y17593 , y17594 , y17595 , y17596 , y17597 , y17598 , y17599 , y17600 , y17601 , y17602 , y17603 , y17604 , y17605 , y17606 , y17607 , y17608 , y17609 , y17610 , y17611 , y17612 , y17613 , y17614 , y17615 , y17616 , y17617 , y17618 , y17619 , y17620 , y17621 , y17622 , y17623 , y17624 , y17625 , y17626 , y17627 , y17628 , y17629 , y17630 , y17631 , y17632 , y17633 , y17634 , y17635 , y17636 , y17637 , y17638 , y17639 , y17640 , y17641 , y17642 , y17643 , y17644 , y17645 , y17646 , y17647 , y17648 , y17649 , y17650 , y17651 , y17652 , y17653 , y17654 , y17655 , y17656 , y17657 , y17658 , y17659 , y17660 , y17661 , y17662 , y17663 , y17664 , y17665 , y17666 , y17667 , y17668 , y17669 , y17670 , y17671 , y17672 , y17673 , y17674 , y17675 , y17676 , y17677 , y17678 , y17679 , y17680 , y17681 , y17682 , y17683 , y17684 , y17685 , y17686 , y17687 , y17688 , y17689 , y17690 , y17691 , y17692 , y17693 , y17694 , y17695 , y17696 , y17697 , y17698 , y17699 , y17700 , y17701 , y17702 , y17703 , y17704 , y17705 , y17706 , y17707 , y17708 , y17709 , y17710 , y17711 , y17712 , y17713 , y17714 , y17715 , y17716 , y17717 , y17718 , y17719 , y17720 , y17721 , y17722 , y17723 , y17724 , y17725 , y17726 , y17727 , y17728 , y17729 , y17730 , y17731 , y17732 , y17733 , y17734 , y17735 , y17736 , y17737 , y17738 , y17739 , y17740 , y17741 , y17742 , y17743 , y17744 , y17745 , y17746 , y17747 , y17748 , y17749 , y17750 , y17751 , y17752 , y17753 , y17754 , y17755 , y17756 , y17757 , y17758 , y17759 , y17760 , y17761 , y17762 , y17763 , y17764 , y17765 , y17766 , y17767 , y17768 , y17769 , y17770 , y17771 , y17772 , y17773 , y17774 , y17775 , y17776 , y17777 , y17778 , y17779 , y17780 , y17781 , y17782 , y17783 , y17784 , y17785 , y17786 , y17787 , y17788 , y17789 , y17790 , y17791 , y17792 , y17793 , y17794 , y17795 , y17796 , y17797 , y17798 , y17799 , y17800 , y17801 , y17802 , y17803 , y17804 , y17805 , y17806 , y17807 , y17808 , y17809 , y17810 , y17811 , y17812 , y17813 , y17814 , y17815 , y17816 , y17817 , y17818 , y17819 , y17820 , y17821 , y17822 , y17823 , y17824 , y17825 , y17826 , y17827 , y17828 , y17829 , y17830 , y17831 , y17832 , y17833 , y17834 , y17835 , y17836 , y17837 , y17838 , y17839 , y17840 , y17841 , y17842 , y17843 , y17844 , y17845 , y17846 , y17847 , y17848 , y17849 , y17850 , y17851 , y17852 , y17853 , y17854 , y17855 , y17856 , y17857 , y17858 , y17859 , y17860 , y17861 , y17862 , y17863 , y17864 , y17865 , y17866 , y17867 , y17868 , y17869 , y17870 , y17871 , y17872 , y17873 , y17874 , y17875 , y17876 , y17877 , y17878 , y17879 , y17880 , y17881 , y17882 , y17883 , y17884 , y17885 , y17886 , y17887 , y17888 , y17889 , y17890 , y17891 , y17892 , y17893 , y17894 , y17895 , y17896 , y17897 , y17898 , y17899 , y17900 , y17901 , y17902 , y17903 , y17904 , y17905 , y17906 , y17907 , y17908 , y17909 , y17910 , y17911 , y17912 , y17913 , y17914 , y17915 , y17916 , y17917 , y17918 , y17919 , y17920 , y17921 , y17922 , y17923 , y17924 , y17925 , y17926 , y17927 , y17928 , y17929 , y17930 , y17931 , y17932 , y17933 , y17934 , y17935 , y17936 , y17937 , y17938 , y17939 , y17940 , y17941 , y17942 , y17943 , y17944 , y17945 , y17946 , y17947 , y17948 , y17949 , y17950 , y17951 , y17952 , y17953 , y17954 , y17955 , y17956 , y17957 , y17958 , y17959 , y17960 , y17961 , y17962 , y17963 , y17964 , y17965 , y17966 , y17967 , y17968 , y17969 , y17970 , y17971 , y17972 , y17973 , y17974 , y17975 , y17976 , y17977 , y17978 , y17979 , y17980 , y17981 , y17982 , y17983 , y17984 , y17985 , y17986 , y17987 , y17988 , y17989 , y17990 , y17991 , y17992 , y17993 , y17994 , y17995 , y17996 , y17997 , y17998 , y17999 , y18000 , y18001 , y18002 , y18003 , y18004 , y18005 , y18006 , y18007 , y18008 , y18009 , y18010 , y18011 , y18012 , y18013 , y18014 , y18015 , y18016 , y18017 , y18018 , y18019 , y18020 , y18021 , y18022 , y18023 , y18024 , y18025 , y18026 , y18027 , y18028 , y18029 , y18030 , y18031 , y18032 , y18033 , y18034 , y18035 , y18036 , y18037 , y18038 , y18039 , y18040 , y18041 , y18042 , y18043 , y18044 , y18045 , y18046 , y18047 , y18048 , y18049 , y18050 , y18051 , y18052 , y18053 , y18054 , y18055 , y18056 , y18057 , y18058 , y18059 , y18060 , y18061 , y18062 , y18063 , y18064 , y18065 , y18066 , y18067 , y18068 , y18069 , y18070 , y18071 , y18072 , y18073 , y18074 , y18075 , y18076 , y18077 , y18078 , y18079 , y18080 , y18081 , y18082 , y18083 , y18084 , y18085 , y18086 , y18087 , y18088 , y18089 , y18090 , y18091 , y18092 , y18093 , y18094 , y18095 , y18096 , y18097 , y18098 , y18099 , y18100 , y18101 , y18102 , y18103 , y18104 , y18105 , y18106 , y18107 , y18108 , y18109 , y18110 , y18111 , y18112 , y18113 , y18114 , y18115 , y18116 , y18117 , y18118 , y18119 , y18120 , y18121 , y18122 , y18123 , y18124 , y18125 , y18126 , y18127 , y18128 , y18129 , y18130 , y18131 , y18132 , y18133 , y18134 , y18135 , y18136 , y18137 , y18138 , y18139 , y18140 , y18141 , y18142 , y18143 , y18144 , y18145 , y18146 , y18147 , y18148 , y18149 , y18150 , y18151 , y18152 , y18153 , y18154 , y18155 , y18156 , y18157 , y18158 , y18159 , y18160 , y18161 , y18162 , y18163 , y18164 , y18165 , y18166 , y18167 , y18168 , y18169 , y18170 , y18171 , y18172 , y18173 , y18174 , y18175 , y18176 , y18177 , y18178 , y18179 , y18180 , y18181 , y18182 , y18183 , y18184 , y18185 , y18186 , y18187 , y18188 , y18189 , y18190 , y18191 , y18192 , y18193 , y18194 , y18195 , y18196 , y18197 , y18198 , y18199 , y18200 , y18201 , y18202 , y18203 , y18204 , y18205 , y18206 , y18207 , y18208 , y18209 , y18210 , y18211 , y18212 , y18213 , y18214 , y18215 , y18216 , y18217 , y18218 , y18219 , y18220 , y18221 , y18222 , y18223 , y18224 , y18225 , y18226 , y18227 , y18228 , y18229 , y18230 , y18231 , y18232 , y18233 , y18234 , y18235 , y18236 , y18237 , y18238 , y18239 , y18240 , y18241 , y18242 , y18243 , y18244 , y18245 , y18246 , y18247 , y18248 , y18249 , y18250 , y18251 , y18252 , y18253 , y18254 , y18255 , y18256 , y18257 , y18258 , y18259 , y18260 , y18261 , y18262 , y18263 , y18264 , y18265 , y18266 , y18267 , y18268 , y18269 , y18270 , y18271 , y18272 , y18273 , y18274 , y18275 , y18276 , y18277 , y18278 , y18279 , y18280 , y18281 , y18282 , y18283 , y18284 , y18285 , y18286 , y18287 , y18288 , y18289 , y18290 , y18291 , y18292 , y18293 , y18294 , y18295 , y18296 , y18297 , y18298 , y18299 , y18300 , y18301 , y18302 , y18303 , y18304 , y18305 , y18306 , y18307 , y18308 , y18309 , y18310 , y18311 , y18312 , y18313 , y18314 , y18315 , y18316 , y18317 , y18318 , y18319 , y18320 , y18321 , y18322 , y18323 , y18324 , y18325 , y18326 , y18327 , y18328 , y18329 , y18330 , y18331 , y18332 , y18333 , y18334 , y18335 , y18336 , y18337 , y18338 , y18339 , y18340 , y18341 , y18342 , y18343 , y18344 , y18345 , y18346 , y18347 , y18348 , y18349 , y18350 , y18351 , y18352 , y18353 , y18354 , y18355 , y18356 , y18357 , y18358 , y18359 , y18360 , y18361 , y18362 , y18363 , y18364 , y18365 , y18366 , y18367 , y18368 , y18369 , y18370 , y18371 , y18372 , y18373 , y18374 , y18375 , y18376 , y18377 , y18378 , y18379 , y18380 , y18381 , y18382 , y18383 , y18384 , y18385 , y18386 , y18387 , y18388 , y18389 , y18390 , y18391 , y18392 , y18393 , y18394 , y18395 , y18396 , y18397 , y18398 , y18399 , y18400 , y18401 , y18402 , y18403 , y18404 , y18405 , y18406 , y18407 , y18408 , y18409 , y18410 , y18411 , y18412 , y18413 , y18414 , y18415 , y18416 , y18417 , y18418 , y18419 , y18420 , y18421 , y18422 , y18423 , y18424 , y18425 , y18426 , y18427 , y18428 , y18429 , y18430 , y18431 , y18432 , y18433 , y18434 , y18435 , y18436 , y18437 , y18438 , y18439 , y18440 , y18441 , y18442 , y18443 , y18444 , y18445 , y18446 , y18447 , y18448 , y18449 , y18450 , y18451 , y18452 , y18453 , y18454 , y18455 , y18456 , y18457 , y18458 , y18459 , y18460 , y18461 , y18462 , y18463 , y18464 , y18465 , y18466 , y18467 , y18468 , y18469 , y18470 , y18471 , y18472 , y18473 , y18474 , y18475 , y18476 , y18477 , y18478 , y18479 , y18480 , y18481 , y18482 , y18483 , y18484 , y18485 , y18486 , y18487 , y18488 , y18489 , y18490 , y18491 , y18492 , y18493 , y18494 , y18495 , y18496 , y18497 , y18498 , y18499 , y18500 , y18501 , y18502 , y18503 , y18504 , y18505 , y18506 , y18507 , y18508 , y18509 , y18510 , y18511 , y18512 , y18513 , y18514 , y18515 , y18516 , y18517 , y18518 , y18519 , y18520 , y18521 , y18522 , y18523 , y18524 , y18525 , y18526 , y18527 , y18528 , y18529 , y18530 , y18531 , y18532 , y18533 , y18534 , y18535 , y18536 , y18537 , y18538 , y18539 , y18540 , y18541 , y18542 , y18543 , y18544 , y18545 , y18546 , y18547 , y18548 , y18549 , y18550 , y18551 , y18552 , y18553 , y18554 , y18555 , y18556 , y18557 , y18558 , y18559 , y18560 , y18561 , y18562 , y18563 , y18564 , y18565 , y18566 , y18567 , y18568 , y18569 , y18570 , y18571 , y18572 , y18573 , y18574 , y18575 , y18576 , y18577 , y18578 , y18579 , y18580 , y18581 , y18582 , y18583 , y18584 , y18585 , y18586 , y18587 , y18588 , y18589 , y18590 , y18591 , y18592 , y18593 , y18594 , y18595 , y18596 , y18597 , y18598 , y18599 , y18600 , y18601 , y18602 , y18603 , y18604 , y18605 , y18606 , y18607 , y18608 , y18609 , y18610 , y18611 , y18612 , y18613 , y18614 , y18615 , y18616 , y18617 , y18618 , y18619 , y18620 , y18621 , y18622 , y18623 , y18624 , y18625 , y18626 , y18627 , y18628 , y18629 , y18630 , y18631 , y18632 , y18633 , y18634 , y18635 , y18636 , y18637 , y18638 , y18639 , y18640 , y18641 , y18642 , y18643 , y18644 , y18645 , y18646 , y18647 , y18648 , y18649 , y18650 , y18651 , y18652 , y18653 , y18654 , y18655 , y18656 , y18657 , y18658 , y18659 , y18660 , y18661 , y18662 , y18663 , y18664 , y18665 , y18666 , y18667 , y18668 , y18669 , y18670 , y18671 , y18672 , y18673 , y18674 , y18675 , y18676 , y18677 , y18678 , y18679 , y18680 , y18681 , y18682 , y18683 , y18684 , y18685 , y18686 , y18687 , y18688 , y18689 , y18690 , y18691 , y18692 , y18693 , y18694 , y18695 , y18696 , y18697 , y18698 , y18699 , y18700 , y18701 , y18702 , y18703 , y18704 , y18705 , y18706 , y18707 , y18708 , y18709 , y18710 , y18711 , y18712 , y18713 , y18714 , y18715 , y18716 , y18717 , y18718 , y18719 , y18720 , y18721 , y18722 , y18723 , y18724 , y18725 , y18726 , y18727 , y18728 , y18729 , y18730 , y18731 , y18732 , y18733 , y18734 , y18735 , y18736 , y18737 , y18738 , y18739 , y18740 , y18741 , y18742 , y18743 , y18744 , y18745 , y18746 , y18747 , y18748 , y18749 , y18750 , y18751 , y18752 , y18753 , y18754 , y18755 , y18756 , y18757 , y18758 , y18759 , y18760 , y18761 , y18762 , y18763 , y18764 , y18765 , y18766 , y18767 , y18768 , y18769 , y18770 , y18771 , y18772 , y18773 , y18774 , y18775 , y18776 , y18777 , y18778 , y18779 , y18780 , y18781 , y18782 , y18783 , y18784 , y18785 , y18786 , y18787 , y18788 , y18789 , y18790 , y18791 , y18792 , y18793 , y18794 , y18795 , y18796 , y18797 , y18798 , y18799 , y18800 , y18801 , y18802 , y18803 , y18804 , y18805 , y18806 , y18807 , y18808 , y18809 , y18810 , y18811 , y18812 , y18813 , y18814 , y18815 , y18816 , y18817 , y18818 , y18819 , y18820 , y18821 , y18822 , y18823 , y18824 , y18825 , y18826 , y18827 , y18828 , y18829 , y18830 , y18831 , y18832 , y18833 , y18834 , y18835 , y18836 , y18837 , y18838 , y18839 , y18840 , y18841 , y18842 , y18843 , y18844 , y18845 , y18846 , y18847 , y18848 , y18849 , y18850 , y18851 , y18852 , y18853 , y18854 , y18855 , y18856 , y18857 , y18858 , y18859 , y18860 , y18861 , y18862 , y18863 , y18864 , y18865 , y18866 , y18867 , y18868 , y18869 , y18870 , y18871 , y18872 , y18873 , y18874 , y18875 , y18876 , y18877 , y18878 , y18879 , y18880 , y18881 , y18882 , y18883 , y18884 , y18885 , y18886 , y18887 , y18888 , y18889 , y18890 , y18891 , y18892 , y18893 , y18894 , y18895 , y18896 , y18897 , y18898 , y18899 , y18900 , y18901 , y18902 , y18903 , y18904 , y18905 , y18906 , y18907 , y18908 , y18909 , y18910 , y18911 , y18912 , y18913 , y18914 , y18915 , y18916 , y18917 , y18918 , y18919 , y18920 , y18921 , y18922 , y18923 , y18924 , y18925 , y18926 , y18927 , y18928 , y18929 , y18930 , y18931 , y18932 , y18933 , y18934 , y18935 , y18936 , y18937 , y18938 , y18939 , y18940 , y18941 , y18942 , y18943 , y18944 , y18945 , y18946 , y18947 , y18948 , y18949 , y18950 , y18951 , y18952 , y18953 , y18954 , y18955 , y18956 , y18957 , y18958 , y18959 , y18960 , y18961 , y18962 , y18963 , y18964 , y18965 , y18966 , y18967 , y18968 , y18969 , y18970 , y18971 , y18972 , y18973 , y18974 , y18975 , y18976 , y18977 , y18978 , y18979 , y18980 , y18981 , y18982 , y18983 , y18984 , y18985 , y18986 , y18987 , y18988 , y18989 , y18990 , y18991 , y18992 , y18993 , y18994 , y18995 , y18996 , y18997 , y18998 , y18999 , y19000 , y19001 , y19002 , y19003 , y19004 , y19005 , y19006 , y19007 , y19008 , y19009 , y19010 , y19011 , y19012 , y19013 , y19014 , y19015 , y19016 , y19017 , y19018 , y19019 , y19020 , y19021 , y19022 , y19023 , y19024 , y19025 , y19026 , y19027 , y19028 , y19029 , y19030 , y19031 , y19032 , y19033 , y19034 , y19035 , y19036 , y19037 , y19038 , y19039 , y19040 , y19041 , y19042 , y19043 , y19044 , y19045 , y19046 , y19047 , y19048 , y19049 , y19050 , y19051 , y19052 , y19053 , y19054 , y19055 , y19056 , y19057 , y19058 , y19059 , y19060 , y19061 , y19062 , y19063 , y19064 , y19065 , y19066 , y19067 , y19068 , y19069 , y19070 , y19071 , y19072 , y19073 , y19074 , y19075 , y19076 , y19077 , y19078 , y19079 , y19080 , y19081 , y19082 , y19083 , y19084 , y19085 , y19086 , y19087 , y19088 , y19089 , y19090 , y19091 , y19092 , y19093 , y19094 , y19095 , y19096 , y19097 , y19098 , y19099 , y19100 , y19101 , y19102 , y19103 , y19104 , y19105 , y19106 , y19107 , y19108 , y19109 , y19110 , y19111 , y19112 , y19113 , y19114 , y19115 , y19116 , y19117 , y19118 , y19119 , y19120 , y19121 , y19122 , y19123 , y19124 , y19125 , y19126 , y19127 , y19128 , y19129 , y19130 , y19131 , y19132 , y19133 , y19134 , y19135 , y19136 , y19137 , y19138 , y19139 , y19140 , y19141 , y19142 , y19143 , y19144 , y19145 , y19146 , y19147 , y19148 , y19149 , y19150 , y19151 , y19152 , y19153 , y19154 , y19155 , y19156 , y19157 , y19158 , y19159 , y19160 , y19161 , y19162 , y19163 , y19164 , y19165 , y19166 , y19167 , y19168 , y19169 , y19170 , y19171 , y19172 , y19173 , y19174 , y19175 , y19176 , y19177 , y19178 , y19179 , y19180 , y19181 , y19182 , y19183 , y19184 , y19185 , y19186 , y19187 , y19188 , y19189 , y19190 , y19191 , y19192 , y19193 , y19194 , y19195 , y19196 , y19197 , y19198 , y19199 , y19200 , y19201 , y19202 , y19203 , y19204 , y19205 , y19206 , y19207 , y19208 , y19209 , y19210 , y19211 , y19212 , y19213 , y19214 , y19215 , y19216 , y19217 , y19218 , y19219 , y19220 , y19221 , y19222 , y19223 , y19224 , y19225 , y19226 , y19227 , y19228 , y19229 , y19230 , y19231 , y19232 , y19233 , y19234 , y19235 , y19236 , y19237 , y19238 , y19239 , y19240 , y19241 , y19242 , y19243 , y19244 , y19245 , y19246 , y19247 , y19248 , y19249 , y19250 , y19251 , y19252 , y19253 , y19254 , y19255 , y19256 , y19257 , y19258 , y19259 , y19260 , y19261 , y19262 , y19263 , y19264 , y19265 , y19266 , y19267 , y19268 , y19269 , y19270 , y19271 , y19272 , y19273 , y19274 , y19275 , y19276 , y19277 , y19278 , y19279 , y19280 , y19281 , y19282 , y19283 , y19284 , y19285 , y19286 , y19287 , y19288 , y19289 , y19290 , y19291 , y19292 , y19293 , y19294 , y19295 , y19296 , y19297 , y19298 , y19299 , y19300 , y19301 , y19302 , y19303 , y19304 , y19305 , y19306 , y19307 , y19308 , y19309 , y19310 , y19311 , y19312 , y19313 , y19314 , y19315 , y19316 , y19317 , y19318 , y19319 , y19320 , y19321 , y19322 , y19323 , y19324 , y19325 , y19326 , y19327 , y19328 , y19329 , y19330 , y19331 , y19332 , y19333 , y19334 , y19335 , y19336 , y19337 , y19338 , y19339 , y19340 , y19341 , y19342 , y19343 , y19344 , y19345 , y19346 , y19347 , y19348 , y19349 , y19350 , y19351 , y19352 , y19353 , y19354 , y19355 , y19356 , y19357 , y19358 , y19359 , y19360 , y19361 , y19362 , y19363 , y19364 , y19365 , y19366 , y19367 , y19368 , y19369 , y19370 , y19371 , y19372 , y19373 , y19374 , y19375 , y19376 , y19377 , y19378 , y19379 , y19380 , y19381 , y19382 , y19383 , y19384 , y19385 , y19386 , y19387 , y19388 , y19389 , y19390 , y19391 , y19392 , y19393 , y19394 , y19395 , y19396 , y19397 , y19398 , y19399 , y19400 , y19401 , y19402 , y19403 , y19404 , y19405 , y19406 , y19407 , y19408 , y19409 , y19410 , y19411 , y19412 , y19413 , y19414 , y19415 , y19416 , y19417 , y19418 , y19419 , y19420 , y19421 , y19422 , y19423 , y19424 , y19425 , y19426 , y19427 , y19428 , y19429 , y19430 , y19431 , y19432 , y19433 , y19434 , y19435 , y19436 , y19437 , y19438 , y19439 , y19440 , y19441 , y19442 , y19443 , y19444 , y19445 , y19446 , y19447 , y19448 , y19449 , y19450 , y19451 , y19452 , y19453 , y19454 , y19455 , y19456 , y19457 , y19458 , y19459 , y19460 , y19461 , y19462 , y19463 , y19464 , y19465 , y19466 , y19467 , y19468 , y19469 , y19470 , y19471 , y19472 , y19473 , y19474 , y19475 , y19476 , y19477 , y19478 , y19479 , y19480 , y19481 , y19482 , y19483 , y19484 , y19485 , y19486 , y19487 , y19488 , y19489 , y19490 , y19491 , y19492 , y19493 , y19494 , y19495 , y19496 , y19497 , y19498 , y19499 , y19500 , y19501 , y19502 , y19503 , y19504 , y19505 , y19506 , y19507 , y19508 , y19509 , y19510 , y19511 , y19512 , y19513 , y19514 , y19515 , y19516 , y19517 , y19518 , y19519 , y19520 , y19521 , y19522 , y19523 , y19524 , y19525 , y19526 , y19527 , y19528 , y19529 , y19530 , y19531 , y19532 , y19533 , y19534 , y19535 , y19536 , y19537 , y19538 , y19539 , y19540 , y19541 , y19542 , y19543 , y19544 , y19545 , y19546 , y19547 , y19548 , y19549 , y19550 , y19551 , y19552 , y19553 , y19554 , y19555 , y19556 , y19557 , y19558 , y19559 , y19560 , y19561 , y19562 , y19563 , y19564 , y19565 , y19566 , y19567 , y19568 , y19569 , y19570 , y19571 , y19572 , y19573 , y19574 , y19575 , y19576 , y19577 , y19578 , y19579 , y19580 , y19581 , y19582 , y19583 , y19584 , y19585 , y19586 , y19587 , y19588 , y19589 , y19590 , y19591 , y19592 , y19593 , y19594 , y19595 , y19596 , y19597 , y19598 , y19599 , y19600 , y19601 , y19602 , y19603 , y19604 , y19605 , y19606 , y19607 , y19608 , y19609 , y19610 , y19611 , y19612 , y19613 , y19614 , y19615 , y19616 , y19617 , y19618 , y19619 , y19620 , y19621 , y19622 , y19623 , y19624 , y19625 , y19626 , y19627 , y19628 , y19629 , y19630 , y19631 , y19632 , y19633 , y19634 , y19635 , y19636 , y19637 , y19638 , y19639 , y19640 , y19641 , y19642 , y19643 , y19644 , y19645 , y19646 , y19647 , y19648 , y19649 , y19650 , y19651 , y19652 , y19653 , y19654 , y19655 , y19656 , y19657 , y19658 , y19659 , y19660 , y19661 , y19662 , y19663 , y19664 , y19665 , y19666 , y19667 , y19668 , y19669 , y19670 , y19671 , y19672 , y19673 , y19674 , y19675 , y19676 , y19677 , y19678 , y19679 , y19680 , y19681 , y19682 , y19683 , y19684 , y19685 , y19686 , y19687 , y19688 , y19689 , y19690 , y19691 , y19692 , y19693 , y19694 , y19695 , y19696 , y19697 , y19698 , y19699 , y19700 , y19701 , y19702 , y19703 , y19704 , y19705 , y19706 , y19707 , y19708 , y19709 , y19710 , y19711 , y19712 , y19713 , y19714 , y19715 , y19716 , y19717 , y19718 , y19719 , y19720 , y19721 , y19722 , y19723 , y19724 , y19725 , y19726 , y19727 , y19728 , y19729 , y19730 , y19731 , y19732 , y19733 , y19734 , y19735 , y19736 , y19737 , y19738 , y19739 , y19740 , y19741 , y19742 , y19743 , y19744 , y19745 , y19746 , y19747 , y19748 , y19749 , y19750 , y19751 , y19752 , y19753 , y19754 , y19755 , y19756 , y19757 , y19758 , y19759 , y19760 , y19761 , y19762 , y19763 , y19764 , y19765 , y19766 , y19767 , y19768 , y19769 , y19770 , y19771 , y19772 , y19773 , y19774 , y19775 , y19776 , y19777 , y19778 , y19779 , y19780 , y19781 , y19782 , y19783 , y19784 , y19785 , y19786 , y19787 , y19788 , y19789 , y19790 , y19791 , y19792 , y19793 , y19794 , y19795 , y19796 , y19797 , y19798 , y19799 , y19800 , y19801 , y19802 , y19803 , y19804 , y19805 , y19806 , y19807 , y19808 , y19809 , y19810 , y19811 , y19812 , y19813 , y19814 , y19815 , y19816 , y19817 , y19818 , y19819 , y19820 , y19821 , y19822 , y19823 , y19824 , y19825 , y19826 , y19827 , y19828 , y19829 , y19830 , y19831 , y19832 , y19833 , y19834 , y19835 , y19836 , y19837 , y19838 , y19839 , y19840 , y19841 , y19842 , y19843 , y19844 , y19845 , y19846 , y19847 , y19848 , y19849 , y19850 , y19851 , y19852 , y19853 , y19854 , y19855 , y19856 , y19857 , y19858 , y19859 , y19860 , y19861 , y19862 , y19863 , y19864 , y19865 , y19866 , y19867 , y19868 , y19869 , y19870 , y19871 , y19872 , y19873 , y19874 , y19875 , y19876 , y19877 , y19878 , y19879 , y19880 , y19881 , y19882 , y19883 , y19884 , y19885 , y19886 , y19887 , y19888 , y19889 , y19890 , y19891 , y19892 , y19893 , y19894 , y19895 , y19896 , y19897 , y19898 , y19899 , y19900 , y19901 , y19902 , y19903 , y19904 , y19905 , y19906 , y19907 , y19908 , y19909 , y19910 , y19911 , y19912 , y19913 , y19914 , y19915 , y19916 , y19917 , y19918 , y19919 , y19920 , y19921 , y19922 , y19923 , y19924 , y19925 , y19926 , y19927 , y19928 , y19929 , y19930 , y19931 , y19932 , y19933 , y19934 , y19935 , y19936 , y19937 , y19938 , y19939 , y19940 , y19941 , y19942 , y19943 , y19944 , y19945 , y19946 , y19947 , y19948 , y19949 , y19950 , y19951 , y19952 , y19953 , y19954 , y19955 , y19956 , y19957 , y19958 , y19959 , y19960 , y19961 , y19962 , y19963 , y19964 , y19965 , y19966 , y19967 , y19968 , y19969 , y19970 , y19971 , y19972 , y19973 , y19974 , y19975 , y19976 , y19977 , y19978 , y19979 , y19980 , y19981 , y19982 , y19983 , y19984 , y19985 , y19986 , y19987 , y19988 , y19989 , y19990 , y19991 , y19992 , y19993 , y19994 , y19995 , y19996 , y19997 , y19998 , y19999 , y20000 , y20001 , y20002 , y20003 , y20004 , y20005 , y20006 , y20007 , y20008 , y20009 , y20010 , y20011 , y20012 , y20013 , y20014 , y20015 , y20016 , y20017 , y20018 , y20019 , y20020 , y20021 , y20022 , y20023 , y20024 , y20025 , y20026 , y20027 , y20028 , y20029 , y20030 , y20031 , y20032 , y20033 , y20034 , y20035 , y20036 , y20037 , y20038 , y20039 , y20040 , y20041 , y20042 , y20043 , y20044 , y20045 , y20046 , y20047 , y20048 , y20049 , y20050 , y20051 , y20052 , y20053 , y20054 , y20055 , y20056 , y20057 , y20058 , y20059 , y20060 , y20061 , y20062 , y20063 , y20064 , y20065 , y20066 , y20067 , y20068 , y20069 , y20070 , y20071 , y20072 , y20073 , y20074 , y20075 , y20076 , y20077 , y20078 , y20079 , y20080 , y20081 , y20082 , y20083 , y20084 , y20085 , y20086 , y20087 , y20088 , y20089 , y20090 , y20091 , y20092 , y20093 , y20094 , y20095 , y20096 , y20097 , y20098 , y20099 , y20100 , y20101 , y20102 , y20103 , y20104 , y20105 , y20106 , y20107 , y20108 , y20109 , y20110 , y20111 , y20112 , y20113 , y20114 , y20115 , y20116 , y20117 , y20118 , y20119 , y20120 , y20121 , y20122 , y20123 , y20124 , y20125 , y20126 , y20127 , y20128 , y20129 , y20130 , y20131 , y20132 , y20133 , y20134 , y20135 , y20136 , y20137 , y20138 , y20139 , y20140 , y20141 , y20142 , y20143 , y20144 , y20145 , y20146 , y20147 , y20148 , y20149 , y20150 , y20151 , y20152 , y20153 , y20154 , y20155 , y20156 , y20157 , y20158 , y20159 , y20160 , y20161 , y20162 , y20163 , y20164 , y20165 , y20166 , y20167 , y20168 , y20169 , y20170 , y20171 , y20172 , y20173 , y20174 , y20175 , y20176 , y20177 , y20178 , y20179 , y20180 , y20181 , y20182 , y20183 , y20184 , y20185 , y20186 , y20187 , y20188 , y20189 , y20190 , y20191 , y20192 , y20193 , y20194 , y20195 , y20196 , y20197 , y20198 , y20199 , y20200 , y20201 , y20202 , y20203 , y20204 , y20205 , y20206 , y20207 , y20208 , y20209 , y20210 , y20211 , y20212 , y20213 , y20214 , y20215 , y20216 , y20217 , y20218 , y20219 , y20220 , y20221 , y20222 , y20223 , y20224 , y20225 , y20226 , y20227 , y20228 , y20229 , y20230 , y20231 , y20232 , y20233 , y20234 , y20235 , y20236 , y20237 , y20238 , y20239 , y20240 , y20241 , y20242 , y20243 , y20244 , y20245 , y20246 , y20247 , y20248 , y20249 , y20250 , y20251 , y20252 , y20253 , y20254 , y20255 , y20256 , y20257 , y20258 , y20259 , y20260 , y20261 , y20262 , y20263 , y20264 , y20265 , y20266 , y20267 , y20268 , y20269 , y20270 , y20271 , y20272 , y20273 , y20274 , y20275 , y20276 , y20277 , y20278 , y20279 , y20280 , y20281 , y20282 , y20283 , y20284 , y20285 , y20286 , y20287 , y20288 , y20289 , y20290 , y20291 , y20292 , y20293 , y20294 , y20295 , y20296 , y20297 , y20298 , y20299 , y20300 , y20301 , y20302 , y20303 , y20304 , y20305 , y20306 , y20307 , y20308 , y20309 , y20310 , y20311 , y20312 , y20313 , y20314 , y20315 , y20316 , y20317 , y20318 , y20319 , y20320 , y20321 , y20322 , y20323 , y20324 , y20325 , y20326 , y20327 , y20328 , y20329 , y20330 , y20331 , y20332 , y20333 , y20334 , y20335 , y20336 , y20337 , y20338 , y20339 , y20340 , y20341 , y20342 , y20343 , y20344 , y20345 , y20346 , y20347 , y20348 , y20349 , y20350 , y20351 , y20352 , y20353 , y20354 , y20355 , y20356 , y20357 , y20358 , y20359 , y20360 , y20361 , y20362 , y20363 , y20364 , y20365 , y20366 , y20367 , y20368 , y20369 , y20370 , y20371 , y20372 , y20373 , y20374 , y20375 , y20376 , y20377 , y20378 , y20379 , y20380 , y20381 , y20382 , y20383 , y20384 , y20385 , y20386 , y20387 , y20388 , y20389 , y20390 , y20391 , y20392 , y20393 , y20394 , y20395 , y20396 , y20397 , y20398 , y20399 , y20400 , y20401 , y20402 , y20403 , y20404 , y20405 , y20406 , y20407 , y20408 , y20409 , y20410 , y20411 , y20412 , y20413 , y20414 , y20415 , y20416 , y20417 , y20418 , y20419 , y20420 , y20421 , y20422 , y20423 , y20424 , y20425 , y20426 , y20427 , y20428 , y20429 , y20430 , y20431 , y20432 , y20433 , y20434 , y20435 , y20436 , y20437 , y20438 , y20439 , y20440 , y20441 , y20442 , y20443 , y20444 , y20445 , y20446 , y20447 , y20448 , y20449 , y20450 , y20451 , y20452 , y20453 , y20454 , y20455 , y20456 , y20457 , y20458 , y20459 , y20460 , y20461 , y20462 , y20463 , y20464 , y20465 , y20466 , y20467 , y20468 , y20469 , y20470 , y20471 , y20472 , y20473 , y20474 , y20475 , y20476 , y20477 , y20478 , y20479 , y20480 , y20481 , y20482 , y20483 , y20484 , y20485 , y20486 , y20487 , y20488 , y20489 , y20490 , y20491 , y20492 , y20493 , y20494 , y20495 , y20496 , y20497 , y20498 , y20499 , y20500 , y20501 , y20502 , y20503 , y20504 , y20505 , y20506 , y20507 , y20508 , y20509 , y20510 , y20511 , y20512 , y20513 , y20514 , y20515 , y20516 , y20517 , y20518 , y20519 , y20520 , y20521 , y20522 , y20523 , y20524 , y20525 , y20526 , y20527 , y20528 , y20529 , y20530 , y20531 , y20532 , y20533 , y20534 , y20535 , y20536 , y20537 , y20538 , y20539 , y20540 , y20541 , y20542 , y20543 , y20544 , y20545 , y20546 , y20547 , y20548 , y20549 , y20550 , y20551 , y20552 , y20553 , y20554 , y20555 , y20556 , y20557 , y20558 , y20559 , y20560 , y20561 , y20562 , y20563 , y20564 , y20565 , y20566 , y20567 , y20568 , y20569 , y20570 , y20571 , y20572 , y20573 , y20574 , y20575 , y20576 , y20577 , y20578 , y20579 , y20580 , y20581 , y20582 , y20583 , y20584 , y20585 , y20586 , y20587 , y20588 , y20589 , y20590 , y20591 , y20592 , y20593 , y20594 , y20595 , y20596 , y20597 , y20598 , y20599 , y20600 , y20601 , y20602 , y20603 , y20604 , y20605 , y20606 , y20607 , y20608 , y20609 , y20610 , y20611 , y20612 , y20613 , y20614 , y20615 , y20616 , y20617 , y20618 , y20619 , y20620 , y20621 , y20622 , y20623 , y20624 , y20625 , y20626 , y20627 , y20628 , y20629 , y20630 , y20631 , y20632 , y20633 , y20634 , y20635 , y20636 , y20637 , y20638 , y20639 , y20640 , y20641 , y20642 , y20643 , y20644 , y20645 , y20646 , y20647 , y20648 , y20649 , y20650 , y20651 , y20652 , y20653 , y20654 , y20655 , y20656 , y20657 , y20658 , y20659 , y20660 , y20661 , y20662 , y20663 , y20664 , y20665 , y20666 , y20667 , y20668 , y20669 , y20670 , y20671 , y20672 , y20673 , y20674 , y20675 , y20676 , y20677 , y20678 , y20679 , y20680 , y20681 , y20682 , y20683 , y20684 , y20685 , y20686 , y20687 , y20688 , y20689 , y20690 , y20691 , y20692 , y20693 , y20694 , y20695 , y20696 , y20697 , y20698 , y20699 , y20700 , y20701 , y20702 , y20703 , y20704 , y20705 , y20706 , y20707 , y20708 , y20709 , y20710 , y20711 , y20712 , y20713 , y20714 , y20715 , y20716 , y20717 , y20718 , y20719 , y20720 , y20721 , y20722 , y20723 , y20724 , y20725 , y20726 , y20727 , y20728 , y20729 , y20730 , y20731 , y20732 , y20733 , y20734 , y20735 , y20736 , y20737 , y20738 , y20739 , y20740 , y20741 , y20742 , y20743 , y20744 , y20745 , y20746 , y20747 , y20748 , y20749 , y20750 , y20751 , y20752 , y20753 , y20754 , y20755 , y20756 , y20757 , y20758 , y20759 , y20760 , y20761 , y20762 , y20763 , y20764 , y20765 , y20766 , y20767 , y20768 , y20769 , y20770 , y20771 , y20772 , y20773 , y20774 , y20775 , y20776 , y20777 , y20778 , y20779 , y20780 , y20781 , y20782 , y20783 , y20784 , y20785 , y20786 , y20787 , y20788 , y20789 , y20790 , y20791 , y20792 , y20793 , y20794 , y20795 , y20796 , y20797 , y20798 , y20799 , y20800 , y20801 , y20802 , y20803 , y20804 , y20805 , y20806 , y20807 , y20808 , y20809 , y20810 , y20811 , y20812 , y20813 , y20814 , y20815 , y20816 , y20817 , y20818 , y20819 , y20820 , y20821 , y20822 , y20823 , y20824 , y20825 , y20826 , y20827 , y20828 , y20829 , y20830 , y20831 , y20832 , y20833 , y20834 , y20835 , y20836 , y20837 , y20838 , y20839 , y20840 , y20841 , y20842 , y20843 , y20844 , y20845 , y20846 , y20847 , y20848 , y20849 , y20850 , y20851 , y20852 , y20853 , y20854 , y20855 , y20856 , y20857 , y20858 , y20859 , y20860 , y20861 , y20862 , y20863 , y20864 , y20865 , y20866 , y20867 , y20868 , y20869 , y20870 , y20871 , y20872 , y20873 , y20874 , y20875 , y20876 , y20877 , y20878 , y20879 , y20880 , y20881 , y20882 , y20883 , y20884 , y20885 , y20886 , y20887 , y20888 , y20889 , y20890 , y20891 , y20892 , y20893 , y20894 , y20895 , y20896 , y20897 , y20898 , y20899 , y20900 , y20901 , y20902 , y20903 , y20904 , y20905 , y20906 , y20907 , y20908 , y20909 , y20910 , y20911 , y20912 , y20913 , y20914 , y20915 , y20916 , y20917 , y20918 , y20919 , y20920 , y20921 , y20922 , y20923 , y20924 , y20925 , y20926 , y20927 , y20928 , y20929 , y20930 , y20931 , y20932 , y20933 , y20934 , y20935 , y20936 , y20937 , y20938 , y20939 , y20940 , y20941 , y20942 , y20943 , y20944 , y20945 , y20946 , y20947 , y20948 , y20949 , y20950 , y20951 , y20952 , y20953 , y20954 , y20955 , y20956 , y20957 , y20958 , y20959 , y20960 , y20961 , y20962 , y20963 , y20964 , y20965 , y20966 , y20967 , y20968 , y20969 , y20970 , y20971 , y20972 , y20973 , y20974 , y20975 , y20976 , y20977 , y20978 , y20979 , y20980 , y20981 , y20982 , y20983 , y20984 , y20985 , y20986 , y20987 , y20988 , y20989 , y20990 , y20991 , y20992 , y20993 , y20994 , y20995 , y20996 , y20997 , y20998 , y20999 , y21000 , y21001 , y21002 , y21003 , y21004 , y21005 , y21006 , y21007 , y21008 , y21009 , y21010 , y21011 , y21012 , y21013 , y21014 , y21015 , y21016 , y21017 , y21018 , y21019 , y21020 , y21021 , y21022 , y21023 , y21024 , y21025 , y21026 , y21027 , y21028 , y21029 , y21030 , y21031 , y21032 , y21033 , y21034 , y21035 , y21036 , y21037 , y21038 , y21039 , y21040 , y21041 , y21042 , y21043 , y21044 , y21045 , y21046 , y21047 , y21048 , y21049 , y21050 , y21051 , y21052 , y21053 , y21054 , y21055 , y21056 , y21057 , y21058 , y21059 , y21060 , y21061 , y21062 , y21063 , y21064 , y21065 , y21066 , y21067 , y21068 , y21069 , y21070 , y21071 , y21072 , y21073 , y21074 , y21075 , y21076 , y21077 , y21078 , y21079 , y21080 , y21081 , y21082 , y21083 , y21084 , y21085 , y21086 , y21087 , y21088 , y21089 , y21090 , y21091 , y21092 , y21093 , y21094 , y21095 , y21096 , y21097 , y21098 , y21099 , y21100 , y21101 , y21102 , y21103 , y21104 , y21105 , y21106 , y21107 , y21108 , y21109 , y21110 , y21111 , y21112 , y21113 , y21114 , y21115 , y21116 , y21117 , y21118 , y21119 , y21120 , y21121 , y21122 , y21123 , y21124 , y21125 , y21126 , y21127 , y21128 , y21129 , y21130 , y21131 , y21132 , y21133 , y21134 , y21135 , y21136 , y21137 , y21138 , y21139 , y21140 , y21141 , y21142 , y21143 , y21144 , y21145 , y21146 , y21147 , y21148 , y21149 , y21150 , y21151 , y21152 , y21153 , y21154 , y21155 , y21156 , y21157 , y21158 , y21159 , y21160 , y21161 , y21162 , y21163 , y21164 , y21165 , y21166 , y21167 , y21168 , y21169 , y21170 , y21171 , y21172 , y21173 , y21174 , y21175 , y21176 , y21177 , y21178 , y21179 , y21180 , y21181 , y21182 , y21183 , y21184 , y21185 , y21186 , y21187 , y21188 , y21189 , y21190 , y21191 , y21192 , y21193 , y21194 , y21195 , y21196 , y21197 , y21198 , y21199 , y21200 , y21201 , y21202 , y21203 , y21204 , y21205 , y21206 , y21207 , y21208 , y21209 , y21210 , y21211 , y21212 , y21213 , y21214 , y21215 , y21216 , y21217 , y21218 , y21219 , y21220 , y21221 , y21222 , y21223 , y21224 , y21225 , y21226 , y21227 , y21228 , y21229 , y21230 , y21231 , y21232 , y21233 , y21234 , y21235 , y21236 , y21237 , y21238 , y21239 , y21240 , y21241 , y21242 , y21243 , y21244 , y21245 , y21246 , y21247 , y21248 , y21249 , y21250 , y21251 , y21252 , y21253 , y21254 , y21255 , y21256 , y21257 , y21258 , y21259 , y21260 , y21261 , y21262 , y21263 , y21264 , y21265 , y21266 , y21267 , y21268 , y21269 , y21270 , y21271 , y21272 , y21273 , y21274 , y21275 , y21276 , y21277 , y21278 , y21279 , y21280 , y21281 , y21282 , y21283 , y21284 , y21285 , y21286 , y21287 , y21288 , y21289 , y21290 , y21291 , y21292 , y21293 , y21294 , y21295 , y21296 , y21297 , y21298 , y21299 , y21300 , y21301 , y21302 , y21303 , y21304 , y21305 , y21306 , y21307 , y21308 , y21309 , y21310 , y21311 , y21312 , y21313 , y21314 , y21315 , y21316 , y21317 , y21318 , y21319 , y21320 , y21321 , y21322 , y21323 , y21324 , y21325 , y21326 , y21327 , y21328 , y21329 , y21330 , y21331 , y21332 , y21333 , y21334 , y21335 , y21336 , y21337 , y21338 , y21339 ;
  wire n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , n46643 , n46644 , n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , n46674 , n46675 , n46676 , n46677 , n46678 , n46679 , n46680 , n46681 , n46682 , n46683 , n46684 , n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , n46711 , n46712 , n46713 , n46714 , n46715 , n46716 , n46717 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , n46725 , n46726 , n46727 , n46728 , n46729 , n46730 , n46731 , n46732 , n46733 , n46734 , n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , n46751 , n46752 , n46753 , n46754 , n46755 , n46756 , n46757 , n46758 , n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , n46765 , n46766 , n46767 , n46768 , n46769 , n46770 , n46771 , n46772 , n46773 , n46774 , n46775 , n46776 , n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , n46785 , n46786 , n46787 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , n46795 , n46796 , n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , n46805 , n46806 , n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , n46815 , n46816 , n46817 , n46818 , n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , n46835 , n46836 , n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , n46845 , n46846 , n46847 , n46848 , n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , n46855 , n46856 , n46857 , n46858 , n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , n46865 , n46866 , n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , n46895 , n46896 , n46897 , n46898 , n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , n46905 , n46906 , n46907 , n46908 , n46909 , n46910 , n46911 , n46912 , n46913 , n46914 , n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , n46924 , n46925 , n46926 , n46927 , n46928 , n46929 , n46930 , n46931 , n46932 , n46933 , n46934 , n46935 , n46936 , n46937 , n46938 , n46939 , n46940 , n46941 , n46942 , n46943 , n46944 , n46945 , n46946 , n46947 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , n46954 , n46955 , n46956 , n46957 , n46958 , n46959 , n46960 , n46961 , n46962 , n46963 , n46964 , n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , n46974 , n46975 , n46976 , n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , n46985 , n46986 , n46987 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , n46995 , n46996 , n46997 , n46998 , n46999 , n47000 , n47001 , n47002 , n47003 , n47004 , n47005 , n47006 , n47007 , n47008 , n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , n47015 , n47016 , n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , n47025 , n47026 , n47027 , n47028 , n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , n47035 , n47036 , n47037 , n47038 , n47039 , n47040 , n47041 , n47042 , n47043 , n47044 , n47045 , n47046 , n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n47053 , n47054 , n47055 , n47056 , n47057 , n47058 , n47059 , n47060 , n47061 , n47062 , n47063 , n47064 , n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , n47071 , n47072 , n47073 , n47074 , n47075 , n47076 , n47077 , n47078 , n47079 , n47080 , n47081 , n47082 , n47083 , n47084 , n47085 , n47086 , n47087 , n47088 , n47089 , n47090 , n47091 , n47092 , n47093 , n47094 , n47095 , n47096 , n47097 , n47098 , n47099 , n47100 , n47101 , n47102 , n47103 , n47104 , n47105 , n47106 , n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n47113 , n47114 , n47115 , n47116 , n47117 , n47118 , n47119 , n47120 , n47121 , n47122 , n47123 , n47124 , n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , n47131 , n47132 , n47133 , n47134 , n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , n47141 , n47142 , n47143 , n47144 , n47145 , n47146 , n47147 , n47148 , n47149 , n47150 , n47151 , n47152 , n47153 , n47154 , n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n47163 , n47164 , n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , n47185 , n47186 , n47187 , n47188 , n47189 , n47190 , n47191 , n47192 , n47193 , n47194 , n47195 , n47196 , n47197 , n47198 , n47199 , n47200 , n47201 , n47202 , n47203 , n47204 , n47205 , n47206 , n47207 , n47208 , n47209 , n47210 , n47211 , n47212 , n47213 , n47214 , n47215 , n47216 , n47217 , n47218 , n47219 , n47220 , n47221 , n47222 , n47223 , n47224 , n47225 , n47226 , n47227 , n47228 , n47229 , n47230 , n47231 , n47232 , n47233 , n47234 , n47235 , n47236 , n47237 , n47238 , n47239 , n47240 , n47241 , n47242 , n47243 , n47244 , n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , n47251 , n47252 , n47253 , n47254 , n47255 , n47256 , n47257 , n47258 , n47259 , n47260 , n47261 , n47262 , n47263 , n47264 , n47265 , n47266 , n47267 , n47268 , n47269 , n47270 , n47271 , n47272 , n47273 , n47274 , n47275 , n47276 , n47277 , n47278 , n47279 , n47280 , n47281 , n47282 , n47283 , n47284 , n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , n47291 , n47292 , n47293 , n47294 , n47295 , n47296 , n47297 , n47298 , n47299 , n47300 , n47301 , n47302 , n47303 , n47304 , n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , n47325 , n47326 , n47327 , n47328 , n47329 , n47330 , n47331 , n47332 , n47333 , n47334 , n47335 , n47336 , n47337 , n47338 , n47339 , n47340 , n47341 , n47342 , n47343 , n47344 , n47345 , n47346 , n47347 , n47348 , n47349 , n47350 , n47351 , n47352 , n47353 , n47354 , n47355 , n47356 , n47357 , n47358 , n47359 , n47360 , n47361 , n47362 , n47363 , n47364 , n47365 , n47366 , n47367 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , n47375 , n47376 , n47377 , n47378 , n47379 , n47380 , n47381 , n47382 , n47383 , n47384 , n47385 , n47386 , n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n47393 , n47394 , n47395 , n47396 , n47397 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , n47404 , n47405 , n47406 , n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , n47414 , n47415 , n47416 , n47417 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , n47424 , n47425 , n47426 , n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , n47435 , n47436 , n47437 , n47438 , n47439 , n47440 , n47441 , n47442 , n47443 , n47444 , n47445 , n47446 , n47447 , n47448 , n47449 , n47450 , n47451 , n47452 , n47453 , n47454 , n47455 , n47456 , n47457 , n47458 , n47459 , n47460 , n47461 , n47462 , n47463 , n47464 , n47465 , n47466 , n47467 , n47468 , n47469 , n47470 , n47471 , n47472 , n47473 , n47474 , n47475 , n47476 , n47477 , n47478 , n47479 , n47480 , n47481 , n47482 , n47483 , n47484 , n47485 , n47486 , n47487 , n47488 , n47489 , n47490 , n47491 , n47492 , n47493 , n47494 , n47495 , n47496 , n47497 , n47498 , n47499 , n47500 , n47501 , n47502 , n47503 , n47504 , n47505 , n47506 , n47507 , n47508 , n47509 , n47510 , n47511 , n47512 , n47513 , n47514 , n47515 , n47516 , n47517 , n47518 , n47519 , n47520 , n47521 , n47522 , n47523 , n47524 , n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , n47535 , n47536 , n47537 , n47538 , n47539 , n47540 , n47541 , n47542 , n47543 , n47544 , n47545 , n47546 , n47547 , n47548 , n47549 , n47550 , n47551 , n47552 , n47553 , n47554 , n47555 , n47556 , n47557 , n47558 , n47559 , n47560 , n47561 , n47562 , n47563 , n47564 , n47565 , n47566 , n47567 , n47568 , n47569 , n47570 , n47571 , n47572 , n47573 , n47574 , n47575 , n47576 , n47577 , n47578 , n47579 , n47580 , n47581 , n47582 , n47583 , n47584 , n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , n47591 , n47592 , n47593 , n47594 , n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , n47601 , n47602 , n47603 , n47604 , n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , n47611 , n47612 , n47613 , n47614 , n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , n47621 , n47622 , n47623 , n47624 , n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , n47641 , n47642 , n47643 , n47644 , n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , n47651 , n47652 , n47653 , n47654 , n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , n47661 , n47662 , n47663 , n47664 , n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , n47671 , n47672 , n47673 , n47674 , n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , n47691 , n47692 , n47693 , n47694 , n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , n47701 , n47702 , n47703 , n47704 , n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , n47711 , n47712 , n47713 , n47714 , n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , n47721 , n47722 , n47723 , n47724 , n47725 , n47726 , n47727 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , n47734 , n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , n47741 , n47742 , n47743 , n47744 , n47745 , n47746 , n47747 , n47748 , n47749 , n47750 , n47751 , n47752 , n47753 , n47754 , n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , n47765 , n47766 , n47767 , n47768 , n47769 , n47770 , n47771 , n47772 , n47773 , n47774 , n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , n47791 , n47792 , n47793 , n47794 , n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , n47801 , n47802 , n47803 , n47804 , n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , n47811 , n47812 , n47813 , n47814 , n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , n47821 , n47822 , n47823 , n47824 , n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , n47831 , n47832 , n47833 , n47834 , n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n47843 , n47844 , n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , n47861 , n47862 , n47863 , n47864 , n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , n47871 , n47872 , n47873 , n47874 , n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , n47881 , n47882 , n47883 , n47884 , n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , n47891 , n47892 , n47893 , n47894 , n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , n47901 , n47902 , n47903 , n47904 , n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , n47911 , n47912 , n47913 , n47914 , n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , n47921 , n47922 , n47923 , n47924 , n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , n47931 , n47932 , n47933 , n47934 , n47935 , n47936 , n47937 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , n47944 , n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , n47951 , n47952 , n47953 , n47954 , n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , n47981 , n47982 , n47983 , n47984 , n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , n47991 , n47992 , n47993 , n47994 , n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , n48001 , n48002 , n48003 , n48004 , n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , n48011 , n48012 , n48013 , n48014 , n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , n48021 , n48022 , n48023 , n48024 , n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , n48031 , n48032 , n48033 , n48034 , n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n48043 , n48044 , n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , n48051 , n48052 , n48053 , n48054 , n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , n48061 , n48062 , n48063 , n48064 , n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , n48071 , n48072 , n48073 , n48074 , n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , n48081 , n48082 , n48083 , n48084 , n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , n48101 , n48102 , n48103 , n48104 , n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , n48111 , n48112 , n48113 , n48114 , n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , n48121 , n48122 , n48123 , n48124 , n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , n48134 , n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , n48141 , n48142 , n48143 , n48144 , n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , n48151 , n48152 , n48153 , n48154 , n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , n48161 , n48162 , n48163 , n48164 , n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , n48191 , n48192 , n48193 , n48194 , n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , n48204 , n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n48213 , n48214 , n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , n48221 , n48222 , n48223 , n48224 , n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , n48231 , n48232 , n48233 , n48234 , n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , n48241 , n48242 , n48243 , n48244 , n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , n48251 , n48252 , n48253 , n48254 , n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , n48261 , n48262 , n48263 , n48264 , n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , n48271 , n48272 , n48273 , n48274 , n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , n48281 , n48282 , n48283 , n48284 , n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , n48291 , n48292 , n48293 , n48294 , n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , n48301 , n48302 , n48303 , n48304 , n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n48313 , n48314 , n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n48323 , n48324 , n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , n48331 , n48332 , n48333 , n48334 , n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , n48341 , n48342 , n48343 , n48344 , n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , n48351 , n48352 , n48353 , n48354 , n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , n48361 , n48362 , n48363 , n48364 , n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , n48371 , n48372 , n48373 , n48374 , n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , n48381 , n48382 , n48383 , n48384 , n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , n48394 , n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , n48401 , n48402 , n48403 , n48404 , n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , n48411 , n48412 , n48413 , n48414 , n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , n48421 , n48422 , n48423 , n48424 , n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n48433 , n48434 , n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , n48441 , n48442 , n48443 , n48444 , n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48453 , n48454 , n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , n48461 , n48462 , n48463 , n48464 , n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , n48471 , n48472 , n48473 , n48474 , n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n48493 , n48494 , n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , n48501 , n48502 , n48503 , n48504 , n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , n48511 , n48512 , n48513 , n48514 , n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , n48521 , n48522 , n48523 , n48524 , n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , n48531 , n48532 , n48533 , n48534 , n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , n48541 , n48542 , n48543 , n48544 , n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , n48551 , n48552 , n48553 , n48554 , n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , n48561 , n48562 , n48563 , n48564 , n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , n48571 , n48572 , n48573 , n48574 , n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , n48581 , n48582 , n48583 , n48584 , n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , n48591 , n48592 , n48593 , n48594 , n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , n48601 , n48602 , n48603 , n48604 , n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , n48611 , n48612 , n48613 , n48614 , n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , n48621 , n48622 , n48623 , n48624 , n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , n48651 , n48652 , n48653 , n48654 , n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n48663 , n48664 , n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , n48671 , n48672 , n48673 , n48674 , n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , n48681 , n48682 , n48683 , n48684 , n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n48693 , n48694 , n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , n48701 , n48702 , n48703 , n48704 , n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , n48711 , n48712 , n48713 , n48714 , n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , n48731 , n48732 , n48733 , n48734 , n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48753 , n48754 , n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , n48761 , n48762 , n48763 , n48764 , n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , n48774 , n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , n48781 , n48782 , n48783 , n48784 , n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , n48791 , n48792 , n48793 , n48794 , n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , n48804 , n48805 , n48806 , n48807 , n48808 , n48809 , n48810 , n48811 , n48812 , n48813 , n48814 , n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , n48821 , n48822 , n48823 , n48824 , n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , n48834 , n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , n48841 , n48842 , n48843 , n48844 , n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , n48851 , n48852 , n48853 , n48854 , n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 , n48864 , n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , n48881 , n48882 , n48883 , n48884 , n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , n48901 , n48902 , n48903 , n48904 , n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , n48921 , n48922 , n48923 , n48924 , n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , n48941 , n48942 , n48943 , n48944 , n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , n48961 , n48962 , n48963 , n48964 , n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , n48981 , n48982 , n48983 , n48984 , n48985 , n48986 , n48987 , n48988 , n48989 , n48990 , n48991 , n48992 , n48993 , n48994 , n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , n49001 , n49002 , n49003 , n49004 , n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , n49011 , n49012 , n49013 , n49014 , n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , n49024 , n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , n49051 , n49052 , n49053 , n49054 , n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , n49061 , n49062 , n49063 , n49064 , n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n49073 , n49074 , n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , n49081 , n49082 , n49083 , n49084 , n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , n49091 , n49092 , n49093 , n49094 , n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , n49101 , n49102 , n49103 , n49104 , n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , n49111 , n49112 , n49113 , n49114 , n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , n49124 , n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , n49131 , n49132 , n49133 , n49134 , n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , n49141 , n49142 , n49143 , n49144 , n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n49153 , n49154 , n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , n49161 , n49162 , n49163 , n49164 , n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , n49171 , n49172 , n49173 , n49174 , n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , n49194 , n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n49213 , n49214 , n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , n49221 , n49222 , n49223 , n49224 , n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , n49231 , n49232 , n49233 , n49234 , n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , n49241 , n49242 , n49243 , n49244 , n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , n49251 , n49252 , n49253 , n49254 , n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , n49261 , n49262 , n49263 , n49264 , n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , n49281 , n49282 , n49283 , n49284 , n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , n49294 , n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , n49301 , n49302 , n49303 , n49304 , n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , n49311 , n49312 , n49313 , n49314 , n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , n49321 , n49322 , n49323 , n49324 , n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , n49331 , n49332 , n49333 , n49334 , n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , n49351 , n49352 , n49353 , n49354 , n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , n49391 , n49392 , n49393 , n49394 , n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , n49411 , n49412 , n49413 , n49414 , n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , n49421 , n49422 , n49423 , n49424 , n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , n49431 , n49432 , n49433 , n49434 , n49435 , n49436 , n49437 , n49438 , n49439 , n49440 , n49441 , n49442 , n49443 , n49444 , n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , n49451 , n49452 , n49453 , n49454 , n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , n49461 , n49462 , n49463 , n49464 , n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , n49471 , n49472 , n49473 , n49474 , n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , n49481 , n49482 , n49483 , n49484 , n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , n49491 , n49492 , n49493 , n49494 , n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , n49501 , n49502 , n49503 , n49504 , n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , n49511 , n49512 , n49513 , n49514 , n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , n49521 , n49522 , n49523 , n49524 , n49525 , n49526 , n49527 , n49528 , n49529 ;
  assign n256 = x69 ^ x44 ^ x33 ;
  assign n257 = x227 ^ x87 ^ x69 ;
  assign n258 = x169 & x252 ;
  assign n259 = n258 ^ x87 ^ 1'b0 ;
  assign n260 = x209 ^ x153 ^ x110 ;
  assign n261 = x85 & x180 ;
  assign n262 = n261 ^ x64 ^ 1'b0 ;
  assign n263 = ( x5 & ~x11 ) | ( x5 & x161 ) | ( ~x11 & x161 ) ;
  assign n264 = x253 ^ x28 ^ x6 ;
  assign n265 = x251 ^ x53 ^ 1'b0 ;
  assign n266 = x163 & n265 ;
  assign n267 = x86 & x171 ;
  assign n268 = n267 ^ x50 ^ 1'b0 ;
  assign n269 = x252 ^ x251 ^ x244 ;
  assign n270 = ( x159 & n257 ) | ( x159 & n269 ) | ( n257 & n269 ) ;
  assign n271 = ( x151 & x225 ) | ( x151 & n259 ) | ( x225 & n259 ) ;
  assign n272 = x207 & x235 ;
  assign n273 = ~x211 & n272 ;
  assign n274 = x174 & ~n273 ;
  assign n275 = ~x180 & n274 ;
  assign n276 = x36 & x236 ;
  assign n277 = n276 ^ x125 ^ 1'b0 ;
  assign n278 = x69 ^ x36 ^ 1'b0 ;
  assign n279 = x152 & n278 ;
  assign n280 = n279 ^ x125 ^ x29 ;
  assign n281 = x6 & x215 ;
  assign n282 = ~x13 & n281 ;
  assign n283 = x21 & x74 ;
  assign n284 = ~x90 & n283 ;
  assign n285 = x90 & x248 ;
  assign n286 = n285 ^ x211 ^ 1'b0 ;
  assign n287 = ( x215 & ~x223 ) | ( x215 & n286 ) | ( ~x223 & n286 ) ;
  assign n288 = x166 ^ x94 ^ x56 ;
  assign n289 = n268 | n288 ;
  assign n290 = x152 | n289 ;
  assign n291 = x84 ^ x64 ^ 1'b0 ;
  assign n292 = ~n282 & n291 ;
  assign n293 = ( x122 & ~x156 ) | ( x122 & n284 ) | ( ~x156 & n284 ) ;
  assign n294 = x30 & ~x237 ;
  assign n295 = x95 ^ x81 ^ 1'b0 ;
  assign n297 = x237 ^ x134 ^ x0 ;
  assign n296 = x53 & x109 ;
  assign n298 = n297 ^ n296 ^ 1'b0 ;
  assign n299 = n284 ^ x198 ^ 1'b0 ;
  assign n300 = x249 & ~n299 ;
  assign n301 = x32 & x214 ;
  assign n302 = n301 ^ x129 ^ 1'b0 ;
  assign n303 = x1 & n302 ;
  assign n304 = x223 ^ x123 ^ x61 ;
  assign n305 = ( x146 & ~x252 ) | ( x146 & n304 ) | ( ~x252 & n304 ) ;
  assign n306 = x49 & ~n305 ;
  assign n307 = ~x225 & n306 ;
  assign n308 = n307 ^ x157 ^ x71 ;
  assign n309 = x13 & x28 ;
  assign n310 = n309 ^ x74 ^ 1'b0 ;
  assign n311 = x63 & x139 ;
  assign n312 = n311 ^ x252 ^ 1'b0 ;
  assign n313 = x80 & ~n312 ;
  assign n314 = ~n308 & n313 ;
  assign n315 = x59 & x157 ;
  assign n316 = ~x179 & n315 ;
  assign n317 = ( ~x47 & x216 ) | ( ~x47 & n316 ) | ( x216 & n316 ) ;
  assign n318 = ( x100 & ~x160 ) | ( x100 & x193 ) | ( ~x160 & x193 ) ;
  assign n319 = x76 ^ x2 ^ 1'b0 ;
  assign n320 = x232 & n319 ;
  assign n321 = x178 & n271 ;
  assign n322 = ~n320 & n321 ;
  assign n324 = x143 & x182 ;
  assign n325 = n324 ^ x33 ^ 1'b0 ;
  assign n326 = ( x9 & ~x213 ) | ( x9 & n325 ) | ( ~x213 & n325 ) ;
  assign n323 = ( ~x36 & x114 ) | ( ~x36 & x188 ) | ( x114 & x188 ) ;
  assign n327 = n326 ^ n323 ^ 1'b0 ;
  assign n328 = x169 ^ x57 ^ 1'b0 ;
  assign n329 = x117 & n328 ;
  assign n330 = x250 & ~n329 ;
  assign n331 = x114 & x144 ;
  assign n332 = ~x165 & n331 ;
  assign n333 = x243 ^ x159 ^ x69 ;
  assign n334 = n332 & ~n333 ;
  assign n335 = x160 ^ x52 ^ 1'b0 ;
  assign n343 = x164 ^ x58 ^ x37 ;
  assign n344 = n343 ^ x88 ^ x83 ;
  assign n336 = x196 ^ x166 ^ 1'b0 ;
  assign n337 = x139 & n336 ;
  assign n338 = x173 ^ x26 ^ x5 ;
  assign n339 = n338 ^ x207 ^ x79 ;
  assign n340 = x159 & n339 ;
  assign n341 = n340 ^ n269 ^ 1'b0 ;
  assign n342 = n337 & n341 ;
  assign n345 = n344 ^ n342 ^ 1'b0 ;
  assign n346 = n345 ^ x252 ^ 1'b0 ;
  assign n347 = x168 & ~n346 ;
  assign n348 = x17 & x101 ;
  assign n349 = ~x165 & n348 ;
  assign n350 = n349 ^ n307 ^ 1'b0 ;
  assign n351 = n271 ^ x108 ^ x37 ;
  assign n352 = n284 ^ x205 ^ x186 ;
  assign n353 = x216 & n279 ;
  assign n354 = ~n352 & n353 ;
  assign n361 = x54 & x76 ;
  assign n362 = ~x223 & n361 ;
  assign n355 = n259 ^ x165 ^ 1'b0 ;
  assign n356 = x72 & ~n355 ;
  assign n357 = x8 & n356 ;
  assign n358 = n357 ^ x98 ^ 1'b0 ;
  assign n359 = n358 ^ x180 ^ 1'b0 ;
  assign n360 = x81 & ~n359 ;
  assign n363 = n362 ^ n360 ^ x32 ;
  assign n364 = x81 ^ x66 ^ 1'b0 ;
  assign n365 = x25 & n364 ;
  assign n366 = ( x79 & x132 ) | ( x79 & ~x230 ) | ( x132 & ~x230 ) ;
  assign n373 = x97 & x148 ;
  assign n374 = n373 ^ n343 ^ 1'b0 ;
  assign n367 = x88 & x181 ;
  assign n368 = n367 ^ x172 ^ 1'b0 ;
  assign n369 = x249 ^ x56 ^ x43 ;
  assign n370 = n368 | n369 ;
  assign n371 = x148 | n370 ;
  assign n372 = x246 & n371 ;
  assign n375 = n374 ^ n372 ^ 1'b0 ;
  assign n383 = x168 & x207 ;
  assign n384 = n383 ^ x65 ^ 1'b0 ;
  assign n376 = x23 & x219 ;
  assign n377 = ~x227 & n376 ;
  assign n378 = n332 ^ x20 ^ 1'b0 ;
  assign n379 = x156 & ~x200 ;
  assign n380 = x29 & ~n379 ;
  assign n381 = n378 & n380 ;
  assign n382 = ( x19 & ~n377 ) | ( x19 & n381 ) | ( ~n377 & n381 ) ;
  assign n385 = n384 ^ n382 ^ n337 ;
  assign n386 = ( x134 & x212 ) | ( x134 & ~x234 ) | ( x212 & ~x234 ) ;
  assign n387 = n386 ^ x1 ^ 1'b0 ;
  assign n388 = x48 & x156 ;
  assign n389 = ~n387 & n388 ;
  assign n390 = x105 ^ x91 ^ 1'b0 ;
  assign n391 = n264 ^ x24 ^ 1'b0 ;
  assign n392 = x142 ^ x140 ^ 1'b0 ;
  assign n393 = x211 & n392 ;
  assign n394 = ( x126 & x208 ) | ( x126 & ~x228 ) | ( x208 & ~x228 ) ;
  assign n395 = x23 & n394 ;
  assign n396 = n395 ^ x235 ^ 1'b0 ;
  assign n397 = x13 & x14 ;
  assign n398 = n397 ^ x246 ^ 1'b0 ;
  assign n399 = ( x45 & ~x64 ) | ( x45 & x156 ) | ( ~x64 & x156 ) ;
  assign n400 = x139 & x237 ;
  assign n401 = ~n399 & n400 ;
  assign n402 = ( ~x169 & x220 ) | ( ~x169 & x223 ) | ( x220 & x223 ) ;
  assign n403 = ( ~x3 & x165 ) | ( ~x3 & n343 ) | ( x165 & n343 ) ;
  assign n404 = x86 ^ x56 ^ 1'b0 ;
  assign n405 = x224 & n404 ;
  assign n406 = n405 ^ x148 ^ 1'b0 ;
  assign n407 = x43 & n406 ;
  assign n408 = x208 & x224 ;
  assign n409 = n408 ^ x238 ^ 1'b0 ;
  assign n410 = ( x11 & ~x127 ) | ( x11 & n409 ) | ( ~x127 & n409 ) ;
  assign n411 = ( ~x92 & x229 ) | ( ~x92 & n410 ) | ( x229 & n410 ) ;
  assign n412 = x84 | n411 ;
  assign n413 = x197 ^ x136 ^ x83 ;
  assign n414 = x234 ^ x80 ^ 1'b0 ;
  assign n415 = x180 & n414 ;
  assign n416 = n415 ^ x35 ^ 1'b0 ;
  assign n417 = ~n302 & n416 ;
  assign n418 = x183 & x197 ;
  assign n419 = ~x154 & n418 ;
  assign n420 = x144 & ~n419 ;
  assign n421 = n420 ^ x133 ^ 1'b0 ;
  assign n426 = x179 ^ x124 ^ x13 ;
  assign n427 = n426 ^ x170 ^ 1'b0 ;
  assign n428 = n427 ^ x236 ^ x224 ;
  assign n423 = ( x37 & ~x185 ) | ( x37 & n386 ) | ( ~x185 & n386 ) ;
  assign n422 = x47 & x71 ;
  assign n424 = n423 ^ n422 ^ 1'b0 ;
  assign n425 = x30 & ~n424 ;
  assign n429 = n428 ^ n425 ^ 1'b0 ;
  assign n430 = ~n421 & n429 ;
  assign n431 = x89 & x151 ;
  assign n432 = n431 ^ x187 ^ 1'b0 ;
  assign n433 = x21 & x180 ;
  assign n434 = ( ~n326 & n432 ) | ( ~n326 & n433 ) | ( n432 & n433 ) ;
  assign n435 = ( x81 & ~x178 ) | ( x81 & x230 ) | ( ~x178 & x230 ) ;
  assign n436 = ( x217 & ~x231 ) | ( x217 & n435 ) | ( ~x231 & n435 ) ;
  assign n437 = n293 ^ x163 ^ 1'b0 ;
  assign n438 = n362 | n437 ;
  assign n439 = x177 & ~n317 ;
  assign n440 = ~x234 & n439 ;
  assign n441 = ~n438 & n440 ;
  assign n442 = ( ~n377 & n436 ) | ( ~n377 & n441 ) | ( n436 & n441 ) ;
  assign n446 = x100 ^ x81 ^ 1'b0 ;
  assign n447 = x198 & n446 ;
  assign n448 = x201 & n447 ;
  assign n449 = n448 ^ x247 ^ 1'b0 ;
  assign n443 = x77 ^ x35 ^ 1'b0 ;
  assign n444 = x11 & n443 ;
  assign n445 = n444 ^ n271 ^ x101 ;
  assign n450 = n449 ^ n445 ^ x215 ;
  assign n451 = n449 ^ x216 ^ x56 ;
  assign n452 = x27 & n451 ;
  assign n453 = ~x144 & n452 ;
  assign n454 = x139 ^ x107 ^ 1'b0 ;
  assign n455 = n271 ^ x47 ^ x8 ;
  assign n456 = n455 ^ n385 ^ 1'b0 ;
  assign n457 = x19 & ~n456 ;
  assign n458 = x57 & x168 ;
  assign n459 = ~x187 & n458 ;
  assign n460 = ~n287 & n459 ;
  assign n461 = ( x97 & x108 ) | ( x97 & n445 ) | ( x108 & n445 ) ;
  assign n462 = ( x117 & n460 ) | ( x117 & ~n461 ) | ( n460 & ~n461 ) ;
  assign n463 = x29 & ~n334 ;
  assign n464 = ~x86 & n463 ;
  assign n466 = x51 & x57 ;
  assign n467 = n466 ^ x228 ^ 1'b0 ;
  assign n468 = x223 ^ x163 ^ x114 ;
  assign n469 = ~n467 & n468 ;
  assign n470 = n469 ^ x207 ^ 1'b0 ;
  assign n471 = x232 & ~n470 ;
  assign n465 = x151 & ~n332 ;
  assign n472 = n471 ^ n465 ^ 1'b0 ;
  assign n473 = n472 ^ n354 ^ 1'b0 ;
  assign n474 = x159 & n473 ;
  assign n475 = x79 & n474 ;
  assign n476 = x199 ^ x194 ^ x107 ;
  assign n477 = x168 & ~n334 ;
  assign n478 = n362 & n477 ;
  assign n479 = ( x209 & n476 ) | ( x209 & ~n478 ) | ( n476 & ~n478 ) ;
  assign n480 = x180 ^ x75 ^ 1'b0 ;
  assign n481 = x149 & n480 ;
  assign n482 = x78 & ~n481 ;
  assign n483 = n482 ^ n320 ^ x206 ;
  assign n484 = n286 ^ x66 ^ 1'b0 ;
  assign n485 = x230 & ~n484 ;
  assign n486 = x192 ^ x181 ^ 1'b0 ;
  assign n487 = x96 & n486 ;
  assign n488 = x250 & n487 ;
  assign n489 = n488 ^ x7 ^ 1'b0 ;
  assign n492 = x106 & x207 ;
  assign n493 = n492 ^ x111 ^ 1'b0 ;
  assign n490 = ( ~x10 & x188 ) | ( ~x10 & n432 ) | ( x188 & n432 ) ;
  assign n494 = n490 ^ n310 ^ 1'b0 ;
  assign n495 = ~n493 & n494 ;
  assign n491 = n445 | n490 ;
  assign n496 = n495 ^ n491 ^ 1'b0 ;
  assign n497 = n300 & ~n343 ;
  assign n498 = ~n451 & n497 ;
  assign n499 = n498 ^ x78 ^ 1'b0 ;
  assign n500 = ( n489 & n496 ) | ( n489 & ~n499 ) | ( n496 & ~n499 ) ;
  assign n501 = n407 ^ x74 ^ x12 ;
  assign n502 = x12 & ~n498 ;
  assign n503 = n502 ^ x2 ^ 1'b0 ;
  assign n504 = x160 ^ x146 ^ 1'b0 ;
  assign n505 = x128 & n504 ;
  assign n510 = x54 ^ x9 ^ 1'b0 ;
  assign n511 = ~n332 & n510 ;
  assign n506 = x235 & ~n277 ;
  assign n507 = n506 ^ x44 ^ 1'b0 ;
  assign n508 = x83 & ~n507 ;
  assign n509 = ~n356 & n508 ;
  assign n512 = n511 ^ n509 ^ 1'b0 ;
  assign n513 = n479 ^ x162 ^ 1'b0 ;
  assign n514 = n513 ^ n339 ^ x108 ;
  assign n515 = ( x119 & ~x148 ) | ( x119 & n450 ) | ( ~x148 & n450 ) ;
  assign n516 = ( x71 & ~x135 ) | ( x71 & x207 ) | ( ~x135 & x207 ) ;
  assign n517 = n469 ^ x139 ^ x48 ;
  assign n518 = n517 ^ n447 ^ x184 ;
  assign n526 = x182 & n308 ;
  assign n527 = n526 ^ x190 ^ 1'b0 ;
  assign n519 = x162 ^ x100 ^ 1'b0 ;
  assign n523 = n284 & n341 ;
  assign n520 = x193 ^ x44 ^ x16 ;
  assign n521 = n520 ^ n320 ^ 1'b0 ;
  assign n522 = x100 & ~n521 ;
  assign n524 = n523 ^ n522 ^ 1'b0 ;
  assign n525 = n519 | n524 ;
  assign n528 = n527 ^ n525 ^ n427 ;
  assign n529 = n356 & n528 ;
  assign n530 = n529 ^ x96 ^ 1'b0 ;
  assign n531 = ( x29 & ~x47 ) | ( x29 & x106 ) | ( ~x47 & x106 ) ;
  assign n532 = n399 & n531 ;
  assign n533 = n532 ^ x240 ^ 1'b0 ;
  assign n535 = ( x10 & ~x241 ) | ( x10 & n326 ) | ( ~x241 & n326 ) ;
  assign n534 = x223 & n339 ;
  assign n536 = n535 ^ n534 ^ 1'b0 ;
  assign n537 = ( x49 & x87 ) | ( x49 & ~x243 ) | ( x87 & ~x243 ) ;
  assign n538 = x233 ^ x179 ^ x31 ;
  assign n539 = ( x179 & x223 ) | ( x179 & n326 ) | ( x223 & n326 ) ;
  assign n540 = ( ~x183 & n538 ) | ( ~x183 & n539 ) | ( n538 & n539 ) ;
  assign n541 = n537 & ~n540 ;
  assign n542 = n541 ^ x107 ^ 1'b0 ;
  assign n543 = x137 & x161 ;
  assign n544 = n543 ^ x44 ^ 1'b0 ;
  assign n545 = ( ~x61 & x202 ) | ( ~x61 & n544 ) | ( x202 & n544 ) ;
  assign n546 = n270 | n545 ;
  assign n547 = x100 | n546 ;
  assign n548 = x216 & n547 ;
  assign n549 = ~x156 & n548 ;
  assign n550 = x28 & ~n298 ;
  assign n551 = ~n269 & n407 ;
  assign n552 = n550 & n551 ;
  assign n553 = x54 & ~n469 ;
  assign n554 = ~x9 & n553 ;
  assign n555 = n554 ^ x48 ^ 1'b0 ;
  assign n556 = x191 & ~n555 ;
  assign n557 = ( x46 & x68 ) | ( x46 & ~x105 ) | ( x68 & ~x105 ) ;
  assign n558 = x240 & n557 ;
  assign n559 = n558 ^ x247 ^ 1'b0 ;
  assign n560 = n426 | n545 ;
  assign n561 = n339 ^ x195 ^ x82 ;
  assign n562 = n561 ^ x27 ^ x11 ;
  assign n563 = ( x174 & n287 ) | ( x174 & n562 ) | ( n287 & n562 ) ;
  assign n564 = ~n335 & n563 ;
  assign n565 = n564 ^ n356 ^ 1'b0 ;
  assign n566 = n565 ^ n302 ^ 1'b0 ;
  assign n567 = x62 & n566 ;
  assign n568 = x8 & x19 ;
  assign n569 = ~x88 & n568 ;
  assign n570 = x146 ^ x98 ^ 1'b0 ;
  assign n571 = ~n569 & n570 ;
  assign n572 = n559 ^ x176 ^ 1'b0 ;
  assign n573 = ~x206 & x211 ;
  assign n574 = ( ~x149 & n343 ) | ( ~x149 & n573 ) | ( n343 & n573 ) ;
  assign n575 = ( n320 & n333 ) | ( n320 & n467 ) | ( n333 & n467 ) ;
  assign n576 = n575 ^ n297 ^ x138 ;
  assign n577 = n398 | n576 ;
  assign n578 = x144 & n402 ;
  assign n579 = n302 ^ n298 ^ 1'b0 ;
  assign n580 = n360 & ~n579 ;
  assign n581 = ~n424 & n580 ;
  assign n582 = n581 ^ n499 ^ 1'b0 ;
  assign n587 = n462 ^ n337 ^ 1'b0 ;
  assign n583 = x27 & x124 ;
  assign n584 = ~x233 & n583 ;
  assign n585 = n308 ^ x2 ^ 1'b0 ;
  assign n586 = ~n584 & n585 ;
  assign n588 = n587 ^ n586 ^ x147 ;
  assign n589 = x104 & ~x158 ;
  assign n590 = n589 ^ n318 ^ 1'b0 ;
  assign n591 = n511 & n590 ;
  assign n592 = x215 ^ x49 ^ 1'b0 ;
  assign n593 = x178 & n592 ;
  assign n594 = n593 ^ n394 ^ 1'b0 ;
  assign n595 = x89 & n594 ;
  assign n596 = x192 ^ x181 ^ x34 ;
  assign n597 = n415 & n596 ;
  assign n598 = n476 | n561 ;
  assign n599 = n598 ^ x196 ^ 1'b0 ;
  assign n600 = ~n517 & n599 ;
  assign n601 = n540 ^ x184 ^ 1'b0 ;
  assign n602 = x110 & ~n601 ;
  assign n603 = ( ~x67 & x142 ) | ( ~x67 & n602 ) | ( x142 & n602 ) ;
  assign n604 = ~x17 & x190 ;
  assign n605 = x81 & ~n378 ;
  assign n606 = n396 & n605 ;
  assign n607 = x203 & x227 ;
  assign n608 = n607 ^ x249 ^ 1'b0 ;
  assign n609 = n379 | n608 ;
  assign n610 = n609 ^ n288 ^ 1'b0 ;
  assign n611 = n308 & ~n453 ;
  assign n612 = n611 ^ x146 ^ 1'b0 ;
  assign n613 = x243 ^ x116 ^ 1'b0 ;
  assign n614 = x151 & n613 ;
  assign n615 = n614 ^ n266 ^ x204 ;
  assign n616 = n615 ^ x96 ^ 1'b0 ;
  assign n617 = n616 ^ n475 ^ 1'b0 ;
  assign n618 = n330 ^ n266 ^ 1'b0 ;
  assign n619 = n445 | n618 ;
  assign n620 = n430 | n619 ;
  assign n621 = x246 & x252 ;
  assign n622 = ~n396 & n621 ;
  assign n623 = n622 ^ x91 ^ 1'b0 ;
  assign n624 = x71 ^ x44 ^ 1'b0 ;
  assign n625 = x189 & n624 ;
  assign n626 = ~n264 & n625 ;
  assign n627 = n626 ^ n316 ^ 1'b0 ;
  assign n628 = n394 & n627 ;
  assign n629 = n623 & n628 ;
  assign n630 = n481 ^ x43 ^ 1'b0 ;
  assign n631 = ( x103 & ~x223 ) | ( x103 & n333 ) | ( ~x223 & n333 ) ;
  assign n632 = n631 ^ x156 ^ 1'b0 ;
  assign n633 = ( ~x7 & n320 ) | ( ~x7 & n632 ) | ( n320 & n632 ) ;
  assign n634 = n633 ^ n294 ^ 1'b0 ;
  assign n635 = x48 & ~n634 ;
  assign n636 = x66 & ~n445 ;
  assign n637 = n636 ^ n312 ^ 1'b0 ;
  assign n638 = ~n562 & n637 ;
  assign n639 = n630 ^ x231 ^ 1'b0 ;
  assign n640 = x40 & ~n385 ;
  assign n641 = x119 & ~n604 ;
  assign n642 = n641 ^ x16 ^ 1'b0 ;
  assign n643 = n266 & n399 ;
  assign n644 = ~x2 & n643 ;
  assign n645 = n569 ^ n399 ^ x229 ;
  assign n646 = n645 ^ x223 ^ 1'b0 ;
  assign n647 = ~n644 & n646 ;
  assign n648 = n415 & n647 ;
  assign n649 = n642 & n648 ;
  assign n650 = x154 & x178 ;
  assign n651 = n650 ^ x3 ^ 1'b0 ;
  assign n652 = n363 ^ x63 ^ 1'b0 ;
  assign n653 = x174 ^ x25 ^ 1'b0 ;
  assign n654 = x178 & n653 ;
  assign n655 = n394 & ~n654 ;
  assign n656 = ( ~n472 & n576 ) | ( ~n472 & n655 ) | ( n576 & n655 ) ;
  assign n659 = x61 | n312 ;
  assign n657 = n493 ^ n481 ^ 1'b0 ;
  assign n658 = x148 & ~n657 ;
  assign n660 = n659 ^ n658 ^ 1'b0 ;
  assign n670 = n308 ^ x87 ^ 1'b0 ;
  assign n671 = n562 & n670 ;
  assign n661 = n485 ^ n307 ^ x55 ;
  assign n666 = x190 & x231 ;
  assign n667 = ~x177 & n666 ;
  assign n662 = x216 & x219 ;
  assign n663 = ~n614 & n662 ;
  assign n664 = x15 & ~n663 ;
  assign n665 = n664 ^ x163 ^ 1'b0 ;
  assign n668 = n667 ^ n665 ^ x61 ;
  assign n669 = ( ~n297 & n661 ) | ( ~n297 & n668 ) | ( n661 & n668 ) ;
  assign n672 = n671 ^ n669 ^ x60 ;
  assign n673 = n365 ^ x21 ^ 1'b0 ;
  assign n695 = n535 ^ x55 ^ 1'b0 ;
  assign n696 = n667 | n695 ;
  assign n674 = x217 & x232 ;
  assign n675 = n674 ^ x52 ^ 1'b0 ;
  assign n676 = n675 ^ n275 ^ x47 ;
  assign n677 = n676 ^ x250 ^ x198 ;
  assign n678 = n677 ^ n523 ^ x70 ;
  assign n679 = ( x195 & n467 ) | ( x195 & n678 ) | ( n467 & n678 ) ;
  assign n680 = ( x0 & x127 ) | ( x0 & ~n679 ) | ( x127 & ~n679 ) ;
  assign n690 = ~x83 & n292 ;
  assign n691 = n690 ^ n593 ^ n390 ;
  assign n681 = x129 ^ x24 ^ 1'b0 ;
  assign n682 = x16 & n681 ;
  assign n683 = n268 ^ x105 ^ 1'b0 ;
  assign n684 = n338 | n683 ;
  assign n685 = x51 & ~n684 ;
  assign n686 = ~n682 & n685 ;
  assign n687 = n560 ^ n487 ^ 1'b0 ;
  assign n688 = n686 | n687 ;
  assign n689 = x41 & ~n688 ;
  assign n692 = n691 ^ n689 ^ 1'b0 ;
  assign n693 = n680 & ~n692 ;
  assign n694 = n398 & n693 ;
  assign n697 = n696 ^ n694 ^ x146 ;
  assign n698 = n374 & n610 ;
  assign n699 = ~n428 & n698 ;
  assign n700 = n339 ^ x211 ^ 1'b0 ;
  assign n701 = ~n554 & n700 ;
  assign n702 = n603 & ~n701 ;
  assign n703 = ( n533 & ~n604 ) | ( n533 & n697 ) | ( ~n604 & n697 ) ;
  assign n704 = n430 ^ n390 ^ x18 ;
  assign n705 = x233 & n704 ;
  assign n706 = ~n536 & n705 ;
  assign n707 = n523 ^ x34 ^ 1'b0 ;
  assign n708 = n478 | n707 ;
  assign n712 = x130 & ~n256 ;
  assign n713 = n712 ^ x109 ^ 1'b0 ;
  assign n709 = ( x78 & x113 ) | ( x78 & ~x163 ) | ( x113 & ~x163 ) ;
  assign n710 = n709 ^ x72 ^ 1'b0 ;
  assign n711 = ( x35 & n569 ) | ( x35 & ~n710 ) | ( n569 & ~n710 ) ;
  assign n714 = n713 ^ n711 ^ 1'b0 ;
  assign n715 = ~n708 & n714 ;
  assign n716 = n316 | n428 ;
  assign n717 = ( x219 & ~n472 ) | ( x219 & n608 ) | ( ~n472 & n608 ) ;
  assign n718 = ( n715 & ~n716 ) | ( n715 & n717 ) | ( ~n716 & n717 ) ;
  assign n719 = x50 & x165 ;
  assign n720 = n297 & n719 ;
  assign n721 = x242 & n308 ;
  assign n722 = n720 & n721 ;
  assign n723 = ( x182 & n615 ) | ( x182 & ~n722 ) | ( n615 & ~n722 ) ;
  assign n724 = n450 ^ n407 ^ 1'b0 ;
  assign n725 = n436 & ~n724 ;
  assign n726 = n725 ^ x227 ^ 1'b0 ;
  assign n727 = ~n620 & n726 ;
  assign n728 = n669 & n715 ;
  assign n729 = n728 ^ x196 ^ 1'b0 ;
  assign n730 = x125 ^ x112 ^ 1'b0 ;
  assign n731 = ~n302 & n730 ;
  assign n732 = x122 & x127 ;
  assign n733 = n493 & n732 ;
  assign n734 = n273 | n733 ;
  assign n735 = n731 | n734 ;
  assign n736 = n735 ^ n696 ^ 1'b0 ;
  assign n737 = x9 & ~x247 ;
  assign n738 = x54 & n737 ;
  assign n739 = x112 & ~n469 ;
  assign n740 = n544 & n739 ;
  assign n741 = ( ~x169 & x223 ) | ( ~x169 & n663 ) | ( x223 & n663 ) ;
  assign n742 = n469 | n741 ;
  assign n743 = n742 ^ n512 ^ 1'b0 ;
  assign n744 = n743 ^ x211 ^ 1'b0 ;
  assign n745 = x133 & n744 ;
  assign n746 = x75 ^ x40 ^ 1'b0 ;
  assign n747 = ~n333 & n746 ;
  assign n748 = n747 ^ n717 ^ 1'b0 ;
  assign n749 = x151 & n747 ;
  assign n750 = n749 ^ x153 ^ 1'b0 ;
  assign n751 = n750 ^ n547 ^ 1'b0 ;
  assign n752 = x14 & ~n751 ;
  assign n753 = ~n651 & n752 ;
  assign n754 = n753 ^ n644 ^ 1'b0 ;
  assign n755 = x116 & ~n472 ;
  assign n756 = n755 ^ x43 ^ 1'b0 ;
  assign n757 = x245 ^ x198 ^ 1'b0 ;
  assign n758 = n757 ^ x128 ^ 1'b0 ;
  assign n759 = ~n756 & n758 ;
  assign n760 = x72 & x143 ;
  assign n761 = n760 ^ x114 ^ 1'b0 ;
  assign n762 = n375 | n761 ;
  assign n763 = n310 & ~n762 ;
  assign n764 = n759 & ~n763 ;
  assign n765 = x176 ^ x55 ^ 1'b0 ;
  assign n766 = x243 & n765 ;
  assign n767 = x242 & n766 ;
  assign n768 = n767 ^ n325 ^ 1'b0 ;
  assign n769 = n768 ^ n609 ^ x241 ;
  assign n770 = n297 | n398 ;
  assign n771 = n770 ^ x111 ^ 1'b0 ;
  assign n772 = n771 ^ x239 ^ 1'b0 ;
  assign n773 = n600 & n772 ;
  assign n774 = ( x93 & n501 ) | ( x93 & n773 ) | ( n501 & n773 ) ;
  assign n776 = x111 & x247 ;
  assign n777 = ~x126 & n776 ;
  assign n775 = ~n287 & n288 ;
  assign n778 = n777 ^ n775 ^ n538 ;
  assign n779 = x91 & n778 ;
  assign n780 = ~x251 & n779 ;
  assign n781 = x24 & x113 ;
  assign n782 = n527 & n781 ;
  assign n783 = ( n582 & n780 ) | ( n582 & n782 ) | ( n780 & n782 ) ;
  assign n786 = x30 & x244 ;
  assign n787 = n786 ^ n593 ^ 1'b0 ;
  assign n784 = n580 ^ n442 ^ 1'b0 ;
  assign n785 = x168 & n784 ;
  assign n788 = n787 ^ n785 ^ 1'b0 ;
  assign n789 = x9 & ~n788 ;
  assign n790 = n789 ^ x166 ^ 1'b0 ;
  assign n791 = n294 ^ x137 ^ 1'b0 ;
  assign n792 = x73 & n791 ;
  assign n793 = n792 ^ n354 ^ 1'b0 ;
  assign n794 = n435 & ~n793 ;
  assign n795 = n621 ^ x102 ^ x84 ;
  assign n796 = x153 & n402 ;
  assign n797 = n795 & n796 ;
  assign n798 = n615 ^ n571 ^ 1'b0 ;
  assign n799 = n424 | n798 ;
  assign n800 = n799 ^ n391 ^ 1'b0 ;
  assign n801 = ( ~x109 & n271 ) | ( ~x109 & n539 ) | ( n271 & n539 ) ;
  assign n802 = ~x104 & n801 ;
  assign n803 = n802 ^ n774 ^ 1'b0 ;
  assign n804 = n663 ^ n369 ^ x191 ;
  assign n805 = n660 ^ x22 ^ 1'b0 ;
  assign n806 = n805 ^ x158 ^ 1'b0 ;
  assign n807 = x248 ^ x20 ^ 1'b0 ;
  assign n808 = n807 ^ n735 ^ n307 ;
  assign n809 = x85 & ~n344 ;
  assign n810 = n334 | n444 ;
  assign n811 = ( ~n312 & n672 ) | ( ~n312 & n810 ) | ( n672 & n810 ) ;
  assign n812 = x126 & ~n362 ;
  assign n813 = n812 ^ n562 ^ 1'b0 ;
  assign n814 = ( x160 & ~n673 ) | ( x160 & n813 ) | ( ~n673 & n813 ) ;
  assign n815 = ( ~x84 & x149 ) | ( ~x84 & n358 ) | ( x149 & n358 ) ;
  assign n816 = n815 ^ n807 ^ x149 ;
  assign n817 = n386 | n816 ;
  assign n818 = n766 ^ n708 ^ n472 ;
  assign n819 = x57 & x188 ;
  assign n820 = ~x82 & n819 ;
  assign n821 = ( x209 & n818 ) | ( x209 & n820 ) | ( n818 & n820 ) ;
  assign n822 = n821 ^ n615 ^ 1'b0 ;
  assign n823 = ~n307 & n822 ;
  assign n824 = ( x1 & x50 ) | ( x1 & n343 ) | ( x50 & n343 ) ;
  assign n825 = n733 ^ n269 ^ x146 ;
  assign n826 = ( x39 & ~n824 ) | ( x39 & n825 ) | ( ~n824 & n825 ) ;
  assign n827 = n467 ^ n290 ^ x102 ;
  assign n828 = ( x14 & n356 ) | ( x14 & ~n827 ) | ( n356 & ~n827 ) ;
  assign n829 = n828 ^ n562 ^ x159 ;
  assign n830 = n829 ^ n678 ^ 1'b0 ;
  assign n831 = n826 | n830 ;
  assign n832 = n430 ^ x115 ^ x108 ;
  assign n833 = n401 | n826 ;
  assign n834 = n442 | n833 ;
  assign n835 = x28 & ~x60 ;
  assign n836 = n835 ^ x48 ^ 1'b0 ;
  assign n837 = n834 & ~n836 ;
  assign n838 = ( ~x11 & x61 ) | ( ~x11 & x154 ) | ( x61 & x154 ) ;
  assign n839 = n838 ^ n631 ^ x112 ;
  assign n840 = ~n837 & n839 ;
  assign n841 = ( x118 & x175 ) | ( x118 & n469 ) | ( x175 & n469 ) ;
  assign n842 = x234 ^ x42 ^ 1'b0 ;
  assign n843 = x229 & n842 ;
  assign n844 = n843 ^ n386 ^ x54 ;
  assign n845 = n844 ^ x100 ^ 1'b0 ;
  assign n846 = n428 & ~n476 ;
  assign n847 = n846 ^ n471 ^ 1'b0 ;
  assign n848 = n729 | n847 ;
  assign n849 = x105 & x158 ;
  assign n850 = ~x56 & n849 ;
  assign n851 = n733 ^ n625 ^ x206 ;
  assign n852 = n851 ^ n259 ^ x183 ;
  assign n853 = n852 ^ n519 ^ x29 ;
  assign n854 = n472 & n853 ;
  assign n855 = n507 | n854 ;
  assign n856 = n850 & ~n855 ;
  assign n857 = x102 & ~x171 ;
  assign n858 = x46 & n593 ;
  assign n859 = n858 ^ x194 ^ 1'b0 ;
  assign n860 = n859 ^ n672 ^ n567 ;
  assign n861 = ( x99 & x250 ) | ( x99 & n493 ) | ( x250 & n493 ) ;
  assign n862 = x35 & n292 ;
  assign n863 = n862 ^ x45 ^ 1'b0 ;
  assign n864 = ( ~x204 & n417 ) | ( ~x204 & n444 ) | ( n417 & n444 ) ;
  assign n867 = n273 | n490 ;
  assign n868 = n867 ^ x175 ^ 1'b0 ;
  assign n869 = n868 ^ x43 ^ 1'b0 ;
  assign n870 = x247 & n869 ;
  assign n871 = x222 & n407 ;
  assign n872 = ~n870 & n871 ;
  assign n865 = n539 ^ n474 ^ 1'b0 ;
  assign n866 = x10 & n865 ;
  assign n873 = n872 ^ n866 ^ 1'b0 ;
  assign n877 = ( x218 & ~n500 ) | ( x218 & n844 ) | ( ~n500 & n844 ) ;
  assign n874 = ( x96 & ~x220 ) | ( x96 & n300 ) | ( ~x220 & n300 ) ;
  assign n875 = n386 ^ x180 ^ 1'b0 ;
  assign n876 = n874 & n875 ;
  assign n878 = n877 ^ n876 ^ 1'b0 ;
  assign n879 = ( x110 & n403 ) | ( x110 & ~n878 ) | ( n403 & ~n878 ) ;
  assign n883 = n386 ^ x160 ^ 1'b0 ;
  assign n880 = x227 & ~n859 ;
  assign n881 = n880 ^ x194 ^ 1'b0 ;
  assign n882 = x176 & ~n881 ;
  assign n884 = n883 ^ n882 ^ 1'b0 ;
  assign n885 = ( n612 & ~n627 ) | ( n612 & n771 ) | ( ~n627 & n771 ) ;
  assign n886 = x185 & ~n519 ;
  assign n887 = n886 ^ n710 ^ 1'b0 ;
  assign n888 = ( x8 & x38 ) | ( x8 & ~n387 ) | ( x38 & ~n387 ) ;
  assign n889 = n888 ^ n509 ^ 1'b0 ;
  assign n890 = n344 & ~n889 ;
  assign n891 = n847 ^ n433 ^ x15 ;
  assign n892 = ( ~x149 & n459 ) | ( ~x149 & n483 ) | ( n459 & n483 ) ;
  assign n893 = n474 & ~n892 ;
  assign n894 = ~n352 & n893 ;
  assign n896 = x158 & ~n264 ;
  assign n897 = n896 ^ n511 ^ 1'b0 ;
  assign n898 = ( x60 & ~n425 ) | ( x60 & n897 ) | ( ~n425 & n897 ) ;
  assign n899 = x208 & ~n898 ;
  assign n900 = n899 ^ x8 ^ 1'b0 ;
  assign n895 = n468 & n704 ;
  assign n901 = n900 ^ n895 ^ n402 ;
  assign n902 = ~x20 & n659 ;
  assign n903 = x231 & n287 ;
  assign n904 = n903 ^ n326 ^ x24 ;
  assign n905 = n904 ^ n844 ^ x53 ;
  assign n907 = ( x172 & ~x193 ) | ( x172 & x207 ) | ( ~x193 & x207 ) ;
  assign n906 = ( x250 & n523 ) | ( x250 & n593 ) | ( n523 & n593 ) ;
  assign n908 = n907 ^ n906 ^ 1'b0 ;
  assign n909 = ~n256 & n908 ;
  assign n910 = x203 & ~n797 ;
  assign n911 = n910 ^ n423 ^ 1'b0 ;
  assign n912 = x249 & n341 ;
  assign n913 = n911 & n912 ;
  assign n914 = n841 ^ n832 ^ x186 ;
  assign n915 = n827 ^ n792 ^ n789 ;
  assign n916 = n490 | n915 ;
  assign n917 = n916 ^ n696 ^ 1'b0 ;
  assign n919 = x112 & x250 ;
  assign n920 = ~x216 & n919 ;
  assign n921 = n468 | n920 ;
  assign n918 = x146 & x247 ;
  assign n922 = n921 ^ n918 ^ 1'b0 ;
  assign n923 = x239 & ~n922 ;
  assign n924 = x127 & x134 ;
  assign n925 = ~x154 & n924 ;
  assign n926 = n405 | n925 ;
  assign n927 = n926 ^ n288 ^ x133 ;
  assign n928 = x215 ^ x13 ^ 1'b0 ;
  assign n929 = ( ~n308 & n709 ) | ( ~n308 & n928 ) | ( n709 & n928 ) ;
  assign n930 = n756 ^ n363 ^ 1'b0 ;
  assign n931 = n851 & ~n930 ;
  assign n934 = n733 ^ n363 ^ 1'b0 ;
  assign n935 = n544 | n934 ;
  assign n937 = n290 & ~n384 ;
  assign n938 = ~x9 & n937 ;
  assign n936 = ( ~x84 & x220 ) | ( ~x84 & x245 ) | ( x220 & x245 ) ;
  assign n939 = n938 ^ n936 ^ n358 ;
  assign n940 = n935 | n939 ;
  assign n941 = n500 | n940 ;
  assign n942 = x156 & n941 ;
  assign n943 = ~n805 & n942 ;
  assign n932 = ~x88 & n294 ;
  assign n933 = n932 ^ n870 ^ n270 ;
  assign n944 = n943 ^ n933 ^ x185 ;
  assign n945 = n269 ^ x227 ^ 1'b0 ;
  assign n953 = n658 ^ x157 ^ 1'b0 ;
  assign n954 = ~n293 & n953 ;
  assign n955 = n954 ^ n401 ^ 1'b0 ;
  assign n948 = x115 & x128 ;
  assign n949 = ~n360 & n948 ;
  assign n950 = n949 ^ n655 ^ x183 ;
  assign n946 = x32 & ~n615 ;
  assign n947 = ~n557 & n946 ;
  assign n951 = n950 ^ n947 ^ x166 ;
  assign n952 = n951 ^ n921 ^ x65 ;
  assign n956 = n955 ^ n952 ^ x27 ;
  assign n957 = x91 & n341 ;
  assign n958 = ( ~n652 & n820 ) | ( ~n652 & n945 ) | ( n820 & n945 ) ;
  assign n959 = ( ~n351 & n669 ) | ( ~n351 & n692 ) | ( n669 & n692 ) ;
  assign n960 = x64 ^ x50 ^ 1'b0 ;
  assign n961 = x113 & n960 ;
  assign n962 = n959 & ~n961 ;
  assign n963 = x203 & ~n303 ;
  assign n964 = ~x177 & n963 ;
  assign n965 = n303 | n964 ;
  assign n966 = x136 | n965 ;
  assign n967 = n415 ^ x154 ^ x34 ;
  assign n968 = n967 ^ x87 ^ 1'b0 ;
  assign n969 = x15 & n968 ;
  assign n970 = ~n966 & n969 ;
  assign n971 = n304 ^ x144 ^ 1'b0 ;
  assign n972 = ~n312 & n423 ;
  assign n973 = n316 & n972 ;
  assign n974 = n973 ^ n485 ^ x140 ;
  assign n975 = ~n561 & n974 ;
  assign n976 = ~n971 & n975 ;
  assign n977 = n444 & n851 ;
  assign n978 = ~x35 & n977 ;
  assign n979 = n729 & ~n978 ;
  assign n980 = ( x118 & n527 ) | ( x118 & n817 ) | ( n527 & n817 ) ;
  assign n981 = ( ~x29 & x108 ) | ( ~x29 & x152 ) | ( x108 & x152 ) ;
  assign n982 = n981 ^ n341 ^ 1'b0 ;
  assign n983 = n783 ^ x238 ^ 1'b0 ;
  assign n985 = n588 ^ x195 ^ 1'b0 ;
  assign n986 = ~n478 & n985 ;
  assign n987 = n639 ^ n338 ^ 1'b0 ;
  assign n988 = n528 & n987 ;
  assign n989 = ~n986 & n988 ;
  assign n984 = x98 & ~n476 ;
  assign n990 = n989 ^ n984 ^ 1'b0 ;
  assign n991 = n256 | n341 ;
  assign n992 = n713 ^ n305 ^ x139 ;
  assign n993 = n992 ^ x216 ^ x129 ;
  assign n996 = n669 ^ x65 ^ 1'b0 ;
  assign n997 = n953 & n996 ;
  assign n994 = n747 ^ n461 ^ n297 ;
  assign n995 = ~n287 & n994 ;
  assign n998 = n997 ^ n995 ^ 1'b0 ;
  assign n999 = n453 ^ x250 ^ 1'b0 ;
  assign n1000 = x41 & ~n999 ;
  assign n1001 = x182 & ~n349 ;
  assign n1002 = ~n266 & n1001 ;
  assign n1003 = n351 ^ x166 ^ 1'b0 ;
  assign n1004 = n1002 | n1003 ;
  assign n1005 = ( x162 & n560 ) | ( x162 & n1004 ) | ( n560 & n1004 ) ;
  assign n1006 = ( ~n998 & n1000 ) | ( ~n998 & n1005 ) | ( n1000 & n1005 ) ;
  assign n1007 = ( x34 & ~x172 ) | ( x34 & n447 ) | ( ~x172 & n447 ) ;
  assign n1008 = n883 & n1007 ;
  assign n1009 = n1008 ^ x16 ^ 1'b0 ;
  assign n1010 = n1009 ^ n986 ^ 1'b0 ;
  assign n1011 = x179 & n391 ;
  assign n1012 = ( x34 & ~x207 ) | ( x34 & n1011 ) | ( ~x207 & n1011 ) ;
  assign n1013 = ( x173 & n307 ) | ( x173 & n317 ) | ( n307 & n317 ) ;
  assign n1014 = n1013 ^ n825 ^ 1'b0 ;
  assign n1015 = ~n1012 & n1014 ;
  assign n1016 = ( ~x233 & x254 ) | ( ~x233 & n802 ) | ( x254 & n802 ) ;
  assign n1017 = ~n1005 & n1016 ;
  assign n1018 = n1017 ^ n432 ^ 1'b0 ;
  assign n1019 = n773 ^ n487 ^ x147 ;
  assign n1024 = x225 ^ x95 ^ x5 ;
  assign n1025 = ( x178 & ~x254 ) | ( x178 & n1024 ) | ( ~x254 & n1024 ) ;
  assign n1020 = n428 ^ n351 ^ 1'b0 ;
  assign n1021 = n268 | n1020 ;
  assign n1022 = n1021 ^ x142 ^ 1'b0 ;
  assign n1023 = n262 & ~n1022 ;
  assign n1026 = n1025 ^ n1023 ^ 1'b0 ;
  assign n1027 = n485 & n754 ;
  assign n1028 = n1027 ^ x45 ^ 1'b0 ;
  assign n1030 = n1023 ^ n651 ^ 1'b0 ;
  assign n1029 = x4 & x192 ;
  assign n1031 = n1030 ^ n1029 ^ 1'b0 ;
  assign n1033 = x34 & x237 ;
  assign n1034 = ~x59 & n1033 ;
  assign n1032 = ~x40 & x192 ;
  assign n1035 = n1034 ^ n1032 ^ x216 ;
  assign n1036 = n757 ^ n533 ^ 1'b0 ;
  assign n1037 = n967 | n1036 ;
  assign n1038 = n838 ^ n515 ^ 1'b0 ;
  assign n1039 = ( ~x121 & x246 ) | ( ~x121 & n831 ) | ( x246 & n831 ) ;
  assign n1044 = ~x131 & n537 ;
  assign n1045 = ( ~x34 & x61 ) | ( ~x34 & n1044 ) | ( x61 & n1044 ) ;
  assign n1046 = ( n270 & n307 ) | ( n270 & ~n1045 ) | ( n307 & ~n1045 ) ;
  assign n1040 = x111 & n697 ;
  assign n1041 = n981 ^ x225 ^ 1'b0 ;
  assign n1042 = n386 & ~n1041 ;
  assign n1043 = ( n981 & ~n1040 ) | ( n981 & n1042 ) | ( ~n1040 & n1042 ) ;
  assign n1047 = n1046 ^ n1043 ^ n890 ;
  assign n1048 = n606 ^ n290 ^ x141 ;
  assign n1049 = n1048 ^ n827 ^ 1'b0 ;
  assign n1050 = ~n894 & n1049 ;
  assign n1051 = x56 & n550 ;
  assign n1052 = n474 & ~n831 ;
  assign n1053 = n1052 ^ n503 ^ 1'b0 ;
  assign n1054 = ~n1026 & n1053 ;
  assign n1055 = n310 | n991 ;
  assign n1056 = x93 & ~n814 ;
  assign n1057 = n1056 ^ n411 ^ 1'b0 ;
  assign n1059 = n800 ^ n419 ^ 1'b0 ;
  assign n1060 = x117 & n1059 ;
  assign n1058 = ( ~x0 & x58 ) | ( ~x0 & n823 ) | ( x58 & n823 ) ;
  assign n1061 = n1060 ^ n1058 ^ 1'b0 ;
  assign n1066 = n432 ^ x77 ^ 1'b0 ;
  assign n1067 = x246 | n1066 ;
  assign n1062 = x237 ^ x132 ^ x123 ;
  assign n1063 = n1062 ^ n349 ^ x171 ;
  assign n1064 = x68 & x238 ;
  assign n1065 = ~n1063 & n1064 ;
  assign n1068 = n1067 ^ n1065 ^ 1'b0 ;
  assign n1069 = x93 ^ x49 ^ x11 ;
  assign n1070 = n1069 ^ n344 ^ 1'b0 ;
  assign n1071 = n1068 | n1070 ;
  assign n1072 = n1022 ^ n748 ^ 1'b0 ;
  assign n1073 = n556 & ~n1072 ;
  assign n1074 = x38 & x219 ;
  assign n1075 = n264 | n620 ;
  assign n1076 = n1075 ^ n503 ^ 1'b0 ;
  assign n1077 = ( n413 & n725 ) | ( n413 & ~n1028 ) | ( n725 & ~n1028 ) ;
  assign n1083 = ( x119 & n428 ) | ( x119 & ~n539 ) | ( n428 & ~n539 ) ;
  assign n1081 = n432 ^ n262 ^ x246 ;
  assign n1078 = x43 & n294 ;
  assign n1079 = ~n423 & n1078 ;
  assign n1080 = n1079 ^ x242 ^ x200 ;
  assign n1082 = n1081 ^ n1080 ^ x252 ;
  assign n1084 = n1083 ^ n1082 ^ n983 ;
  assign n1089 = x136 & ~n286 ;
  assign n1090 = n381 & n1089 ;
  assign n1085 = x227 & ~n967 ;
  assign n1086 = ~x252 & n1085 ;
  assign n1087 = x49 & n853 ;
  assign n1088 = n1086 & n1087 ;
  assign n1091 = n1090 ^ n1088 ^ 1'b0 ;
  assign n1092 = n655 ^ n440 ^ 1'b0 ;
  assign n1093 = x244 & ~n1092 ;
  assign n1094 = ( x253 & ~n514 ) | ( x253 & n1093 ) | ( ~n514 & n1093 ) ;
  assign n1095 = n845 & n1094 ;
  assign n1096 = n1091 & n1095 ;
  assign n1097 = n320 ^ x203 ^ 1'b0 ;
  assign n1098 = n339 & n1097 ;
  assign n1099 = x241 & n953 ;
  assign n1100 = ~x69 & n1099 ;
  assign n1101 = n675 ^ n485 ^ 1'b0 ;
  assign n1102 = x209 & ~n1101 ;
  assign n1103 = ~n515 & n1102 ;
  assign n1104 = n1103 ^ n1035 ^ n923 ;
  assign n1105 = n986 ^ x58 ^ 1'b0 ;
  assign n1106 = n625 ^ x201 ^ x39 ;
  assign n1107 = n764 & n810 ;
  assign n1108 = ~n1106 & n1107 ;
  assign n1109 = n1105 | n1108 ;
  assign n1110 = x167 | n1109 ;
  assign n1111 = x210 & n460 ;
  assign n1115 = n766 ^ x29 ^ x16 ;
  assign n1112 = x81 & x195 ;
  assign n1113 = ~x88 & n1112 ;
  assign n1114 = n582 & ~n1113 ;
  assign n1116 = n1115 ^ n1114 ^ 1'b0 ;
  assign n1117 = n931 ^ n816 ^ 1'b0 ;
  assign n1118 = n549 | n1117 ;
  assign n1119 = x243 ^ x127 ^ 1'b0 ;
  assign n1120 = ~n269 & n1119 ;
  assign n1121 = ~n1021 & n1120 ;
  assign n1122 = n1121 ^ x10 ^ 1'b0 ;
  assign n1123 = n1122 ^ n958 ^ n701 ;
  assign n1124 = x89 & ~x159 ;
  assign n1125 = x40 & x172 ;
  assign n1126 = n1125 ^ x37 ^ 1'b0 ;
  assign n1127 = x27 & n690 ;
  assign n1128 = ~n682 & n1127 ;
  assign n1130 = x39 & n941 ;
  assign n1131 = ~x36 & n1130 ;
  assign n1129 = ( x61 & ~x168 ) | ( x61 & n403 ) | ( ~x168 & n403 ) ;
  assign n1132 = n1131 ^ n1129 ^ 1'b0 ;
  assign n1135 = x83 & x180 ;
  assign n1136 = n307 & n1135 ;
  assign n1137 = n1136 ^ x26 ^ 1'b0 ;
  assign n1138 = n1012 | n1137 ;
  assign n1133 = ( n612 & n952 ) | ( n612 & n1025 ) | ( n952 & n1025 ) ;
  assign n1134 = n1133 ^ n738 ^ 1'b0 ;
  assign n1139 = n1138 ^ n1134 ^ 1'b0 ;
  assign n1140 = n1132 & ~n1139 ;
  assign n1141 = ( n627 & n1128 ) | ( n627 & n1140 ) | ( n1128 & n1140 ) ;
  assign n1142 = ( ~n356 & n1126 ) | ( ~n356 & n1141 ) | ( n1126 & n1141 ) ;
  assign n1143 = n1124 | n1142 ;
  assign n1144 = n620 & ~n1143 ;
  assign n1145 = ~x24 & n457 ;
  assign n1147 = n295 & n462 ;
  assign n1148 = n1147 ^ x235 ^ 1'b0 ;
  assign n1146 = x151 & n768 ;
  assign n1149 = n1148 ^ n1146 ^ 1'b0 ;
  assign n1150 = ( n489 & n1021 ) | ( n489 & n1149 ) | ( n1021 & n1149 ) ;
  assign n1151 = x241 ^ x68 ^ x59 ;
  assign n1152 = n750 & ~n1151 ;
  assign n1153 = n326 | n1129 ;
  assign n1154 = n385 | n1153 ;
  assign n1158 = n415 & ~n973 ;
  assign n1159 = n1158 ^ x105 ^ 1'b0 ;
  assign n1160 = x158 & n1159 ;
  assign n1161 = ~x195 & n1160 ;
  assign n1155 = n511 ^ n459 ^ x198 ;
  assign n1156 = n1155 ^ x183 ^ x74 ;
  assign n1157 = n709 & ~n1156 ;
  assign n1162 = n1161 ^ n1157 ^ 1'b0 ;
  assign n1163 = n800 | n1066 ;
  assign n1164 = n560 & ~n1163 ;
  assign n1165 = n897 ^ n264 ^ 1'b0 ;
  assign n1166 = ~n684 & n1165 ;
  assign n1167 = n804 ^ n444 ^ 1'b0 ;
  assign n1168 = n362 | n1167 ;
  assign n1169 = n1166 & ~n1168 ;
  assign n1170 = n1164 & n1169 ;
  assign n1171 = x119 & ~n850 ;
  assign n1172 = ~x126 & n1171 ;
  assign n1173 = ( x58 & ~x207 ) | ( x58 & n300 ) | ( ~x207 & n300 ) ;
  assign n1174 = ~n256 & n1173 ;
  assign n1175 = n595 & n1174 ;
  assign n1176 = ( x232 & n1172 ) | ( x232 & ~n1175 ) | ( n1172 & ~n1175 ) ;
  assign n1177 = n950 ^ x58 ^ 1'b0 ;
  assign n1178 = n462 & n1177 ;
  assign n1179 = ( x205 & n263 ) | ( x205 & n859 ) | ( n263 & n859 ) ;
  assign n1180 = x133 & n1179 ;
  assign n1181 = n612 & n1180 ;
  assign n1182 = n1178 & ~n1181 ;
  assign n1183 = ~n479 & n582 ;
  assign n1184 = n1182 & n1183 ;
  assign n1185 = n1184 ^ n813 ^ 1'b0 ;
  assign n1188 = x99 & x228 ;
  assign n1189 = n273 & n1188 ;
  assign n1186 = n1175 ^ n335 ^ 1'b0 ;
  assign n1187 = x127 & ~n1186 ;
  assign n1190 = n1189 ^ n1187 ^ n735 ;
  assign n1191 = x186 & n298 ;
  assign n1192 = ~x254 & n1191 ;
  assign n1193 = n642 | n1192 ;
  assign n1194 = n774 | n1193 ;
  assign n1195 = n976 ^ n787 ^ 1'b0 ;
  assign n1196 = ~n861 & n1195 ;
  assign n1197 = n387 ^ x21 ^ 1'b0 ;
  assign n1198 = n474 ^ x8 ^ 1'b0 ;
  assign n1199 = x34 & n1198 ;
  assign n1200 = ( ~n366 & n1197 ) | ( ~n366 & n1199 ) | ( n1197 & n1199 ) ;
  assign n1201 = x58 & x251 ;
  assign n1202 = ( x37 & ~x186 ) | ( x37 & n447 ) | ( ~x186 & n447 ) ;
  assign n1203 = x156 | n684 ;
  assign n1204 = n451 ^ n401 ^ 1'b0 ;
  assign n1205 = ( n1202 & n1203 ) | ( n1202 & n1204 ) | ( n1203 & n1204 ) ;
  assign n1206 = n600 ^ n378 ^ x159 ;
  assign n1207 = n1206 ^ n803 ^ 1'b0 ;
  assign n1208 = n906 & n1207 ;
  assign n1209 = ~n485 & n1208 ;
  assign n1210 = x24 & ~n1209 ;
  assign n1211 = n1210 ^ n344 ^ 1'b0 ;
  assign n1212 = n907 ^ x89 ^ 1'b0 ;
  assign n1213 = n436 & n1212 ;
  assign n1214 = ~n496 & n1213 ;
  assign n1215 = x38 & ~n1214 ;
  assign n1216 = n1004 & n1215 ;
  assign n1217 = n1216 ^ n1022 ^ n597 ;
  assign n1218 = n604 ^ n586 ^ 1'b0 ;
  assign n1219 = n1172 | n1218 ;
  assign n1220 = x223 ^ x88 ^ x84 ;
  assign n1221 = n1220 ^ x224 ^ 1'b0 ;
  assign n1222 = n560 | n1221 ;
  assign n1223 = x62 & ~n1222 ;
  assign n1224 = n1223 ^ n527 ^ 1'b0 ;
  assign n1225 = n990 ^ n608 ^ x83 ;
  assign n1228 = n861 ^ n394 ^ x251 ;
  assign n1229 = ( n270 & n575 ) | ( n270 & ~n1228 ) | ( n575 & ~n1228 ) ;
  assign n1230 = n716 & ~n1229 ;
  assign n1231 = ~x69 & n1230 ;
  assign n1226 = ( ~x181 & n323 ) | ( ~x181 & n947 ) | ( n323 & n947 ) ;
  assign n1227 = n1226 ^ x5 ^ 1'b0 ;
  assign n1232 = n1231 ^ n1227 ^ n1068 ;
  assign n1233 = n561 | n1086 ;
  assign n1234 = n496 | n1233 ;
  assign n1235 = ~n817 & n961 ;
  assign n1236 = ~n1234 & n1235 ;
  assign n1237 = n763 ^ n642 ^ 1'b0 ;
  assign n1238 = n1237 ^ n803 ^ 1'b0 ;
  assign n1239 = n951 & n1238 ;
  assign n1240 = n902 ^ n659 ^ 1'b0 ;
  assign n1243 = n990 & ~n1032 ;
  assign n1241 = ( n275 & n474 ) | ( n275 & n710 ) | ( n474 & n710 ) ;
  assign n1242 = ~n1022 & n1241 ;
  assign n1244 = n1243 ^ n1242 ^ 1'b0 ;
  assign n1245 = n333 | n878 ;
  assign n1246 = n1245 ^ x130 ^ 1'b0 ;
  assign n1247 = ( x142 & n599 ) | ( x142 & n1151 ) | ( n599 & n1151 ) ;
  assign n1248 = n440 | n1247 ;
  assign n1249 = n837 ^ x216 ^ 1'b0 ;
  assign n1250 = ( x228 & n574 ) | ( x228 & ~n1249 ) | ( n574 & ~n1249 ) ;
  assign n1251 = n1079 ^ n938 ^ x224 ;
  assign n1252 = ( ~n347 & n481 ) | ( ~n347 & n667 ) | ( n481 & n667 ) ;
  assign n1253 = ( x102 & n365 ) | ( x102 & n608 ) | ( n365 & n608 ) ;
  assign n1254 = ( n270 & n1252 ) | ( n270 & n1253 ) | ( n1252 & n1253 ) ;
  assign n1255 = n490 | n1254 ;
  assign n1256 = n1251 & ~n1255 ;
  assign n1257 = n1151 ^ n580 ^ n432 ;
  assign n1258 = n384 & ~n1257 ;
  assign n1259 = ~n1256 & n1258 ;
  assign n1260 = n1259 ^ n964 ^ 1'b0 ;
  assign n1261 = n562 ^ n343 ^ x50 ;
  assign n1262 = ( ~n853 & n877 ) | ( ~n853 & n1261 ) | ( n877 & n1261 ) ;
  assign n1263 = n1262 ^ n649 ^ 1'b0 ;
  assign n1264 = x141 & ~n1263 ;
  assign n1265 = n1264 ^ n961 ^ n606 ;
  assign n1266 = n316 | n824 ;
  assign n1267 = n1266 ^ n1185 ^ n841 ;
  assign n1268 = x206 ^ x49 ^ 1'b0 ;
  assign n1269 = x136 & n1268 ;
  assign n1270 = ( x120 & ~n495 ) | ( x120 & n1269 ) | ( ~n495 & n1269 ) ;
  assign n1271 = n389 ^ x134 ^ x8 ;
  assign n1272 = n1271 ^ x74 ^ x52 ;
  assign n1273 = n1022 & ~n1272 ;
  assign n1274 = x245 & n1273 ;
  assign n1284 = n279 & ~n667 ;
  assign n1281 = n684 ^ n460 ^ n350 ;
  assign n1279 = n1106 ^ x97 ^ 1'b0 ;
  assign n1280 = n290 & ~n1279 ;
  assign n1282 = n1281 ^ n1280 ^ 1'b0 ;
  assign n1283 = n1134 & n1282 ;
  assign n1275 = n275 ^ x48 ^ 1'b0 ;
  assign n1276 = n702 & n870 ;
  assign n1277 = n1275 & n1276 ;
  assign n1278 = ~n1041 & n1277 ;
  assign n1285 = n1284 ^ n1283 ^ n1278 ;
  assign n1286 = ( n460 & n1274 ) | ( n460 & ~n1285 ) | ( n1274 & ~n1285 ) ;
  assign n1287 = n344 & n827 ;
  assign n1288 = ~n266 & n1287 ;
  assign n1289 = n1288 ^ n782 ^ x106 ;
  assign n1290 = n1289 ^ n1024 ^ x213 ;
  assign n1291 = n1290 ^ n1226 ^ n923 ;
  assign n1292 = ~n795 & n1211 ;
  assign n1293 = x57 ^ x39 ^ 1'b0 ;
  assign n1294 = x131 & n1293 ;
  assign n1295 = n352 & n1294 ;
  assign n1296 = n1295 ^ n1289 ^ n1115 ;
  assign n1297 = n535 | n920 ;
  assign n1298 = n1296 & ~n1297 ;
  assign n1299 = n262 | n994 ;
  assign n1300 = n1299 ^ n1189 ^ n790 ;
  assign n1301 = n1299 ^ n660 ^ 1'b0 ;
  assign n1303 = n381 ^ x196 ^ 1'b0 ;
  assign n1304 = n287 | n1303 ;
  assign n1305 = n752 & ~n847 ;
  assign n1306 = n1304 & n1305 ;
  assign n1302 = x149 & ~n1002 ;
  assign n1307 = n1306 ^ n1302 ^ n1227 ;
  assign n1308 = ( x73 & ~x226 ) | ( x73 & n516 ) | ( ~x226 & n516 ) ;
  assign n1309 = ( x200 & n939 ) | ( x200 & n1128 ) | ( n939 & n1128 ) ;
  assign n1310 = n718 ^ n275 ^ 1'b0 ;
  assign n1311 = n1310 ^ n876 ^ 1'b0 ;
  assign n1312 = ~n1309 & n1311 ;
  assign n1313 = x78 & x184 ;
  assign n1314 = ~n393 & n1313 ;
  assign n1315 = n374 ^ n280 ^ 1'b0 ;
  assign n1316 = n1314 | n1315 ;
  assign n1317 = n1316 ^ n1077 ^ 1'b0 ;
  assign n1318 = n1312 & ~n1317 ;
  assign n1320 = n535 ^ x57 ^ 1'b0 ;
  assign n1319 = ( x47 & n554 ) | ( x47 & n952 ) | ( n554 & n952 ) ;
  assign n1321 = n1320 ^ n1319 ^ n859 ;
  assign n1322 = x13 & ~n562 ;
  assign n1323 = n1322 ^ n600 ^ 1'b0 ;
  assign n1324 = ~x245 & n778 ;
  assign n1325 = n1323 | n1324 ;
  assign n1326 = n1325 ^ n610 ^ n606 ;
  assign n1327 = n500 ^ n433 ^ 1'b0 ;
  assign n1328 = x143 & n741 ;
  assign n1329 = ( x107 & x111 ) | ( x107 & n1328 ) | ( x111 & n1328 ) ;
  assign n1330 = ~n333 & n851 ;
  assign n1331 = ~x236 & n1330 ;
  assign n1332 = n803 | n1331 ;
  assign n1333 = x251 & ~n813 ;
  assign n1334 = n1333 ^ x162 ^ 1'b0 ;
  assign n1335 = n1334 ^ n1048 ^ 1'b0 ;
  assign n1336 = n1024 ^ x163 ^ x55 ;
  assign n1337 = n1336 ^ x176 ^ 1'b0 ;
  assign n1338 = x24 & x97 ;
  assign n1339 = n1189 & n1338 ;
  assign n1340 = n1131 ^ n857 ^ 1'b0 ;
  assign n1341 = ~n826 & n1340 ;
  assign n1342 = ~n1339 & n1341 ;
  assign n1343 = n1342 ^ n1181 ^ 1'b0 ;
  assign n1344 = ~n282 & n460 ;
  assign n1345 = n817 & n1344 ;
  assign n1346 = ~n552 & n1308 ;
  assign n1347 = n1346 ^ x118 ^ 1'b0 ;
  assign n1348 = x247 & ~n1088 ;
  assign n1349 = n1348 ^ n1086 ^ 1'b0 ;
  assign n1350 = ( x32 & ~x173 ) | ( x32 & n1229 ) | ( ~x173 & n1229 ) ;
  assign n1351 = ( ~x63 & x126 ) | ( ~x63 & x157 ) | ( x126 & x157 ) ;
  assign n1352 = n1351 ^ n656 ^ 1'b0 ;
  assign n1353 = ( ~x9 & x112 ) | ( ~x9 & n441 ) | ( x112 & n441 ) ;
  assign n1354 = x148 | n421 ;
  assign n1355 = ~n1353 & n1354 ;
  assign n1356 = n1355 ^ n557 ^ 1'b0 ;
  assign n1357 = ( ~x23 & n1352 ) | ( ~x23 & n1356 ) | ( n1352 & n1356 ) ;
  assign n1358 = n1220 ^ n704 ^ 1'b0 ;
  assign n1359 = n1226 | n1358 ;
  assign n1360 = n944 | n1359 ;
  assign n1361 = n710 ^ n403 ^ 1'b0 ;
  assign n1362 = n600 & ~n1361 ;
  assign n1363 = n1362 ^ x135 ^ 1'b0 ;
  assign n1364 = n947 ^ n490 ^ 1'b0 ;
  assign n1365 = x218 ^ x122 ^ x35 ;
  assign n1366 = x190 | n1365 ;
  assign n1367 = n459 & n1284 ;
  assign n1368 = n1367 ^ n1090 ^ n1022 ;
  assign n1369 = n286 & n1368 ;
  assign n1370 = ( n1332 & ~n1366 ) | ( n1332 & n1369 ) | ( ~n1366 & n1369 ) ;
  assign n1371 = n1370 ^ n300 ^ 1'b0 ;
  assign n1372 = n277 | n1371 ;
  assign n1374 = ~n559 & n1024 ;
  assign n1375 = n630 | n1374 ;
  assign n1376 = n454 | n1375 ;
  assign n1373 = ~n944 & n952 ;
  assign n1377 = n1376 ^ n1373 ^ 1'b0 ;
  assign n1378 = n1220 ^ x157 ^ x101 ;
  assign n1379 = ( x239 & ~n487 ) | ( x239 & n974 ) | ( ~n487 & n974 ) ;
  assign n1380 = x146 & n1105 ;
  assign n1381 = n1379 & ~n1380 ;
  assign n1382 = ~x109 & n1381 ;
  assign n1383 = n824 | n911 ;
  assign n1384 = ~n1382 & n1383 ;
  assign n1385 = ~n1247 & n1384 ;
  assign n1386 = ( x98 & n1035 ) | ( x98 & n1248 ) | ( n1035 & n1248 ) ;
  assign n1387 = n668 | n1040 ;
  assign n1388 = n978 ^ x134 ^ 1'b0 ;
  assign n1389 = n1388 ^ n1252 ^ 1'b0 ;
  assign n1390 = n1389 ^ n915 ^ 1'b0 ;
  assign n1391 = n496 & n547 ;
  assign n1392 = ~n1390 & n1391 ;
  assign n1393 = n1392 ^ x81 ^ x11 ;
  assign n1394 = n389 | n1393 ;
  assign n1395 = ( x55 & ~x135 ) | ( x55 & n686 ) | ( ~x135 & n686 ) ;
  assign n1396 = n1395 ^ n1012 ^ 1'b0 ;
  assign n1397 = x76 & n1396 ;
  assign n1398 = n1397 ^ n914 ^ 1'b0 ;
  assign n1399 = n303 & n654 ;
  assign n1400 = n1398 & n1399 ;
  assign n1401 = n550 & n1400 ;
  assign n1402 = n1295 ^ n911 ^ x204 ;
  assign n1403 = n906 ^ n876 ^ 1'b0 ;
  assign n1404 = n1294 ^ n509 ^ 1'b0 ;
  assign n1405 = x121 & ~n1404 ;
  assign n1406 = ( ~x34 & x196 ) | ( ~x34 & n499 ) | ( x196 & n499 ) ;
  assign n1407 = ~n733 & n1406 ;
  assign n1408 = n1407 ^ x241 ^ 1'b0 ;
  assign n1409 = n1405 & n1408 ;
  assign n1410 = x137 | n325 ;
  assign n1411 = n964 ^ n609 ^ 1'b0 ;
  assign n1412 = ~n343 & n1411 ;
  assign n1413 = n1412 ^ n522 ^ 1'b0 ;
  assign n1414 = n1281 & n1413 ;
  assign n1415 = n1410 & n1414 ;
  assign n1416 = x7 & ~n314 ;
  assign n1417 = x180 & x246 ;
  assign n1418 = n1417 ^ n493 ^ 1'b0 ;
  assign n1419 = n931 & n1418 ;
  assign n1420 = ~x45 & n1419 ;
  assign n1421 = n715 ^ x194 ^ 1'b0 ;
  assign n1422 = x35 & n1421 ;
  assign n1423 = n1422 ^ n694 ^ n660 ;
  assign n1424 = n680 & n1423 ;
  assign n1425 = x245 & ~n573 ;
  assign n1426 = n327 & ~n1275 ;
  assign n1427 = n1425 & n1426 ;
  assign n1428 = n717 & ~n1427 ;
  assign n1429 = ~n764 & n1428 ;
  assign n1430 = ~x67 & n1179 ;
  assign n1431 = n1422 ^ n441 ^ 1'b0 ;
  assign n1432 = x104 & ~n1431 ;
  assign n1433 = ( n482 & ~n1304 ) | ( n482 & n1432 ) | ( ~n1304 & n1432 ) ;
  assign n1434 = n1270 & ~n1433 ;
  assign n1438 = x88 ^ x78 ^ 1'b0 ;
  assign n1439 = ( x51 & ~n478 ) | ( x51 & n1438 ) | ( ~n478 & n1438 ) ;
  assign n1440 = ~x56 & n1439 ;
  assign n1437 = n1108 | n1214 ;
  assign n1441 = n1440 ^ n1437 ^ 1'b0 ;
  assign n1435 = n1019 ^ n951 ^ 1'b0 ;
  assign n1436 = n750 | n1435 ;
  assign n1442 = n1441 ^ n1436 ^ 1'b0 ;
  assign n1443 = n638 | n958 ;
  assign n1444 = n1443 ^ x183 ^ 1'b0 ;
  assign n1445 = x194 & x229 ;
  assign n1446 = n1445 ^ x174 ^ 1'b0 ;
  assign n1447 = n782 | n1446 ;
  assign n1452 = ( x146 & n708 ) | ( x146 & n920 ) | ( n708 & n920 ) ;
  assign n1448 = ( ~x143 & x194 ) | ( ~x143 & n1004 ) | ( x194 & n1004 ) ;
  assign n1449 = x100 & ~n1448 ;
  assign n1450 = n1449 ^ x207 ^ 1'b0 ;
  assign n1451 = n1450 ^ n1034 ^ 1'b0 ;
  assign n1453 = n1452 ^ n1451 ^ n806 ;
  assign n1454 = ( ~x144 & x154 ) | ( ~x144 & n1390 ) | ( x154 & n1390 ) ;
  assign n1460 = n499 & ~n1228 ;
  assign n1455 = n615 ^ x172 ^ x110 ;
  assign n1456 = n1455 ^ n642 ^ 1'b0 ;
  assign n1457 = n322 | n1456 ;
  assign n1458 = n1457 ^ n1366 ^ x10 ;
  assign n1459 = x218 & n1458 ;
  assign n1461 = n1460 ^ n1459 ^ 1'b0 ;
  assign n1462 = ~n381 & n1461 ;
  assign n1463 = n1462 ^ x154 ^ 1'b0 ;
  assign n1464 = n391 ^ x51 ^ 1'b0 ;
  assign n1465 = n440 | n1464 ;
  assign n1466 = n356 & ~n1465 ;
  assign n1467 = n1466 ^ n287 ^ 1'b0 ;
  assign n1468 = n1335 ^ x227 ^ x30 ;
  assign n1469 = ~n1434 & n1468 ;
  assign n1470 = n1467 & n1469 ;
  assign n1471 = n1395 ^ n623 ^ 1'b0 ;
  assign n1472 = n997 & n1471 ;
  assign n1473 = n945 ^ x18 ^ 1'b0 ;
  assign n1474 = n1472 & n1473 ;
  assign n1475 = n351 | n1418 ;
  assign n1476 = ( n616 & n1474 ) | ( n616 & n1475 ) | ( n1474 & n1475 ) ;
  assign n1477 = x251 & ~n672 ;
  assign n1478 = n1477 ^ n1314 ^ 1'b0 ;
  assign n1479 = ( ~x139 & n562 ) | ( ~x139 & n824 ) | ( n562 & n824 ) ;
  assign n1480 = n282 & ~n1126 ;
  assign n1481 = ( n1032 & ~n1479 ) | ( n1032 & n1480 ) | ( ~n1479 & n1480 ) ;
  assign n1482 = ~x146 & n394 ;
  assign n1483 = n363 & ~n835 ;
  assign n1484 = n1483 ^ n1022 ^ 1'b0 ;
  assign n1485 = x247 & n1484 ;
  assign n1486 = n1485 ^ n438 ^ 1'b0 ;
  assign n1487 = ~n297 & n978 ;
  assign n1488 = n335 | n1487 ;
  assign n1489 = n1488 ^ n878 ^ 1'b0 ;
  assign n1491 = n378 | n515 ;
  assign n1492 = n1491 ^ n615 ^ 1'b0 ;
  assign n1490 = x76 & n1175 ;
  assign n1493 = n1492 ^ n1490 ^ 1'b0 ;
  assign n1494 = n841 ^ n747 ^ 1'b0 ;
  assign n1495 = n935 ^ x237 ^ 1'b0 ;
  assign n1496 = ( x141 & x251 ) | ( x141 & ~n1495 ) | ( x251 & ~n1495 ) ;
  assign n1499 = ( x196 & ~n976 ) | ( x196 & n1251 ) | ( ~n976 & n1251 ) ;
  assign n1497 = n1007 ^ x48 ^ x14 ;
  assign n1498 = n288 | n1497 ;
  assign n1500 = n1499 ^ n1498 ^ 1'b0 ;
  assign n1501 = n1500 ^ n462 ^ 1'b0 ;
  assign n1502 = n1496 & ~n1501 ;
  assign n1503 = ~n1444 & n1502 ;
  assign n1504 = n292 ^ x198 ^ 1'b0 ;
  assign n1505 = n584 & ~n1504 ;
  assign n1506 = n487 ^ x203 ^ x106 ;
  assign n1507 = n1372 | n1506 ;
  assign n1508 = x46 | n1507 ;
  assign n1509 = n1141 & n1295 ;
  assign n1510 = n1509 ^ n286 ^ 1'b0 ;
  assign n1511 = n507 ^ x125 ^ 1'b0 ;
  assign n1512 = n552 | n1511 ;
  assign n1513 = n757 & n1512 ;
  assign n1514 = n825 & n1513 ;
  assign n1515 = n1514 ^ n909 ^ n436 ;
  assign n1516 = n1515 ^ n713 ^ n394 ;
  assign n1517 = n1239 & n1275 ;
  assign n1518 = n1508 & n1517 ;
  assign n1519 = n1518 ^ n1031 ^ 1'b0 ;
  assign n1520 = n385 & ~n1136 ;
  assign n1521 = ~x27 & n1520 ;
  assign n1522 = n1521 ^ n763 ^ 1'b0 ;
  assign n1523 = n838 ^ x37 ^ 1'b0 ;
  assign n1524 = n1523 ^ n1175 ^ x63 ;
  assign n1525 = n511 ^ n479 ^ 1'b0 ;
  assign n1526 = x242 & n621 ;
  assign n1527 = n1526 ^ n768 ^ 1'b0 ;
  assign n1528 = n872 | n1527 ;
  assign n1529 = x167 | n1528 ;
  assign n1530 = ( x212 & n920 ) | ( x212 & ~n1050 ) | ( n920 & ~n1050 ) ;
  assign n1531 = n1530 ^ n1094 ^ 1'b0 ;
  assign n1532 = n857 | n1531 ;
  assign n1536 = n394 ^ x84 ^ 1'b0 ;
  assign n1537 = n464 & n1536 ;
  assign n1533 = ( n423 & n1192 ) | ( n423 & ~n1299 ) | ( n1192 & ~n1299 ) ;
  assign n1534 = n287 & ~n1533 ;
  assign n1535 = n426 | n1534 ;
  assign n1538 = n1537 ^ n1535 ^ 1'b0 ;
  assign n1539 = n630 | n949 ;
  assign n1540 = x241 | n1539 ;
  assign n1541 = x169 & ~n1199 ;
  assign n1542 = ( n471 & n808 ) | ( n471 & n1541 ) | ( n808 & n1541 ) ;
  assign n1543 = x51 & ~n450 ;
  assign n1544 = x126 & n337 ;
  assign n1545 = n1544 ^ n677 ^ 1'b0 ;
  assign n1546 = n295 ^ x238 ^ 1'b0 ;
  assign n1547 = x43 & n1546 ;
  assign n1548 = ( n599 & n1406 ) | ( n599 & ~n1547 ) | ( n1406 & ~n1547 ) ;
  assign n1549 = n385 & ~n1548 ;
  assign n1550 = ( ~n445 & n1028 ) | ( ~n445 & n1549 ) | ( n1028 & n1549 ) ;
  assign n1551 = n1550 ^ n981 ^ 1'b0 ;
  assign n1552 = ~n1545 & n1551 ;
  assign n1553 = n1322 ^ n1275 ^ 1'b0 ;
  assign n1554 = n735 & ~n1553 ;
  assign n1555 = n300 & ~n1018 ;
  assign n1556 = ~n840 & n866 ;
  assign n1557 = ~x133 & n1556 ;
  assign n1558 = n1115 ^ n959 ^ n619 ;
  assign n1559 = n1558 ^ n890 ^ 1'b0 ;
  assign n1560 = n362 | n1090 ;
  assign n1561 = x89 | n1560 ;
  assign n1562 = n1561 ^ n1479 ^ n1247 ;
  assign n1563 = n971 & ~n1562 ;
  assign n1564 = n425 & n1302 ;
  assign n1565 = n1460 ^ x68 ^ 1'b0 ;
  assign n1566 = ~n623 & n1565 ;
  assign n1567 = n1511 ^ n438 ^ x101 ;
  assign n1568 = n1567 ^ x82 ^ 1'b0 ;
  assign n1569 = n1566 & n1568 ;
  assign n1570 = ( n761 & ~n771 ) | ( n761 & n792 ) | ( ~n771 & n792 ) ;
  assign n1571 = n955 ^ n825 ^ x10 ;
  assign n1572 = ( x26 & n970 ) | ( x26 & ~n1450 ) | ( n970 & ~n1450 ) ;
  assign n1573 = n1571 & ~n1572 ;
  assign n1574 = ( n1448 & n1561 ) | ( n1448 & n1573 ) | ( n1561 & n1573 ) ;
  assign n1575 = x135 & n931 ;
  assign n1576 = n1575 ^ n677 ^ 1'b0 ;
  assign n1577 = n913 ^ n505 ^ 1'b0 ;
  assign n1578 = n1576 | n1577 ;
  assign n1579 = n876 ^ n665 ^ x10 ;
  assign n1580 = n1579 ^ n813 ^ x225 ;
  assign n1581 = ~n1321 & n1580 ;
  assign n1582 = n1581 ^ x223 ^ 1'b0 ;
  assign n1583 = ( x4 & n783 ) | ( x4 & ~n802 ) | ( n783 & ~n802 ) ;
  assign n1584 = n1093 ^ n787 ^ x118 ;
  assign n1585 = x20 & ~n1584 ;
  assign n1586 = x82 & ~x168 ;
  assign n1587 = n317 | n1586 ;
  assign n1588 = n1587 ^ n1071 ^ 1'b0 ;
  assign n1589 = n1320 | n1588 ;
  assign n1590 = n704 | n1589 ;
  assign n1591 = x127 & n1590 ;
  assign n1592 = n501 & n1591 ;
  assign n1593 = x36 | n401 ;
  assign n1594 = n320 ^ x67 ^ 1'b0 ;
  assign n1595 = n1593 | n1594 ;
  assign n1596 = n768 ^ x220 ^ x75 ;
  assign n1597 = ( ~n894 & n902 ) | ( ~n894 & n1596 ) | ( n902 & n1596 ) ;
  assign n1598 = n467 & ~n1335 ;
  assign n1599 = ~n928 & n1302 ;
  assign n1600 = ~n953 & n1599 ;
  assign n1603 = n668 ^ x5 ^ 1'b0 ;
  assign n1604 = ( ~n549 & n1383 ) | ( ~n549 & n1603 ) | ( n1383 & n1603 ) ;
  assign n1601 = n503 ^ x200 ^ 1'b0 ;
  assign n1602 = n597 | n1601 ;
  assign n1605 = n1604 ^ n1602 ^ 1'b0 ;
  assign n1606 = n1605 ^ n1382 ^ x254 ;
  assign n1607 = ~x189 & n531 ;
  assign n1608 = x106 & ~n1334 ;
  assign n1609 = n1607 & n1608 ;
  assign n1610 = ~n262 & n415 ;
  assign n1611 = n1610 ^ n637 ^ 1'b0 ;
  assign n1612 = x190 & ~n1611 ;
  assign n1613 = n1612 ^ n469 ^ 1'b0 ;
  assign n1614 = x211 & n1271 ;
  assign n1615 = n1172 & n1614 ;
  assign n1616 = ( n843 & ~n1613 ) | ( n843 & n1615 ) | ( ~n1613 & n1615 ) ;
  assign n1617 = n1616 ^ n1271 ^ n944 ;
  assign n1618 = n1172 | n1617 ;
  assign n1619 = n654 & ~n1332 ;
  assign n1620 = n1619 ^ n1252 ^ 1'b0 ;
  assign n1621 = n1359 ^ x4 ^ 1'b0 ;
  assign n1622 = n1511 & ~n1621 ;
  assign n1623 = ~n1427 & n1622 ;
  assign n1624 = n750 & n1623 ;
  assign n1625 = n638 | n1290 ;
  assign n1626 = n1244 & ~n1625 ;
  assign n1627 = n1626 ^ n600 ^ 1'b0 ;
  assign n1628 = n1352 & ~n1627 ;
  assign n1629 = n860 ^ n513 ^ n441 ;
  assign n1630 = n567 & n1629 ;
  assign n1634 = n675 ^ x109 ^ x9 ;
  assign n1635 = n1634 ^ n1069 ^ n335 ;
  assign n1631 = n537 & ~n1288 ;
  assign n1632 = n1323 & n1631 ;
  assign n1633 = x131 | n1632 ;
  assign n1636 = n1635 ^ n1633 ^ n550 ;
  assign n1637 = ( n1103 & n1266 ) | ( n1103 & n1636 ) | ( n1266 & n1636 ) ;
  assign n1638 = ( n454 & n599 ) | ( n454 & n897 ) | ( n599 & n897 ) ;
  assign n1652 = ~n596 & n673 ;
  assign n1653 = ~n1098 & n1652 ;
  assign n1646 = x197 ^ x168 ^ 1'b0 ;
  assign n1647 = ~n316 & n1646 ;
  assign n1648 = x236 & x242 ;
  assign n1649 = n1648 ^ x73 ^ 1'b0 ;
  assign n1650 = n1647 & n1649 ;
  assign n1643 = ~x13 & x31 ;
  assign n1639 = ( ~x48 & x61 ) | ( ~x48 & x92 ) | ( x61 & x92 ) ;
  assign n1640 = n403 & n1639 ;
  assign n1641 = n1561 ^ n580 ^ 1'b0 ;
  assign n1642 = ~n1640 & n1641 ;
  assign n1644 = n1643 ^ n1642 ^ 1'b0 ;
  assign n1645 = n794 & n1644 ;
  assign n1651 = n1650 ^ n1645 ^ 1'b0 ;
  assign n1654 = n1653 ^ n1651 ^ 1'b0 ;
  assign n1655 = n1638 & n1654 ;
  assign n1656 = x183 ^ x10 ^ 1'b0 ;
  assign n1657 = n655 & n1656 ;
  assign n1658 = n1657 ^ n1289 ^ 1'b0 ;
  assign n1659 = x22 | n623 ;
  assign n1660 = x139 & n435 ;
  assign n1661 = ~n1659 & n1660 ;
  assign n1662 = x30 & x76 ;
  assign n1663 = n947 & n1662 ;
  assign n1664 = ( n874 & ~n1410 ) | ( n874 & n1663 ) | ( ~n1410 & n1663 ) ;
  assign n1665 = n1318 ^ n1166 ^ 1'b0 ;
  assign n1666 = n925 ^ n853 ^ x65 ;
  assign n1667 = n1665 & ~n1666 ;
  assign n1668 = ~n1066 & n1650 ;
  assign n1669 = n1668 ^ n602 ^ 1'b0 ;
  assign n1670 = n1669 ^ n982 ^ 1'b0 ;
  assign n1671 = n688 | n1670 ;
  assign n1672 = n1475 ^ x129 ^ 1'b0 ;
  assign n1673 = ~n396 & n445 ;
  assign n1674 = n1673 ^ n1038 ^ x110 ;
  assign n1675 = n1674 ^ n1366 ^ 1'b0 ;
  assign n1676 = ~n441 & n1351 ;
  assign n1677 = n1676 ^ n645 ^ 1'b0 ;
  assign n1678 = n1677 ^ x216 ^ 1'b0 ;
  assign n1679 = n1678 ^ n1019 ^ 1'b0 ;
  assign n1680 = x157 & n1679 ;
  assign n1681 = ~n807 & n1680 ;
  assign n1682 = n1681 ^ x54 ^ 1'b0 ;
  assign n1683 = n1653 | n1672 ;
  assign n1684 = n1155 | n1683 ;
  assign n1685 = n1044 ^ x179 ^ 1'b0 ;
  assign n1686 = x215 & ~n1685 ;
  assign n1687 = ~n393 & n1686 ;
  assign n1688 = n1687 ^ n1316 ^ x32 ;
  assign n1689 = n335 | n1131 ;
  assign n1690 = x167 & n623 ;
  assign n1691 = ( ~n1504 & n1678 ) | ( ~n1504 & n1690 ) | ( n1678 & n1690 ) ;
  assign n1692 = x24 & ~n1691 ;
  assign n1693 = n1689 & n1692 ;
  assign n1694 = ( x216 & n816 ) | ( x216 & n1693 ) | ( n816 & n1693 ) ;
  assign n1695 = ~x219 & n678 ;
  assign n1696 = n1316 | n1559 ;
  assign n1697 = n308 ^ x137 ^ 1'b0 ;
  assign n1698 = x25 & n1697 ;
  assign n1699 = ~n467 & n839 ;
  assign n1700 = ~n1698 & n1699 ;
  assign n1701 = x48 & n1700 ;
  assign n1702 = n1701 ^ n913 ^ 1'b0 ;
  assign n1703 = x206 ^ x41 ^ 1'b0 ;
  assign n1704 = x74 & ~n1703 ;
  assign n1705 = n1704 ^ n1691 ^ 1'b0 ;
  assign n1718 = n1365 ^ x81 ^ x65 ;
  assign n1717 = n708 ^ n656 ^ n415 ;
  assign n1710 = n377 ^ x149 ^ 1'b0 ;
  assign n1711 = n633 | n1710 ;
  assign n1712 = n1711 ^ n1009 ^ 1'b0 ;
  assign n1713 = ~n1356 & n1712 ;
  assign n1706 = x228 & ~n686 ;
  assign n1707 = ~x85 & n1706 ;
  assign n1708 = x150 & ~n1707 ;
  assign n1709 = n1708 ^ n647 ^ 1'b0 ;
  assign n1714 = n1713 ^ n1709 ^ 1'b0 ;
  assign n1715 = x55 & ~n1714 ;
  assign n1716 = ( n671 & n913 ) | ( n671 & n1715 ) | ( n913 & n1715 ) ;
  assign n1719 = n1718 ^ n1717 ^ n1716 ;
  assign n1720 = n737 ^ x151 ^ 1'b0 ;
  assign n1721 = n1720 ^ n756 ^ 1'b0 ;
  assign n1722 = n1090 | n1721 ;
  assign n1723 = n398 | n997 ;
  assign n1724 = ( ~x61 & x112 ) | ( ~x61 & n493 ) | ( x112 & n493 ) ;
  assign n1725 = n898 ^ n425 ^ x241 ;
  assign n1726 = n1725 ^ n1068 ^ 1'b0 ;
  assign n1727 = n1724 | n1726 ;
  assign n1728 = n987 ^ n352 ^ 1'b0 ;
  assign n1729 = n921 ^ n694 ^ n552 ;
  assign n1741 = n1729 ^ n1068 ^ x254 ;
  assign n1730 = n1729 ^ x41 ^ 1'b0 ;
  assign n1731 = ~n519 & n1730 ;
  assign n1732 = ( n1173 & n1304 ) | ( n1173 & n1731 ) | ( n1304 & n1731 ) ;
  assign n1733 = n257 ^ x74 ^ 1'b0 ;
  assign n1734 = n717 ^ x8 ^ 1'b0 ;
  assign n1735 = x233 & n729 ;
  assign n1736 = n1734 & n1735 ;
  assign n1737 = n1736 ^ x93 ^ 1'b0 ;
  assign n1738 = n1733 | n1737 ;
  assign n1739 = n1738 ^ n407 ^ 1'b0 ;
  assign n1740 = ( n1415 & n1732 ) | ( n1415 & ~n1739 ) | ( n1732 & ~n1739 ) ;
  assign n1742 = n1741 ^ n1740 ^ 1'b0 ;
  assign n1743 = x89 & n1484 ;
  assign n1744 = n1743 ^ x214 ^ 1'b0 ;
  assign n1745 = n680 & n961 ;
  assign n1746 = n1228 & n1745 ;
  assign n1747 = n794 & ~n1289 ;
  assign n1748 = n1747 ^ n599 ^ 1'b0 ;
  assign n1749 = n1711 ^ n1386 ^ 1'b0 ;
  assign n1751 = ( x8 & ~n759 ) | ( x8 & n1406 ) | ( ~n759 & n1406 ) ;
  assign n1750 = ( n326 & ~n461 ) | ( n326 & n926 ) | ( ~n461 & n926 ) ;
  assign n1752 = n1751 ^ n1750 ^ n1164 ;
  assign n1754 = n444 & ~n818 ;
  assign n1753 = n603 & n1301 ;
  assign n1755 = n1754 ^ n1753 ^ 1'b0 ;
  assign n1756 = n783 | n1356 ;
  assign n1757 = n440 & ~n1756 ;
  assign n1758 = n1140 & n1757 ;
  assign n1759 = n667 | n1002 ;
  assign n1760 = n1759 ^ n1319 ^ 1'b0 ;
  assign n1761 = ( x183 & n1576 ) | ( x183 & n1760 ) | ( n1576 & n1760 ) ;
  assign n1762 = n271 & ~n489 ;
  assign n1763 = ~n953 & n1762 ;
  assign n1764 = n1145 | n1763 ;
  assign n1765 = n1764 ^ n733 ^ 1'b0 ;
  assign n1766 = ( n531 & n773 ) | ( n531 & n1750 ) | ( n773 & n1750 ) ;
  assign n1767 = n1766 ^ n1120 ^ 1'b0 ;
  assign n1768 = n679 & n1767 ;
  assign n1770 = n381 ^ x122 ^ x89 ;
  assign n1769 = ( n672 & ~n845 ) | ( n672 & n1352 ) | ( ~n845 & n1352 ) ;
  assign n1771 = n1770 ^ n1769 ^ 1'b0 ;
  assign n1772 = n1010 | n1771 ;
  assign n1773 = ( ~n256 & n1768 ) | ( ~n256 & n1772 ) | ( n1768 & n1772 ) ;
  assign n1774 = n936 ^ n785 ^ 1'b0 ;
  assign n1775 = n1774 ^ n256 ^ 1'b0 ;
  assign n1777 = x121 & n256 ;
  assign n1778 = n1777 ^ n507 ^ 1'b0 ;
  assign n1779 = n1594 ^ n939 ^ 1'b0 ;
  assign n1780 = n1778 & ~n1779 ;
  assign n1776 = n1579 ^ x157 ^ 1'b0 ;
  assign n1781 = n1780 ^ n1776 ^ 1'b0 ;
  assign n1783 = x148 & ~n1353 ;
  assign n1784 = ~n341 & n1783 ;
  assign n1785 = n385 & ~n1784 ;
  assign n1786 = n1785 ^ x52 ^ 1'b0 ;
  assign n1782 = x55 & ~n335 ;
  assign n1787 = n1786 ^ n1782 ^ 1'b0 ;
  assign n1788 = n1781 & ~n1787 ;
  assign n1789 = ( n642 & n994 ) | ( n642 & n1247 ) | ( n994 & n1247 ) ;
  assign n1790 = n1031 ^ x59 ^ 1'b0 ;
  assign n1791 = n1789 & n1790 ;
  assign n1792 = n344 ^ x65 ^ 1'b0 ;
  assign n1793 = x200 & n1792 ;
  assign n1794 = n1793 ^ x98 ^ 1'b0 ;
  assign n1798 = x218 & ~n780 ;
  assign n1799 = n464 & n1798 ;
  assign n1800 = ( ~n260 & n1452 ) | ( ~n260 & n1799 ) | ( n1452 & n1799 ) ;
  assign n1795 = ( x98 & x205 ) | ( x98 & n377 ) | ( x205 & n377 ) ;
  assign n1796 = n1094 & n1795 ;
  assign n1797 = n1796 ^ n369 ^ 1'b0 ;
  assign n1801 = n1800 ^ n1797 ^ 1'b0 ;
  assign n1802 = n1794 & ~n1801 ;
  assign n1803 = n1802 ^ n903 ^ n513 ;
  assign n1804 = x120 & ~n1803 ;
  assign n1805 = n1804 ^ n1376 ^ n1160 ;
  assign n1806 = ( x127 & ~n1791 ) | ( x127 & n1805 ) | ( ~n1791 & n1805 ) ;
  assign n1807 = ~n615 & n787 ;
  assign n1808 = n1807 ^ n872 ^ 1'b0 ;
  assign n1809 = ~n1803 & n1808 ;
  assign n1810 = n1285 ^ x178 ^ 1'b0 ;
  assign n1811 = n1810 ^ x10 ^ 1'b0 ;
  assign n1812 = n1809 & n1811 ;
  assign n1826 = x217 & n727 ;
  assign n1827 = ~x36 & n1826 ;
  assign n1828 = n1827 ^ n764 ^ 1'b0 ;
  assign n1829 = ( n806 & n1701 ) | ( n806 & n1828 ) | ( n1701 & n1828 ) ;
  assign n1813 = n1720 ^ n994 ^ 1'b0 ;
  assign n1814 = x123 & n820 ;
  assign n1815 = n586 & n1814 ;
  assign n1816 = n1815 ^ n1432 ^ 1'b0 ;
  assign n1817 = n1729 ^ n496 ^ x187 ;
  assign n1818 = ( n1813 & ~n1816 ) | ( n1813 & n1817 ) | ( ~n1816 & n1817 ) ;
  assign n1819 = x64 & n966 ;
  assign n1820 = ~x208 & n1819 ;
  assign n1821 = n1647 ^ n535 ^ x18 ;
  assign n1822 = x196 & n1821 ;
  assign n1823 = n1820 & n1822 ;
  assign n1824 = n1590 & ~n1823 ;
  assign n1825 = ~n1818 & n1824 ;
  assign n1830 = n1829 ^ n1825 ^ 1'b0 ;
  assign n1834 = n1086 ^ x48 ^ 1'b0 ;
  assign n1835 = n1222 | n1834 ;
  assign n1832 = n735 & n820 ;
  assign n1833 = n345 | n1832 ;
  assign n1836 = n1835 ^ n1833 ^ 1'b0 ;
  assign n1831 = ( ~x26 & n500 ) | ( ~x26 & n606 ) | ( n500 & n606 ) ;
  assign n1837 = n1836 ^ n1831 ^ 1'b0 ;
  assign n1838 = ~n894 & n1837 ;
  assign n1839 = n715 ^ n485 ^ 1'b0 ;
  assign n1840 = ~n259 & n1839 ;
  assign n1842 = n263 & ~n556 ;
  assign n1841 = n704 & n1579 ;
  assign n1843 = n1842 ^ n1841 ^ 1'b0 ;
  assign n1844 = n1843 ^ n1039 ^ x188 ;
  assign n1845 = ( ~n1439 & n1840 ) | ( ~n1439 & n1844 ) | ( n1840 & n1844 ) ;
  assign n1846 = n1606 ^ n644 ^ 1'b0 ;
  assign n1847 = n433 & ~n1846 ;
  assign n1848 = n967 ^ n885 ^ 1'b0 ;
  assign n1849 = ( ~n854 & n1068 ) | ( ~n854 & n1154 ) | ( n1068 & n1154 ) ;
  assign n1850 = x188 & n410 ;
  assign n1851 = n1521 ^ n877 ^ n839 ;
  assign n1852 = n1850 & n1851 ;
  assign n1853 = ~x138 & n537 ;
  assign n1854 = x149 & n1853 ;
  assign n1855 = n708 & n1854 ;
  assign n1856 = ( x4 & n1011 ) | ( x4 & ~n1855 ) | ( n1011 & ~n1855 ) ;
  assign n1857 = n1856 ^ n499 ^ 1'b0 ;
  assign n1858 = n638 | n1857 ;
  assign n1859 = n1858 ^ n1271 ^ 1'b0 ;
  assign n1860 = ( ~x12 & x133 ) | ( ~x12 & n514 ) | ( x133 & n514 ) ;
  assign n1861 = n962 & n1860 ;
  assign n1862 = n1861 ^ x71 ^ 1'b0 ;
  assign n1863 = n347 & n1220 ;
  assign n1864 = n561 | n1863 ;
  assign n1865 = n1021 & ~n1864 ;
  assign n1866 = n1288 | n1829 ;
  assign n1867 = n1067 | n1866 ;
  assign n1868 = ~n1865 & n1867 ;
  assign n1869 = ~n868 & n1868 ;
  assign n1870 = n375 & ~n1869 ;
  assign n1871 = n444 ^ n403 ^ n351 ;
  assign n1872 = x242 ^ x223 ^ 1'b0 ;
  assign n1873 = x103 & n1872 ;
  assign n1874 = n1873 ^ n572 ^ 1'b0 ;
  assign n1875 = n1874 ^ x70 ^ x1 ;
  assign n1876 = ~n1871 & n1875 ;
  assign n1877 = ~n852 & n1876 ;
  assign n1878 = n1665 & ~n1877 ;
  assign n1879 = n1878 ^ x16 ^ 1'b0 ;
  assign n1880 = x160 ^ x139 ^ 1'b0 ;
  assign n1881 = n1880 ^ n1126 ^ x32 ;
  assign n1882 = n1881 ^ n1548 ^ x112 ;
  assign n1883 = n1585 ^ x79 ^ 1'b0 ;
  assign n1884 = n1116 & ~n1883 ;
  assign n1885 = ~n1754 & n1884 ;
  assign n1886 = n1525 ^ x252 ^ 1'b0 ;
  assign n1887 = x46 & ~n349 ;
  assign n1888 = ~n292 & n1887 ;
  assign n1889 = x57 & ~n928 ;
  assign n1890 = n1888 & n1889 ;
  assign n1891 = n825 ^ x227 ^ 1'b0 ;
  assign n1892 = ~n490 & n1891 ;
  assign n1893 = n1892 ^ x178 ^ 1'b0 ;
  assign n1894 = n1118 ^ n509 ^ 1'b0 ;
  assign n1895 = ~n1893 & n1894 ;
  assign n1896 = n1890 | n1895 ;
  assign n1898 = n1795 ^ n1562 ^ 1'b0 ;
  assign n1897 = x194 & n444 ;
  assign n1899 = n1898 ^ n1897 ^ 1'b0 ;
  assign n1900 = ~n816 & n1649 ;
  assign n1901 = n1286 | n1900 ;
  assign n1902 = n1899 | n1901 ;
  assign n1903 = ~n854 & n1458 ;
  assign n1904 = n1903 ^ n1440 ^ 1'b0 ;
  assign n1905 = n387 & n1904 ;
  assign n1906 = n1905 ^ x144 ^ 1'b0 ;
  assign n1907 = ( x242 & n1361 ) | ( x242 & ~n1906 ) | ( n1361 & ~n1906 ) ;
  assign n1908 = n1795 ^ n1514 ^ 1'b0 ;
  assign n1909 = ( x46 & n665 ) | ( x46 & ~n939 ) | ( n665 & ~n939 ) ;
  assign n1910 = n1909 ^ n1190 ^ 1'b0 ;
  assign n1911 = n1910 ^ n1836 ^ 1'b0 ;
  assign n1912 = n1908 | n1911 ;
  assign n1913 = n936 | n1071 ;
  assign n1917 = n881 ^ x160 ^ 1'b0 ;
  assign n1918 = n1113 | n1917 ;
  assign n1919 = ( ~n609 & n943 ) | ( ~n609 & n1918 ) | ( n943 & n1918 ) ;
  assign n1920 = n1329 & ~n1919 ;
  assign n1921 = ~n627 & n1920 ;
  assign n1914 = x94 & ~x241 ;
  assign n1915 = x85 & ~n1914 ;
  assign n1916 = n1915 ^ x51 ^ 1'b0 ;
  assign n1922 = n1921 ^ n1916 ^ x202 ;
  assign n1923 = n898 ^ n861 ^ n387 ;
  assign n1924 = ~n1835 & n1923 ;
  assign n1925 = n1924 ^ x71 ^ 1'b0 ;
  assign n1926 = n478 | n1925 ;
  assign n1927 = n1926 ^ n371 ^ 1'b0 ;
  assign n1928 = n951 ^ n743 ^ n409 ;
  assign n1929 = n1910 & n1928 ;
  assign n1930 = n1929 ^ n1523 ^ 1'b0 ;
  assign n1931 = x133 ^ x66 ^ 1'b0 ;
  assign n1932 = n460 | n1532 ;
  assign n1933 = ~n1931 & n1932 ;
  assign n1934 = n1718 ^ n1700 ^ n1011 ;
  assign n1935 = n297 & ~n1934 ;
  assign n1936 = n936 & ~n1935 ;
  assign n1937 = n1202 & ~n1936 ;
  assign n1938 = n1632 ^ n393 ^ 1'b0 ;
  assign n1939 = ( x38 & ~n591 ) | ( x38 & n1938 ) | ( ~n591 & n1938 ) ;
  assign n1940 = ~n375 & n1939 ;
  assign n1941 = x159 & n1031 ;
  assign n1944 = n405 ^ x139 ^ 1'b0 ;
  assign n1942 = n262 ^ x102 ^ 1'b0 ;
  assign n1943 = n716 & ~n1942 ;
  assign n1945 = n1944 ^ n1943 ^ 1'b0 ;
  assign n1946 = n1941 & ~n1945 ;
  assign n1947 = x186 & ~n314 ;
  assign n1948 = n1947 ^ n1723 ^ 1'b0 ;
  assign n1949 = n911 & n1451 ;
  assign n1950 = n1949 ^ n1292 ^ n260 ;
  assign n1951 = n427 ^ x25 ^ 1'b0 ;
  assign n1952 = n936 & n1413 ;
  assign n1953 = n1952 ^ n1442 ^ 1'b0 ;
  assign n1954 = x74 & n853 ;
  assign n1955 = n1954 ^ n1553 ^ 1'b0 ;
  assign n1956 = n1867 ^ n554 ^ n298 ;
  assign n1957 = n1550 ^ n371 ^ 1'b0 ;
  assign n1958 = n382 & n1957 ;
  assign n1959 = ( n1019 & n1881 ) | ( n1019 & n1958 ) | ( n1881 & n1958 ) ;
  assign n1960 = n1956 & ~n1959 ;
  assign n1961 = n1955 & n1960 ;
  assign n1962 = ( n300 & n795 ) | ( n300 & n1057 ) | ( n795 & n1057 ) ;
  assign n1963 = n1962 ^ x145 ^ 1'b0 ;
  assign n1964 = n1076 ^ n801 ^ 1'b0 ;
  assign n1968 = n1809 ^ n1035 ^ 1'b0 ;
  assign n1965 = n824 & ~n1174 ;
  assign n1966 = ~n580 & n1965 ;
  assign n1967 = n1079 & ~n1966 ;
  assign n1969 = n1968 ^ n1967 ^ 1'b0 ;
  assign n1970 = n1803 ^ n1251 ^ 1'b0 ;
  assign n1971 = ~x72 & n1970 ;
  assign n1972 = n1971 ^ n1064 ^ 1'b0 ;
  assign n1974 = n627 & n1067 ;
  assign n1975 = ~n1793 & n1974 ;
  assign n1976 = x105 | n1148 ;
  assign n1977 = ~n1975 & n1976 ;
  assign n1978 = n1977 ^ n1329 ^ 1'b0 ;
  assign n1973 = x192 & ~n297 ;
  assign n1979 = n1978 ^ n1973 ^ 1'b0 ;
  assign n1980 = n1979 ^ n417 ^ 1'b0 ;
  assign n1981 = n405 ^ x116 ^ x70 ;
  assign n1982 = n314 | n1981 ;
  assign n1983 = n1982 ^ n1331 ^ 1'b0 ;
  assign n1984 = n1179 ^ x150 ^ 1'b0 ;
  assign n1985 = n1573 | n1984 ;
  assign n1986 = n794 & ~n1037 ;
  assign n1987 = n1986 ^ n914 ^ 1'b0 ;
  assign n1988 = x17 & ~n1987 ;
  assign n1989 = n1988 ^ n1174 ^ 1'b0 ;
  assign n1990 = n1989 ^ x140 ^ 1'b0 ;
  assign n1991 = n1985 | n1990 ;
  assign n1992 = ~n1002 & n1312 ;
  assign n1993 = n1759 & n1992 ;
  assign n1994 = n1993 ^ n1806 ^ n1597 ;
  assign n1995 = n1616 ^ n1274 ^ n923 ;
  assign n1996 = ( ~x234 & x239 ) | ( ~x234 & n1995 ) | ( x239 & n1995 ) ;
  assign n1997 = ~n1669 & n1996 ;
  assign n1998 = ~n1031 & n1997 ;
  assign n1999 = n1189 ^ x172 ^ x45 ;
  assign n2000 = n794 & n1622 ;
  assign n2001 = n1142 & n2000 ;
  assign n2002 = x110 & x213 ;
  assign n2003 = n2001 & n2002 ;
  assign n2004 = n907 ^ n498 ^ x202 ;
  assign n2005 = n2004 ^ n667 ^ 1'b0 ;
  assign n2006 = n1787 | n2005 ;
  assign n2007 = n2006 ^ n1040 ^ n974 ;
  assign n2008 = x123 & ~n523 ;
  assign n2009 = n2008 ^ n870 ^ 1'b0 ;
  assign n2011 = n522 & n1253 ;
  assign n2012 = ~n823 & n2011 ;
  assign n2010 = n1150 | n1335 ;
  assign n2013 = n2012 ^ n2010 ^ 1'b0 ;
  assign n2014 = n2009 | n2013 ;
  assign n2015 = n757 | n2014 ;
  assign n2016 = n2015 ^ n1882 ^ 1'b0 ;
  assign n2017 = n1759 ^ n1647 ^ 1'b0 ;
  assign n2018 = x197 & n1319 ;
  assign n2019 = ~n2017 & n2018 ;
  assign n2020 = ~n565 & n593 ;
  assign n2021 = n2020 ^ n316 ^ 1'b0 ;
  assign n2022 = n2021 ^ n1174 ^ n1104 ;
  assign n2023 = ( n1846 & n2019 ) | ( n1846 & ~n2022 ) | ( n2019 & ~n2022 ) ;
  assign n2024 = n1702 ^ n322 ^ 1'b0 ;
  assign n2025 = ( n512 & n967 ) | ( n512 & ~n1918 ) | ( n967 & ~n1918 ) ;
  assign n2026 = n1111 ^ x198 ^ 1'b0 ;
  assign n2027 = ~n1314 & n1629 ;
  assign n2028 = ~n516 & n2027 ;
  assign n2029 = n2028 ^ n973 ^ 1'b0 ;
  assign n2030 = ~n280 & n2029 ;
  assign n2031 = ~n1345 & n2030 ;
  assign n2032 = ~x169 & n2031 ;
  assign n2033 = ( n756 & n947 ) | ( n756 & ~n2032 ) | ( n947 & ~n2032 ) ;
  assign n2034 = n690 ^ n310 ^ 1'b0 ;
  assign n2035 = n1659 & ~n2034 ;
  assign n2036 = n282 ^ x77 ^ 1'b0 ;
  assign n2037 = n1312 & ~n2036 ;
  assign n2038 = n1863 & n2037 ;
  assign n2039 = n293 & n415 ;
  assign n2040 = n2039 ^ n1161 ^ 1'b0 ;
  assign n2041 = ~n1309 & n2040 ;
  assign n2042 = ( n1944 & n2038 ) | ( n1944 & n2041 ) | ( n2038 & n2041 ) ;
  assign n2043 = n2042 ^ n1750 ^ 1'b0 ;
  assign n2044 = x4 & ~n513 ;
  assign n2045 = n2044 ^ x72 ^ 1'b0 ;
  assign n2046 = n1173 | n2045 ;
  assign n2047 = n2046 ^ n706 ^ x71 ;
  assign n2048 = n337 & n2047 ;
  assign n2049 = n1314 ^ n557 ^ n270 ;
  assign n2050 = ( ~x99 & n785 ) | ( ~x99 & n2049 ) | ( n785 & n2049 ) ;
  assign n2052 = x186 & ~n1677 ;
  assign n2053 = x213 & n1281 ;
  assign n2054 = n1012 & n2053 ;
  assign n2055 = n606 ^ n302 ^ 1'b0 ;
  assign n2056 = ( n2052 & n2054 ) | ( n2052 & ~n2055 ) | ( n2054 & ~n2055 ) ;
  assign n2051 = n2017 ^ n415 ^ 1'b0 ;
  assign n2057 = n2056 ^ n2051 ^ n1628 ;
  assign n2058 = n1200 ^ n754 ^ x25 ;
  assign n2059 = ~n2057 & n2058 ;
  assign n2060 = n1388 & ~n1651 ;
  assign n2061 = n440 & n2060 ;
  assign n2062 = n2061 ^ n691 ^ 1'b0 ;
  assign n2063 = n1736 ^ n1005 ^ 1'b0 ;
  assign n2064 = n1439 & n2063 ;
  assign n2065 = n1312 & n2064 ;
  assign n2066 = ~n627 & n2065 ;
  assign n2067 = ~x154 & n602 ;
  assign n2068 = ~x21 & n596 ;
  assign n2069 = n644 | n1687 ;
  assign n2070 = n2069 ^ n856 ^ 1'b0 ;
  assign n2071 = n557 | n1669 ;
  assign n2072 = n2071 ^ n1318 ^ 1'b0 ;
  assign n2073 = ~n2070 & n2072 ;
  assign n2074 = ~n2068 & n2073 ;
  assign n2075 = n2067 & n2074 ;
  assign n2076 = n2066 | n2075 ;
  assign n2077 = n1285 & ~n2076 ;
  assign n2078 = n567 & n810 ;
  assign n2079 = ~n317 & n890 ;
  assign n2080 = n1690 & n2079 ;
  assign n2081 = n1778 | n2080 ;
  assign n2082 = n2078 & ~n2081 ;
  assign n2083 = n297 ^ x47 ^ 1'b0 ;
  assign n2084 = ~n1987 & n2083 ;
  assign n2085 = n2084 ^ x153 ^ 1'b0 ;
  assign n2086 = n2012 ^ x135 ^ 1'b0 ;
  assign n2087 = x207 ^ x143 ^ 1'b0 ;
  assign n2088 = x163 & n2087 ;
  assign n2089 = ( n711 & ~n986 ) | ( n711 & n2088 ) | ( ~n986 & n2088 ) ;
  assign n2090 = n2089 ^ n1615 ^ n440 ;
  assign n2091 = x56 & ~n1447 ;
  assign n2092 = ~n2090 & n2091 ;
  assign n2093 = n2092 ^ n1231 ^ 1'b0 ;
  assign n2094 = ~n280 & n2093 ;
  assign n2095 = n1096 | n1606 ;
  assign n2096 = n339 & n1781 ;
  assign n2097 = n2096 ^ n1274 ^ 1'b0 ;
  assign n2098 = n2097 ^ x91 ^ 1'b0 ;
  assign n2099 = n561 | n1768 ;
  assign n2100 = n2099 ^ n1856 ^ 1'b0 ;
  assign n2101 = x77 & ~n419 ;
  assign n2102 = n2101 ^ x196 ^ 1'b0 ;
  assign n2103 = ( n338 & n576 ) | ( n338 & ~n2102 ) | ( n576 & ~n2102 ) ;
  assign n2110 = x233 | n1314 ;
  assign n2105 = n795 ^ n531 ^ x31 ;
  assign n2104 = n612 | n967 ;
  assign n2106 = n2105 ^ n2104 ^ 1'b0 ;
  assign n2107 = ( n635 & n903 ) | ( n635 & ~n2106 ) | ( n903 & ~n2106 ) ;
  assign n2108 = n1853 ^ n487 ^ 1'b0 ;
  assign n2109 = ~n2107 & n2108 ;
  assign n2111 = n2110 ^ n2109 ^ 1'b0 ;
  assign n2112 = n356 & ~n1110 ;
  assign n2113 = n2112 ^ n1904 ^ n1580 ;
  assign n2114 = n1567 ^ x158 ^ 1'b0 ;
  assign n2115 = n1684 & n2097 ;
  assign n2116 = ~n425 & n2115 ;
  assign n2119 = n1644 ^ n885 ^ n436 ;
  assign n2117 = n1553 ^ n1023 ^ n453 ;
  assign n2118 = n2117 ^ n588 ^ x15 ;
  assign n2120 = n2119 ^ n2118 ^ 1'b0 ;
  assign n2121 = n956 | n2120 ;
  assign n2122 = x58 & n2121 ;
  assign n2123 = n2122 ^ n2088 ^ 1'b0 ;
  assign n2124 = n1068 ^ n545 ^ x191 ;
  assign n2125 = ( n449 & n715 ) | ( n449 & ~n1607 ) | ( n715 & ~n1607 ) ;
  assign n2126 = ( x246 & ~n1310 ) | ( x246 & n1829 ) | ( ~n1310 & n1829 ) ;
  assign n2127 = n859 | n2126 ;
  assign n2128 = n2127 ^ n704 ^ 1'b0 ;
  assign n2129 = n2125 & n2128 ;
  assign n2130 = ~n536 & n2129 ;
  assign n2131 = ( x67 & n2124 ) | ( x67 & n2130 ) | ( n2124 & n2130 ) ;
  assign n2132 = n629 | n825 ;
  assign n2133 = n2132 ^ n632 ^ 1'b0 ;
  assign n2134 = n467 | n2133 ;
  assign n2135 = n2134 ^ n273 ^ 1'b0 ;
  assign n2136 = x21 & n312 ;
  assign n2137 = ( x146 & n493 ) | ( x146 & n2136 ) | ( n493 & n2136 ) ;
  assign n2138 = ~n1131 & n2137 ;
  assign n2139 = x246 & ~n811 ;
  assign n2140 = n545 & n2139 ;
  assign n2141 = ( n729 & ~n990 ) | ( n729 & n2125 ) | ( ~n990 & n2125 ) ;
  assign n2142 = n2141 ^ n790 ^ n638 ;
  assign n2143 = x73 & ~n1370 ;
  assign n2144 = ~n1543 & n2143 ;
  assign n2145 = n843 ^ n614 ^ 1'b0 ;
  assign n2146 = ~n1362 & n2145 ;
  assign n2147 = ( n572 & ~n825 ) | ( n572 & n1479 ) | ( ~n825 & n1479 ) ;
  assign n2148 = n2147 ^ n402 ^ 1'b0 ;
  assign n2149 = n1285 & n2148 ;
  assign n2150 = n807 & n2149 ;
  assign n2151 = n284 | n1425 ;
  assign n2152 = n1836 ^ n1123 ^ 1'b0 ;
  assign n2153 = n2151 | n2152 ;
  assign n2154 = n1643 & ~n2153 ;
  assign n2155 = ( ~n862 & n986 ) | ( ~n862 & n1352 ) | ( n986 & n1352 ) ;
  assign n2156 = n1009 ^ n421 ^ 1'b0 ;
  assign n2157 = ~n638 & n2156 ;
  assign n2158 = n1264 & n2157 ;
  assign n2159 = n2158 ^ n1644 ^ 1'b0 ;
  assign n2160 = n1713 ^ n576 ^ 1'b0 ;
  assign n2161 = ~n1122 & n1460 ;
  assign n2162 = n2161 ^ n1435 ^ 1'b0 ;
  assign n2163 = x179 & ~n782 ;
  assign n2164 = ~n771 & n2163 ;
  assign n2165 = x127 ^ x71 ^ 1'b0 ;
  assign n2166 = n2165 ^ n1034 ^ 1'b0 ;
  assign n2167 = ~n2164 & n2166 ;
  assign n2168 = n382 & n2167 ;
  assign n2169 = ~n2162 & n2168 ;
  assign n2170 = n503 | n2169 ;
  assign n2171 = n2160 & ~n2170 ;
  assign n2172 = n1069 ^ n807 ^ x13 ;
  assign n2173 = n496 & n947 ;
  assign n2174 = n1328 & ~n1993 ;
  assign n2175 = n436 & n2174 ;
  assign n2176 = n2175 ^ n679 ^ 1'b0 ;
  assign n2177 = n1243 ^ x134 ^ 1'b0 ;
  assign n2178 = n1561 & n2177 ;
  assign n2179 = x83 & ~n1620 ;
  assign n2181 = n873 & ~n1757 ;
  assign n2182 = n2181 ^ n1744 ^ 1'b0 ;
  assign n2180 = ~n288 & n1082 ;
  assign n2183 = n2182 ^ n2180 ^ 1'b0 ;
  assign n2184 = n1643 ^ x128 ^ 1'b0 ;
  assign n2185 = x162 | n2184 ;
  assign n2186 = x107 | n2185 ;
  assign n2187 = n655 ^ x218 ^ 1'b0 ;
  assign n2188 = ~n967 & n2187 ;
  assign n2189 = ( n413 & ~n1600 ) | ( n413 & n2188 ) | ( ~n1600 & n2188 ) ;
  assign n2190 = x30 & ~n609 ;
  assign n2191 = n2190 ^ x101 ^ 1'b0 ;
  assign n2192 = ( x149 & n262 ) | ( x149 & ~n2191 ) | ( n262 & ~n2191 ) ;
  assign n2193 = n2192 ^ n1296 ^ n571 ;
  assign n2194 = ~x103 & n399 ;
  assign n2195 = n2136 & ~n2194 ;
  assign n2196 = ~n2193 & n2195 ;
  assign n2197 = n1360 ^ n421 ^ 1'b0 ;
  assign n2198 = ~n848 & n1174 ;
  assign n2199 = ~n352 & n2198 ;
  assign n2200 = n619 | n2199 ;
  assign n2201 = n407 & ~n1525 ;
  assign n2203 = x146 ^ x27 ^ 1'b0 ;
  assign n2204 = x246 & ~n2203 ;
  assign n2205 = ( ~x129 & n403 ) | ( ~x129 & n2204 ) | ( n403 & n2204 ) ;
  assign n2202 = n282 ^ x117 ^ 1'b0 ;
  assign n2206 = n2205 ^ n2202 ^ 1'b0 ;
  assign n2207 = x109 & n2206 ;
  assign n2208 = ( n686 & n2201 ) | ( n686 & n2207 ) | ( n2201 & n2207 ) ;
  assign n2209 = ( ~n2073 & n2200 ) | ( ~n2073 & n2208 ) | ( n2200 & n2208 ) ;
  assign n2210 = n490 ^ x225 ^ x186 ;
  assign n2211 = x229 & n2210 ;
  assign n2212 = n2211 ^ x5 ^ 1'b0 ;
  assign n2213 = x149 & ~x162 ;
  assign n2214 = n2213 ^ x198 ^ 1'b0 ;
  assign n2215 = ( n399 & n1472 ) | ( n399 & n2214 ) | ( n1472 & n2214 ) ;
  assign n2216 = ( n1236 & ~n2212 ) | ( n1236 & n2215 ) | ( ~n2212 & n2215 ) ;
  assign n2217 = n2216 ^ x93 ^ 1'b0 ;
  assign n2218 = n1616 ^ n270 ^ 1'b0 ;
  assign n2219 = n1873 & n2218 ;
  assign n2223 = n1622 ^ x74 ^ x70 ;
  assign n2220 = n545 ^ x196 ^ 1'b0 ;
  assign n2221 = n1687 ^ x36 ^ 1'b0 ;
  assign n2222 = ( n2090 & n2220 ) | ( n2090 & n2221 ) | ( n2220 & n2221 ) ;
  assign n2224 = n2223 ^ n2222 ^ 1'b0 ;
  assign n2225 = n630 | n2224 ;
  assign n2226 = ~x230 & n1478 ;
  assign n2228 = n1209 ^ n717 ^ 1'b0 ;
  assign n2227 = ( x193 & n501 ) | ( x193 & ~n1243 ) | ( n501 & ~n1243 ) ;
  assign n2229 = n2228 ^ n2227 ^ 1'b0 ;
  assign n2230 = n1500 ^ n472 ^ x117 ;
  assign n2231 = ~n710 & n2230 ;
  assign n2232 = n704 & ~n1005 ;
  assign n2233 = n2232 ^ n1144 ^ 1'b0 ;
  assign n2237 = x139 & ~n1533 ;
  assign n2238 = ~x214 & n2237 ;
  assign n2239 = n2238 ^ n1647 ^ 1'b0 ;
  assign n2240 = x144 & ~n2239 ;
  assign n2236 = x73 & n396 ;
  assign n2241 = n2240 ^ n2236 ^ 1'b0 ;
  assign n2242 = n1965 & n2241 ;
  assign n2234 = n654 ^ n449 ^ 1'b0 ;
  assign n2235 = n440 | n2234 ;
  assign n2243 = n2242 ^ n2235 ^ 1'b0 ;
  assign n2246 = n586 ^ x137 ^ 1'b0 ;
  assign n2247 = ~n894 & n2246 ;
  assign n2244 = ( x65 & n847 ) | ( x65 & ~n1100 ) | ( n847 & ~n1100 ) ;
  assign n2245 = n2244 ^ n1842 ^ n578 ;
  assign n2248 = n2247 ^ n2245 ^ n1295 ;
  assign n2249 = ~n1136 & n1776 ;
  assign n2250 = n809 & n2249 ;
  assign n2251 = ~n1120 & n1140 ;
  assign n2252 = x17 & ~n2251 ;
  assign n2253 = n2252 ^ n474 ^ 1'b0 ;
  assign n2254 = ~n1256 & n1499 ;
  assign n2255 = ~n1271 & n2254 ;
  assign n2261 = n1644 & n1886 ;
  assign n2256 = n635 ^ n287 ^ 1'b0 ;
  assign n2257 = x188 | n1784 ;
  assign n2258 = n2256 & ~n2257 ;
  assign n2259 = ~n952 & n2258 ;
  assign n2260 = ( x90 & ~n537 ) | ( x90 & n2259 ) | ( ~n537 & n2259 ) ;
  assign n2262 = n2261 ^ n2260 ^ n2068 ;
  assign n2263 = n740 & ~n1172 ;
  assign n2264 = n1802 ^ n514 ^ 1'b0 ;
  assign n2265 = n2264 ^ n990 ^ 1'b0 ;
  assign n2266 = ~n1013 & n2265 ;
  assign n2267 = n2266 ^ n1432 ^ x219 ;
  assign n2268 = ( n863 & n1328 ) | ( n863 & ~n2267 ) | ( n1328 & ~n2267 ) ;
  assign n2269 = n562 ^ x120 ^ 1'b0 ;
  assign n2270 = n1055 & n2269 ;
  assign n2271 = n1814 & n1853 ;
  assign n2272 = n2271 ^ n545 ^ 1'b0 ;
  assign n2273 = n1262 & n2272 ;
  assign n2274 = ~n1732 & n2273 ;
  assign n2275 = n1216 ^ n829 ^ n457 ;
  assign n2276 = x6 & ~n322 ;
  assign n2277 = n925 & n2276 ;
  assign n2278 = n2277 ^ n1131 ^ 1'b0 ;
  assign n2279 = n1523 ^ n1047 ^ n323 ;
  assign n2280 = ~n1880 & n2279 ;
  assign n2281 = n2280 ^ n1545 ^ 1'b0 ;
  assign n2282 = n2278 & ~n2281 ;
  assign n2283 = n2242 ^ n1468 ^ 1'b0 ;
  assign n2284 = ( x157 & n2038 ) | ( x157 & ~n2283 ) | ( n2038 & ~n2283 ) ;
  assign n2285 = n308 & ~n1367 ;
  assign n2286 = n1360 & n2285 ;
  assign n2287 = n2286 ^ n1978 ^ x129 ;
  assign n2292 = n1363 ^ n837 ^ 1'b0 ;
  assign n2293 = ( n1402 & n1877 ) | ( n1402 & n2292 ) | ( n1877 & n2292 ) ;
  assign n2288 = x49 & n495 ;
  assign n2289 = ~n428 & n2288 ;
  assign n2290 = n2289 ^ n847 ^ x77 ;
  assign n2291 = x198 | n2290 ;
  assign n2294 = n2293 ^ n2291 ^ 1'b0 ;
  assign n2295 = n2294 ^ n1934 ^ n1780 ;
  assign n2301 = ~x82 & n986 ;
  assign n2297 = n821 ^ n401 ^ 1'b0 ;
  assign n2296 = ~n468 & n920 ;
  assign n2298 = n2297 ^ n2296 ^ 1'b0 ;
  assign n2299 = ~n1447 & n2298 ;
  assign n2300 = n287 & n2299 ;
  assign n2302 = n2301 ^ n2300 ^ 1'b0 ;
  assign n2303 = n968 & n1201 ;
  assign n2304 = n2303 ^ n1757 ^ 1'b0 ;
  assign n2305 = n1521 ^ n1478 ^ 1'b0 ;
  assign n2306 = n1269 ^ n1257 ^ 1'b0 ;
  assign n2307 = ( n1377 & n1970 ) | ( n1377 & n2306 ) | ( n1970 & n2306 ) ;
  assign n2308 = n1025 ^ n915 ^ 1'b0 ;
  assign n2313 = ( n1289 & n1537 ) | ( n1289 & ~n2036 ) | ( n1537 & ~n2036 ) ;
  assign n2309 = x250 & ~n684 ;
  assign n2310 = n2309 ^ n403 ^ 1'b0 ;
  assign n2311 = n2310 ^ n835 ^ n752 ;
  assign n2312 = n1308 & ~n2311 ;
  assign n2314 = n2313 ^ n2312 ^ n1257 ;
  assign n2315 = n1891 ^ x142 ^ x8 ;
  assign n2316 = n2220 | n2315 ;
  assign n2317 = n1674 & ~n2316 ;
  assign n2318 = n1804 ^ x46 ^ 1'b0 ;
  assign n2319 = n1018 & ~n2318 ;
  assign n2320 = n1272 ^ n623 ^ 1'b0 ;
  assign n2321 = n1962 & n2320 ;
  assign n2322 = x238 & n794 ;
  assign n2323 = n2322 ^ n852 ^ 1'b0 ;
  assign n2324 = n2323 ^ n533 ^ 1'b0 ;
  assign n2325 = n1424 & n2324 ;
  assign n2326 = n2325 ^ n318 ^ x56 ;
  assign n2327 = n2326 ^ n932 ^ 1'b0 ;
  assign n2328 = n2321 & n2327 ;
  assign n2329 = n1463 ^ n741 ^ x23 ;
  assign n2330 = x209 | n520 ;
  assign n2331 = n2330 ^ x207 ^ 1'b0 ;
  assign n2332 = n1723 & n2205 ;
  assign n2333 = n2099 ^ n487 ^ 1'b0 ;
  assign n2334 = n1025 | n1561 ;
  assign n2335 = n2334 ^ n992 ^ 1'b0 ;
  assign n2336 = x187 & ~n2335 ;
  assign n2337 = n571 & ~n1252 ;
  assign n2338 = n840 & n2337 ;
  assign n2339 = n2338 ^ n574 ^ 1'b0 ;
  assign n2340 = ~n396 & n2339 ;
  assign n2341 = n1675 ^ n665 ^ 1'b0 ;
  assign n2342 = n1172 ^ n697 ^ n256 ;
  assign n2343 = n645 & n1154 ;
  assign n2344 = n750 & n2343 ;
  assign n2345 = x191 & x201 ;
  assign n2346 = n1803 & n2345 ;
  assign n2347 = n1772 & ~n2174 ;
  assign n2348 = x186 ^ x64 ^ 1'b0 ;
  assign n2349 = n2348 ^ n333 ^ 1'b0 ;
  assign n2350 = ( n783 & ~n2294 ) | ( n783 & n2349 ) | ( ~n2294 & n2349 ) ;
  assign n2351 = n479 ^ x27 ^ 1'b0 ;
  assign n2352 = n277 & n2351 ;
  assign n2353 = n939 | n1090 ;
  assign n2354 = n795 & ~n2353 ;
  assign n2355 = n872 & n1965 ;
  assign n2356 = n2355 ^ n814 ^ n678 ;
  assign n2357 = ( n522 & n587 ) | ( n522 & ~n1550 ) | ( n587 & ~n1550 ) ;
  assign n2358 = n1806 | n2313 ;
  assign n2359 = n866 ^ n631 ^ 1'b0 ;
  assign n2360 = x222 ^ x159 ^ 1'b0 ;
  assign n2361 = n1820 ^ n440 ^ 1'b0 ;
  assign n2362 = n2360 & n2361 ;
  assign n2363 = n898 & n1031 ;
  assign n2364 = n1820 ^ n1032 ^ 1'b0 ;
  assign n2365 = n747 & n2364 ;
  assign n2366 = n600 & ~n642 ;
  assign n2367 = n2366 ^ n1632 ^ 1'b0 ;
  assign n2368 = n2365 & n2367 ;
  assign n2369 = n2368 ^ n2066 ^ 1'b0 ;
  assign n2370 = ( x182 & n468 ) | ( x182 & n476 ) | ( n468 & n476 ) ;
  assign n2371 = n2370 ^ n733 ^ 1'b0 ;
  assign n2372 = ~n1356 & n2371 ;
  assign n2373 = ~n783 & n2372 ;
  assign n2374 = x43 & ~n1064 ;
  assign n2375 = n671 & n1620 ;
  assign n2376 = n970 ^ n678 ^ 1'b0 ;
  assign n2377 = n2376 ^ n2256 ^ 1'b0 ;
  assign n2378 = ~n1136 & n2377 ;
  assign n2379 = n2378 ^ n2248 ^ n750 ;
  assign n2380 = n1547 ^ n850 ^ 1'b0 ;
  assign n2381 = n2379 | n2380 ;
  assign n2382 = n1653 ^ n1603 ^ 1'b0 ;
  assign n2383 = ~n525 & n2382 ;
  assign n2384 = n2383 ^ n1051 ^ 1'b0 ;
  assign n2385 = n2381 | n2384 ;
  assign n2386 = n1176 | n1658 ;
  assign n2387 = n877 ^ n549 ^ 1'b0 ;
  assign n2388 = n2387 ^ n691 ^ 1'b0 ;
  assign n2389 = n675 & ~n2388 ;
  assign n2390 = n1545 | n1564 ;
  assign n2391 = n511 ^ x202 ^ x176 ;
  assign n2393 = n2301 ^ n1298 ^ 1'b0 ;
  assign n2394 = n2024 | n2393 ;
  assign n2392 = n1058 & ~n1257 ;
  assign n2395 = n2394 ^ n2392 ^ 1'b0 ;
  assign n2396 = n2304 & ~n2395 ;
  assign n2397 = n2261 & ~n2387 ;
  assign n2403 = n2301 ^ n1611 ^ n327 ;
  assign n2404 = ~n358 & n2403 ;
  assign n2405 = n2404 ^ n1022 ^ 1'b0 ;
  assign n2398 = n625 & ~n1600 ;
  assign n2399 = n694 & n2398 ;
  assign n2400 = n1389 ^ x156 ^ 1'b0 ;
  assign n2401 = n1970 & n2400 ;
  assign n2402 = ~n2399 & n2401 ;
  assign n2406 = n2405 ^ n2402 ^ 1'b0 ;
  assign n2407 = n1308 ^ n1168 ^ 1'b0 ;
  assign n2408 = n961 & ~n1131 ;
  assign n2409 = ( n829 & n994 ) | ( n829 & ~n2408 ) | ( n994 & ~n2408 ) ;
  assign n2410 = x129 & n2367 ;
  assign n2411 = n2410 ^ n1671 ^ 1'b0 ;
  assign n2417 = n809 | n2047 ;
  assign n2418 = n1275 | n2417 ;
  assign n2415 = x119 & ~n338 ;
  assign n2416 = n2415 ^ n686 ^ 1'b0 ;
  assign n2419 = n2418 ^ n2416 ^ x75 ;
  assign n2412 = n1302 ^ n902 ^ x124 ;
  assign n2413 = ~n1131 & n2412 ;
  assign n2414 = n2413 ^ n302 ^ 1'b0 ;
  assign n2420 = n2419 ^ n2414 ^ 1'b0 ;
  assign n2421 = n2370 | n2420 ;
  assign n2422 = n1351 ^ n1216 ^ 1'b0 ;
  assign n2423 = n2422 ^ n2397 ^ x218 ;
  assign n2424 = x28 & ~n1504 ;
  assign n2425 = n665 & n2424 ;
  assign n2426 = n1690 | n2425 ;
  assign n2427 = ~n668 & n2426 ;
  assign n2428 = x167 & n952 ;
  assign n2429 = n2428 ^ x254 ^ 1'b0 ;
  assign n2430 = n2429 ^ n1156 ^ n1039 ;
  assign n2431 = n1858 | n2430 ;
  assign n2432 = n827 & n1647 ;
  assign n2433 = n1062 & n2432 ;
  assign n2436 = x35 & x97 ;
  assign n2437 = n2436 ^ n979 ^ 1'b0 ;
  assign n2434 = x247 & ~n259 ;
  assign n2435 = n2434 ^ n1644 ^ 1'b0 ;
  assign n2438 = n2437 ^ n2435 ^ 1'b0 ;
  assign n2439 = ~n2019 & n2438 ;
  assign n2440 = ( ~n2406 & n2433 ) | ( ~n2406 & n2439 ) | ( n2433 & n2439 ) ;
  assign n2441 = n1004 ^ x136 ^ 1'b0 ;
  assign n2442 = n1154 & ~n2441 ;
  assign n2443 = ~n1416 & n2442 ;
  assign n2444 = n2443 ^ n559 ^ n436 ;
  assign n2445 = ( n1005 & n1374 ) | ( n1005 & n2444 ) | ( n1374 & n2444 ) ;
  assign n2446 = ~n293 & n671 ;
  assign n2447 = n2446 ^ n1024 ^ 1'b0 ;
  assign n2448 = x248 ^ x1 ^ 1'b0 ;
  assign n2449 = n2448 ^ n2372 ^ n1812 ;
  assign n2450 = ( n454 & ~n2447 ) | ( n454 & n2449 ) | ( ~n2447 & n2449 ) ;
  assign n2451 = ~n710 & n1149 ;
  assign n2452 = ( x245 & n525 ) | ( x245 & ~n1174 ) | ( n525 & ~n1174 ) ;
  assign n2453 = n485 & n2452 ;
  assign n2454 = n2453 ^ n363 ^ 1'b0 ;
  assign n2455 = n1232 ^ n933 ^ 1'b0 ;
  assign n2456 = n616 & ~n2455 ;
  assign n2457 = n260 ^ x115 ^ 1'b0 ;
  assign n2458 = n2456 & ~n2457 ;
  assign n2459 = n2370 ^ x118 ^ 1'b0 ;
  assign n2460 = n369 | n2459 ;
  assign n2461 = x150 | n2460 ;
  assign n2462 = ( x207 & ~n2458 ) | ( x207 & n2461 ) | ( ~n2458 & n2461 ) ;
  assign n2463 = ( ~n1162 & n2454 ) | ( ~n1162 & n2462 ) | ( n2454 & n2462 ) ;
  assign n2464 = ( ~n417 & n993 ) | ( ~n417 & n2441 ) | ( n993 & n2441 ) ;
  assign n2465 = n2464 ^ n1579 ^ n1460 ;
  assign n2466 = ( x107 & n615 ) | ( x107 & ~n1178 ) | ( n615 & ~n1178 ) ;
  assign n2467 = n1873 & ~n2466 ;
  assign n2468 = n2467 ^ n2054 ^ 1'b0 ;
  assign n2469 = n2468 ^ n2435 ^ 1'b0 ;
  assign n2470 = n459 ^ x209 ^ 1'b0 ;
  assign n2471 = n992 | n2470 ;
  assign n2472 = n1329 & n2471 ;
  assign n2473 = ( n544 & n1713 ) | ( n544 & ~n2351 ) | ( n1713 & ~n2351 ) ;
  assign n2474 = n655 ^ n329 ^ 1'b0 ;
  assign n2475 = x198 & n2474 ;
  assign n2476 = n680 & ~n2475 ;
  assign n2477 = n1173 & n2476 ;
  assign n2478 = n2477 ^ n1838 ^ 1'b0 ;
  assign n2479 = ( x246 & ~n993 ) | ( x246 & n2128 ) | ( ~n993 & n2128 ) ;
  assign n2482 = x171 & n1559 ;
  assign n2480 = x78 & n953 ;
  assign n2481 = n831 & n2480 ;
  assign n2483 = n2482 ^ n2481 ^ 1'b0 ;
  assign n2484 = n1021 | n2483 ;
  assign n2485 = n715 & n1208 ;
  assign n2486 = ~n1225 & n2485 ;
  assign n2487 = n1567 ^ n941 ^ n843 ;
  assign n2488 = x42 & n2487 ;
  assign n2489 = ( n472 & ~n927 ) | ( n472 & n1048 ) | ( ~n927 & n1048 ) ;
  assign n2490 = ( n589 & n2488 ) | ( n589 & ~n2489 ) | ( n2488 & ~n2489 ) ;
  assign n2491 = n2490 ^ x158 ^ x15 ;
  assign n2492 = n2491 ^ n2376 ^ 1'b0 ;
  assign n2493 = n457 & ~n2492 ;
  assign n2494 = n1356 ^ n701 ^ 1'b0 ;
  assign n2495 = n514 ^ x12 ^ 1'b0 ;
  assign n2496 = x154 & n2495 ;
  assign n2497 = n2496 ^ n1846 ^ 1'b0 ;
  assign n2498 = n1243 & ~n2497 ;
  assign n2499 = n2067 ^ n1582 ^ n795 ;
  assign n2500 = n1383 ^ n645 ^ 1'b0 ;
  assign n2503 = x199 & n1000 ;
  assign n2504 = n287 & n2503 ;
  assign n2505 = n2504 ^ n1380 ^ n1113 ;
  assign n2501 = n848 ^ x239 ^ 1'b0 ;
  assign n2502 = n478 | n2501 ;
  assign n2506 = n2505 ^ n2502 ^ n303 ;
  assign n2512 = ~n317 & n599 ;
  assign n2513 = n2370 & n2512 ;
  assign n2507 = ( ~x58 & n1013 ) | ( ~x58 & n1116 ) | ( n1013 & n1116 ) ;
  assign n2508 = x163 & ~n2507 ;
  assign n2509 = n286 & n2508 ;
  assign n2510 = n2509 ^ n1440 ^ 1'b0 ;
  assign n2511 = n2510 ^ n2294 ^ n818 ;
  assign n2514 = n2513 ^ n2511 ^ 1'b0 ;
  assign n2515 = ~n2443 & n2514 ;
  assign n2516 = n2372 ^ n1044 ^ 1'b0 ;
  assign n2522 = n870 ^ x155 ^ x27 ;
  assign n2523 = n1615 & ~n2522 ;
  assign n2521 = n481 & n990 ;
  assign n2524 = n2523 ^ n2521 ^ 1'b0 ;
  assign n2517 = x37 & ~x201 ;
  assign n2518 = ( n589 & ~n990 ) | ( n589 & n2126 ) | ( ~n990 & n2126 ) ;
  assign n2519 = n2517 & ~n2518 ;
  assign n2520 = n860 & n2519 ;
  assign n2525 = n2524 ^ n2520 ^ 1'b0 ;
  assign n2526 = n675 | n2525 ;
  assign n2527 = n1220 ^ n897 ^ n451 ;
  assign n2528 = ~n493 & n627 ;
  assign n2529 = n2528 ^ n773 ^ 1'b0 ;
  assign n2530 = n2496 ^ n671 ^ 1'b0 ;
  assign n2531 = n993 & n2530 ;
  assign n2532 = ( n704 & n1160 ) | ( n704 & ~n2531 ) | ( n1160 & ~n2531 ) ;
  assign n2533 = n516 & n2532 ;
  assign n2534 = n2529 & n2533 ;
  assign n2535 = ~n403 & n1472 ;
  assign n2536 = n1501 & n2535 ;
  assign n2537 = n2117 & ~n2536 ;
  assign n2538 = n334 & n2537 ;
  assign n2539 = ( x239 & n925 ) | ( x239 & ~n2045 ) | ( n925 & ~n2045 ) ;
  assign n2540 = n2539 ^ n362 ^ 1'b0 ;
  assign n2541 = n970 | n2540 ;
  assign n2542 = n2389 ^ n2339 ^ 1'b0 ;
  assign n2545 = ~n259 & n953 ;
  assign n2546 = n729 & n2545 ;
  assign n2547 = n2546 ^ n1843 ^ n513 ;
  assign n2543 = n1267 ^ n1071 ^ 1'b0 ;
  assign n2544 = ~n1908 & n2543 ;
  assign n2548 = n2547 ^ n2544 ^ 1'b0 ;
  assign n2549 = ( n623 & ~n1794 ) | ( n623 & n2119 ) | ( ~n1794 & n2119 ) ;
  assign n2550 = n1108 ^ n338 ^ 1'b0 ;
  assign n2551 = x206 & n2550 ;
  assign n2552 = ~n668 & n2551 ;
  assign n2553 = n468 & n2552 ;
  assign n2554 = ~n736 & n1789 ;
  assign n2555 = n2553 & n2554 ;
  assign n2556 = x70 & ~n286 ;
  assign n2557 = n2556 ^ x232 ^ 1'b0 ;
  assign n2558 = n2557 ^ n2370 ^ n901 ;
  assign n2559 = ~n338 & n2558 ;
  assign n2560 = n377 & n2559 ;
  assign n2561 = n399 ^ x47 ^ 1'b0 ;
  assign n2562 = ~n515 & n2561 ;
  assign n2563 = n1309 ^ n1022 ^ n671 ;
  assign n2564 = n2562 & ~n2563 ;
  assign n2565 = n2560 & n2564 ;
  assign n2566 = n2453 ^ n1252 ^ n888 ;
  assign n2567 = n402 | n2566 ;
  assign n2568 = n2567 ^ n474 ^ n338 ;
  assign n2569 = n326 | n1047 ;
  assign n2570 = n820 & ~n2569 ;
  assign n2571 = ~x7 & x70 ;
  assign n2572 = n2571 ^ n1206 ^ n351 ;
  assign n2573 = ~n2570 & n2572 ;
  assign n2574 = n1534 & n2017 ;
  assign n2575 = ( n441 & n447 ) | ( n441 & n803 ) | ( n447 & n803 ) ;
  assign n2576 = ~n1350 & n2575 ;
  assign n2577 = n2574 & n2576 ;
  assign n2578 = n2427 ^ n1830 ^ 1'b0 ;
  assign n2579 = x43 & ~n1442 ;
  assign n2580 = n2579 ^ n547 ^ 1'b0 ;
  assign n2584 = n280 & n1639 ;
  assign n2581 = n1761 ^ x215 ^ 1'b0 ;
  assign n2582 = n1270 & n2581 ;
  assign n2583 = n2582 ^ n1948 ^ n964 ;
  assign n2585 = n2584 ^ n2583 ^ n1176 ;
  assign n2586 = n1091 & n1185 ;
  assign n2589 = n562 & ~n2021 ;
  assign n2587 = ~n1603 & n2030 ;
  assign n2588 = ~x125 & n2587 ;
  assign n2590 = n2589 ^ n2588 ^ n1503 ;
  assign n2591 = x161 & ~n2507 ;
  assign n2592 = n2591 ^ n1324 ^ 1'b0 ;
  assign n2593 = ~n1133 & n1522 ;
  assign n2594 = n2593 ^ n1898 ^ 1'b0 ;
  assign n2595 = ( n1467 & ~n2592 ) | ( n1467 & n2594 ) | ( ~n2592 & n2594 ) ;
  assign n2596 = n769 ^ n396 ^ 1'b0 ;
  assign n2597 = x51 & ~n2596 ;
  assign n2598 = ~n2426 & n2597 ;
  assign n2599 = ~n763 & n1873 ;
  assign n2600 = n2599 ^ n304 ^ 1'b0 ;
  assign n2601 = n2600 ^ n1322 ^ 1'b0 ;
  assign n2602 = n595 ^ n509 ^ 1'b0 ;
  assign n2603 = n318 & ~n2602 ;
  assign n2604 = n2603 ^ n1004 ^ 1'b0 ;
  assign n2605 = n2601 | n2604 ;
  assign n2606 = n2605 ^ n1877 ^ 1'b0 ;
  assign n2607 = n358 | n2606 ;
  assign n2608 = n649 | n1484 ;
  assign n2609 = ~n1010 & n1349 ;
  assign n2610 = ~n402 & n2609 ;
  assign n2611 = ( n874 & ~n1050 ) | ( n874 & n2610 ) | ( ~n1050 & n2610 ) ;
  assign n2612 = n2611 ^ n1399 ^ 1'b0 ;
  assign n2613 = n2608 & ~n2612 ;
  assign n2614 = ~n785 & n1571 ;
  assign n2615 = n1962 ^ n1650 ^ n1174 ;
  assign n2616 = ( n467 & n1116 ) | ( n467 & n2615 ) | ( n1116 & n2615 ) ;
  assign n2619 = x111 | n949 ;
  assign n2617 = n926 & ~n2422 ;
  assign n2618 = n2617 ^ n678 ^ 1'b0 ;
  assign n2620 = n2619 ^ n2618 ^ 1'b0 ;
  assign n2621 = n711 | n2620 ;
  assign n2622 = ( n467 & n522 ) | ( n467 & n967 ) | ( n522 & n967 ) ;
  assign n2623 = n2151 | n2622 ;
  assign n2624 = n2621 & ~n2623 ;
  assign n2625 = n2624 ^ x116 ^ 1'b0 ;
  assign n2626 = n1750 | n2625 ;
  assign n2627 = n2616 | n2626 ;
  assign n2628 = n1110 & ~n2627 ;
  assign n2632 = n327 & ~n545 ;
  assign n2633 = n1596 & n2632 ;
  assign n2629 = n679 ^ x240 ^ 1'b0 ;
  assign n2630 = ~n675 & n2629 ;
  assign n2631 = x140 & n2630 ;
  assign n2634 = n2633 ^ n2631 ^ 1'b0 ;
  assign n2635 = n522 & ~n2634 ;
  assign n2636 = ( n1603 & n2136 ) | ( n1603 & n2635 ) | ( n2136 & n2635 ) ;
  assign n2637 = n387 ^ x114 ^ 1'b0 ;
  assign n2638 = n2637 ^ n1877 ^ n1571 ;
  assign n2639 = ( n1618 & n1752 ) | ( n1618 & n2638 ) | ( n1752 & n2638 ) ;
  assign n2640 = ( n1200 & n2590 ) | ( n1200 & n2639 ) | ( n2590 & n2639 ) ;
  assign n2641 = n1291 ^ n763 ^ 1'b0 ;
  assign n2642 = x14 & ~n2641 ;
  assign n2643 = ( n1943 & ~n2025 ) | ( n1943 & n2642 ) | ( ~n2025 & n2642 ) ;
  assign n2644 = ( n363 & ~n574 ) | ( n363 & n1553 ) | ( ~n574 & n1553 ) ;
  assign n2645 = ~n2013 & n2644 ;
  assign n2646 = x51 & x125 ;
  assign n2647 = ~n2645 & n2646 ;
  assign n2648 = n2370 ^ n720 ^ x164 ;
  assign n2649 = n2648 ^ n1804 ^ 1'b0 ;
  assign n2650 = ~n2471 & n2649 ;
  assign n2651 = n1548 ^ n862 ^ 1'b0 ;
  assign n2652 = n1034 | n2651 ;
  assign n2653 = n2652 ^ n1540 ^ 1'b0 ;
  assign n2654 = ( x111 & ~n633 ) | ( x111 & n1309 ) | ( ~n633 & n1309 ) ;
  assign n2655 = n725 ^ x51 ^ 1'b0 ;
  assign n2656 = ~n507 & n2655 ;
  assign n2657 = ( ~n1202 & n1935 ) | ( ~n1202 & n2656 ) | ( n1935 & n2656 ) ;
  assign n2658 = n2657 ^ n1002 ^ x78 ;
  assign n2659 = n1107 ^ n806 ^ 1'b0 ;
  assign n2660 = n1425 | n2659 ;
  assign n2661 = ( x73 & ~n2648 ) | ( x73 & n2660 ) | ( ~n2648 & n2660 ) ;
  assign n2662 = n1430 & n2141 ;
  assign n2663 = ~n2085 & n2662 ;
  assign n2664 = n1617 | n2553 ;
  assign n2665 = n2664 ^ n1323 ^ 1'b0 ;
  assign n2666 = n2665 ^ n678 ^ 1'b0 ;
  assign n2667 = x70 & ~n2666 ;
  assign n2668 = ~n498 & n528 ;
  assign n2669 = ~n981 & n2668 ;
  assign n2670 = ( ~n303 & n990 ) | ( ~n303 & n2669 ) | ( n990 & n2669 ) ;
  assign n2671 = x73 | n509 ;
  assign n2672 = n1665 ^ n725 ^ 1'b0 ;
  assign n2674 = n873 ^ n835 ^ 1'b0 ;
  assign n2675 = n2674 ^ n1511 ^ 1'b0 ;
  assign n2673 = x169 & n1838 ;
  assign n2676 = n2675 ^ n2673 ^ 1'b0 ;
  assign n2677 = n1272 ^ n690 ^ n584 ;
  assign n2678 = n2677 ^ n1224 ^ n841 ;
  assign n2679 = ( x69 & x113 ) | ( x69 & ~n1082 ) | ( x113 & ~n1082 ) ;
  assign n2680 = n587 & n2679 ;
  assign n2681 = n2678 & ~n2680 ;
  assign n2682 = ~n2676 & n2681 ;
  assign n2683 = n982 & n2682 ;
  assign n2686 = ~n815 & n1158 ;
  assign n2687 = n2686 ^ n449 ^ 1'b0 ;
  assign n2684 = n931 & ~n1038 ;
  assign n2685 = n2684 ^ n617 ^ 1'b0 ;
  assign n2688 = n2687 ^ n2685 ^ n2571 ;
  assign n2689 = x250 & n2679 ;
  assign n2690 = n2689 ^ n2005 ^ 1'b0 ;
  assign n2691 = n1530 | n2690 ;
  assign n2692 = n1873 ^ n1228 ^ x6 ;
  assign n2693 = ~n1366 & n2692 ;
  assign n2694 = n2225 ^ n1715 ^ 1'b0 ;
  assign n2695 = n2541 | n2694 ;
  assign n2696 = ~n490 & n2383 ;
  assign n2697 = ~n1999 & n2696 ;
  assign n2698 = x217 & n266 ;
  assign n2699 = ~n2204 & n2698 ;
  assign n2700 = n1635 ^ n576 ^ 1'b0 ;
  assign n2701 = n2700 ^ n1775 ^ n1772 ;
  assign n2702 = n2699 | n2701 ;
  assign n2703 = n2121 ^ n256 ^ 1'b0 ;
  assign n2705 = x132 & ~n284 ;
  assign n2704 = n993 & ~n2126 ;
  assign n2706 = n2705 ^ n2704 ^ 1'b0 ;
  assign n2707 = n2706 ^ n671 ^ 1'b0 ;
  assign n2708 = n1615 | n2707 ;
  assign n2709 = n1410 ^ n1197 ^ x252 ;
  assign n2710 = ~n2061 & n2709 ;
  assign n2711 = n2710 ^ n347 ^ 1'b0 ;
  assign n2712 = n998 | n1517 ;
  assign n2713 = x171 & n1285 ;
  assign n2714 = n1508 | n2016 ;
  assign n2715 = ( n389 & n1304 ) | ( n389 & ~n1611 ) | ( n1304 & ~n1611 ) ;
  assign n2716 = n716 & ~n1374 ;
  assign n2717 = n2716 ^ n2259 ^ 1'b0 ;
  assign n2718 = x240 & n520 ;
  assign n2719 = ~n507 & n2718 ;
  assign n2720 = ~n2717 & n2719 ;
  assign n2721 = n1622 ^ n1360 ^ 1'b0 ;
  assign n2722 = n528 & ~n2243 ;
  assign n2723 = n2138 ^ n1077 ^ 1'b0 ;
  assign n2724 = n903 ^ x227 ^ 1'b0 ;
  assign n2725 = n870 & n1141 ;
  assign n2726 = n2724 & n2725 ;
  assign n2727 = n2726 ^ n2310 ^ n1299 ;
  assign n2728 = n2687 ^ n2577 ^ 1'b0 ;
  assign n2729 = n2172 & n2728 ;
  assign n2736 = n1719 ^ n922 ^ 1'b0 ;
  assign n2730 = n704 ^ n300 ^ x51 ;
  assign n2731 = ( x44 & ~n711 ) | ( x44 & n2730 ) | ( ~n711 & n2730 ) ;
  assign n2732 = n1622 & n2731 ;
  assign n2733 = n2732 ^ n850 ^ 1'b0 ;
  assign n2734 = x104 & ~n2733 ;
  assign n2735 = ( ~n1023 & n1682 ) | ( ~n1023 & n2734 ) | ( n1682 & n2734 ) ;
  assign n2737 = n2736 ^ n2735 ^ 1'b0 ;
  assign n2738 = n998 ^ n952 ^ n813 ;
  assign n2739 = x30 & n805 ;
  assign n2740 = n1805 & n2739 ;
  assign n2741 = n821 ^ x24 ^ 1'b0 ;
  assign n2742 = n2740 | n2741 ;
  assign n2743 = n2656 ^ x133 ^ 1'b0 ;
  assign n2744 = ~n2742 & n2743 ;
  assign n2745 = n2744 ^ n702 ^ 1'b0 ;
  assign n2746 = n1781 & n2745 ;
  assign n2747 = ~n2738 & n2746 ;
  assign n2748 = n2747 ^ n2500 ^ 1'b0 ;
  assign n2749 = n2035 & ~n2151 ;
  assign n2750 = ~n1776 & n2749 ;
  assign n2751 = n1474 ^ n1284 ^ 1'b0 ;
  assign n2752 = n790 & n2751 ;
  assign n2753 = ~n1106 & n2752 ;
  assign n2754 = n740 & n2753 ;
  assign n2755 = n752 & n2754 ;
  assign n2756 = n1187 ^ x34 ^ x9 ;
  assign n2757 = n1018 & ~n1353 ;
  assign n2758 = n2756 & n2757 ;
  assign n2759 = n2758 ^ n1232 ^ 1'b0 ;
  assign n2760 = ( n1727 & ~n1774 ) | ( n1727 & n2482 ) | ( ~n1774 & n2482 ) ;
  assign n2761 = n2760 ^ n1585 ^ 1'b0 ;
  assign n2762 = n2735 | n2761 ;
  assign n2763 = n2001 ^ n1289 ^ 1'b0 ;
  assign n2764 = ( n621 & ~n802 ) | ( n621 & n818 ) | ( ~n802 & n818 ) ;
  assign n2765 = n1962 & ~n2764 ;
  assign n2766 = ~n2763 & n2765 ;
  assign n2767 = n686 | n1615 ;
  assign n2768 = n1821 ^ n877 ^ 1'b0 ;
  assign n2769 = x109 & n2768 ;
  assign n2770 = ( n297 & ~n722 ) | ( n297 & n2769 ) | ( ~n722 & n2769 ) ;
  assign n2771 = n371 & ~n2770 ;
  assign n2772 = ( n1324 & n2767 ) | ( n1324 & n2771 ) | ( n2767 & n2771 ) ;
  assign n2773 = n2439 & ~n2772 ;
  assign n2774 = n2773 ^ n584 ^ 1'b0 ;
  assign n2775 = n1395 ^ n1309 ^ 1'b0 ;
  assign n2776 = n974 & n2775 ;
  assign n2777 = n2776 ^ n394 ^ 1'b0 ;
  assign n2778 = n509 ^ x83 ^ 1'b0 ;
  assign n2779 = x34 & ~n2221 ;
  assign n2780 = n752 | n1689 ;
  assign n2781 = ~n956 & n2780 ;
  assign n2782 = ( x80 & n1232 ) | ( x80 & ~n1605 ) | ( n1232 & ~n1605 ) ;
  assign n2786 = ~x209 & n884 ;
  assign n2783 = ( ~n1116 & n1734 ) | ( ~n1116 & n2110 ) | ( n1734 & n2110 ) ;
  assign n2784 = ( x24 & n2441 ) | ( x24 & ~n2783 ) | ( n2441 & ~n2783 ) ;
  assign n2785 = x95 & n2784 ;
  assign n2787 = n2786 ^ n2785 ^ 1'b0 ;
  assign n2788 = ( n2520 & ~n2782 ) | ( n2520 & n2787 ) | ( ~n2782 & n2787 ) ;
  assign n2789 = x58 & x242 ;
  assign n2790 = n2789 ^ x87 ^ 1'b0 ;
  assign n2791 = ( x217 & n847 ) | ( x217 & n2790 ) | ( n847 & n2790 ) ;
  assign n2792 = x171 & x254 ;
  assign n2793 = n2792 ^ n407 ^ 1'b0 ;
  assign n2794 = n1667 & n2793 ;
  assign n2797 = x56 & n462 ;
  assign n2798 = n2797 ^ n1372 ^ 1'b0 ;
  assign n2799 = n2798 ^ n1969 ^ x156 ;
  assign n2795 = n1394 & n2634 ;
  assign n2796 = n2795 ^ n736 ^ 1'b0 ;
  assign n2800 = n2799 ^ n2796 ^ n1569 ;
  assign n2801 = x54 & ~n750 ;
  assign n2802 = n1425 & n2801 ;
  assign n2803 = n629 ^ x98 ^ 1'b0 ;
  assign n2804 = n2802 | n2803 ;
  assign n2805 = n723 ^ x156 ^ 1'b0 ;
  assign n2806 = x246 & n2805 ;
  assign n2807 = n1385 | n2806 ;
  assign n2808 = x235 & ~n1022 ;
  assign n2809 = n2637 ^ x77 ^ 1'b0 ;
  assign n2810 = n2809 ^ n2639 ^ 1'b0 ;
  assign n2811 = n2808 & ~n2810 ;
  assign n2812 = ( ~n445 & n2529 ) | ( ~n445 & n2811 ) | ( n2529 & n2811 ) ;
  assign n2813 = x146 & n586 ;
  assign n2814 = n2813 ^ n1999 ^ 1'b0 ;
  assign n2815 = n333 | n2814 ;
  assign n2816 = n952 | n2815 ;
  assign n2817 = n2816 ^ n2702 ^ n591 ;
  assign n2818 = ~n944 & n1420 ;
  assign n2826 = n1007 ^ n600 ^ 1'b0 ;
  assign n2824 = ( x134 & x227 ) | ( x134 & n343 ) | ( x227 & n343 ) ;
  assign n2822 = n1774 ^ n1182 ^ 1'b0 ;
  assign n2821 = n1817 ^ n1604 ^ n1353 ;
  assign n2820 = ~n1148 & n1179 ;
  assign n2823 = n2822 ^ n2821 ^ n2820 ;
  assign n2819 = n2601 ^ n1592 ^ 1'b0 ;
  assign n2825 = n2824 ^ n2823 ^ n2819 ;
  assign n2827 = n2826 ^ n2825 ^ n1328 ;
  assign n2828 = n2401 & ~n2577 ;
  assign n2829 = x74 & x107 ;
  assign n2830 = n2829 ^ n312 ^ 1'b0 ;
  assign n2831 = x91 & ~n1658 ;
  assign n2832 = n1197 & n2678 ;
  assign n2834 = x100 & n599 ;
  assign n2835 = ~x160 & n2834 ;
  assign n2833 = n1382 ^ n343 ^ 1'b0 ;
  assign n2836 = n2835 ^ n2833 ^ 1'b0 ;
  assign n2837 = n811 ^ n677 ^ x142 ;
  assign n2838 = ( ~n1200 & n1644 ) | ( ~n1200 & n2118 ) | ( n1644 & n2118 ) ;
  assign n2839 = n617 & ~n2838 ;
  assign n2840 = n1504 & n2839 ;
  assign n2841 = n593 & n2840 ;
  assign n2844 = n1236 & n2299 ;
  assign n2842 = n1063 & n1479 ;
  assign n2843 = n2842 ^ n1405 ^ 1'b0 ;
  assign n2845 = n2844 ^ n2843 ^ n441 ;
  assign n2846 = n658 ^ n575 ^ 1'b0 ;
  assign n2847 = n1865 ^ n593 ^ 1'b0 ;
  assign n2848 = x6 & ~n2847 ;
  assign n2849 = n2848 ^ x26 ^ 1'b0 ;
  assign n2850 = n1727 ^ n1711 ^ 1'b0 ;
  assign n2851 = n891 ^ n885 ^ x192 ;
  assign n2852 = n2851 ^ n1231 ^ 1'b0 ;
  assign n2853 = n2852 ^ n2769 ^ 1'b0 ;
  assign n2854 = ( x103 & n415 ) | ( x103 & ~n2268 ) | ( n415 & ~n2268 ) ;
  assign n2855 = x5 & ~n2513 ;
  assign n2856 = n2855 ^ x146 ^ 1'b0 ;
  assign n2857 = n2856 ^ n596 ^ 1'b0 ;
  assign n2858 = n1729 & n2510 ;
  assign n2859 = ~x178 & n2858 ;
  assign n2860 = n1717 ^ n1352 ^ x239 ;
  assign n2861 = n2859 | n2860 ;
  assign n2862 = n2645 ^ n454 ^ 1'b0 ;
  assign n2863 = ~n554 & n2862 ;
  assign n2864 = n1327 | n1576 ;
  assign n2865 = n2864 ^ x198 ^ 1'b0 ;
  assign n2870 = n701 & ~n947 ;
  assign n2871 = n2870 ^ n1273 ^ 1'b0 ;
  assign n2872 = n2679 & n2871 ;
  assign n2873 = n2872 ^ n544 ^ 1'b0 ;
  assign n2866 = n673 ^ n630 ^ 1'b0 ;
  assign n2867 = n1152 & ~n2866 ;
  assign n2868 = n549 | n2867 ;
  assign n2869 = x149 & n2868 ;
  assign n2874 = n2873 ^ n2869 ^ 1'b0 ;
  assign n2877 = x202 | n1746 ;
  assign n2875 = x89 & ~n1067 ;
  assign n2876 = n1543 & n2875 ;
  assign n2878 = n2877 ^ n2876 ^ 1'b0 ;
  assign n2879 = ~n2447 & n2878 ;
  assign n2880 = n327 & ~n2679 ;
  assign n2881 = ~n1744 & n1780 ;
  assign n2882 = n2174 & n2881 ;
  assign n2883 = ~n2880 & n2882 ;
  assign n2884 = n1286 ^ n317 ^ 1'b0 ;
  assign n2885 = n1784 ^ n623 ^ 1'b0 ;
  assign n2886 = n2884 | n2885 ;
  assign n2887 = ( n763 & n1380 ) | ( n763 & ~n2699 ) | ( n1380 & ~n2699 ) ;
  assign n2889 = x183 & ~n1472 ;
  assign n2890 = n2889 ^ n287 ^ 1'b0 ;
  assign n2891 = n2890 ^ n1989 ^ n407 ;
  assign n2892 = n1350 & n2891 ;
  assign n2888 = ( x58 & n1552 ) | ( x58 & ~n2229 ) | ( n1552 & ~n2229 ) ;
  assign n2893 = n2892 ^ n2888 ^ 1'b0 ;
  assign n2896 = n386 & n959 ;
  assign n2897 = ~x15 & n2896 ;
  assign n2894 = n1179 ^ n464 ^ x153 ;
  assign n2895 = ( n1966 & n2140 ) | ( n1966 & n2894 ) | ( n2140 & n2894 ) ;
  assign n2898 = n2897 ^ n2895 ^ 1'b0 ;
  assign n2899 = ~n2338 & n2898 ;
  assign n2900 = n1452 ^ n1134 ^ 1'b0 ;
  assign n2901 = n479 & n2900 ;
  assign n2902 = n2901 ^ n2615 ^ 1'b0 ;
  assign n2903 = ~n1816 & n2902 ;
  assign n2904 = n2903 ^ n1579 ^ x159 ;
  assign n2905 = ~n1722 & n2904 ;
  assign n2906 = ~n2899 & n2905 ;
  assign n2907 = n2370 ^ n314 ^ 1'b0 ;
  assign n2908 = ( n440 & ~n1661 ) | ( n440 & n2907 ) | ( ~n1661 & n2907 ) ;
  assign n2909 = ~n1930 & n2908 ;
  assign n2910 = ( ~n1907 & n2174 ) | ( ~n1907 & n2610 ) | ( n2174 & n2610 ) ;
  assign n2911 = n2468 ^ n1451 ^ n656 ;
  assign n2912 = ( x105 & n1100 ) | ( x105 & n1423 ) | ( n1100 & n1423 ) ;
  assign n2913 = x120 & ~n1118 ;
  assign n2914 = n2913 ^ x50 ^ 1'b0 ;
  assign n2915 = n2912 | n2914 ;
  assign n2916 = n1723 ^ n423 ^ 1'b0 ;
  assign n2917 = ( n1222 & n2915 ) | ( n1222 & n2916 ) | ( n2915 & n2916 ) ;
  assign n2918 = n1090 & n1605 ;
  assign n2919 = n2918 ^ n2155 ^ 1'b0 ;
  assign n2920 = n2041 | n2919 ;
  assign n2921 = n2920 ^ n591 ^ 1'b0 ;
  assign n2922 = n2921 ^ n1415 ^ 1'b0 ;
  assign n2923 = n2705 ^ x154 ^ 1'b0 ;
  assign n2924 = x121 & n2923 ;
  assign n2925 = ( x57 & n2378 ) | ( x57 & n2775 ) | ( n2378 & n2775 ) ;
  assign n2926 = n2925 ^ n926 ^ 1'b0 ;
  assign n2927 = n2924 & n2926 ;
  assign n2928 = x17 & ~n1562 ;
  assign n2929 = n2928 ^ n457 ^ 1'b0 ;
  assign n2930 = n981 & ~n2929 ;
  assign n2931 = n2930 ^ x55 ^ 1'b0 ;
  assign n2932 = ( ~n720 & n1728 ) | ( ~n720 & n2931 ) | ( n1728 & n2931 ) ;
  assign n2933 = ~n2441 & n2932 ;
  assign n2934 = n2933 ^ n973 ^ 1'b0 ;
  assign n2935 = x116 & x216 ;
  assign n2936 = n2935 ^ x14 ^ 1'b0 ;
  assign n2937 = n2936 ^ x91 ^ 1'b0 ;
  assign n2938 = n1644 ^ x135 ^ 1'b0 ;
  assign n2939 = n715 & n1995 ;
  assign n2940 = n1496 ^ n1423 ^ x161 ;
  assign n2941 = n2939 & ~n2940 ;
  assign n2942 = n2941 ^ n2107 ^ 1'b0 ;
  assign n2943 = n2942 ^ n2179 ^ n921 ;
  assign n2945 = ~x2 & n1970 ;
  assign n2944 = n1672 | n2118 ;
  assign n2946 = n2945 ^ n2944 ^ 1'b0 ;
  assign n2947 = x68 & n1860 ;
  assign n2948 = n2947 ^ n1956 ^ 1'b0 ;
  assign n2949 = n768 & ~n1505 ;
  assign n2950 = ~n2006 & n2949 ;
  assign n2951 = n1213 & ~n2950 ;
  assign n2952 = x122 & x228 ;
  assign n2953 = n2952 ^ x216 ^ 1'b0 ;
  assign n2954 = ~n1890 & n2953 ;
  assign n2955 = n1022 & ~n1047 ;
  assign n2956 = n468 ^ x188 ^ 1'b0 ;
  assign n2957 = n2955 & ~n2956 ;
  assign n2958 = n2957 ^ n1231 ^ 1'b0 ;
  assign n2959 = n978 | n2958 ;
  assign n2961 = n268 & n805 ;
  assign n2960 = ~n1685 & n2871 ;
  assign n2962 = n2961 ^ n2960 ^ 1'b0 ;
  assign n2966 = n561 & ~n2100 ;
  assign n2963 = n1175 & n2448 ;
  assign n2964 = n2963 ^ n971 ^ 1'b0 ;
  assign n2965 = n1965 & ~n2964 ;
  assign n2967 = n2966 ^ n2965 ^ 1'b0 ;
  assign n2968 = x195 & n1998 ;
  assign n2971 = n1579 ^ n904 ^ 1'b0 ;
  assign n2969 = n2892 ^ n1538 ^ 1'b0 ;
  assign n2970 = n1667 & ~n2969 ;
  assign n2972 = n2971 ^ n2970 ^ 1'b0 ;
  assign n2977 = n2019 ^ n1702 ^ n260 ;
  assign n2975 = n1150 ^ n549 ^ 1'b0 ;
  assign n2976 = ~n500 & n2975 ;
  assign n2973 = n559 | n1211 ;
  assign n2974 = n2973 ^ n1696 ^ 1'b0 ;
  assign n2978 = n2977 ^ n2976 ^ n2974 ;
  assign n2979 = x199 & ~n2727 ;
  assign n2980 = n1922 & n2979 ;
  assign n2982 = n614 ^ x164 ^ 1'b0 ;
  assign n2983 = ~n699 & n2982 ;
  assign n2984 = ( n1082 & n1258 ) | ( n1082 & ~n2983 ) | ( n1258 & ~n2983 ) ;
  assign n2981 = x86 & n966 ;
  assign n2985 = n2984 ^ n2981 ^ 1'b0 ;
  assign n2986 = x77 & n335 ;
  assign n2987 = n2986 ^ n2522 ^ n363 ;
  assign n2988 = ~n619 & n2987 ;
  assign n2989 = n349 & n2988 ;
  assign n2990 = n2989 ^ n1671 ^ x113 ;
  assign n2991 = n438 ^ x177 ^ x23 ;
  assign n2992 = x145 & ~n2991 ;
  assign n2993 = ( ~n2257 & n2571 ) | ( ~n2257 & n2992 ) | ( n2571 & n2992 ) ;
  assign n2994 = n314 | n386 ;
  assign n2995 = ( x230 & ~n1909 ) | ( x230 & n2994 ) | ( ~n1909 & n2994 ) ;
  assign n2996 = n409 | n2995 ;
  assign n2997 = ~x125 & n2996 ;
  assign n2998 = ( n1164 & ~n1592 ) | ( n1164 & n1703 ) | ( ~n1592 & n1703 ) ;
  assign n2999 = x150 & ~n1597 ;
  assign n3000 = n2999 ^ n2680 ^ 1'b0 ;
  assign n3004 = ( n305 & ~n384 ) | ( n305 & n1208 ) | ( ~n384 & n1208 ) ;
  assign n3003 = n318 & n434 ;
  assign n3005 = n3004 ^ n3003 ^ 1'b0 ;
  assign n3006 = n1484 & ~n3005 ;
  assign n3007 = n1978 & n3006 ;
  assign n3001 = n2585 ^ n2216 ^ 1'b0 ;
  assign n3002 = ~n2275 & n3001 ;
  assign n3008 = n3007 ^ n3002 ^ 1'b0 ;
  assign n3009 = x162 | n3008 ;
  assign n3010 = n3009 ^ n1024 ^ 1'b0 ;
  assign n3011 = n2230 ^ n417 ^ x166 ;
  assign n3012 = n642 ^ n635 ^ 1'b0 ;
  assign n3013 = n3012 ^ n1655 ^ 1'b0 ;
  assign n3014 = n1740 | n3013 ;
  assign n3015 = ( n577 & n1840 ) | ( n577 & ~n2523 ) | ( n1840 & ~n2523 ) ;
  assign n3016 = n2538 | n3015 ;
  assign n3017 = n3016 ^ n1264 ^ n672 ;
  assign n3021 = x88 | n857 ;
  assign n3018 = n1118 | n1219 ;
  assign n3019 = n600 | n3018 ;
  assign n3020 = n1633 & n3019 ;
  assign n3022 = n3021 ^ n3020 ^ 1'b0 ;
  assign n3023 = ( n917 & n1980 ) | ( n917 & n3022 ) | ( n1980 & n3022 ) ;
  assign n3032 = n300 | n333 ;
  assign n3024 = x212 & ~n1941 ;
  assign n3028 = x58 & ~n2513 ;
  assign n3029 = n3028 ^ n609 ^ 1'b0 ;
  assign n3025 = ( x113 & n1172 ) | ( x113 & n1229 ) | ( n1172 & n1229 ) ;
  assign n3026 = n888 & ~n3025 ;
  assign n3027 = ~x179 & n3026 ;
  assign n3030 = n3029 ^ n3027 ^ n1389 ;
  assign n3031 = n3024 & n3030 ;
  assign n3033 = n3032 ^ n3031 ^ 1'b0 ;
  assign n3034 = ( x231 & n347 ) | ( x231 & n992 ) | ( n347 & n992 ) ;
  assign n3035 = n3034 ^ n1253 ^ 1'b0 ;
  assign n3036 = ~n264 & n3035 ;
  assign n3038 = n1733 ^ x90 ^ 1'b0 ;
  assign n3039 = n1495 & ~n3038 ;
  assign n3037 = ( n369 & n951 ) | ( n369 & ~n1173 ) | ( n951 & ~n1173 ) ;
  assign n3040 = n3039 ^ n3037 ^ n1046 ;
  assign n3041 = n2287 | n3040 ;
  assign n3042 = n3041 ^ n2188 ^ 1'b0 ;
  assign n3043 = n1071 | n2274 ;
  assign n3044 = n845 | n3043 ;
  assign n3045 = n1769 | n1843 ;
  assign n3047 = n1321 | n1836 ;
  assign n3046 = ( x133 & ~n371 ) | ( x133 & n1084 ) | ( ~n371 & n1084 ) ;
  assign n3048 = n3047 ^ n3046 ^ 1'b0 ;
  assign n3049 = ~n3045 & n3048 ;
  assign n3050 = ( n817 & ~n1647 ) | ( n817 & n3049 ) | ( ~n1647 & n3049 ) ;
  assign n3051 = ( n2465 & n2713 ) | ( n2465 & ~n3050 ) | ( n2713 & ~n3050 ) ;
  assign n3062 = n1251 | n1597 ;
  assign n3061 = ( x78 & n663 ) | ( x78 & ~n1226 ) | ( n663 & ~n1226 ) ;
  assign n3058 = n1243 & n2871 ;
  assign n3059 = n3058 ^ n2191 ^ 1'b0 ;
  assign n3056 = n1266 | n1855 ;
  assign n3053 = ~x163 & n1547 ;
  assign n3054 = ~n967 & n3053 ;
  assign n3055 = n1274 | n3054 ;
  assign n3057 = n3056 ^ n3055 ^ 1'b0 ;
  assign n3052 = ~x7 & n1480 ;
  assign n3060 = n3059 ^ n3057 ^ n3052 ;
  assign n3063 = n3062 ^ n3061 ^ n3060 ;
  assign n3064 = n2308 ^ n2145 ^ n1639 ;
  assign n3065 = n1423 ^ n565 ^ 1'b0 ;
  assign n3067 = x102 | n1151 ;
  assign n3068 = n591 & ~n3067 ;
  assign n3069 = n3068 ^ n294 ^ 1'b0 ;
  assign n3070 = ~n884 & n3069 ;
  assign n3066 = n1821 ^ n1364 ^ n1314 ;
  assign n3071 = n3070 ^ n3066 ^ 1'b0 ;
  assign n3072 = ~n1144 & n1226 ;
  assign n3073 = n2313 ^ n1213 ^ n1009 ;
  assign n3074 = n3073 ^ n1744 ^ 1'b0 ;
  assign n3075 = ( n2135 & n3072 ) | ( n2135 & ~n3074 ) | ( n3072 & ~n3074 ) ;
  assign n3077 = x110 & n339 ;
  assign n3078 = ~x115 & n3077 ;
  assign n3076 = n2028 | n2809 ;
  assign n3079 = n3078 ^ n3076 ^ 1'b0 ;
  assign n3080 = ( ~n790 & n1149 ) | ( ~n790 & n1763 ) | ( n1149 & n1763 ) ;
  assign n3081 = n884 ^ n326 ^ 1'b0 ;
  assign n3082 = x73 & ~n3081 ;
  assign n3083 = n3082 ^ x171 ^ 1'b0 ;
  assign n3084 = n3083 ^ n2351 ^ 1'b0 ;
  assign n3085 = n341 & ~n3084 ;
  assign n3086 = n1120 & ~n1377 ;
  assign n3087 = ( n2921 & n3085 ) | ( n2921 & n3086 ) | ( n3085 & n3086 ) ;
  assign n3088 = ~n2444 & n3087 ;
  assign n3089 = n3088 ^ n2938 ^ 1'b0 ;
  assign n3090 = ~n3080 & n3089 ;
  assign n3092 = ~n1251 & n2088 ;
  assign n3093 = n3092 ^ n1133 ^ 1'b0 ;
  assign n3094 = n1763 | n3093 ;
  assign n3091 = ( x193 & n752 ) | ( x193 & ~n2210 ) | ( n752 & ~n2210 ) ;
  assign n3095 = n3094 ^ n3091 ^ 1'b0 ;
  assign n3096 = n1441 ^ n1164 ^ 1'b0 ;
  assign n3097 = ~n587 & n945 ;
  assign n3104 = x153 & n1357 ;
  assign n3098 = n1649 | n1989 ;
  assign n3099 = n3098 ^ n385 ^ 1'b0 ;
  assign n3100 = n688 & n862 ;
  assign n3101 = n3100 ^ n1545 ^ 1'b0 ;
  assign n3102 = n3099 & ~n3101 ;
  assign n3103 = ~n1687 & n3102 ;
  assign n3105 = n3104 ^ n3103 ^ 1'b0 ;
  assign n3106 = n1076 & n3105 ;
  assign n3107 = n2136 ^ n270 ^ 1'b0 ;
  assign n3108 = n377 ^ x70 ^ 1'b0 ;
  assign n3109 = n2524 ^ n2441 ^ x171 ;
  assign n3110 = x54 & n1763 ;
  assign n3111 = n3109 & ~n3110 ;
  assign n3112 = n2840 & n3111 ;
  assign n3113 = ~n1540 & n1634 ;
  assign n3114 = n3113 ^ n1593 ^ 1'b0 ;
  assign n3115 = ~n302 & n3114 ;
  assign n3118 = n673 & ~n1700 ;
  assign n3119 = n2730 & n3118 ;
  assign n3120 = n3119 ^ n3037 ^ n901 ;
  assign n3116 = n1019 | n1107 ;
  assign n3117 = n1320 & ~n3116 ;
  assign n3121 = n3120 ^ n3117 ^ n2119 ;
  assign n3122 = n647 & n939 ;
  assign n3123 = n1536 | n3122 ;
  assign n3124 = n1776 & ~n3123 ;
  assign n3125 = n3124 ^ n412 ^ 1'b0 ;
  assign n3126 = n1880 ^ n1131 ^ 1'b0 ;
  assign n3127 = x70 & n3126 ;
  assign n3128 = n310 & n3127 ;
  assign n3129 = n476 | n3128 ;
  assign n3130 = n3129 ^ n292 ^ 1'b0 ;
  assign n3131 = ~n1672 & n3130 ;
  assign n3132 = ~n3099 & n3131 ;
  assign n3133 = ~n1038 & n3132 ;
  assign n3134 = ~n2615 & n2806 ;
  assign n3135 = ~n2193 & n3134 ;
  assign n3136 = n3135 ^ n906 ^ n800 ;
  assign n3137 = n350 & n371 ;
  assign n3138 = n500 & n3137 ;
  assign n3139 = n531 & n3138 ;
  assign n3140 = n1090 ^ x212 ^ 1'b0 ;
  assign n3141 = ~n1136 & n1861 ;
  assign n3142 = ~n3140 & n3141 ;
  assign n3143 = n2052 | n3142 ;
  assign n3144 = n3143 ^ n1202 ^ 1'b0 ;
  assign n3146 = n941 | n2900 ;
  assign n3145 = n1818 ^ n501 ^ x250 ;
  assign n3147 = n3146 ^ n3145 ^ n1851 ;
  assign n3148 = ~n1906 & n2411 ;
  assign n3149 = ~n1339 & n3004 ;
  assign n3150 = n3149 ^ n651 ^ 1'b0 ;
  assign n3153 = n2215 ^ n354 ^ 1'b0 ;
  assign n3154 = ( x167 & n2471 ) | ( x167 & ~n3153 ) | ( n2471 & ~n3153 ) ;
  assign n3151 = n2009 ^ n967 ^ 1'b0 ;
  assign n3152 = ( n923 & ~n1501 ) | ( n923 & n3151 ) | ( ~n1501 & n3151 ) ;
  assign n3155 = n3154 ^ n3152 ^ n3146 ;
  assign n3158 = x247 & ~n2705 ;
  assign n3159 = ( n706 & ~n2709 ) | ( n706 & n3158 ) | ( ~n2709 & n3158 ) ;
  assign n3156 = n2942 ^ n1644 ^ n1481 ;
  assign n3157 = n3156 ^ n617 ^ n457 ;
  assign n3160 = n3159 ^ n3157 ^ x168 ;
  assign n3161 = n1657 ^ n1651 ^ 1'b0 ;
  assign n3162 = n1225 & ~n3161 ;
  assign n3163 = n3160 & n3162 ;
  assign n3164 = n701 & ~n1042 ;
  assign n3165 = n3164 ^ x124 ^ 1'b0 ;
  assign n3166 = x35 & ~n3165 ;
  assign n3167 = n1504 ^ x103 ^ 1'b0 ;
  assign n3168 = n921 | n3167 ;
  assign n3169 = n1399 ^ n1246 ^ x151 ;
  assign n3170 = n3169 ^ n1979 ^ 1'b0 ;
  assign n3171 = x149 & ~n872 ;
  assign n3172 = ~x230 & n3171 ;
  assign n3173 = n3172 ^ n860 ^ 1'b0 ;
  assign n3174 = n658 & n1398 ;
  assign n3175 = n3174 ^ n2456 ^ 1'b0 ;
  assign n3176 = n1214 & ~n3175 ;
  assign n3177 = n1294 & n2986 ;
  assign n3178 = n3177 ^ n354 ^ 1'b0 ;
  assign n3179 = n3178 ^ n989 ^ 1'b0 ;
  assign n3180 = n1307 | n3179 ;
  assign n3189 = n1220 & ~n1380 ;
  assign n3190 = n3189 ^ n1723 ^ 1'b0 ;
  assign n3187 = n1774 ^ n824 ^ n654 ;
  assign n3182 = x127 & ~n967 ;
  assign n3183 = n3182 ^ x67 ^ 1'b0 ;
  assign n3184 = n1270 & n3183 ;
  assign n3185 = n3184 ^ n1136 ^ 1'b0 ;
  assign n3186 = ~n335 & n3185 ;
  assign n3188 = n3187 ^ n3186 ^ 1'b0 ;
  assign n3191 = n3190 ^ n3188 ^ n1950 ;
  assign n3181 = n1727 ^ n639 ^ 1'b0 ;
  assign n3192 = n3191 ^ n3181 ^ n451 ;
  assign n3193 = n3192 ^ n3185 ^ 1'b0 ;
  assign n3194 = ~n3180 & n3193 ;
  assign n3195 = n1192 ^ x39 ^ 1'b0 ;
  assign n3196 = x202 & ~n3195 ;
  assign n3197 = n1005 ^ n542 ^ x162 ;
  assign n3198 = n464 & n3197 ;
  assign n3199 = n3198 ^ n715 ^ 1'b0 ;
  assign n3200 = n3196 & n3199 ;
  assign n3202 = x199 & ~n859 ;
  assign n3203 = n1164 & n3202 ;
  assign n3201 = n427 | n482 ;
  assign n3204 = n3203 ^ n3201 ^ 1'b0 ;
  assign n3205 = n818 ^ x144 ^ 1'b0 ;
  assign n3206 = n1069 | n3205 ;
  assign n3207 = x147 & ~n3206 ;
  assign n3208 = n1231 | n3207 ;
  assign n3209 = n902 | n3208 ;
  assign n3210 = n3204 & ~n3209 ;
  assign n3211 = n1418 & n3210 ;
  assign n3212 = n1537 ^ x143 ^ 1'b0 ;
  assign n3213 = n3212 ^ n3100 ^ 1'b0 ;
  assign n3214 = x103 & ~n1975 ;
  assign n3215 = n2200 & n3214 ;
  assign n3216 = n803 & n2373 ;
  assign n3217 = n2727 ^ n1674 ^ n1420 ;
  assign n3218 = n861 ^ x246 ^ 1'b0 ;
  assign n3219 = n405 & n3218 ;
  assign n3220 = ( ~n1205 & n1727 ) | ( ~n1205 & n1921 ) | ( n1727 & n1921 ) ;
  assign n3221 = n2778 ^ n1817 ^ 1'b0 ;
  assign n3222 = ~n2693 & n3221 ;
  assign n3223 = ( n1891 & n1893 ) | ( n1891 & n1959 ) | ( n1893 & n1959 ) ;
  assign n3224 = n1290 | n3223 ;
  assign n3225 = n2150 | n3224 ;
  assign n3226 = n1935 ^ n655 ^ 1'b0 ;
  assign n3227 = n3226 ^ n2594 ^ 1'b0 ;
  assign n3228 = n1309 ^ n1004 ^ 1'b0 ;
  assign n3229 = x52 & n3228 ;
  assign n3230 = n341 & n517 ;
  assign n3231 = n3230 ^ x96 ^ 1'b0 ;
  assign n3232 = n1308 & n3231 ;
  assign n3233 = n3232 ^ n2476 ^ x140 ;
  assign n3234 = n3100 ^ n1220 ^ 1'b0 ;
  assign n3235 = ( ~n3073 & n3233 ) | ( ~n3073 & n3234 ) | ( n3233 & n3234 ) ;
  assign n3236 = n3235 ^ n335 ^ 1'b0 ;
  assign n3238 = n1561 | n1930 ;
  assign n3237 = n769 & n1294 ;
  assign n3239 = n3238 ^ n3237 ^ 1'b0 ;
  assign n3240 = n1472 ^ n577 ^ 1'b0 ;
  assign n3241 = x108 & ~n840 ;
  assign n3242 = n3241 ^ n396 ^ 1'b0 ;
  assign n3243 = n3242 ^ n2856 ^ 1'b0 ;
  assign n3244 = n3240 & ~n3243 ;
  assign n3245 = n1329 & n3244 ;
  assign n3247 = n1053 & n1533 ;
  assign n3246 = x184 & n2644 ;
  assign n3248 = n3247 ^ n3246 ^ 1'b0 ;
  assign n3249 = n3248 ^ n3100 ^ 1'b0 ;
  assign n3250 = n1082 & ~n3249 ;
  assign n3254 = n369 | n409 ;
  assign n3255 = ( x137 & n1586 ) | ( x137 & n3254 ) | ( n1586 & n3254 ) ;
  assign n3251 = ~n835 & n1174 ;
  assign n3252 = n2116 & n3251 ;
  assign n3253 = n1343 & ~n3252 ;
  assign n3256 = n3255 ^ n3253 ^ 1'b0 ;
  assign n3257 = x22 & ~n2240 ;
  assign n3258 = n2547 | n2977 ;
  assign n3259 = n3257 | n3258 ;
  assign n3260 = n2917 ^ n2539 ^ 1'b0 ;
  assign n3261 = n905 ^ n599 ^ n425 ;
  assign n3262 = n3261 ^ n2328 ^ n1270 ;
  assign n3263 = ( n351 & n1076 ) | ( n351 & n2046 ) | ( n1076 & n2046 ) ;
  assign n3264 = n591 | n3263 ;
  assign n3265 = n2375 & n3264 ;
  assign n3266 = ~n475 & n3265 ;
  assign n3267 = x30 & ~n1062 ;
  assign n3268 = n3267 ^ n1981 ^ n1452 ;
  assign n3269 = n1296 ^ n1141 ^ 1'b0 ;
  assign n3270 = n2692 ^ n1564 ^ 1'b0 ;
  assign n3271 = n2230 & n3270 ;
  assign n3274 = n330 & n442 ;
  assign n3273 = n614 ^ x174 ^ 1'b0 ;
  assign n3272 = x138 & ~n436 ;
  assign n3275 = n3274 ^ n3273 ^ n3272 ;
  assign n3276 = n3275 ^ n2058 ^ 1'b0 ;
  assign n3277 = n3271 & n3276 ;
  assign n3278 = n2197 & n3277 ;
  assign n3279 = n3269 & n3278 ;
  assign n3280 = n3268 | n3279 ;
  assign n3281 = n3266 & ~n3280 ;
  assign n3282 = n450 & ~n2463 ;
  assign n3283 = ( x95 & n268 ) | ( x95 & n2706 ) | ( n268 & n2706 ) ;
  assign n3284 = n3283 ^ n1319 ^ 1'b0 ;
  assign n3285 = n2284 | n3284 ;
  assign n3286 = n993 & n3081 ;
  assign n3287 = n2868 & ~n3286 ;
  assign n3288 = n3285 & n3287 ;
  assign n3289 = n2216 ^ n1467 ^ n1234 ;
  assign n3290 = n763 | n1987 ;
  assign n3291 = n1148 & ~n3290 ;
  assign n3292 = n3291 ^ n2055 ^ n1604 ;
  assign n3293 = n2970 & n3292 ;
  assign n3294 = ~n3289 & n3293 ;
  assign n3295 = n1789 & ~n1944 ;
  assign n3296 = n3295 ^ n1778 ^ 1'b0 ;
  assign n3297 = n3296 ^ n1080 ^ x218 ;
  assign n3298 = n3085 ^ n514 ^ 1'b0 ;
  assign n3299 = n329 & n3298 ;
  assign n3300 = ( n872 & ~n2680 ) | ( n872 & n3299 ) | ( ~n2680 & n3299 ) ;
  assign n3301 = n3300 ^ n1994 ^ 1'b0 ;
  assign n3302 = ~n2574 & n3301 ;
  assign n3303 = n1319 & ~n2618 ;
  assign n3304 = ~n1705 & n3303 ;
  assign n3305 = n1328 ^ n1006 ^ 1'b0 ;
  assign n3306 = ~n2286 & n3034 ;
  assign n3307 = n3306 ^ n1856 ^ 1'b0 ;
  assign n3308 = ( n277 & n1007 ) | ( n277 & n1304 ) | ( n1007 & n1304 ) ;
  assign n3309 = n2945 & n3308 ;
  assign n3310 = n1179 | n3309 ;
  assign n3311 = ~n3307 & n3310 ;
  assign n3312 = n3305 & n3311 ;
  assign n3313 = x136 & ~n1922 ;
  assign n3314 = n2019 & n3313 ;
  assign n3315 = ~n854 & n2660 ;
  assign n3316 = n1105 ^ n322 ^ 1'b0 ;
  assign n3317 = n3316 ^ x131 ^ 1'b0 ;
  assign n3318 = n1002 | n3317 ;
  assign n3319 = n3318 ^ x13 ^ 1'b0 ;
  assign n3320 = n3315 & ~n3319 ;
  assign n3321 = ~n498 & n900 ;
  assign n3322 = n1108 | n3120 ;
  assign n3323 = x27 & ~n1869 ;
  assign n3324 = n3323 ^ n1362 ^ 1'b0 ;
  assign n3325 = n390 ^ n266 ^ 1'b0 ;
  assign n3326 = n1406 ^ n578 ^ 1'b0 ;
  assign n3327 = n3325 & ~n3326 ;
  assign n3328 = n3327 ^ n533 ^ n421 ;
  assign n3329 = ( x108 & ~n565 ) | ( x108 & n3328 ) | ( ~n565 & n3328 ) ;
  assign n3330 = n2086 ^ x164 ^ 1'b0 ;
  assign n3331 = n3329 & ~n3330 ;
  assign n3332 = n2730 ^ n2088 ^ n587 ;
  assign n3333 = n326 ^ x143 ^ 1'b0 ;
  assign n3334 = ~n3332 & n3333 ;
  assign n3335 = n3334 ^ n3185 ^ 1'b0 ;
  assign n3336 = ( n326 & n539 ) | ( n326 & ~n1452 ) | ( n539 & ~n1452 ) ;
  assign n3337 = x137 ^ x8 ^ 1'b0 ;
  assign n3338 = n1310 & n3337 ;
  assign n3339 = ( n735 & ~n1074 ) | ( n735 & n3338 ) | ( ~n1074 & n3338 ) ;
  assign n3340 = n1083 & n3234 ;
  assign n3341 = ~n3339 & n3340 ;
  assign n3342 = ( n559 & n1634 ) | ( n559 & n2342 ) | ( n1634 & n2342 ) ;
  assign n3343 = n2708 ^ n1042 ^ 1'b0 ;
  assign n3344 = n3237 & n3343 ;
  assign n3345 = n2240 ^ x68 ^ 1'b0 ;
  assign n3346 = x106 & n3345 ;
  assign n3347 = n3346 ^ n1353 ^ 1'b0 ;
  assign n3348 = n3040 | n3347 ;
  assign n3349 = ( n606 & ~n2102 ) | ( n606 & n2674 ) | ( ~n2102 & n2674 ) ;
  assign n3350 = x169 & ~n1850 ;
  assign n3351 = n3350 ^ n1249 ^ 1'b0 ;
  assign n3352 = ( x198 & ~n2005 ) | ( x198 & n3351 ) | ( ~n2005 & n3351 ) ;
  assign n3354 = n1181 ^ n950 ^ 1'b0 ;
  assign n3355 = n1840 & ~n3354 ;
  assign n3356 = n3355 ^ n857 ^ 1'b0 ;
  assign n3353 = ( x84 & ~n403 ) | ( x84 & n850 ) | ( ~n403 & n850 ) ;
  assign n3357 = n3356 ^ n3353 ^ n1650 ;
  assign n3358 = n1214 & ~n3357 ;
  assign n3359 = ( n3349 & n3352 ) | ( n3349 & n3358 ) | ( n3352 & n3358 ) ;
  assign n3360 = n2807 | n3359 ;
  assign n3364 = n2039 ^ n1349 ^ n379 ;
  assign n3365 = n3364 ^ n1266 ^ 1'b0 ;
  assign n3366 = n2705 & ~n3365 ;
  assign n3367 = n3366 ^ n1971 ^ 1'b0 ;
  assign n3368 = n507 | n3367 ;
  assign n3369 = ( x48 & ~n945 ) | ( x48 & n3368 ) | ( ~n945 & n3368 ) ;
  assign n3370 = n3369 ^ n593 ^ 1'b0 ;
  assign n3361 = n476 | n785 ;
  assign n3362 = ~n1993 & n3361 ;
  assign n3363 = n3362 ^ n1023 ^ 1'b0 ;
  assign n3371 = n3370 ^ n3363 ^ n1286 ;
  assign n3377 = n1829 ^ n1069 ^ 1'b0 ;
  assign n3378 = n725 & n3377 ;
  assign n3379 = x4 & ~n3378 ;
  assign n3380 = n1606 ^ n417 ^ 1'b0 ;
  assign n3381 = ~n3379 & n3380 ;
  assign n3375 = n2692 ^ n525 ^ 1'b0 ;
  assign n3372 = n294 & ~n699 ;
  assign n3373 = n3372 ^ n1175 ^ 1'b0 ;
  assign n3374 = n3373 ^ n2656 ^ n2259 ;
  assign n3376 = n3375 ^ n3374 ^ 1'b0 ;
  assign n3382 = n3381 ^ n3376 ^ 1'b0 ;
  assign n3383 = n2886 & n3382 ;
  assign n3384 = ~n310 & n735 ;
  assign n3385 = n449 & n3384 ;
  assign n3386 = n3385 ^ n2200 ^ 1'b0 ;
  assign n3387 = n806 & ~n986 ;
  assign n3388 = n3387 ^ n1302 ^ 1'b0 ;
  assign n3389 = x169 & n3388 ;
  assign n3390 = ( n571 & n1022 ) | ( n571 & n1063 ) | ( n1022 & n1063 ) ;
  assign n3394 = ( x6 & x71 ) | ( x6 & ~x250 ) | ( x71 & ~x250 ) ;
  assign n3391 = ( n1240 & n1709 ) | ( n1240 & n2924 ) | ( n1709 & n2924 ) ;
  assign n3392 = n1252 | n3391 ;
  assign n3393 = n2437 & ~n3392 ;
  assign n3395 = n3394 ^ n3393 ^ 1'b0 ;
  assign n3396 = n3390 | n3395 ;
  assign n3400 = ~n256 & n537 ;
  assign n3397 = n1633 ^ n264 ^ 1'b0 ;
  assign n3398 = n2416 & ~n3397 ;
  assign n3399 = ~n3223 & n3398 ;
  assign n3401 = n3400 ^ n3399 ^ 1'b0 ;
  assign n3402 = ( x90 & n423 ) | ( x90 & n615 ) | ( n423 & n615 ) ;
  assign n3403 = n3402 ^ n1206 ^ 1'b0 ;
  assign n3404 = n545 ^ n338 ^ 1'b0 ;
  assign n3405 = x209 & x220 ;
  assign n3406 = ~x126 & n3405 ;
  assign n3407 = n1388 & ~n3406 ;
  assign n3408 = n1944 & n3407 ;
  assign n3409 = n589 & n3408 ;
  assign n3410 = n3409 ^ n394 ^ x169 ;
  assign n3411 = n1768 & n3410 ;
  assign n3412 = n3411 ^ n419 ^ 1'b0 ;
  assign n3413 = ~n2105 & n2431 ;
  assign n3414 = n1133 | n3413 ;
  assign n3415 = n2603 ^ x108 ^ 1'b0 ;
  assign n3416 = n922 & n3415 ;
  assign n3417 = x88 & ~n3416 ;
  assign n3418 = x158 & n1369 ;
  assign n3419 = n3083 ^ n2107 ^ 1'b0 ;
  assign n3420 = n2268 & n3419 ;
  assign n3421 = ~n1349 & n3420 ;
  assign n3422 = n1595 & n1723 ;
  assign n3423 = x8 & n955 ;
  assign n3424 = ( n604 & n797 ) | ( n604 & n3423 ) | ( n797 & n3423 ) ;
  assign n3425 = n3424 ^ n1069 ^ 1'b0 ;
  assign n3426 = n1045 ^ n257 ^ 1'b0 ;
  assign n3427 = n3426 ^ n2940 ^ 1'b0 ;
  assign n3428 = ~n1690 & n3427 ;
  assign n3429 = n410 & n1261 ;
  assign n3430 = n697 | n3429 ;
  assign n3431 = ( x195 & n764 ) | ( x195 & n3430 ) | ( n764 & n3430 ) ;
  assign n3432 = n2715 ^ n2510 ^ n876 ;
  assign n3433 = ( n1733 & n3431 ) | ( n1733 & n3432 ) | ( n3431 & n3432 ) ;
  assign n3435 = x156 & n2030 ;
  assign n3436 = ~x236 & n3435 ;
  assign n3434 = n3047 & n3159 ;
  assign n3437 = n3436 ^ n3434 ^ n2950 ;
  assign n3438 = n2220 ^ n1351 ^ 1'b0 ;
  assign n3439 = n1787 & ~n3438 ;
  assign n3440 = n3439 ^ n2365 ^ 1'b0 ;
  assign n3441 = n1194 & n3245 ;
  assign n3442 = n3070 & n3441 ;
  assign n3451 = n1758 ^ n517 ^ 1'b0 ;
  assign n3452 = x157 & ~n3451 ;
  assign n3443 = x218 & n704 ;
  assign n3444 = n3443 ^ n859 ^ 1'b0 ;
  assign n3445 = ( ~n268 & n2454 ) | ( ~n268 & n3444 ) | ( n2454 & n3444 ) ;
  assign n3446 = n764 & ~n2048 ;
  assign n3447 = n3332 & n3446 ;
  assign n3448 = n3122 | n3447 ;
  assign n3449 = n3448 ^ n1858 ^ 1'b0 ;
  assign n3450 = n3445 & ~n3449 ;
  assign n3453 = n3452 ^ n3450 ^ 1'b0 ;
  assign n3456 = ( n282 & n588 ) | ( n282 & ~n1288 ) | ( n588 & ~n1288 ) ;
  assign n3454 = ~n450 & n2931 ;
  assign n3455 = n3454 ^ n1787 ^ x219 ;
  assign n3457 = n3456 ^ n3455 ^ 1'b0 ;
  assign n3458 = x160 | n1685 ;
  assign n3460 = n1199 & n1729 ;
  assign n3461 = n3460 ^ x190 ^ 1'b0 ;
  assign n3459 = n820 & ~n1807 ;
  assign n3462 = n3461 ^ n3459 ^ 1'b0 ;
  assign n3463 = ~n1950 & n3462 ;
  assign n3464 = ( ~x213 & n2367 ) | ( ~x213 & n2459 ) | ( n2367 & n2459 ) ;
  assign n3465 = x52 & n417 ;
  assign n3466 = ~n853 & n3465 ;
  assign n3467 = n649 & ~n1966 ;
  assign n3468 = n3467 ^ n1890 ^ 1'b0 ;
  assign n3469 = n2671 & ~n3468 ;
  assign n3470 = x83 & ~n354 ;
  assign n3471 = n3470 ^ x71 ^ 1'b0 ;
  assign n3472 = n1254 & n2208 ;
  assign n3473 = n3471 & ~n3472 ;
  assign n3474 = n3473 ^ n3060 ^ 1'b0 ;
  assign n3475 = n2532 ^ n1035 ^ 1'b0 ;
  assign n3476 = n3475 ^ n1718 ^ 1'b0 ;
  assign n3477 = ~n333 & n402 ;
  assign n3478 = n1328 & n3233 ;
  assign n3479 = n3478 ^ n1871 ^ 1'b0 ;
  assign n3480 = n1579 & n3479 ;
  assign n3481 = ~n487 & n3480 ;
  assign n3482 = n3477 & ~n3481 ;
  assign n3483 = n3482 ^ n623 ^ 1'b0 ;
  assign n3484 = n2515 & ~n3305 ;
  assign n3485 = ~n3483 & n3484 ;
  assign n3486 = n3476 | n3485 ;
  assign n3487 = n3486 ^ n2780 ^ 1'b0 ;
  assign n3488 = n715 | n741 ;
  assign n3491 = n801 & n1197 ;
  assign n3492 = n3491 ^ n552 ^ 1'b0 ;
  assign n3493 = n3492 ^ n3142 ^ 1'b0 ;
  assign n3494 = n322 | n3493 ;
  assign n3489 = n2207 & n2245 ;
  assign n3490 = n3489 ^ n2289 ^ 1'b0 ;
  assign n3495 = n3494 ^ n3490 ^ 1'b0 ;
  assign n3496 = n3488 & ~n3495 ;
  assign n3497 = n3496 ^ n1919 ^ 1'b0 ;
  assign n3498 = n1176 ^ n902 ^ x33 ;
  assign n3499 = n1071 ^ n654 ^ 1'b0 ;
  assign n3500 = n603 & ~n3499 ;
  assign n3501 = n567 & n3500 ;
  assign n3502 = ~n731 & n3501 ;
  assign n3503 = n3502 ^ x82 ^ 1'b0 ;
  assign n3504 = n1262 & ~n3503 ;
  assign n3505 = n3504 ^ n811 ^ 1'b0 ;
  assign n3506 = n2833 & ~n3505 ;
  assign n3507 = ~n3498 & n3506 ;
  assign n3508 = ( ~x68 & n2551 ) | ( ~x68 & n3507 ) | ( n2551 & n3507 ) ;
  assign n3516 = n1985 ^ n725 ^ x218 ;
  assign n3517 = n718 & n3516 ;
  assign n3513 = n958 ^ n625 ^ 1'b0 ;
  assign n3514 = n2045 | n3513 ;
  assign n3509 = n1229 ^ n537 ^ 1'b0 ;
  assign n3510 = n434 & ~n3509 ;
  assign n3511 = n3510 ^ n1709 ^ 1'b0 ;
  assign n3512 = ( x130 & n2222 ) | ( x130 & ~n3511 ) | ( n2222 & ~n3511 ) ;
  assign n3515 = n3514 ^ n3512 ^ n1543 ;
  assign n3518 = n3517 ^ n3515 ^ n974 ;
  assign n3520 = n1615 | n2940 ;
  assign n3521 = n3520 ^ n1602 ^ 1'b0 ;
  assign n3522 = n457 & ~n3521 ;
  assign n3523 = ~n3072 & n3522 ;
  assign n3519 = n1725 ^ x78 ^ 1'b0 ;
  assign n3524 = n3523 ^ n3519 ^ 1'b0 ;
  assign n3525 = n807 | n3524 ;
  assign n3526 = n345 | n2342 ;
  assign n3527 = n3526 ^ n978 ^ 1'b0 ;
  assign n3528 = ( n575 & ~n1022 ) | ( n575 & n2182 ) | ( ~n1022 & n2182 ) ;
  assign n3529 = n3528 ^ n3277 ^ n1848 ;
  assign n3530 = n3425 | n3529 ;
  assign n3531 = n402 & ~n3530 ;
  assign n3537 = x132 & ~n2355 ;
  assign n3538 = n3390 & n3537 ;
  assign n3532 = n1454 ^ n706 ^ 1'b0 ;
  assign n3533 = ( ~n1778 & n3317 ) | ( ~n1778 & n3532 ) | ( n3317 & n3532 ) ;
  assign n3534 = n1955 | n1966 ;
  assign n3535 = n3534 ^ n1144 ^ 1'b0 ;
  assign n3536 = n3533 | n3535 ;
  assign n3539 = n3538 ^ n3536 ^ 1'b0 ;
  assign n3540 = n407 ^ x233 ^ 1'b0 ;
  assign n3541 = ( n514 & ~n915 ) | ( n514 & n1189 ) | ( ~n915 & n1189 ) ;
  assign n3542 = n3541 ^ n1086 ^ n539 ;
  assign n3543 = n632 & ~n1420 ;
  assign n3544 = ( ~n2440 & n3542 ) | ( ~n2440 & n3543 ) | ( n3542 & n3543 ) ;
  assign n3546 = ( x230 & n905 ) | ( x230 & n3289 ) | ( n905 & n3289 ) ;
  assign n3545 = n1701 ^ n644 ^ 1'b0 ;
  assign n3547 = n3546 ^ n3545 ^ n989 ;
  assign n3548 = n593 & ~n741 ;
  assign n3549 = n3548 ^ n2287 ^ 1'b0 ;
  assign n3550 = ~n1383 & n3549 ;
  assign n3555 = n805 & ~n3444 ;
  assign n3551 = x87 & n1673 ;
  assign n3552 = n3551 ^ n2056 ^ x214 ;
  assign n3553 = n2860 & n3552 ;
  assign n3554 = n290 & n3553 ;
  assign n3556 = n3555 ^ n3554 ^ 1'b0 ;
  assign n3557 = n1478 & ~n1719 ;
  assign n3558 = n1453 ^ n1241 ^ 1'b0 ;
  assign n3559 = n3557 & n3558 ;
  assign n3562 = n1222 | n2137 ;
  assign n3563 = n3562 ^ n1203 ^ 1'b0 ;
  assign n3560 = n807 & ~n1133 ;
  assign n3561 = n1685 & n3560 ;
  assign n3564 = n3563 ^ n3561 ^ 1'b0 ;
  assign n3565 = x233 & ~n632 ;
  assign n3566 = n3565 ^ x129 ^ 1'b0 ;
  assign n3567 = ( ~x89 & n1290 ) | ( ~x89 & n2531 ) | ( n1290 & n2531 ) ;
  assign n3568 = ( x45 & x128 ) | ( x45 & n3567 ) | ( x128 & n3567 ) ;
  assign n3569 = n3568 ^ n2416 ^ 1'b0 ;
  assign n3570 = n1644 & n3569 ;
  assign n3571 = n3140 ^ n2080 ^ 1'b0 ;
  assign n3572 = n3571 ^ n639 ^ 1'b0 ;
  assign n3573 = ( n3566 & n3570 ) | ( n3566 & ~n3572 ) | ( n3570 & ~n3572 ) ;
  assign n3574 = n881 | n1440 ;
  assign n3575 = n3574 ^ n973 ^ 1'b0 ;
  assign n3576 = x55 & ~n3575 ;
  assign n3577 = ~x218 & n3576 ;
  assign n3578 = n3577 ^ n288 ^ 1'b0 ;
  assign n3579 = n1280 & n1495 ;
  assign n3580 = n362 & n3579 ;
  assign n3581 = x251 | n3580 ;
  assign n3582 = n1510 & ~n3215 ;
  assign n3583 = n3581 & n3582 ;
  assign n3584 = n1468 ^ n1199 ^ 1'b0 ;
  assign n3585 = ~n2804 & n3584 ;
  assign n3586 = n3065 & n3585 ;
  assign n3587 = ~n3463 & n3586 ;
  assign n3589 = ( x150 & n464 ) | ( x150 & ~n1209 ) | ( n464 & ~n1209 ) ;
  assign n3588 = n952 | n1703 ;
  assign n3590 = n3589 ^ n3588 ^ 1'b0 ;
  assign n3591 = ( x219 & n1880 ) | ( x219 & ~n3590 ) | ( n1880 & ~n3590 ) ;
  assign n3592 = ~n1300 & n1407 ;
  assign n3593 = n1678 & n3592 ;
  assign n3594 = x121 & n807 ;
  assign n3595 = n3594 ^ x65 ^ 1'b0 ;
  assign n3596 = n870 & n2505 ;
  assign n3597 = n3596 ^ n1702 ^ 1'b0 ;
  assign n3598 = ~n2993 & n3597 ;
  assign n3599 = n3598 ^ n1429 ^ 1'b0 ;
  assign n3600 = n1080 | n2425 ;
  assign n3601 = n2635 ^ n1732 ^ 1'b0 ;
  assign n3602 = n2726 | n3601 ;
  assign n3603 = ~n1961 & n3528 ;
  assign n3604 = n3603 ^ n2103 ^ 1'b0 ;
  assign n3606 = x106 & x216 ;
  assign n3607 = ~x124 & n3606 ;
  assign n3605 = n2268 ^ n1595 ^ 1'b0 ;
  assign n3608 = n3607 ^ n3605 ^ n1519 ;
  assign n3612 = n2548 ^ x62 ^ 1'b0 ;
  assign n3610 = n2648 ^ n1080 ^ 1'b0 ;
  assign n3611 = n966 | n3610 ;
  assign n3613 = n3612 ^ n3611 ^ 1'b0 ;
  assign n3609 = n2885 ^ x159 ^ 1'b0 ;
  assign n3614 = n3613 ^ n3609 ^ n3514 ;
  assign n3615 = n1480 | n2009 ;
  assign n3616 = n951 & ~n3615 ;
  assign n3617 = ~n3614 & n3616 ;
  assign n3618 = ~n736 & n3242 ;
  assign n3619 = n3079 & n3618 ;
  assign n3620 = n3053 ^ x53 ^ 1'b0 ;
  assign n3621 = ~n519 & n1058 ;
  assign n3622 = ( n2138 & n3156 ) | ( n2138 & ~n3621 ) | ( n3156 & ~n3621 ) ;
  assign n3623 = n2056 ^ n804 ^ 1'b0 ;
  assign n3624 = x50 & n3623 ;
  assign n3627 = ~n649 & n1639 ;
  assign n3628 = ~n1718 & n3627 ;
  assign n3625 = x91 & ~n1863 ;
  assign n3626 = n1140 & n3625 ;
  assign n3629 = n3628 ^ n3626 ^ 1'b0 ;
  assign n3630 = n1234 ^ n423 ^ 1'b0 ;
  assign n3631 = n2235 ^ n1504 ^ 1'b0 ;
  assign n3632 = n2348 | n3631 ;
  assign n3633 = n3429 ^ n1439 ^ 1'b0 ;
  assign n3634 = n3632 & ~n3633 ;
  assign n3635 = x208 & n3634 ;
  assign n3636 = n3635 ^ n2942 ^ 1'b0 ;
  assign n3637 = ~x68 & n1809 ;
  assign n3638 = n3636 & ~n3637 ;
  assign n3639 = n1043 ^ n1024 ^ n848 ;
  assign n3640 = n394 & ~n3639 ;
  assign n3641 = ~n1661 & n3640 ;
  assign n3642 = ( n647 & n798 ) | ( n647 & ~n1336 ) | ( n798 & ~n1336 ) ;
  assign n3643 = n1374 | n3642 ;
  assign n3644 = n3268 & ~n3643 ;
  assign n3645 = ~n2964 & n3644 ;
  assign n3646 = n2313 & n3645 ;
  assign n3647 = n3203 ^ n1802 ^ n883 ;
  assign n3648 = n2624 & n3647 ;
  assign n3649 = x86 & ~n1302 ;
  assign n3650 = n3649 ^ n3261 ^ 1'b0 ;
  assign n3651 = n2049 | n3650 ;
  assign n3652 = n2784 & ~n3651 ;
  assign n3653 = n1807 | n3385 ;
  assign n3654 = n1126 ^ x205 ^ x162 ;
  assign n3655 = n2816 & n3654 ;
  assign n3656 = n3655 ^ n1522 ^ 1'b0 ;
  assign n3657 = n926 & n3656 ;
  assign n3658 = n3657 ^ n941 ^ 1'b0 ;
  assign n3659 = n2024 ^ n256 ^ 1'b0 ;
  assign n3660 = ( x15 & n2038 ) | ( x15 & ~n3566 ) | ( n2038 & ~n3566 ) ;
  assign n3661 = ~n1962 & n3660 ;
  assign n3662 = n1769 ^ n945 ^ 1'b0 ;
  assign n3663 = ~n2277 & n3184 ;
  assign n3664 = n3663 ^ n2280 ^ 1'b0 ;
  assign n3665 = n617 & ~n3664 ;
  assign n3666 = n3665 ^ n382 ^ 1'b0 ;
  assign n3667 = n853 | n1103 ;
  assign n3668 = n684 & n3115 ;
  assign n3669 = n3668 ^ n2379 ^ 1'b0 ;
  assign n3670 = n982 ^ x244 ^ 1'b0 ;
  assign n3671 = n1299 & ~n3670 ;
  assign n3672 = n3671 ^ n1258 ^ 1'b0 ;
  assign n3673 = n2286 | n3672 ;
  assign n3674 = n3673 ^ n1510 ^ 1'b0 ;
  assign n3675 = n1115 | n3674 ;
  assign n3676 = n2295 ^ n1474 ^ 1'b0 ;
  assign n3681 = n1323 ^ n672 ^ 1'b0 ;
  assign n3677 = x221 & ~n256 ;
  assign n3678 = n3677 ^ n1736 ^ 1'b0 ;
  assign n3679 = ( n1148 & n1636 ) | ( n1148 & n3678 ) | ( n1636 & n3678 ) ;
  assign n3680 = n3679 ^ n826 ^ 1'b0 ;
  assign n3682 = n3681 ^ n3680 ^ 1'b0 ;
  assign n3683 = ~n1724 & n3682 ;
  assign n3684 = ~n3066 & n3683 ;
  assign n3685 = ~n2915 & n3684 ;
  assign n3690 = n2554 & n3047 ;
  assign n3686 = x214 & ~n1091 ;
  assign n3687 = n3615 & n3686 ;
  assign n3688 = n3687 ^ n3015 ^ n318 ;
  assign n3689 = n3688 ^ n2683 ^ 1'b0 ;
  assign n3691 = n3690 ^ n3689 ^ n3458 ;
  assign n3692 = ( n507 & ~n790 ) | ( n507 & n1281 ) | ( ~n790 & n1281 ) ;
  assign n3693 = n3692 ^ n1958 ^ 1'b0 ;
  assign n3694 = n3693 ^ n750 ^ 1'b0 ;
  assign n3695 = ~n715 & n2222 ;
  assign n3696 = n1170 ^ x165 ^ 1'b0 ;
  assign n3697 = n3696 ^ n2939 ^ 1'b0 ;
  assign n3698 = n3695 & n3697 ;
  assign n3699 = n1158 ^ n259 ^ 1'b0 ;
  assign n3700 = x219 & ~n3699 ;
  assign n3701 = ~n2560 & n3700 ;
  assign n3702 = n2880 & n3701 ;
  assign n3703 = n2888 ^ n557 ^ 1'b0 ;
  assign n3704 = ~n1734 & n3703 ;
  assign n3705 = n3310 ^ n2112 ^ 1'b0 ;
  assign n3706 = n3705 ^ n3622 ^ 1'b0 ;
  assign n3707 = n1098 & n3706 ;
  assign n3708 = ( ~n1352 & n1613 ) | ( ~n1352 & n1939 ) | ( n1613 & n1939 ) ;
  assign n3709 = ~n2068 & n3708 ;
  assign n3710 = n3709 ^ n2897 ^ 1'b0 ;
  assign n3711 = n1314 | n1987 ;
  assign n3712 = n3711 ^ n1423 ^ 1'b0 ;
  assign n3713 = n3712 ^ n1248 ^ 1'b0 ;
  assign n3714 = n2760 & n3713 ;
  assign n3715 = ( n623 & ~n3710 ) | ( n623 & n3714 ) | ( ~n3710 & n3714 ) ;
  assign n3716 = ( x177 & ~n757 ) | ( x177 & n803 ) | ( ~n757 & n803 ) ;
  assign n3717 = ( n2032 & ~n3351 ) | ( n2032 & n3716 ) | ( ~n3351 & n3716 ) ;
  assign n3718 = n3148 & n3631 ;
  assign n3719 = ~x26 & n3718 ;
  assign n3720 = n3719 ^ n3192 ^ 1'b0 ;
  assign n3721 = n3717 & ~n3720 ;
  assign n3722 = ~n644 & n2763 ;
  assign n3723 = n2509 ^ n913 ^ n859 ;
  assign n3724 = n3146 & n3723 ;
  assign n3725 = n2742 ^ n2225 ^ n2215 ;
  assign n3726 = n949 | n3176 ;
  assign n3727 = ( ~n403 & n1012 ) | ( ~n403 & n2539 ) | ( n1012 & n2539 ) ;
  assign n3728 = ( ~n1395 & n1921 ) | ( ~n1395 & n3727 ) | ( n1921 & n3727 ) ;
  assign n3729 = ( n1272 & n2961 ) | ( n1272 & n3728 ) | ( n2961 & n3728 ) ;
  assign n3730 = x242 & n3729 ;
  assign n3731 = n591 | n2506 ;
  assign n3737 = ( ~n861 & n922 ) | ( ~n861 & n2929 ) | ( n922 & n2929 ) ;
  assign n3738 = n774 ^ n290 ^ 1'b0 ;
  assign n3739 = n3737 & n3738 ;
  assign n3734 = n2305 ^ n2032 ^ 1'b0 ;
  assign n3735 = n1042 | n3734 ;
  assign n3732 = ~n468 & n863 ;
  assign n3733 = n1496 & ~n3732 ;
  assign n3736 = n3735 ^ n3733 ^ 1'b0 ;
  assign n3740 = n3739 ^ n3736 ^ 1'b0 ;
  assign n3744 = ( x244 & n1649 ) | ( x244 & n3317 ) | ( n1649 & n3317 ) ;
  assign n3741 = n440 | n2523 ;
  assign n3742 = n1703 & ~n3741 ;
  assign n3743 = ( x86 & n2904 ) | ( x86 & n3742 ) | ( n2904 & n3742 ) ;
  assign n3745 = n3744 ^ n3743 ^ 1'b0 ;
  assign n3746 = n3745 ^ n2277 ^ 1'b0 ;
  assign n3747 = n2222 & ~n3746 ;
  assign n3748 = x161 & n385 ;
  assign n3749 = n1853 & n3748 ;
  assign n3750 = n688 ^ x151 ^ x91 ;
  assign n3751 = ( ~n1201 & n3749 ) | ( ~n1201 & n3750 ) | ( n3749 & n3750 ) ;
  assign n3754 = n3633 ^ n1655 ^ 1'b0 ;
  assign n3755 = n1265 & ~n3754 ;
  assign n3752 = n320 & ~n1611 ;
  assign n3753 = n3752 ^ n1179 ^ 1'b0 ;
  assign n3756 = n3755 ^ n3753 ^ n1063 ;
  assign n3757 = n1511 & n1641 ;
  assign n3758 = n3757 ^ n1867 ^ 1'b0 ;
  assign n3759 = n950 ^ n412 ^ n366 ;
  assign n3760 = n3758 | n3759 ;
  assign n3761 = n3760 ^ n1013 ^ 1'b0 ;
  assign n3762 = n3761 ^ n1653 ^ n1416 ;
  assign n3763 = n3535 ^ n2145 ^ 1'b0 ;
  assign n3764 = ( ~n1385 & n3762 ) | ( ~n1385 & n3763 ) | ( n3762 & n3763 ) ;
  assign n3765 = n1742 | n1778 ;
  assign n3766 = n3765 ^ n2297 ^ 1'b0 ;
  assign n3767 = n938 & n3766 ;
  assign n3768 = ( n926 & n1607 ) | ( n926 & n3767 ) | ( n1607 & n3767 ) ;
  assign n3769 = x252 & n774 ;
  assign n3770 = n3769 ^ n1018 ^ 1'b0 ;
  assign n3771 = x5 | n3770 ;
  assign n3772 = n3661 ^ n658 ^ 1'b0 ;
  assign n3773 = x197 & ~n3772 ;
  assign n3775 = n1174 & n2444 ;
  assign n3774 = n3078 ^ n804 ^ x25 ;
  assign n3776 = n3775 ^ n3774 ^ 1'b0 ;
  assign n3777 = n2771 ^ x15 ^ 1'b0 ;
  assign n3778 = n2155 & n3777 ;
  assign n3779 = ~n3776 & n3778 ;
  assign n3780 = n2993 ^ n2197 ^ 1'b0 ;
  assign n3781 = n1739 & ~n3780 ;
  assign n3782 = ( n649 & ~n2444 ) | ( n649 & n2884 ) | ( ~n2444 & n2884 ) ;
  assign n3789 = n1718 ^ n785 ^ 1'b0 ;
  assign n3783 = n358 | n1088 ;
  assign n3784 = n1940 | n3783 ;
  assign n3785 = n1950 | n2355 ;
  assign n3786 = n3784 | n3785 ;
  assign n3787 = n385 & ~n915 ;
  assign n3788 = ~n3786 & n3787 ;
  assign n3790 = n3789 ^ n3788 ^ n1630 ;
  assign n3791 = ( n1037 & ~n2767 ) | ( n1037 & n2825 ) | ( ~n2767 & n2825 ) ;
  assign n3792 = n1442 & n2236 ;
  assign n3793 = n2731 ^ n1320 ^ 1'b0 ;
  assign n3794 = n495 | n3793 ;
  assign n3795 = n3794 ^ x158 ^ 1'b0 ;
  assign n3796 = n3669 ^ n2140 ^ 1'b0 ;
  assign n3797 = n895 | n3047 ;
  assign n3798 = n3254 ^ n2733 ^ x132 ;
  assign n3799 = ~n3797 & n3798 ;
  assign n3800 = n3799 ^ n998 ^ 1'b0 ;
  assign n3801 = x187 & ~n2943 ;
  assign n3802 = n3801 ^ n351 ^ 1'b0 ;
  assign n3803 = n2515 & n3802 ;
  assign n3804 = n3800 & ~n3803 ;
  assign n3805 = n326 | n3804 ;
  assign n3806 = n3805 ^ n384 ^ 1'b0 ;
  assign n3807 = n1048 & n1766 ;
  assign n3808 = n3807 ^ x50 ^ 1'b0 ;
  assign n3809 = n3808 ^ n959 ^ 1'b0 ;
  assign n3810 = n1364 | n3809 ;
  assign n3811 = n589 & n1067 ;
  assign n3812 = ~n1213 & n3811 ;
  assign n3813 = ( ~n298 & n386 ) | ( ~n298 & n413 ) | ( n386 & n413 ) ;
  assign n3814 = ( n838 & n1347 ) | ( n838 & ~n3813 ) | ( n1347 & ~n3813 ) ;
  assign n3815 = n3471 & n3814 ;
  assign n3816 = n3815 ^ n514 ^ 1'b0 ;
  assign n3817 = n3816 ^ n1615 ^ n1343 ;
  assign n3818 = n1069 ^ n608 ^ 1'b0 ;
  assign n3819 = ~n3817 & n3818 ;
  assign n3820 = ( n3810 & ~n3812 ) | ( n3810 & n3819 ) | ( ~n3812 & n3819 ) ;
  assign n3821 = n3820 ^ n1047 ^ x198 ;
  assign n3822 = n1570 | n3413 ;
  assign n3823 = n3822 ^ n1435 ^ 1'b0 ;
  assign n3824 = n310 | n1661 ;
  assign n3825 = n3824 ^ n1632 ^ 1'b0 ;
  assign n3826 = ( ~n3566 & n3632 ) | ( ~n3566 & n3825 ) | ( n3632 & n3825 ) ;
  assign n3827 = ~n3252 & n3826 ;
  assign n3828 = ~n2942 & n3827 ;
  assign n3829 = n3788 | n3828 ;
  assign n3830 = n3657 | n3829 ;
  assign n3831 = ~n1724 & n1736 ;
  assign n3832 = n1412 ^ n292 ^ 1'b0 ;
  assign n3833 = ~n3831 & n3832 ;
  assign n3834 = n3833 ^ n574 ^ 1'b0 ;
  assign n3835 = n859 | n3834 ;
  assign n3836 = ~n1772 & n3835 ;
  assign n3837 = n3526 ^ n3304 ^ 1'b0 ;
  assign n3838 = ~n2049 & n3471 ;
  assign n3839 = n3838 ^ n3408 ^ 1'b0 ;
  assign n3840 = ( x64 & ~n982 ) | ( x64 & n3839 ) | ( ~n982 & n3839 ) ;
  assign n3841 = n1593 & n1999 ;
  assign n3842 = n3841 ^ n1292 ^ 1'b0 ;
  assign n3846 = n1067 & ~n1286 ;
  assign n3847 = n3846 ^ n540 ^ 1'b0 ;
  assign n3843 = ( x196 & ~n1076 ) | ( x196 & n1955 ) | ( ~n1076 & n1955 ) ;
  assign n3844 = ~n1150 & n3843 ;
  assign n3845 = n3844 ^ n305 ^ 1'b0 ;
  assign n3848 = n3847 ^ n3845 ^ 1'b0 ;
  assign n3849 = n2267 ^ n341 ^ 1'b0 ;
  assign n3850 = n1110 ^ n892 ^ 1'b0 ;
  assign n3851 = x71 & ~n3850 ;
  assign n3852 = n3851 ^ n2657 ^ 1'b0 ;
  assign n3853 = n3849 & ~n3852 ;
  assign n3854 = ( ~n1118 & n1734 ) | ( ~n1118 & n3409 ) | ( n1734 & n3409 ) ;
  assign n3855 = ~n2315 & n3854 ;
  assign n3858 = n1474 ^ x174 ^ 1'b0 ;
  assign n3857 = ( n1569 & n2890 ) | ( n1569 & ~n3192 ) | ( n2890 & ~n3192 ) ;
  assign n3856 = n1835 ^ n971 ^ 1'b0 ;
  assign n3859 = n3858 ^ n3857 ^ n3856 ;
  assign n3861 = n344 & ~n1611 ;
  assign n3862 = n269 & n3861 ;
  assign n3863 = x165 & ~n3862 ;
  assign n3864 = n3863 ^ n2730 ^ 1'b0 ;
  assign n3860 = ~n2657 & n3678 ;
  assign n3865 = n3864 ^ n3860 ^ 1'b0 ;
  assign n3866 = ( x132 & n503 ) | ( x132 & n2522 ) | ( n503 & n2522 ) ;
  assign n3867 = n464 | n3866 ;
  assign n3868 = n263 | n3867 ;
  assign n3869 = ( ~n873 & n2346 ) | ( ~n873 & n3868 ) | ( n2346 & n3868 ) ;
  assign n3871 = x47 & ~n1034 ;
  assign n3872 = n1689 & n3871 ;
  assign n3870 = n271 & ~n675 ;
  assign n3873 = n3872 ^ n3870 ^ 1'b0 ;
  assign n3874 = n3873 ^ n1172 ^ 1'b0 ;
  assign n3875 = n1364 & ~n1470 ;
  assign n3876 = x63 & ~n3875 ;
  assign n3877 = ~n2266 & n3876 ;
  assign n3878 = n1208 & ~n1301 ;
  assign n3879 = n2033 | n3878 ;
  assign n3880 = n3877 & ~n3879 ;
  assign n3881 = n2814 ^ n665 ^ n293 ;
  assign n3882 = ~n2553 & n3004 ;
  assign n3883 = ~n1644 & n3882 ;
  assign n3884 = n3883 ^ n1727 ^ 1'b0 ;
  assign n3885 = n3439 & n3884 ;
  assign n3886 = ~n2772 & n3885 ;
  assign n3887 = ~n3881 & n3886 ;
  assign n3888 = n1479 & ~n2840 ;
  assign n3889 = n3888 ^ n1598 ^ 1'b0 ;
  assign n3890 = n2642 & ~n2658 ;
  assign n3891 = ~n1958 & n3890 ;
  assign n3895 = n387 & n3551 ;
  assign n3896 = n3895 ^ n1312 ^ 1'b0 ;
  assign n3897 = n1910 & ~n3896 ;
  assign n3898 = n3897 ^ n665 ^ 1'b0 ;
  assign n3892 = n1082 | n1918 ;
  assign n3893 = n3892 ^ n3165 ^ x81 ;
  assign n3894 = n2279 & ~n3893 ;
  assign n3899 = n3898 ^ n3894 ^ n935 ;
  assign n3900 = n3234 ^ n620 ^ 1'b0 ;
  assign n3901 = ~n902 & n1178 ;
  assign n3902 = n3901 ^ n901 ^ 1'b0 ;
  assign n3903 = n2279 & n3902 ;
  assign n3904 = ~n2705 & n3903 ;
  assign n3905 = ( ~n1103 & n1830 ) | ( ~n1103 & n3369 ) | ( n1830 & n3369 ) ;
  assign n3906 = ~n1555 & n3905 ;
  assign n3907 = n3904 & n3906 ;
  assign n3908 = n409 | n3025 ;
  assign n3909 = n3908 ^ x53 ^ 1'b0 ;
  assign n3910 = ( n275 & n656 ) | ( n275 & n1189 ) | ( n656 & n1189 ) ;
  assign n3911 = n3909 & ~n3910 ;
  assign n3912 = ~n3327 & n3911 ;
  assign n3913 = x81 & ~n533 ;
  assign n3914 = ~n3261 & n3913 ;
  assign n3915 = ( n1021 & n1501 ) | ( n1021 & n3716 ) | ( n1501 & n3716 ) ;
  assign n3916 = n2430 & ~n3915 ;
  assign n3917 = n2287 & n3916 ;
  assign n3918 = n1863 | n3917 ;
  assign n3919 = n3914 & ~n3918 ;
  assign n3922 = ( ~n507 & n540 ) | ( ~n507 & n677 ) | ( n540 & n677 ) ;
  assign n3920 = x21 & ~x159 ;
  assign n3921 = n790 & ~n3920 ;
  assign n3923 = n3922 ^ n3921 ^ 1'b0 ;
  assign n3924 = n1525 & ~n1993 ;
  assign n3925 = n3637 | n3924 ;
  assign n3926 = n398 & ~n3925 ;
  assign n3930 = n428 & ~n1021 ;
  assign n3931 = n3930 ^ x150 ^ 1'b0 ;
  assign n3927 = n273 | n3263 ;
  assign n3928 = n3927 ^ n997 ^ 1'b0 ;
  assign n3929 = ~n3566 & n3928 ;
  assign n3932 = n3931 ^ n3929 ^ 1'b0 ;
  assign n3933 = n2991 ^ n922 ^ 1'b0 ;
  assign n3934 = ~n2028 & n3933 ;
  assign n3935 = ( ~n829 & n1257 ) | ( ~n829 & n3934 ) | ( n1257 & n3934 ) ;
  assign n3936 = ( n644 & ~n1758 ) | ( n644 & n3935 ) | ( ~n1758 & n3935 ) ;
  assign n3937 = n1046 & n3936 ;
  assign n3938 = n3932 & n3937 ;
  assign n3939 = n3938 ^ n1082 ^ x116 ;
  assign n3940 = n2523 | n2626 ;
  assign n3941 = n3940 ^ n3523 ^ n1882 ;
  assign n3942 = n562 & n1132 ;
  assign n3943 = n787 & n3942 ;
  assign n3944 = n3943 ^ n1707 ^ n629 ;
  assign n3946 = n1152 & n3109 ;
  assign n3947 = n3946 ^ n1023 ^ 1'b0 ;
  assign n3948 = n3947 ^ n270 ^ 1'b0 ;
  assign n3945 = n3011 ^ n2054 ^ n1705 ;
  assign n3949 = n3948 ^ n3945 ^ n1695 ;
  assign n3950 = n1893 & n2939 ;
  assign n3951 = x224 & ~n3950 ;
  assign n3952 = n3951 ^ n2287 ^ 1'b0 ;
  assign n3953 = n3144 | n3952 ;
  assign n3954 = n1044 ^ x186 ^ x92 ;
  assign n3955 = n3954 ^ n3391 ^ n1234 ;
  assign n3956 = x52 | n782 ;
  assign n3957 = ~n2157 & n3956 ;
  assign n3958 = n3957 ^ n1494 ^ 1'b0 ;
  assign n3959 = ( n1928 & ~n3955 ) | ( n1928 & n3958 ) | ( ~n3955 & n3958 ) ;
  assign n3960 = n3615 ^ n774 ^ x193 ;
  assign n3962 = n1722 ^ n515 ^ 1'b0 ;
  assign n3961 = n2179 ^ n2032 ^ n1199 ;
  assign n3963 = n3962 ^ n3961 ^ n2786 ;
  assign n3964 = n3893 ^ x41 ^ 1'b0 ;
  assign n3965 = n3015 & n3964 ;
  assign n3966 = n3074 ^ n428 ^ 1'b0 ;
  assign n3967 = n2490 ^ n1393 ^ x48 ;
  assign n3968 = n926 & ~n2387 ;
  assign n3969 = n2977 & n3968 ;
  assign n3970 = n1267 ^ n708 ^ x112 ;
  assign n3971 = n3970 ^ n1989 ^ 1'b0 ;
  assign n3972 = n1444 & n3971 ;
  assign n3973 = ~n3969 & n3972 ;
  assign n3974 = ~x125 & n3973 ;
  assign n3975 = ( ~x49 & n419 ) | ( ~x49 & n1183 ) | ( n419 & n1183 ) ;
  assign n3976 = n563 ^ n363 ^ 1'b0 ;
  assign n3977 = n3975 | n3976 ;
  assign n3978 = ( n3967 & ~n3974 ) | ( n3967 & n3977 ) | ( ~n3974 & n3977 ) ;
  assign n3979 = ~n341 & n2499 ;
  assign n3980 = n3979 ^ n1416 ^ 1'b0 ;
  assign n3984 = n1405 & ~n2244 ;
  assign n3982 = ~n572 & n1269 ;
  assign n3983 = ( n761 & n1737 ) | ( n761 & n3982 ) | ( n1737 & n3982 ) ;
  assign n3981 = n2219 ^ n1806 ^ 1'b0 ;
  assign n3985 = n3984 ^ n3983 ^ n3981 ;
  assign n3986 = n3985 ^ n2679 ^ n1678 ;
  assign n3987 = ( ~x70 & n2744 ) | ( ~x70 & n3010 ) | ( n2744 & n3010 ) ;
  assign n3988 = x236 & ~n2185 ;
  assign n3989 = n3364 & n3988 ;
  assign n3990 = n3814 ^ n3182 ^ 1'b0 ;
  assign n3991 = n2095 ^ n1123 ^ 1'b0 ;
  assign n3992 = n512 & n2517 ;
  assign n3993 = ~n390 & n2678 ;
  assign n3994 = n3993 ^ n464 ^ 1'b0 ;
  assign n3995 = ( n1350 & n3992 ) | ( n1350 & n3994 ) | ( n3992 & n3994 ) ;
  assign n3996 = n2204 ^ n1979 ^ n913 ;
  assign n3997 = ~n3875 & n3996 ;
  assign n3998 = n3997 ^ n3923 ^ n3332 ;
  assign n3999 = n2964 ^ x140 ^ 1'b0 ;
  assign n4000 = n412 & n2656 ;
  assign n4001 = ~n1644 & n4000 ;
  assign n4002 = n1009 | n4001 ;
  assign n4003 = n1486 | n4002 ;
  assign n4004 = ( n1136 & n3237 ) | ( n1136 & n4003 ) | ( n3237 & n4003 ) ;
  assign n4005 = n1778 ^ n1000 ^ 1'b0 ;
  assign n4006 = n604 | n2461 ;
  assign n4007 = n574 ^ x92 ^ 1'b0 ;
  assign n4008 = n4007 ^ n3912 ^ n2445 ;
  assign n4012 = n877 & n1976 ;
  assign n4013 = x202 & n4012 ;
  assign n4014 = n1458 ^ n1359 ^ n804 ;
  assign n4015 = n547 & ~n4014 ;
  assign n4016 = n4015 ^ x47 ^ 1'b0 ;
  assign n4017 = n4013 | n4016 ;
  assign n4018 = x251 | n4017 ;
  assign n4009 = n2566 ^ n2021 ^ 1'b0 ;
  assign n4010 = ~n1503 & n4009 ;
  assign n4011 = n4010 ^ n3165 ^ 1'b0 ;
  assign n4019 = n4018 ^ n4011 ^ n1418 ;
  assign n4020 = ( ~x47 & n684 ) | ( ~x47 & n1000 ) | ( n684 & n1000 ) ;
  assign n4021 = n1976 & n2634 ;
  assign n4022 = n3123 & n4021 ;
  assign n4023 = n4020 | n4022 ;
  assign n4024 = n4023 ^ n3873 ^ 1'b0 ;
  assign n4025 = ~n351 & n1369 ;
  assign n4026 = n4025 ^ n1727 ^ 1'b0 ;
  assign n4027 = n1324 & ~n2809 ;
  assign n4028 = n481 & n1569 ;
  assign n4029 = ~n4027 & n4028 ;
  assign n4030 = n4026 & ~n4029 ;
  assign n4031 = ~n4024 & n4030 ;
  assign n4032 = n1354 & n2762 ;
  assign n4033 = ( n335 & ~n377 ) | ( n335 & n1959 ) | ( ~n377 & n1959 ) ;
  assign n4034 = n4033 ^ n1795 ^ n1392 ;
  assign n4035 = n4034 ^ n2590 ^ 1'b0 ;
  assign n4036 = ~n1617 & n4035 ;
  assign n4037 = ~n1784 & n1843 ;
  assign n4038 = ~n802 & n4037 ;
  assign n4039 = ( n1637 & ~n2936 ) | ( n1637 & n4038 ) | ( ~n2936 & n4038 ) ;
  assign n4040 = n577 | n3408 ;
  assign n4041 = n4040 ^ n825 ^ 1'b0 ;
  assign n4042 = n4041 ^ n2275 ^ 1'b0 ;
  assign n4043 = n2367 & n4042 ;
  assign n4044 = n766 ^ n365 ^ 1'b0 ;
  assign n4045 = x150 & n4044 ;
  assign n4046 = n1363 & ~n4045 ;
  assign n4047 = n4046 ^ n1931 ^ n572 ;
  assign n4048 = ( n2209 & n2240 ) | ( n2209 & ~n3557 ) | ( n2240 & ~n3557 ) ;
  assign n4049 = n3020 ^ n922 ^ n591 ;
  assign n4050 = n823 & ~n1812 ;
  assign n4051 = n257 | n2914 ;
  assign n4052 = n1818 | n4051 ;
  assign n4053 = ( n805 & ~n3310 ) | ( n805 & n4052 ) | ( ~n3310 & n4052 ) ;
  assign n4054 = n4053 ^ n2253 ^ 1'b0 ;
  assign n4055 = x83 & ~n4054 ;
  assign n4056 = n2551 & n3304 ;
  assign n4058 = x226 & n522 ;
  assign n4059 = n1669 & n4058 ;
  assign n4057 = n2583 | n3154 ;
  assign n4060 = n4059 ^ n4057 ^ 1'b0 ;
  assign n4061 = n2548 ^ n1702 ^ x26 ;
  assign n4062 = n2523 ^ n303 ^ 1'b0 ;
  assign n4063 = n1500 & n4062 ;
  assign n4064 = n4063 ^ n2217 ^ 1'b0 ;
  assign n4065 = ~n4061 & n4064 ;
  assign n4066 = ~n740 & n2733 ;
  assign n4067 = ~n294 & n4066 ;
  assign n4068 = ( n1045 & n2242 ) | ( n1045 & n4067 ) | ( n2242 & n4067 ) ;
  assign n4069 = n4068 ^ n1323 ^ n843 ;
  assign n4070 = ( x210 & n1093 ) | ( x210 & n4069 ) | ( n1093 & n4069 ) ;
  assign n4071 = n3271 ^ n1971 ^ x59 ;
  assign n4072 = x214 & n4071 ;
  assign n4073 = n4072 ^ n2733 ^ 1'b0 ;
  assign n4074 = n3599 & n4073 ;
  assign n4078 = n1284 ^ n630 ^ x96 ;
  assign n4079 = ( n2517 & n2860 ) | ( n2517 & ~n4078 ) | ( n2860 & ~n4078 ) ;
  assign n4075 = n1805 ^ n861 ^ 1'b0 ;
  assign n4076 = n2408 & n4075 ;
  assign n4077 = n3510 & n4076 ;
  assign n4080 = n4079 ^ n4077 ^ 1'b0 ;
  assign n4081 = n4080 ^ n2422 ^ 1'b0 ;
  assign n4082 = n3749 ^ n427 ^ 1'b0 ;
  assign n4083 = ~n1229 & n4082 ;
  assign n4084 = n1104 ^ n495 ^ n277 ;
  assign n4085 = n4084 ^ n1262 ^ n824 ;
  assign n4086 = n4085 ^ n1817 ^ 1'b0 ;
  assign n4087 = n2680 ^ n2520 ^ 1'b0 ;
  assign n4088 = n1265 & n4087 ;
  assign n4089 = n1018 ^ n857 ^ 1'b0 ;
  assign n4090 = n2532 ^ n1064 ^ 1'b0 ;
  assign n4091 = n1752 ^ n1671 ^ n629 ;
  assign n4092 = n868 & n3984 ;
  assign n4093 = n4092 ^ n2439 ^ 1'b0 ;
  assign n4094 = n1470 | n3940 ;
  assign n4096 = ~n1828 & n2687 ;
  assign n4097 = n4096 ^ n956 ^ 1'b0 ;
  assign n4095 = n1853 ^ n902 ^ n527 ;
  assign n4098 = n4097 ^ n4095 ^ n3637 ;
  assign n4099 = n4098 ^ n1999 ^ 1'b0 ;
  assign n4100 = n794 & n4099 ;
  assign n4101 = n4100 ^ n4009 ^ 1'b0 ;
  assign n4102 = ~n4094 & n4101 ;
  assign n4103 = n1719 & n4102 ;
  assign n4104 = n3614 ^ n2286 ^ n1653 ;
  assign n4110 = n3494 ^ n994 ^ 1'b0 ;
  assign n4111 = n3932 & ~n4110 ;
  assign n4108 = n710 ^ x65 ^ 1'b0 ;
  assign n4105 = n432 ^ x133 ^ 1'b0 ;
  assign n4106 = n1895 & ~n4105 ;
  assign n4107 = n4106 ^ n2116 ^ 1'b0 ;
  assign n4109 = n4108 ^ n4107 ^ n1582 ;
  assign n4112 = n4111 ^ n4109 ^ 1'b0 ;
  assign n4113 = ( n1208 & n1906 ) | ( n1208 & n2245 ) | ( n1906 & n2245 ) ;
  assign n4114 = n813 & n1120 ;
  assign n4115 = n1031 | n1492 ;
  assign n4116 = n4115 ^ n3494 ^ 1'b0 ;
  assign n4117 = n4114 | n4116 ;
  assign n4118 = ( n640 & n1050 ) | ( n640 & n1809 ) | ( n1050 & n1809 ) ;
  assign n4119 = n2231 ^ n1949 ^ 1'b0 ;
  assign n4120 = n4118 & ~n4119 ;
  assign n4121 = ( n2259 & ~n3944 ) | ( n2259 & n4120 ) | ( ~n3944 & n4120 ) ;
  assign n4122 = n3753 ^ n1671 ^ x0 ;
  assign n4123 = ~n1955 & n4122 ;
  assign n4125 = ~n307 & n837 ;
  assign n4126 = n4125 ^ n1851 ^ 1'b0 ;
  assign n4124 = n1074 ^ n366 ^ n365 ;
  assign n4127 = n4126 ^ n4124 ^ 1'b0 ;
  assign n4128 = n3072 ^ n1628 ^ 1'b0 ;
  assign n4129 = n386 | n1105 ;
  assign n4130 = n3766 ^ n2657 ^ n1312 ;
  assign n4132 = n2441 ^ n1448 ^ 1'b0 ;
  assign n4131 = n358 | n3473 ;
  assign n4133 = n4132 ^ n4131 ^ 1'b0 ;
  assign n4137 = n2724 & ~n3309 ;
  assign n4134 = ~n440 & n3563 ;
  assign n4135 = x114 & n2282 ;
  assign n4136 = n4134 & n4135 ;
  assign n4138 = n4137 ^ n4136 ^ 1'b0 ;
  assign n4139 = n4105 ^ x14 ^ 1'b0 ;
  assign n4140 = n3207 & ~n4139 ;
  assign n4141 = n4140 ^ n3469 ^ n3100 ;
  assign n4142 = x25 & n1220 ;
  assign n4143 = n4142 ^ n345 ^ 1'b0 ;
  assign n4144 = ~n3874 & n4143 ;
  assign n4145 = n2570 & ~n2977 ;
  assign n4146 = ~n1694 & n4145 ;
  assign n4147 = n4146 ^ n769 ^ 1'b0 ;
  assign n4148 = n410 & ~n1727 ;
  assign n4149 = ( n559 & n1647 ) | ( n559 & n2679 ) | ( n1647 & n2679 ) ;
  assign n4150 = x226 & ~n665 ;
  assign n4151 = ( ~n2517 & n4149 ) | ( ~n2517 & n4150 ) | ( n4149 & n4150 ) ;
  assign n4152 = ~n1933 & n4151 ;
  assign n4153 = ~n4148 & n4152 ;
  assign n4154 = n2931 ^ n727 ^ x26 ;
  assign n4155 = n4154 ^ n1179 ^ x147 ;
  assign n4156 = n3842 ^ n2422 ^ n554 ;
  assign n4157 = n3813 ^ n1275 ^ 1'b0 ;
  assign n4158 = ( n4155 & ~n4156 ) | ( n4155 & n4157 ) | ( ~n4156 & n4157 ) ;
  assign n4159 = n489 ^ x105 ^ 1'b0 ;
  assign n4161 = n3122 ^ x246 ^ 1'b0 ;
  assign n4162 = n804 | n4161 ;
  assign n4160 = n1256 | n2897 ;
  assign n4163 = n4162 ^ n4160 ^ 1'b0 ;
  assign n4164 = n4163 ^ n3093 ^ n795 ;
  assign n4165 = n727 & ~n4164 ;
  assign n4166 = n4159 & n4165 ;
  assign n4167 = n2566 | n4166 ;
  assign n4168 = n2549 & ~n4167 ;
  assign n4169 = n478 | n1062 ;
  assign n4170 = n2522 & ~n4169 ;
  assign n4171 = n2916 & ~n4170 ;
  assign n4172 = ~n3100 & n4171 ;
  assign n4173 = n3914 ^ n2329 ^ n599 ;
  assign n4174 = ( n1891 & n2937 ) | ( n1891 & ~n4173 ) | ( n2937 & ~n4173 ) ;
  assign n4175 = n660 & ~n1347 ;
  assign n4176 = n2648 & n4175 ;
  assign n4177 = n925 & ~n4176 ;
  assign n4178 = x54 & n514 ;
  assign n4179 = n992 & n4178 ;
  assign n4180 = n2024 | n4179 ;
  assign n4181 = n1499 & ~n1640 ;
  assign n4182 = n4180 & n4181 ;
  assign n4183 = n1944 | n2766 ;
  assign n4184 = n4183 ^ n1430 ^ 1'b0 ;
  assign n4185 = n3452 & ~n4184 ;
  assign n4186 = n1748 ^ n1331 ^ 1'b0 ;
  assign n4187 = n861 & n4186 ;
  assign n4188 = n1073 & n4187 ;
  assign n4189 = n4188 ^ n3433 ^ 1'b0 ;
  assign n4190 = n1405 ^ x192 ^ 1'b0 ;
  assign n4191 = n4190 ^ n1594 ^ x106 ;
  assign n4192 = n4191 ^ n2822 ^ n684 ;
  assign n4193 = n4192 ^ x45 ^ 1'b0 ;
  assign n4194 = n2496 & ~n4193 ;
  assign n4195 = ~n1537 & n4194 ;
  assign n4196 = n1517 ^ n964 ^ 1'b0 ;
  assign n4197 = n2128 & ~n4196 ;
  assign n4198 = n4197 ^ n2268 ^ 1'b0 ;
  assign n4199 = n2294 ^ n1836 ^ x227 ;
  assign n4202 = n981 ^ x183 ^ 1'b0 ;
  assign n4201 = x115 & ~n967 ;
  assign n4203 = n4202 ^ n4201 ^ 1'b0 ;
  assign n4200 = ~x29 & x37 ;
  assign n4204 = n4203 ^ n4200 ^ 1'b0 ;
  assign n4205 = n467 | n4204 ;
  assign n4206 = n4205 ^ n3461 ^ 1'b0 ;
  assign n4207 = n4206 ^ n4170 ^ n4022 ;
  assign n4208 = n3272 | n4207 ;
  assign n4209 = n4208 ^ x114 ^ 1'b0 ;
  assign n4210 = n2182 ^ n1880 ^ n951 ;
  assign n4211 = n2196 ^ n1393 ^ 1'b0 ;
  assign n4212 = n4210 & ~n4211 ;
  assign n4214 = n3327 ^ n3012 ^ 1'b0 ;
  assign n4213 = n1508 & ~n1636 ;
  assign n4215 = n4214 ^ n4213 ^ 1'b0 ;
  assign n4216 = n1793 ^ x175 ^ 1'b0 ;
  assign n4217 = ( x244 & ~n4215 ) | ( x244 & n4216 ) | ( ~n4215 & n4216 ) ;
  assign n4218 = ~n354 & n3708 ;
  assign n4219 = n4218 ^ n1632 ^ 1'b0 ;
  assign n4220 = ( n1140 & n2831 ) | ( n1140 & n4219 ) | ( n2831 & n4219 ) ;
  assign n4221 = n1716 & n3198 ;
  assign n4222 = n4104 ^ n2868 ^ 1'b0 ;
  assign n4223 = n4221 & ~n4222 ;
  assign n4224 = n1334 ^ x120 ^ 1'b0 ;
  assign n4225 = n4224 ^ n2270 ^ 1'b0 ;
  assign n4226 = n2314 & ~n4225 ;
  assign n4227 = n1881 & n4226 ;
  assign n4228 = n417 & n1541 ;
  assign n4229 = ( n1021 & n1142 ) | ( n1021 & n4228 ) | ( n1142 & n4228 ) ;
  assign n4230 = n1120 & ~n3957 ;
  assign n4231 = n1983 ^ n1746 ^ 1'b0 ;
  assign n4232 = n3199 & n4231 ;
  assign n4233 = n1225 & n4232 ;
  assign n4234 = ( ~x14 & n790 ) | ( ~x14 & n2248 ) | ( n790 & n2248 ) ;
  assign n4235 = n3245 & ~n4234 ;
  assign n4236 = n2140 & n4235 ;
  assign n4237 = n2201 ^ n1835 ^ 1'b0 ;
  assign n4238 = x165 & ~n840 ;
  assign n4239 = n4237 & n4238 ;
  assign n4240 = n4239 ^ n3866 ^ n1206 ;
  assign n4241 = n4240 ^ n3376 ^ x4 ;
  assign n4242 = n1357 & n4095 ;
  assign n4243 = n2585 & ~n4242 ;
  assign n4244 = ( n1081 & n2126 ) | ( n1081 & ~n2394 ) | ( n2126 & ~n2394 ) ;
  assign n4245 = n323 & ~n4244 ;
  assign n4246 = n312 | n1108 ;
  assign n4247 = n2929 & ~n4246 ;
  assign n4248 = n1543 ^ n1394 ^ 1'b0 ;
  assign n4249 = ~n4247 & n4248 ;
  assign n4250 = ~n1429 & n4249 ;
  assign n4251 = n4250 ^ n2133 ^ 1'b0 ;
  assign n4252 = ~n565 & n3002 ;
  assign n4253 = n4252 ^ n4108 ^ 1'b0 ;
  assign n4254 = n4253 ^ n2835 ^ n2102 ;
  assign n4255 = ( n481 & ~n2212 ) | ( n481 & n4254 ) | ( ~n2212 & n4254 ) ;
  assign n4256 = n2451 ^ x25 ^ 1'b0 ;
  assign n4257 = n2894 ^ n1977 ^ n1812 ;
  assign n4258 = n4257 ^ n4177 ^ 1'b0 ;
  assign n4259 = n2675 ^ n769 ^ 1'b0 ;
  assign n4260 = n2526 | n4259 ;
  assign n4261 = n4260 ^ n4180 ^ 1'b0 ;
  assign n4266 = n3056 ^ n2506 ^ 1'b0 ;
  assign n4267 = n3010 | n3283 ;
  assign n4268 = n1115 & ~n4267 ;
  assign n4269 = ~n4266 & n4268 ;
  assign n4262 = ~n2165 & n3072 ;
  assign n4263 = ~n371 & n4262 ;
  assign n4264 = ( n1933 & n4142 ) | ( n1933 & n4263 ) | ( n4142 & n4263 ) ;
  assign n4265 = n4264 ^ n2407 ^ n2057 ;
  assign n4270 = n4269 ^ n4265 ^ n920 ;
  assign n4271 = ( x190 & n955 ) | ( x190 & ~n4270 ) | ( n955 & ~n4270 ) ;
  assign n4272 = x178 & n2551 ;
  assign n4273 = ~x227 & n4272 ;
  assign n4274 = n3151 ^ n1123 ^ n266 ;
  assign n4275 = n774 & n4274 ;
  assign n4276 = n4275 ^ n1347 ^ 1'b0 ;
  assign n4285 = ( ~x28 & n1264 ) | ( ~x28 & n2128 ) | ( n1264 & n2128 ) ;
  assign n4279 = n305 | n349 ;
  assign n4280 = n4279 ^ n512 ^ 1'b0 ;
  assign n4281 = ~n1534 & n4280 ;
  assign n4282 = ~n1907 & n4281 ;
  assign n4277 = n2009 ^ n763 ^ 1'b0 ;
  assign n4278 = n4277 ^ n932 ^ 1'b0 ;
  assign n4283 = n4282 ^ n4278 ^ n3074 ;
  assign n4284 = ~n958 & n4283 ;
  assign n4286 = n4285 ^ n4284 ^ 1'b0 ;
  assign n4287 = n4276 & ~n4286 ;
  assign n4288 = ( n1274 & ~n4162 ) | ( n1274 & n4287 ) | ( ~n4162 & n4287 ) ;
  assign n4289 = ~n316 & n1060 ;
  assign n4290 = n4289 ^ n374 ^ 1'b0 ;
  assign n4291 = n4191 ^ n1369 ^ 1'b0 ;
  assign n4292 = n3361 & n3793 ;
  assign n4293 = n4291 & n4292 ;
  assign n4294 = ( n2414 & n4290 ) | ( n2414 & ~n4293 ) | ( n4290 & ~n4293 ) ;
  assign n4295 = n1505 ^ n807 ^ 1'b0 ;
  assign n4296 = n1136 | n4295 ;
  assign n4297 = n1475 | n4296 ;
  assign n4298 = n4297 ^ n1369 ^ 1'b0 ;
  assign n4299 = x113 & ~n4298 ;
  assign n4300 = n3045 ^ n1585 ^ 1'b0 ;
  assign n4301 = n4300 ^ n1499 ^ n369 ;
  assign n4302 = n1039 | n4114 ;
  assign n4303 = n4302 ^ n2692 ^ n432 ;
  assign n4304 = n2626 ^ n764 ^ n647 ;
  assign n4305 = n3302 & n3899 ;
  assign n4306 = ( n2227 & n4304 ) | ( n2227 & ~n4305 ) | ( n4304 & ~n4305 ) ;
  assign n4307 = ( ~x139 & n3689 ) | ( ~x139 & n4306 ) | ( n3689 & n4306 ) ;
  assign n4308 = n864 & ~n2555 ;
  assign n4309 = n976 | n1755 ;
  assign n4310 = n2389 | n4309 ;
  assign n4311 = n3165 ^ n3062 ^ 1'b0 ;
  assign n4312 = n344 & ~n4311 ;
  assign n4313 = ~n1302 & n4312 ;
  assign n4316 = n1374 ^ n1320 ^ x251 ;
  assign n4314 = ( x87 & n1069 ) | ( x87 & n1919 ) | ( n1069 & n1919 ) ;
  assign n4315 = n3017 & ~n4314 ;
  assign n4317 = n4316 ^ n4315 ^ 1'b0 ;
  assign n4318 = n4132 ^ n957 ^ 1'b0 ;
  assign n4319 = n4318 ^ n1994 ^ 1'b0 ;
  assign n4320 = n1006 & ~n4319 ;
  assign n4321 = n4317 & n4320 ;
  assign n4322 = ~n1045 & n1478 ;
  assign n4323 = n3447 ^ n1890 ^ n1077 ;
  assign n4324 = n1588 | n4323 ;
  assign n4325 = n3928 ^ n300 ^ 1'b0 ;
  assign n4326 = ~n535 & n4325 ;
  assign n4327 = n986 ^ n360 ^ 1'b0 ;
  assign n4328 = ~n832 & n4327 ;
  assign n4329 = ~n4326 & n4328 ;
  assign n4330 = n4329 ^ n4024 ^ 1'b0 ;
  assign n4331 = n2444 ^ n1936 ^ 1'b0 ;
  assign n4332 = ~n1972 & n4331 ;
  assign n4333 = n1789 & n4332 ;
  assign n4334 = n1900 ^ n1298 ^ 1'b0 ;
  assign n4335 = n419 | n1655 ;
  assign n4336 = n1891 | n4335 ;
  assign n4342 = n691 ^ x76 ^ 1'b0 ;
  assign n4343 = n3204 ^ n3128 ^ n2878 ;
  assign n4344 = n1172 | n4343 ;
  assign n4345 = n4342 & ~n4344 ;
  assign n4337 = n505 & n1895 ;
  assign n4338 = ~n1079 & n4337 ;
  assign n4339 = n1744 ^ x155 ^ 1'b0 ;
  assign n4340 = n1327 | n4339 ;
  assign n4341 = ( n860 & ~n4338 ) | ( n860 & n4340 ) | ( ~n4338 & n4340 ) ;
  assign n4346 = n4345 ^ n4341 ^ n4277 ;
  assign n4347 = n351 | n4210 ;
  assign n4349 = n381 | n1750 ;
  assign n4350 = n4349 ^ x28 ^ 1'b0 ;
  assign n4351 = n4350 ^ n1731 ^ 1'b0 ;
  assign n4348 = n1403 & n4300 ;
  assign n4352 = n4351 ^ n4348 ^ 1'b0 ;
  assign n4353 = n1733 ^ n487 ^ 1'b0 ;
  assign n4354 = n1552 & n4353 ;
  assign n4355 = ~n2890 & n4354 ;
  assign n4356 = n1132 & n4355 ;
  assign n4357 = ( ~n1641 & n1848 ) | ( ~n1641 & n4356 ) | ( n1848 & n4356 ) ;
  assign n4358 = n989 | n4357 ;
  assign n4359 = n2680 & ~n4358 ;
  assign n4360 = n1636 | n4090 ;
  assign n4361 = n2344 & ~n4360 ;
  assign n4362 = n4304 ^ n3625 ^ 1'b0 ;
  assign n4363 = n3417 & n4362 ;
  assign n4364 = n490 | n2297 ;
  assign n4365 = ( ~x129 & x160 ) | ( ~x129 & x240 ) | ( x160 & x240 ) ;
  assign n4366 = n4365 ^ n1570 ^ 1'b0 ;
  assign n4367 = n3257 & ~n4366 ;
  assign n4368 = n2676 & n4084 ;
  assign n4369 = ~n4367 & n4368 ;
  assign n4370 = n4369 ^ n2644 ^ n667 ;
  assign n4371 = n2386 ^ n1374 ^ 1'b0 ;
  assign n4372 = n4371 ^ n1427 ^ 1'b0 ;
  assign n4373 = n1040 ^ n708 ^ 1'b0 ;
  assign n4374 = n4345 & ~n4373 ;
  assign n4377 = n1493 ^ n1450 ^ 1'b0 ;
  assign n4378 = n936 & ~n4377 ;
  assign n4375 = n540 | n2024 ;
  assign n4376 = n2435 & ~n4375 ;
  assign n4379 = n4378 ^ n4376 ^ n352 ;
  assign n4380 = n1225 ^ n766 ^ 1'b0 ;
  assign n4381 = ~n3254 & n4380 ;
  assign n4382 = ~n1124 & n4381 ;
  assign n4383 = n4382 ^ n1534 ^ 1'b0 ;
  assign n4384 = n1129 | n1377 ;
  assign n4385 = n4384 ^ n1647 ^ 1'b0 ;
  assign n4386 = n4383 & n4385 ;
  assign n4387 = n402 & n1956 ;
  assign n4388 = ~n3564 & n4387 ;
  assign n4389 = ~n273 & n967 ;
  assign n4391 = n1479 & n1751 ;
  assign n4390 = ~n1168 & n1775 ;
  assign n4392 = n4391 ^ n4390 ^ n4123 ;
  assign n4393 = n2162 ^ n1467 ^ 1'b0 ;
  assign n4394 = n4392 | n4393 ;
  assign n4395 = ( x94 & n1566 ) | ( x94 & n3649 ) | ( n1566 & n3649 ) ;
  assign n4396 = n433 & n4395 ;
  assign n4397 = n3938 ^ x66 ^ 1'b0 ;
  assign n4398 = n3985 ^ n2667 ^ x148 ;
  assign n4399 = n3659 & n4398 ;
  assign n4400 = n4399 ^ n1262 ^ 1'b0 ;
  assign n4401 = n2873 & ~n3165 ;
  assign n4402 = n4401 ^ n3500 ^ 1'b0 ;
  assign n4403 = n3982 & ~n4402 ;
  assign n4404 = ~n706 & n4403 ;
  assign n4405 = n1602 ^ n1098 ^ n771 ;
  assign n4406 = n2319 & ~n3656 ;
  assign n4407 = n4406 ^ n1030 ^ 1'b0 ;
  assign n4408 = n4405 & n4407 ;
  assign n4409 = ~n4207 & n4408 ;
  assign n4410 = n3128 & n4409 ;
  assign n4411 = n3825 & ~n4410 ;
  assign n4413 = n3409 ^ n2352 ^ 1'b0 ;
  assign n4412 = n1818 & n4088 ;
  assign n4414 = n4413 ^ n4412 ^ 1'b0 ;
  assign n4415 = n921 ^ n652 ^ 1'b0 ;
  assign n4416 = x128 & ~n4415 ;
  assign n4417 = n4416 ^ n1874 ^ n1405 ;
  assign n4418 = n1399 & n4417 ;
  assign n4419 = n3210 & n4418 ;
  assign n4420 = n632 | n3679 ;
  assign n4421 = n931 | n4420 ;
  assign n4422 = ~n377 & n4421 ;
  assign n4423 = n2362 ^ n735 ^ x165 ;
  assign n4424 = n4423 ^ n4290 ^ n759 ;
  assign n4425 = ( x234 & n1296 ) | ( x234 & ~n1993 ) | ( n1296 & ~n1993 ) ;
  assign n4426 = n4425 ^ n2107 ^ x43 ;
  assign n4427 = n2993 ^ n939 ^ 1'b0 ;
  assign n4428 = n1655 ^ n1231 ^ n1083 ;
  assign n4429 = n4428 ^ n892 ^ 1'b0 ;
  assign n4430 = n1175 & ~n4429 ;
  assign n4431 = n4430 ^ n3646 ^ 1'b0 ;
  assign n4432 = ( n2111 & ~n4287 ) | ( n2111 & n4431 ) | ( ~n4287 & n4431 ) ;
  assign n4433 = n768 | n4432 ;
  assign n4434 = n1843 ^ x90 ^ 1'b0 ;
  assign n4435 = n888 & ~n2370 ;
  assign n4436 = n4435 ^ n501 ^ 1'b0 ;
  assign n4437 = n1176 | n4436 ;
  assign n4438 = n1164 | n2932 ;
  assign n4439 = n1040 ^ n854 ^ x93 ;
  assign n4440 = n1365 | n1900 ;
  assign n4441 = n1644 | n4440 ;
  assign n4442 = x215 & n2310 ;
  assign n4443 = n4442 ^ n2868 ^ 1'b0 ;
  assign n4444 = ( x146 & n4441 ) | ( x146 & n4443 ) | ( n4441 & n4443 ) ;
  assign n4445 = x104 & ~n1961 ;
  assign n4446 = n4445 ^ n338 ^ 1'b0 ;
  assign n4447 = ~n2931 & n3661 ;
  assign n4448 = n2667 ^ n1863 ^ n821 ;
  assign n4449 = ( ~x78 & n1091 ) | ( ~x78 & n2306 ) | ( n1091 & n2306 ) ;
  assign n4450 = n3269 & ~n4449 ;
  assign n4451 = n3572 ^ n3122 ^ 1'b0 ;
  assign n4453 = n3165 ^ n2214 ^ x234 ;
  assign n4454 = n4453 ^ n3737 ^ 1'b0 ;
  assign n4452 = n425 & n2147 ;
  assign n4455 = n4454 ^ n4452 ^ 1'b0 ;
  assign n4456 = n4455 ^ n460 ^ 1'b0 ;
  assign n4457 = ( n2255 & ~n3676 ) | ( n2255 & n4456 ) | ( ~n3676 & n4456 ) ;
  assign n4458 = x210 | n1081 ;
  assign n4459 = x42 & ~n4458 ;
  assign n4460 = n464 & n4459 ;
  assign n4461 = ~n1828 & n4460 ;
  assign n4462 = n2165 & ~n3990 ;
  assign n4464 = n3393 ^ n335 ^ 1'b0 ;
  assign n4463 = ~n1789 & n3194 ;
  assign n4465 = n4464 ^ n4463 ^ 1'b0 ;
  assign n4466 = n2312 ^ n1956 ^ 1'b0 ;
  assign n4467 = ~n1989 & n4466 ;
  assign n4468 = n2601 | n4467 ;
  assign n4469 = n3470 ^ n1111 ^ x127 ;
  assign n4470 = n606 ^ x130 ^ 1'b0 ;
  assign n4471 = n4469 | n4470 ;
  assign n4472 = ~n1028 & n4471 ;
  assign n4473 = n4134 ^ n3966 ^ 1'b0 ;
  assign n4474 = n658 & ~n1962 ;
  assign n4479 = n300 & ~n1179 ;
  assign n4475 = ( ~n1320 & n2724 ) | ( ~n1320 & n3188 ) | ( n2724 & n3188 ) ;
  assign n4476 = n530 & n2064 ;
  assign n4477 = ~n609 & n4476 ;
  assign n4478 = n4475 | n4477 ;
  assign n4480 = n4479 ^ n4478 ^ 1'b0 ;
  assign n4481 = n4474 | n4480 ;
  assign n4482 = ( x162 & n1107 ) | ( x162 & ~n3797 ) | ( n1107 & ~n3797 ) ;
  assign n4483 = n4482 ^ n3704 ^ 1'b0 ;
  assign n4484 = ~n3907 & n4483 ;
  assign n4485 = n1446 ^ n387 ^ 1'b0 ;
  assign n4486 = n4024 ^ n413 ^ 1'b0 ;
  assign n4487 = n2236 & ~n4486 ;
  assign n4488 = n1522 & ~n4229 ;
  assign n4489 = n4479 & n4488 ;
  assign n4490 = ( ~n2314 & n4203 ) | ( ~n2314 & n4303 ) | ( n4203 & n4303 ) ;
  assign n4496 = x251 & n652 ;
  assign n4497 = n4496 ^ n2883 ^ 1'b0 ;
  assign n4498 = n2231 & ~n4497 ;
  assign n4491 = n1693 | n3523 ;
  assign n4492 = n4491 ^ n811 ^ 1'b0 ;
  assign n4493 = n4492 ^ n1024 ^ 1'b0 ;
  assign n4494 = ~n1465 & n4493 ;
  assign n4495 = n4494 ^ n3016 ^ 1'b0 ;
  assign n4499 = n4498 ^ n4495 ^ n3531 ;
  assign n4500 = n2297 ^ n1409 ^ n256 ;
  assign n4501 = ~n1462 & n4500 ;
  assign n4502 = n854 ^ n438 ^ 1'b0 ;
  assign n4503 = n4502 ^ n4455 ^ x3 ;
  assign n4504 = ~n4501 & n4503 ;
  assign n4505 = n4504 ^ n2885 ^ 1'b0 ;
  assign n4506 = ( x243 & ~n2317 ) | ( x243 & n3188 ) | ( ~n2317 & n3188 ) ;
  assign n4507 = n3364 ^ n432 ^ 1'b0 ;
  assign n4508 = x36 & n4507 ;
  assign n4509 = ~n892 & n3102 ;
  assign n4510 = n3069 & n4509 ;
  assign n4511 = n802 & ~n817 ;
  assign n4512 = n4511 ^ n3858 ^ 1'b0 ;
  assign n4513 = n4510 | n4512 ;
  assign n4514 = n4513 ^ n1932 ^ 1'b0 ;
  assign n4515 = n4514 ^ n4121 ^ 1'b0 ;
  assign n4516 = n539 & n3533 ;
  assign n4517 = ( n2332 & ~n3339 ) | ( n2332 & n4516 ) | ( ~n3339 & n4516 ) ;
  assign n4518 = n2297 ^ n1677 ^ 1'b0 ;
  assign n4519 = ~n4215 & n4518 ;
  assign n4520 = n3425 ^ n2986 ^ 1'b0 ;
  assign n4521 = n4519 & ~n4520 ;
  assign n4522 = n1156 | n4521 ;
  assign n4523 = n2596 & n4522 ;
  assign n4524 = n892 | n1677 ;
  assign n4525 = n4524 ^ n3742 ^ 1'b0 ;
  assign n4526 = n2301 ^ n1671 ^ 1'b0 ;
  assign n4527 = ~n4373 & n4526 ;
  assign n4528 = n1497 ^ n354 ^ 1'b0 ;
  assign n4529 = ( n1570 & n1845 ) | ( n1570 & ~n4528 ) | ( n1845 & ~n4528 ) ;
  assign n4530 = ~n1002 & n1657 ;
  assign n4531 = ~n1120 & n4530 ;
  assign n4532 = ( ~n3328 & n4529 ) | ( ~n3328 & n4531 ) | ( n4529 & n4531 ) ;
  assign n4533 = n3343 ^ n1450 ^ 1'b0 ;
  assign n4534 = n2338 | n4166 ;
  assign n4535 = n3982 | n4534 ;
  assign n4536 = x57 | n4535 ;
  assign n4537 = ~n3640 & n4008 ;
  assign n4538 = n1511 ^ n845 ^ 1'b0 ;
  assign n4539 = ( ~n2033 & n2247 ) | ( ~n2033 & n2386 ) | ( n2247 & n2386 ) ;
  assign n4540 = n2193 ^ n1972 ^ n1638 ;
  assign n4541 = n4540 ^ n2983 ^ 1'b0 ;
  assign n4542 = ( ~n4538 & n4539 ) | ( ~n4538 & n4541 ) | ( n4539 & n4541 ) ;
  assign n4543 = n1015 | n1870 ;
  assign n4544 = n4543 ^ n1846 ^ 1'b0 ;
  assign n4545 = n1655 & ~n3108 ;
  assign n4546 = n4545 ^ n3593 ^ 1'b0 ;
  assign n4547 = n4546 ^ n3502 ^ x4 ;
  assign n4548 = ~n575 & n3369 ;
  assign n4549 = n2236 & n4078 ;
  assign n4550 = n4549 ^ n3184 ^ 1'b0 ;
  assign n4551 = x70 & ~n2740 ;
  assign n4552 = n4551 ^ n4266 ^ 1'b0 ;
  assign n4553 = n4469 ^ n2908 ^ n409 ;
  assign n4554 = ~n464 & n3155 ;
  assign n4555 = ~n3418 & n4554 ;
  assign n4557 = n2983 ^ n1326 ^ n302 ;
  assign n4558 = ( n1765 & ~n3182 ) | ( n1765 & n4557 ) | ( ~n3182 & n4557 ) ;
  assign n4556 = n1806 & ~n2706 ;
  assign n4559 = n4558 ^ n4556 ^ 1'b0 ;
  assign n4560 = ~n4400 & n4559 ;
  assign n4561 = n4560 ^ n3222 ^ 1'b0 ;
  assign n4562 = x62 & ~n1079 ;
  assign n4563 = n572 & n4562 ;
  assign n4564 = n4563 ^ n1424 ^ x234 ;
  assign n4565 = n3470 ^ n2182 ^ 1'b0 ;
  assign n4566 = x69 & n4565 ;
  assign n4567 = ~n4564 & n4566 ;
  assign n4576 = n1794 ^ n1729 ^ 1'b0 ;
  assign n4577 = ~n1406 & n4576 ;
  assign n4573 = n1045 ^ x37 ^ 1'b0 ;
  assign n4574 = n982 & ~n4573 ;
  assign n4575 = n4574 ^ n2283 ^ n1145 ;
  assign n4568 = n2205 | n3172 ;
  assign n4569 = n1325 | n4568 ;
  assign n4570 = ( ~x174 & n2167 ) | ( ~x174 & n4569 ) | ( n2167 & n4569 ) ;
  assign n4571 = n4570 ^ n1390 ^ 1'b0 ;
  assign n4572 = n1760 & n4571 ;
  assign n4578 = n4577 ^ n4575 ^ n4572 ;
  assign n4579 = n3786 ^ n329 ^ 1'b0 ;
  assign n4580 = n1422 & ~n4579 ;
  assign n4581 = n1140 ^ n615 ^ n284 ;
  assign n4582 = n1879 | n4581 ;
  assign n4583 = n4247 & ~n4582 ;
  assign n4584 = n2989 | n4583 ;
  assign n4585 = n2953 & ~n4584 ;
  assign n4586 = n2394 | n4585 ;
  assign n4587 = n3883 & ~n4586 ;
  assign n4588 = ( n434 & n694 ) | ( n434 & n1447 ) | ( n694 & n1447 ) ;
  assign n4589 = ( ~x24 & n2653 ) | ( ~x24 & n4588 ) | ( n2653 & n4588 ) ;
  assign n4590 = n3758 ^ n2642 ^ n2509 ;
  assign n4591 = n4590 ^ n2701 ^ 1'b0 ;
  assign n4592 = n671 & n4591 ;
  assign n4593 = ( x137 & n449 ) | ( x137 & n1732 ) | ( n449 & n1732 ) ;
  assign n4594 = n4593 ^ n602 ^ 1'b0 ;
  assign n4595 = n678 & n4594 ;
  assign n4596 = ~n4592 & n4595 ;
  assign n4597 = n4596 ^ n1718 ^ 1'b0 ;
  assign n4598 = ~n1989 & n2090 ;
  assign n4599 = n512 & n4598 ;
  assign n4600 = n4599 ^ n3881 ^ 1'b0 ;
  assign n4601 = ( n1401 & n2636 ) | ( n1401 & ~n4476 ) | ( n2636 & ~n4476 ) ;
  assign n4602 = n1206 & ~n2205 ;
  assign n4603 = x43 & ~n4602 ;
  assign n4604 = x69 ^ x50 ^ 1'b0 ;
  assign n4605 = n4604 ^ n903 ^ 1'b0 ;
  assign n4606 = n4603 & ~n4605 ;
  assign n4608 = n655 & ~n1273 ;
  assign n4609 = n4608 ^ n614 ^ 1'b0 ;
  assign n4610 = n4609 ^ n1438 ^ 1'b0 ;
  assign n4611 = ~n1013 & n4610 ;
  assign n4607 = x65 & n1280 ;
  assign n4612 = n4611 ^ n4607 ^ 1'b0 ;
  assign n4613 = n4612 ^ n4350 ^ 1'b0 ;
  assign n4614 = x10 & ~n4613 ;
  assign n4615 = n4614 ^ n2759 ^ 1'b0 ;
  assign n4616 = x231 | n4615 ;
  assign n4618 = n264 | n483 ;
  assign n4617 = n511 & n572 ;
  assign n4619 = n4618 ^ n4617 ^ n737 ;
  assign n4620 = x150 ^ x148 ^ 1'b0 ;
  assign n4621 = n1718 & ~n4620 ;
  assign n4622 = ~n1257 & n2125 ;
  assign n4623 = n4622 ^ n2088 ^ 1'b0 ;
  assign n4624 = n1394 ^ x219 ^ 1'b0 ;
  assign n4625 = n2994 & n4624 ;
  assign n4626 = ( n4621 & n4623 ) | ( n4621 & ~n4625 ) | ( n4623 & ~n4625 ) ;
  assign n4627 = n3356 & ~n4626 ;
  assign n4628 = n4619 & n4627 ;
  assign n4629 = n351 | n1757 ;
  assign n4630 = n3248 & ~n4629 ;
  assign n4631 = n1004 ^ n333 ^ 1'b0 ;
  assign n4632 = n1398 & n4631 ;
  assign n4633 = n4531 & n4632 ;
  assign n4634 = ~n706 & n2468 ;
  assign n4635 = ~n2642 & n4634 ;
  assign n4636 = n4635 ^ n3948 ^ 1'b0 ;
  assign n4637 = n2636 | n4636 ;
  assign n4638 = n878 & ~n4317 ;
  assign n4639 = n559 & ~n640 ;
  assign n4640 = n1902 ^ n1380 ^ 1'b0 ;
  assign n4641 = n4639 | n4640 ;
  assign n4642 = n4641 ^ n4273 ^ 1'b0 ;
  assign n4645 = n3564 ^ n2974 ^ 1'b0 ;
  assign n4643 = x131 & n394 ;
  assign n4644 = ~x100 & n4643 ;
  assign n4646 = n4645 ^ n4644 ^ 1'b0 ;
  assign n4649 = x39 & n1388 ;
  assign n4650 = n4649 ^ n417 ^ 1'b0 ;
  assign n4651 = n2443 | n4650 ;
  assign n4647 = n2860 ^ n1418 ^ 1'b0 ;
  assign n4648 = n3254 | n4647 ;
  assign n4652 = n4651 ^ n4648 ^ x117 ;
  assign n4653 = n2365 ^ x233 ^ 1'b0 ;
  assign n4654 = n4653 ^ n668 ^ n270 ;
  assign n4655 = n929 & ~n2133 ;
  assign n4656 = ~n1908 & n4493 ;
  assign n4657 = n4655 & n4656 ;
  assign n4658 = n4654 | n4657 ;
  assign n4659 = n1176 & ~n4658 ;
  assign n4663 = n3532 ^ n1136 ^ 1'b0 ;
  assign n4664 = x27 & n4663 ;
  assign n4660 = n4118 ^ n1452 ^ 1'b0 ;
  assign n4661 = n982 & n4660 ;
  assign n4662 = ( n2884 & n3950 ) | ( n2884 & ~n4661 ) | ( n3950 & ~n4661 ) ;
  assign n4665 = n4664 ^ n4662 ^ 1'b0 ;
  assign n4666 = n2626 | n4665 ;
  assign n4667 = n3708 ^ n676 ^ 1'b0 ;
  assign n4668 = n1750 ^ n669 ^ 1'b0 ;
  assign n4669 = n1387 & ~n1724 ;
  assign n4670 = n4669 ^ x119 ^ 1'b0 ;
  assign n4671 = n4668 | n4670 ;
  assign n4672 = n4667 & ~n4671 ;
  assign n4673 = n750 & ~n884 ;
  assign n4674 = n1657 & ~n4673 ;
  assign n4675 = ~n3200 & n4674 ;
  assign n4676 = n4675 ^ n2292 ^ n1742 ;
  assign n4677 = n4280 ^ n2820 ^ n1435 ;
  assign n4678 = n4355 ^ n1131 ^ 1'b0 ;
  assign n4679 = n1527 ^ n1172 ^ n530 ;
  assign n4680 = ~n569 & n4679 ;
  assign n4681 = n4680 ^ n1527 ^ 1'b0 ;
  assign n4682 = n375 & ~n4139 ;
  assign n4683 = n4682 ^ n1357 ^ 1'b0 ;
  assign n4684 = n625 & n4683 ;
  assign n4685 = n4684 ^ n549 ^ 1'b0 ;
  assign n4686 = ~n4681 & n4685 ;
  assign n4694 = ( ~n2358 & n3190 ) | ( ~n2358 & n3409 ) | ( n3190 & n3409 ) ;
  assign n4689 = ~n1457 & n3172 ;
  assign n4690 = n1934 ^ n1886 ^ 1'b0 ;
  assign n4691 = ~n561 & n4690 ;
  assign n4692 = n4691 ^ n866 ^ 1'b0 ;
  assign n4693 = ( ~n3817 & n4689 ) | ( ~n3817 & n4692 ) | ( n4689 & n4692 ) ;
  assign n4695 = n4694 ^ n4693 ^ n945 ;
  assign n4687 = n1409 & n1768 ;
  assign n4688 = n4687 ^ n1040 ^ 1'b0 ;
  assign n4696 = n4695 ^ n4688 ^ 1'b0 ;
  assign n4697 = n2700 | n3859 ;
  assign n4698 = n4648 ^ n3059 ^ 1'b0 ;
  assign n4699 = x7 & n1770 ;
  assign n4700 = ~n884 & n4699 ;
  assign n4701 = n3990 ^ n2760 ^ 1'b0 ;
  assign n4702 = n2680 ^ n1148 ^ 1'b0 ;
  assign n4703 = n4018 & n4702 ;
  assign n4704 = n4564 ^ n1103 ^ 1'b0 ;
  assign n4705 = n4422 & ~n4704 ;
  assign n4706 = n4705 ^ n2458 ^ 1'b0 ;
  assign n4707 = ~n1919 & n4706 ;
  assign n4708 = n4041 ^ n2310 ^ 1'b0 ;
  assign n4709 = n3054 | n4708 ;
  assign n4710 = n4439 & ~n4709 ;
  assign n4711 = n4710 ^ n1258 ^ 1'b0 ;
  assign n4712 = n1604 & n2023 ;
  assign n4713 = n2844 ^ n1327 ^ n1174 ;
  assign n4714 = n4713 ^ n3775 ^ 1'b0 ;
  assign n4715 = n4528 ^ n4475 ^ n1880 ;
  assign n4716 = ~n921 & n1201 ;
  assign n4717 = n4716 ^ n3009 ^ 1'b0 ;
  assign n4718 = n2048 | n3060 ;
  assign n4719 = n2016 & ~n4718 ;
  assign n4720 = n4719 ^ x240 ^ 1'b0 ;
  assign n4721 = n4720 ^ n1611 ^ 1'b0 ;
  assign n4722 = ~n2506 & n4721 ;
  assign n4723 = n1694 & n2439 ;
  assign n4724 = n4469 & ~n4723 ;
  assign n4725 = n2890 ^ n2611 ^ 1'b0 ;
  assign n4726 = n4725 ^ n2454 ^ 1'b0 ;
  assign n4728 = ~n2326 & n3100 ;
  assign n4729 = ~n1561 & n4728 ;
  assign n4727 = ~n398 & n2201 ;
  assign n4730 = n4729 ^ n4727 ^ 1'b0 ;
  assign n4731 = ( n3112 & ~n4726 ) | ( n3112 & n4730 ) | ( ~n4726 & n4730 ) ;
  assign n4732 = n4065 ^ n1257 ^ 1'b0 ;
  assign n4733 = n1336 & ~n4732 ;
  assign n4734 = x2 & n3459 ;
  assign n4735 = ( n1751 & ~n4588 ) | ( n1751 & n4734 ) | ( ~n4588 & n4734 ) ;
  assign n4736 = ( n2030 & n3100 ) | ( n2030 & n4369 ) | ( n3100 & n4369 ) ;
  assign n4737 = n4736 ^ n4273 ^ 1'b0 ;
  assign n4738 = x62 & ~n4737 ;
  assign n4739 = n2939 ^ n1935 ^ n273 ;
  assign n4740 = n4739 ^ n1853 ^ 1'b0 ;
  assign n4741 = ~n1390 & n4740 ;
  assign n4742 = n1148 | n4741 ;
  assign n4743 = n4742 ^ n3056 ^ 1'b0 ;
  assign n4744 = ( x214 & n1641 ) | ( x214 & ~n4743 ) | ( n1641 & ~n4743 ) ;
  assign n4745 = n2456 ^ n852 ^ 1'b0 ;
  assign n4754 = n3580 | n3770 ;
  assign n4755 = ~n850 & n4754 ;
  assign n4746 = n1809 ^ n723 ^ 1'b0 ;
  assign n4751 = n1002 ^ n877 ^ n679 ;
  assign n4747 = n729 & ~n970 ;
  assign n4748 = n3213 | n4747 ;
  assign n4749 = n4748 ^ n3175 ^ 1'b0 ;
  assign n4750 = n3698 & ~n4749 ;
  assign n4752 = n4751 ^ n4750 ^ 1'b0 ;
  assign n4753 = n4746 & ~n4752 ;
  assign n4756 = n4755 ^ n4753 ^ 1'b0 ;
  assign n4757 = n3015 ^ n2346 ^ 1'b0 ;
  assign n4758 = n4397 | n4757 ;
  assign n4759 = ( n287 & ~n337 ) | ( n287 & n973 ) | ( ~n337 & n973 ) ;
  assign n4760 = n4759 ^ n1617 ^ n1481 ;
  assign n4761 = n2186 & ~n4760 ;
  assign n4762 = n4761 ^ x180 ^ 1'b0 ;
  assign n4763 = n1940 & ~n4762 ;
  assign n4764 = n1961 ^ x192 ^ 1'b0 ;
  assign n4765 = n2543 & n4764 ;
  assign n4766 = ~n4763 & n4765 ;
  assign n4767 = n1647 & ~n1995 ;
  assign n4768 = ( ~n617 & n3029 ) | ( ~n617 & n4767 ) | ( n3029 & n4767 ) ;
  assign n4769 = n2987 & ~n4768 ;
  assign n4770 = n487 | n3692 ;
  assign n4771 = ( n1935 & n4350 ) | ( n1935 & ~n4564 ) | ( n4350 & ~n4564 ) ;
  assign n4772 = n4770 | n4771 ;
  assign n4773 = n4769 | n4772 ;
  assign n4774 = x58 & n1174 ;
  assign n4775 = n4774 ^ n1521 ^ 1'b0 ;
  assign n4776 = n476 | n4775 ;
  assign n4777 = n1387 & ~n4776 ;
  assign n4780 = n1450 | n3308 ;
  assign n4778 = n1504 & n2733 ;
  assign n4779 = ~n1765 & n4778 ;
  assign n4781 = n4780 ^ n4779 ^ 1'b0 ;
  assign n4782 = n423 & ~n4781 ;
  assign n4783 = ~n4777 & n4782 ;
  assign n4784 = n4388 ^ n1803 ^ n1458 ;
  assign n4785 = ( x151 & ~x159 ) | ( x151 & n1211 ) | ( ~x159 & n1211 ) ;
  assign n4788 = n259 & ~n596 ;
  assign n4786 = n971 & ~n2767 ;
  assign n4787 = n4786 ^ n3833 ^ 1'b0 ;
  assign n4789 = n4788 ^ n4787 ^ 1'b0 ;
  assign n4790 = ( n1951 & ~n4785 ) | ( n1951 & n4789 ) | ( ~n4785 & n4789 ) ;
  assign n4791 = x182 | n3220 ;
  assign n4792 = ( n715 & n2574 ) | ( n715 & ~n4791 ) | ( n2574 & ~n4791 ) ;
  assign n4793 = n326 & n1540 ;
  assign n4794 = n4793 ^ n2978 ^ 1'b0 ;
  assign n4795 = n4679 & n4794 ;
  assign n4796 = n1956 & n4795 ;
  assign n4797 = n4796 ^ n2274 ^ 1'b0 ;
  assign n4798 = n1295 & ~n1602 ;
  assign n4799 = n1275 & n4798 ;
  assign n4800 = n4631 & ~n4799 ;
  assign n4801 = n4800 ^ n2688 ^ 1'b0 ;
  assign n4802 = n1716 & ~n4801 ;
  assign n4803 = n4802 ^ n4004 ^ 1'b0 ;
  assign n4804 = n391 & ~n2411 ;
  assign n4805 = n1323 ^ n1102 ^ n921 ;
  assign n4806 = n690 & n4805 ;
  assign n4807 = n774 & n4806 ;
  assign n4808 = n4189 | n4525 ;
  assign n4809 = n4808 ^ n2513 ^ 1'b0 ;
  assign n4810 = n1795 & ~n1823 ;
  assign n4811 = n4810 ^ n3263 ^ 1'b0 ;
  assign n4812 = n4811 ^ x124 ^ 1'b0 ;
  assign n4813 = x70 ^ x48 ^ 1'b0 ;
  assign n4814 = n1369 & n4813 ;
  assign n4815 = n3751 ^ n904 ^ 1'b0 ;
  assign n4816 = n4814 & n4815 ;
  assign n4821 = x190 & n580 ;
  assign n4822 = n4821 ^ n531 ^ 1'b0 ;
  assign n4823 = x124 | n4822 ;
  assign n4820 = x165 & n2210 ;
  assign n4824 = n4823 ^ n4820 ^ 1'b0 ;
  assign n4825 = n4824 ^ n3708 ^ 1'b0 ;
  assign n4817 = ~n1717 & n3277 ;
  assign n4818 = n4185 ^ n3436 ^ n1855 ;
  assign n4819 = ~n4817 & n4818 ;
  assign n4826 = n4825 ^ n4819 ^ 1'b0 ;
  assign n4827 = ~n994 & n4013 ;
  assign n4828 = n4078 ^ x42 ^ 1'b0 ;
  assign n4829 = n2019 | n4828 ;
  assign n4830 = n4829 ^ n2800 ^ 1'b0 ;
  assign n4831 = n298 & ~n1110 ;
  assign n4832 = n4830 & n4831 ;
  assign n4833 = n3521 ^ n468 ^ 1'b0 ;
  assign n4834 = n337 & ~n4803 ;
  assign n4835 = ~n1641 & n4834 ;
  assign n4836 = ( n1252 & n2204 ) | ( n1252 & n3328 ) | ( n2204 & n3328 ) ;
  assign n4837 = n1994 & ~n2075 ;
  assign n4838 = ~n3376 & n4837 ;
  assign n4839 = n2667 & n4838 ;
  assign n4840 = ~n3625 & n4839 ;
  assign n4841 = n2456 ^ x4 ^ 1'b0 ;
  assign n4842 = n3885 & n4841 ;
  assign n4843 = n1814 & n4842 ;
  assign n4844 = n4843 ^ n3255 ^ 1'b0 ;
  assign n4845 = ( ~x139 & n1194 ) | ( ~x139 & n2301 ) | ( n1194 & n2301 ) ;
  assign n4846 = n1741 & n4845 ;
  assign n4847 = n3641 & n4846 ;
  assign n4848 = ~n3839 & n4083 ;
  assign n4849 = n2376 ^ x150 ^ 1'b0 ;
  assign n4850 = n3375 & n4849 ;
  assign n4851 = n427 & n4850 ;
  assign n4852 = n2039 & ~n4851 ;
  assign n4853 = ~n2781 & n4129 ;
  assign n4854 = n2502 & n4853 ;
  assign n4855 = n1985 & n2308 ;
  assign n4856 = ~n325 & n2147 ;
  assign n4857 = n4856 ^ n2321 ^ 1'b0 ;
  assign n4858 = ~x108 & n3325 ;
  assign n4860 = x188 & ~n2522 ;
  assign n4861 = n619 & n4860 ;
  assign n4859 = n257 | n3975 ;
  assign n4862 = n4861 ^ n4859 ^ 1'b0 ;
  assign n4863 = ( ~n987 & n4858 ) | ( ~n987 & n4862 ) | ( n4858 & n4862 ) ;
  assign n4864 = n1266 & ~n3005 ;
  assign n4865 = n1307 & n4864 ;
  assign n4866 = n3197 & n4653 ;
  assign n4867 = n720 & n4866 ;
  assign n4868 = ~n4865 & n4867 ;
  assign n4869 = ( n4857 & n4863 ) | ( n4857 & n4868 ) | ( n4863 & n4868 ) ;
  assign n4870 = ( x135 & ~n829 ) | ( x135 & n4869 ) | ( ~n829 & n4869 ) ;
  assign n4871 = n4269 ^ n1719 ^ 1'b0 ;
  assign n4872 = n3242 & ~n4871 ;
  assign n4873 = n2277 | n2618 ;
  assign n4874 = n4873 ^ n415 ^ 1'b0 ;
  assign n4875 = ( ~x92 & n1825 ) | ( ~x92 & n4874 ) | ( n1825 & n4874 ) ;
  assign n4879 = n4067 ^ x50 ^ 1'b0 ;
  assign n4876 = n1106 ^ n1039 ^ 1'b0 ;
  assign n4877 = n807 & ~n1504 ;
  assign n4878 = ~n4876 & n4877 ;
  assign n4880 = n4879 ^ n4878 ^ 1'b0 ;
  assign n4881 = ~n4875 & n4880 ;
  assign n4882 = ~n1511 & n1540 ;
  assign n4883 = n4882 ^ n4019 ^ 1'b0 ;
  assign n4884 = ~x84 & x235 ;
  assign n4885 = ~n1765 & n3962 ;
  assign n4886 = n4884 & n4885 ;
  assign n4887 = n3922 ^ x77 ^ 1'b0 ;
  assign n4888 = n671 & n4887 ;
  assign n4889 = ( n947 & ~n2425 ) | ( n947 & n4888 ) | ( ~n2425 & n4888 ) ;
  assign n4890 = n4659 ^ n3190 ^ n1715 ;
  assign n4894 = ~n1882 & n4421 ;
  assign n4895 = n4894 ^ n1345 ^ 1'b0 ;
  assign n4896 = n2331 & n4895 ;
  assign n4891 = n3743 ^ n1368 ^ n925 ;
  assign n4892 = ~n3963 & n4764 ;
  assign n4893 = ~n4891 & n4892 ;
  assign n4897 = n4896 ^ n4893 ^ 1'b0 ;
  assign n4898 = n1727 & ~n4897 ;
  assign n4899 = n2171 ^ n1515 ^ n1442 ;
  assign n4900 = n2583 ^ n1374 ^ 1'b0 ;
  assign n4901 = ~n4899 & n4900 ;
  assign n4902 = n957 | n3568 ;
  assign n4903 = n4902 ^ n574 ^ 1'b0 ;
  assign n4904 = n428 & ~n4903 ;
  assign n4905 = ~n1804 & n4904 ;
  assign n4906 = ~n4901 & n4905 ;
  assign n4909 = n1567 & n3943 ;
  assign n4908 = x142 & ~n469 ;
  assign n4910 = n4909 ^ n4908 ^ 1'b0 ;
  assign n4911 = n4910 ^ n3909 ^ n857 ;
  assign n4907 = ~n1084 & n1439 ;
  assign n4912 = n4911 ^ n4907 ^ 1'b0 ;
  assign n4913 = ( x31 & n1549 ) | ( x31 & n3581 ) | ( n1549 & n3581 ) ;
  assign n4914 = n2601 | n4296 ;
  assign n4915 = n4913 | n4914 ;
  assign n4916 = n1372 & n4915 ;
  assign n4917 = n3078 ^ x95 ^ 1'b0 ;
  assign n4918 = n386 & ~n3163 ;
  assign n4919 = ~n2769 & n4918 ;
  assign n4920 = ( n845 & n853 ) | ( n845 & ~n1979 ) | ( n853 & ~n1979 ) ;
  assign n4921 = n2295 | n2680 ;
  assign n4922 = n2118 & ~n4921 ;
  assign n4923 = x254 & ~n2819 ;
  assign n4924 = ~n1838 & n4923 ;
  assign n4925 = n1176 | n4924 ;
  assign n4926 = n4922 & ~n4925 ;
  assign n4927 = ~n4888 & n4926 ;
  assign n4928 = n1265 & n4469 ;
  assign n4929 = n4928 ^ n3949 ^ n3585 ;
  assign n4940 = ~n378 & n3226 ;
  assign n4932 = x158 & n599 ;
  assign n4933 = n4932 ^ n1379 ^ x215 ;
  assign n4934 = n3786 & ~n4933 ;
  assign n4935 = ( x49 & ~n1232 ) | ( x49 & n3370 ) | ( ~n1232 & n3370 ) ;
  assign n4936 = ~n4651 & n4935 ;
  assign n4937 = ~n3439 & n4936 ;
  assign n4938 = ( ~n4078 & n4934 ) | ( ~n4078 & n4937 ) | ( n4934 & n4937 ) ;
  assign n4930 = ( n398 & n827 ) | ( n398 & n1271 ) | ( n827 & n1271 ) ;
  assign n4931 = n4930 ^ x146 ^ 1'b0 ;
  assign n4939 = n4938 ^ n4931 ^ n1741 ;
  assign n4941 = n4940 ^ n4939 ^ n4572 ;
  assign n4942 = n1046 | n4475 ;
  assign n4943 = n476 & ~n4942 ;
  assign n4944 = n2052 ^ n1899 ^ 1'b0 ;
  assign n4945 = n1585 & n4944 ;
  assign n4946 = n4945 ^ n2648 ^ 1'b0 ;
  assign n4947 = ( n1232 & ~n3194 ) | ( n1232 & n4946 ) | ( ~n3194 & n4946 ) ;
  assign n4951 = x55 & n1970 ;
  assign n4952 = n4951 ^ n720 ^ 1'b0 ;
  assign n4948 = ~n1700 & n3150 ;
  assign n4949 = n4948 ^ n4614 ^ 1'b0 ;
  assign n4950 = ~n2786 & n4949 ;
  assign n4953 = n4952 ^ n4950 ^ x45 ;
  assign n4954 = n945 | n4523 ;
  assign n4955 = n4353 | n4672 ;
  assign n4956 = n1082 & n2603 ;
  assign n4957 = n2674 & n4956 ;
  assign n4958 = n4957 ^ n4318 ^ n800 ;
  assign n4959 = n4958 ^ n1320 ^ 1'b0 ;
  assign n4960 = ( n2280 & ~n4395 ) | ( n2280 & n4959 ) | ( ~n4395 & n4959 ) ;
  assign n4961 = n4960 ^ n1296 ^ n731 ;
  assign n4966 = n3817 ^ x25 ^ 1'b0 ;
  assign n4967 = n2001 | n4966 ;
  assign n4968 = n1576 & ~n4967 ;
  assign n4975 = ~x48 & n1284 ;
  assign n4969 = ~n482 & n861 ;
  assign n4970 = n4969 ^ n813 ^ 1'b0 ;
  assign n4971 = n4970 ^ n517 ^ x104 ;
  assign n4972 = n1225 & ~n4971 ;
  assign n4973 = n4972 ^ x123 ^ 1'b0 ;
  assign n4974 = n2335 | n4973 ;
  assign n4976 = n4975 ^ n4974 ^ 1'b0 ;
  assign n4977 = n4968 | n4976 ;
  assign n4962 = n2401 ^ n2024 ^ 1'b0 ;
  assign n4963 = n501 | n4962 ;
  assign n4964 = ~n887 & n4053 ;
  assign n4965 = n4963 & n4964 ;
  assign n4978 = n4977 ^ n4965 ^ n1533 ;
  assign n4979 = ~n1096 & n2630 ;
  assign n4980 = n1900 | n4979 ;
  assign n4981 = ~n1141 & n4980 ;
  assign n4982 = n2102 & n4614 ;
  assign n4983 = ( x121 & ~n287 ) | ( x121 & n4982 ) | ( ~n287 & n4982 ) ;
  assign n4984 = n4983 ^ n4824 ^ 1'b0 ;
  assign n4985 = n4111 ^ n1120 ^ n706 ;
  assign n4986 = ( n1376 & n4468 ) | ( n1376 & ~n4985 ) | ( n4468 & ~n4985 ) ;
  assign n4987 = n507 & ~n2315 ;
  assign n4988 = ( n787 & n1728 ) | ( n787 & n4316 ) | ( n1728 & n4316 ) ;
  assign n4989 = n1649 | n4988 ;
  assign n4990 = n2899 & n4274 ;
  assign n4991 = ~n2304 & n4990 ;
  assign n4992 = n4991 ^ n1258 ^ 1'b0 ;
  assign n4993 = n2802 ^ n2025 ^ n1859 ;
  assign n4996 = ( n807 & n1496 ) | ( n807 & n3679 ) | ( n1496 & n3679 ) ;
  assign n4997 = n333 | n4996 ;
  assign n4998 = n4997 ^ n1252 ^ 1'b0 ;
  assign n4999 = ~n1671 & n4998 ;
  assign n4994 = ~n2937 & n3140 ;
  assign n4995 = n4994 ^ n3994 ^ n1971 ;
  assign n5000 = n4999 ^ n4995 ^ 1'b0 ;
  assign n5001 = n4993 | n5000 ;
  assign n5005 = n649 | n825 ;
  assign n5006 = n5005 ^ x115 ^ 1'b0 ;
  assign n5002 = n1044 ^ n813 ^ 1'b0 ;
  assign n5003 = x225 | n5002 ;
  assign n5004 = n257 & ~n5003 ;
  assign n5007 = n5006 ^ n5004 ^ n1416 ;
  assign n5008 = n365 & ~n2165 ;
  assign n5009 = n3567 & n5008 ;
  assign n5010 = x39 & ~n804 ;
  assign n5011 = n5010 ^ n1272 ^ 1'b0 ;
  assign n5012 = n3751 ^ n2373 ^ n898 ;
  assign n5013 = n3893 & ~n5012 ;
  assign n5014 = n5013 ^ n2121 ^ 1'b0 ;
  assign n5015 = n5011 | n5014 ;
  assign n5016 = n3105 ^ n478 ^ 1'b0 ;
  assign n5017 = n1933 | n5016 ;
  assign n5018 = n5017 ^ x142 ^ 1'b0 ;
  assign n5019 = n3207 & n4389 ;
  assign n5020 = n335 & n5019 ;
  assign n5021 = ( n1041 & ~n2321 ) | ( n1041 & n2416 ) | ( ~n2321 & n2416 ) ;
  assign n5022 = ~n1132 & n5021 ;
  assign n5023 = n476 | n2657 ;
  assign n5024 = n5023 ^ n2954 ^ 1'b0 ;
  assign n5025 = n5024 ^ n2929 ^ n1594 ;
  assign n5026 = n785 & n968 ;
  assign n5027 = ~n1715 & n5026 ;
  assign n5028 = x66 & ~n766 ;
  assign n5029 = n1734 ^ n1596 ^ 1'b0 ;
  assign n5030 = ~n5028 & n5029 ;
  assign n5031 = ~n5027 & n5030 ;
  assign n5032 = ( n332 & n2411 ) | ( n332 & n5031 ) | ( n2411 & n5031 ) ;
  assign n5036 = ~n469 & n785 ;
  assign n5037 = n5036 ^ n2822 ^ 1'b0 ;
  assign n5038 = ( ~x152 & n3526 ) | ( ~x152 & n5037 ) | ( n3526 & n5037 ) ;
  assign n5033 = n4909 ^ n262 ^ 1'b0 ;
  assign n5034 = n5033 ^ n3910 ^ n1182 ;
  assign n5035 = n3455 & n5034 ;
  assign n5039 = n5038 ^ n5035 ^ 1'b0 ;
  assign n5042 = n701 & n1524 ;
  assign n5043 = n5042 ^ n1789 ^ 1'b0 ;
  assign n5040 = n1836 | n1989 ;
  assign n5041 = n5040 ^ n2980 ^ 1'b0 ;
  assign n5044 = n5043 ^ n5041 ^ n1746 ;
  assign n5045 = n533 & n3476 ;
  assign n5046 = n4528 | n5045 ;
  assign n5047 = n1347 & ~n5046 ;
  assign n5048 = ~n2280 & n4422 ;
  assign n5049 = n3481 & n5048 ;
  assign n5051 = n3735 ^ n2816 ^ 1'b0 ;
  assign n5052 = n1861 & ~n5051 ;
  assign n5053 = n5052 ^ n2484 ^ 1'b0 ;
  assign n5050 = ( ~n635 & n1760 ) | ( ~n635 & n2097 ) | ( n1760 & n2097 ) ;
  assign n5054 = n5053 ^ n5050 ^ 1'b0 ;
  assign n5055 = n3708 | n5054 ;
  assign n5056 = n1946 & n2893 ;
  assign n5057 = n3181 ^ n1482 ^ 1'b0 ;
  assign n5058 = ( n1013 & n2196 ) | ( n1013 & n5057 ) | ( n2196 & n5057 ) ;
  assign n5059 = ~n2202 & n5058 ;
  assign n5060 = ( ~n3978 & n4391 ) | ( ~n3978 & n5059 ) | ( n4391 & n5059 ) ;
  assign n5061 = n5060 ^ n2067 ^ 1'b0 ;
  assign n5062 = ~n5056 & n5061 ;
  assign n5071 = n1196 ^ n997 ^ x57 ;
  assign n5072 = n5071 ^ n3182 ^ n2348 ;
  assign n5063 = n3156 ^ n2717 ^ 1'b0 ;
  assign n5064 = n2764 | n5063 ;
  assign n5065 = n3178 | n5064 ;
  assign n5066 = n1424 ^ x33 ^ 1'b0 ;
  assign n5067 = n5066 ^ n2251 ^ 1'b0 ;
  assign n5068 = n5067 ^ n3952 ^ 1'b0 ;
  assign n5069 = n1409 & n5068 ;
  assign n5070 = ( n2379 & n5065 ) | ( n2379 & ~n5069 ) | ( n5065 & ~n5069 ) ;
  assign n5073 = n5072 ^ n5070 ^ n3796 ;
  assign n5074 = n1486 & n4938 ;
  assign n5075 = ~n3953 & n5074 ;
  assign n5076 = n5075 ^ n1791 ^ 1'b0 ;
  assign n5077 = n3593 & n3970 ;
  assign n5078 = ( n402 & ~n706 ) | ( n402 & n1510 ) | ( ~n706 & n1510 ) ;
  assign n5079 = n5078 ^ n3732 ^ 1'b0 ;
  assign n5080 = n1251 | n4341 ;
  assign n5081 = n3112 & ~n5080 ;
  assign n5085 = x234 & ~n3054 ;
  assign n5086 = n5085 ^ n1133 ^ 1'b0 ;
  assign n5087 = ~n2370 & n5086 ;
  assign n5082 = n1875 ^ n1843 ^ 1'b0 ;
  assign n5083 = ~n1700 & n5082 ;
  assign n5084 = ~n881 & n5083 ;
  assign n5088 = n5087 ^ n5084 ^ 1'b0 ;
  assign n5089 = n3506 | n5088 ;
  assign n5090 = n5089 ^ n4922 ^ 1'b0 ;
  assign n5091 = ( n362 & n1368 ) | ( n362 & n1938 ) | ( n1368 & n1938 ) ;
  assign n5092 = n5091 ^ n1142 ^ 1'b0 ;
  assign n5093 = n3517 & ~n5092 ;
  assign n5094 = ~x208 & n789 ;
  assign n5095 = n1515 & n5094 ;
  assign n5096 = n2543 & n4130 ;
  assign n5097 = ~n3781 & n5096 ;
  assign n5099 = n1684 & n1759 ;
  assign n5098 = ( n1113 & n1820 ) | ( n1113 & n3452 ) | ( n1820 & n3452 ) ;
  assign n5100 = n5099 ^ n5098 ^ 1'b0 ;
  assign n5101 = ~n5097 & n5100 ;
  assign n5102 = n635 | n829 ;
  assign n5103 = n462 & ~n764 ;
  assign n5104 = n5103 ^ n2990 ^ 1'b0 ;
  assign n5105 = n3843 ^ n1388 ^ 1'b0 ;
  assign n5106 = ( ~n1361 & n2373 ) | ( ~n1361 & n5105 ) | ( n2373 & n5105 ) ;
  assign n5107 = n5106 ^ n3940 ^ x146 ;
  assign n5108 = ( n2369 & ~n3630 ) | ( n2369 & n5107 ) | ( ~n3630 & n5107 ) ;
  assign n5109 = ( n358 & n1260 ) | ( n358 & ~n1429 ) | ( n1260 & ~n1429 ) ;
  assign n5110 = n922 | n5109 ;
  assign n5111 = ( n3425 & n4673 ) | ( n3425 & n5110 ) | ( n4673 & n5110 ) ;
  assign n5112 = ~n3025 & n3575 ;
  assign n5113 = n913 | n3813 ;
  assign n5114 = n1774 & ~n5113 ;
  assign n5115 = n5112 & ~n5114 ;
  assign n5116 = n363 | n5115 ;
  assign n5117 = n5111 & ~n5116 ;
  assign n5118 = n945 & ~n4611 ;
  assign n5119 = ~n632 & n5118 ;
  assign n5120 = n1199 & ~n3080 ;
  assign n5121 = n921 & n5120 ;
  assign n5122 = n317 | n1595 ;
  assign n5123 = n385 | n5122 ;
  assign n5124 = n1880 | n5123 ;
  assign n5125 = n2515 & ~n3817 ;
  assign n5126 = n5125 ^ n887 ^ 1'b0 ;
  assign n5127 = x155 & n2667 ;
  assign n5128 = n5127 ^ n3024 ^ 1'b0 ;
  assign n5129 = ~n4971 & n5128 ;
  assign n5130 = n1389 ^ n945 ^ 1'b0 ;
  assign n5131 = x28 & n5130 ;
  assign n5132 = n1666 ^ n1511 ^ 1'b0 ;
  assign n5133 = n3632 & n5132 ;
  assign n5134 = n3007 & n5133 ;
  assign n5135 = n4623 & n5134 ;
  assign n5136 = n1956 & ~n3294 ;
  assign n5137 = n5136 ^ n2381 ^ 1'b0 ;
  assign n5146 = n3471 ^ n2844 ^ 1'b0 ;
  assign n5147 = ~n1955 & n4595 ;
  assign n5148 = ~n5146 & n5147 ;
  assign n5138 = n356 ^ x18 ^ 1'b0 ;
  assign n5139 = n5138 ^ n4085 ^ n1760 ;
  assign n5140 = n2831 & n5139 ;
  assign n5141 = n5140 ^ n1624 ^ 1'b0 ;
  assign n5142 = n2142 ^ n2131 ^ 1'b0 ;
  assign n5143 = n3333 & ~n5142 ;
  assign n5144 = ( n2676 & ~n5141 ) | ( n2676 & n5143 ) | ( ~n5141 & n5143 ) ;
  assign n5145 = x242 & n5144 ;
  assign n5149 = n5148 ^ n5145 ^ 1'b0 ;
  assign n5156 = n517 | n606 ;
  assign n5157 = n2394 | n5156 ;
  assign n5150 = n4958 & ~n4982 ;
  assign n5151 = n5150 ^ n2816 ^ 1'b0 ;
  assign n5152 = ~n1786 & n2709 ;
  assign n5153 = n5152 ^ n1288 ^ 1'b0 ;
  assign n5154 = n1666 & n5153 ;
  assign n5155 = n5151 & n5154 ;
  assign n5158 = n5157 ^ n5155 ^ n2358 ;
  assign n5159 = n1564 | n4020 ;
  assign n5160 = n275 & n874 ;
  assign n5161 = n5160 ^ n2032 ^ 1'b0 ;
  assign n5162 = ~n5159 & n5161 ;
  assign n5163 = x159 & ~n2885 ;
  assign n5164 = n4306 & n5163 ;
  assign n5165 = ~n5162 & n5164 ;
  assign n5170 = n1787 ^ n1069 ^ n898 ;
  assign n5169 = ( ~n677 & n4416 ) | ( ~n677 & n4435 ) | ( n4416 & n4435 ) ;
  assign n5171 = n5170 ^ n5169 ^ n2058 ;
  assign n5166 = ~n1611 & n2113 ;
  assign n5167 = ~n2510 & n5166 ;
  assign n5168 = n1399 & ~n5167 ;
  assign n5172 = n5171 ^ n5168 ^ 1'b0 ;
  assign n5173 = n5172 ^ n4192 ^ n1393 ;
  assign n5174 = n1828 & n2257 ;
  assign n5175 = n3219 & ~n5174 ;
  assign n5185 = n1797 ^ n866 ^ 1'b0 ;
  assign n5184 = n580 & n2157 ;
  assign n5186 = n5185 ^ n5184 ^ 1'b0 ;
  assign n5176 = n1308 & ~n2449 ;
  assign n5177 = ~n1884 & n5176 ;
  assign n5180 = ~n256 & n4024 ;
  assign n5181 = n5180 ^ n1123 ^ 1'b0 ;
  assign n5178 = n2733 ^ n1480 ^ 1'b0 ;
  assign n5179 = n5178 ^ n1284 ^ n828 ;
  assign n5182 = n5181 ^ n5179 ^ 1'b0 ;
  assign n5183 = ~n5177 & n5182 ;
  assign n5187 = n5186 ^ n5183 ^ 1'b0 ;
  assign n5188 = n4681 ^ n410 ^ 1'b0 ;
  assign n5189 = n4342 ^ n2687 ^ 1'b0 ;
  assign n5190 = ~n5188 & n5189 ;
  assign n5191 = n5190 ^ n2682 ^ 1'b0 ;
  assign n5195 = n706 & ~n4004 ;
  assign n5192 = n1574 | n3436 ;
  assign n5193 = n3019 | n5192 ;
  assign n5194 = x131 & n5193 ;
  assign n5196 = n5195 ^ n5194 ^ 1'b0 ;
  assign n5197 = n5196 ^ n1902 ^ 1'b0 ;
  assign n5198 = n1427 ^ n1299 ^ 1'b0 ;
  assign n5199 = n1644 | n2695 ;
  assign n5200 = ~n2754 & n5199 ;
  assign n5201 = ~n1162 & n5200 ;
  assign n5202 = n2830 ^ n1510 ^ 1'b0 ;
  assign n5203 = ~n3889 & n5202 ;
  assign n5204 = n2727 & ~n5203 ;
  assign n5205 = n2767 | n3349 ;
  assign n5206 = n5205 ^ n3273 ^ 1'b0 ;
  assign n5207 = n1543 & n5206 ;
  assign n5208 = n5207 ^ n3731 ^ n2782 ;
  assign n5209 = ( n4193 & n5166 ) | ( n4193 & ~n5208 ) | ( n5166 & ~n5208 ) ;
  assign n5210 = n861 & ~n1406 ;
  assign n5211 = n5210 ^ n3873 ^ 1'b0 ;
  assign n5212 = ~n3813 & n4690 ;
  assign n5213 = n5211 & n5212 ;
  assign n5214 = n3328 & n5213 ;
  assign n5215 = ~n3640 & n5214 ;
  assign n5216 = n2572 ^ n1959 ^ 1'b0 ;
  assign n5217 = n2897 | n5216 ;
  assign n5218 = n5217 ^ n4920 ^ 1'b0 ;
  assign n5219 = n2352 | n5218 ;
  assign n5220 = n1754 ^ n1634 ^ 1'b0 ;
  assign n5221 = n974 & n5220 ;
  assign n5222 = n5221 ^ n627 ^ 1'b0 ;
  assign n5223 = n4148 & n5222 ;
  assign n5224 = n968 & n3727 ;
  assign n5225 = ~n1120 & n5224 ;
  assign n5226 = x182 | n5225 ;
  assign n5227 = ~n800 & n5226 ;
  assign n5228 = ~n2369 & n5227 ;
  assign n5229 = n4029 ^ n263 ^ 1'b0 ;
  assign n5230 = n2191 & n5229 ;
  assign n5231 = n1399 & ~n5230 ;
  assign n5232 = ~n5131 & n5231 ;
  assign n5233 = n1776 & ~n2024 ;
  assign n5234 = n1976 & n3308 ;
  assign n5235 = n4105 ^ n3310 ^ 1'b0 ;
  assign n5236 = ( n5233 & ~n5234 ) | ( n5233 & n5235 ) | ( ~n5234 & n5235 ) ;
  assign n5237 = n1916 ^ n304 ^ 1'b0 ;
  assign n5238 = n3744 ^ n2618 ^ 1'b0 ;
  assign n5239 = ( n1713 & n5237 ) | ( n1713 & n5238 ) | ( n5237 & n5238 ) ;
  assign n5240 = n2934 ^ n1187 ^ 1'b0 ;
  assign n5241 = n2240 & ~n5240 ;
  assign n5242 = n4982 & n5241 ;
  assign n5243 = n2856 | n4723 ;
  assign n5244 = n5243 ^ n487 ^ 1'b0 ;
  assign n5255 = n1120 ^ n704 ^ 1'b0 ;
  assign n5256 = n2800 & ~n5255 ;
  assign n5257 = n4237 & n5256 ;
  assign n5245 = n740 | n1222 ;
  assign n5246 = n1976 ^ n1300 ^ 1'b0 ;
  assign n5247 = ~n1129 & n1269 ;
  assign n5248 = ~x152 & n5247 ;
  assign n5249 = ( n2278 & n2660 ) | ( n2278 & n5248 ) | ( n2660 & n5248 ) ;
  assign n5250 = n428 & ~n1142 ;
  assign n5251 = n5250 ^ n1503 ^ 1'b0 ;
  assign n5252 = n729 & n5251 ;
  assign n5253 = n5249 & n5252 ;
  assign n5254 = ( n5245 & n5246 ) | ( n5245 & n5253 ) | ( n5246 & n5253 ) ;
  assign n5258 = n5257 ^ n5254 ^ n2511 ;
  assign n5259 = n3872 ^ n1877 ^ 1'b0 ;
  assign n5260 = ~n2042 & n2720 ;
  assign n5261 = ~n5259 & n5260 ;
  assign n5262 = n5261 ^ n1202 ^ 1'b0 ;
  assign n5263 = n2123 ^ n1543 ^ n856 ;
  assign n5264 = n286 & n1514 ;
  assign n5265 = ( n405 & ~n768 ) | ( n405 & n5264 ) | ( ~n768 & n5264 ) ;
  assign n5266 = ~n5263 & n5265 ;
  assign n5267 = n1390 ^ x141 ^ 1'b0 ;
  assign n5268 = n5267 ^ n1976 ^ 1'b0 ;
  assign n5269 = ~n4321 & n5268 ;
  assign n5270 = ( n2030 & n5058 ) | ( n2030 & ~n5269 ) | ( n5058 & ~n5269 ) ;
  assign n5271 = n3948 & ~n5270 ;
  assign n5272 = ~n5266 & n5271 ;
  assign n5273 = n318 & ~n1557 ;
  assign n5274 = n5273 ^ n3373 ^ 1'b0 ;
  assign n5275 = n1435 & n2110 ;
  assign n5276 = n2900 | n3277 ;
  assign n5277 = ( n2491 & ~n5275 ) | ( n2491 & n5276 ) | ( ~n5275 & n5276 ) ;
  assign n5278 = n5277 ^ n935 ^ 1'b0 ;
  assign n5279 = n5274 & n5278 ;
  assign n5280 = n5155 ^ n300 ^ 1'b0 ;
  assign n5281 = x71 & ~n5280 ;
  assign n5289 = ( n493 & n2752 ) | ( n493 & ~n4858 ) | ( n2752 & ~n4858 ) ;
  assign n5282 = n3608 & ~n3950 ;
  assign n5283 = n2449 & n5282 ;
  assign n5284 = x34 & n1452 ;
  assign n5285 = ~n1324 & n5284 ;
  assign n5286 = n4561 | n5285 ;
  assign n5287 = n5286 ^ n3704 ^ 1'b0 ;
  assign n5288 = ~n5283 & n5287 ;
  assign n5290 = n5289 ^ n5288 ^ n2120 ;
  assign n5291 = n4777 ^ n1093 ^ 1'b0 ;
  assign n5292 = ~n2713 & n4574 ;
  assign n5293 = n2676 ^ n1406 ^ 1'b0 ;
  assign n5294 = n1084 | n5293 ;
  assign n5295 = n2677 | n4767 ;
  assign n5296 = n5294 & ~n5295 ;
  assign n5297 = n1980 ^ n1249 ^ 1'b0 ;
  assign n5298 = n5296 | n5297 ;
  assign n5299 = n2041 ^ n390 ^ 1'b0 ;
  assign n5300 = n5298 | n5299 ;
  assign n5301 = n514 & n686 ;
  assign n5302 = n5301 ^ n2692 ^ n1435 ;
  assign n5303 = x55 & ~n2650 ;
  assign n5304 = n5303 ^ n1032 ^ 1'b0 ;
  assign n5305 = n5302 | n5304 ;
  assign n5306 = n1496 ^ n780 ^ 1'b0 ;
  assign n5307 = n4746 ^ n1723 ^ n1586 ;
  assign n5308 = ( n3394 & n5153 ) | ( n3394 & ~n5307 ) | ( n5153 & ~n5307 ) ;
  assign n5310 = n4151 ^ n1543 ^ n737 ;
  assign n5309 = n288 | n4342 ;
  assign n5311 = n5310 ^ n5309 ^ 1'b0 ;
  assign n5312 = n5311 ^ n4451 ^ 1'b0 ;
  assign n5313 = n1262 & ~n5312 ;
  assign n5314 = n1711 | n1802 ;
  assign n5315 = n5314 ^ n3286 ^ 1'b0 ;
  assign n5316 = n3998 & ~n5315 ;
  assign n5317 = n2191 ^ n1265 ^ x170 ;
  assign n5318 = n2120 & n5317 ;
  assign n5319 = n282 | n5318 ;
  assign n5320 = n5319 ^ n3607 ^ 1'b0 ;
  assign n5321 = n5320 ^ n614 ^ 1'b0 ;
  assign n5322 = ~n4257 & n5321 ;
  assign n5323 = ( ~n577 & n1226 ) | ( ~n577 & n3810 ) | ( n1226 & n3810 ) ;
  assign n5324 = n5323 ^ n3683 ^ n2360 ;
  assign n5325 = n2874 | n5324 ;
  assign n5326 = n2454 ^ n2094 ^ 1'b0 ;
  assign n5327 = n1647 & ~n2509 ;
  assign n5328 = ( n625 & n2433 ) | ( n625 & n5327 ) | ( n2433 & n5327 ) ;
  assign n5329 = n5328 ^ n4086 ^ 1'b0 ;
  assign n5330 = n5326 & ~n5329 ;
  assign n5331 = n1164 ^ x116 ^ x84 ;
  assign n5332 = n2193 & n5331 ;
  assign n5333 = n5332 ^ n5115 ^ 1'b0 ;
  assign n5334 = x139 ^ x85 ^ 1'b0 ;
  assign n5335 = ( ~x246 & n1257 ) | ( ~x246 & n5334 ) | ( n1257 & n5334 ) ;
  assign n5336 = n1999 & n4535 ;
  assign n5337 = n5336 ^ n5057 ^ 1'b0 ;
  assign n5338 = n3145 ^ n725 ^ 1'b0 ;
  assign n5339 = n2916 & n5338 ;
  assign n5340 = ~n4034 & n5339 ;
  assign n5341 = n5340 ^ n2054 ^ 1'b0 ;
  assign n5342 = ( n2939 & n5337 ) | ( n2939 & ~n5341 ) | ( n5337 & ~n5341 ) ;
  assign n5343 = n2826 ^ n1067 ^ 1'b0 ;
  assign n5344 = n3408 | n5343 ;
  assign n5345 = ~n663 & n5344 ;
  assign n5346 = x83 & n3400 ;
  assign n5347 = n5346 ^ n2884 ^ 1'b0 ;
  assign n5348 = n2070 | n3190 ;
  assign n5349 = n2618 & ~n5348 ;
  assign n5351 = n1347 ^ n1106 ^ n576 ;
  assign n5352 = n4353 & n5351 ;
  assign n5353 = ~x194 & n5352 ;
  assign n5354 = n2638 & ~n5353 ;
  assign n5355 = n275 & n5354 ;
  assign n5356 = n4618 & ~n5355 ;
  assign n5350 = n2567 & ~n2651 ;
  assign n5357 = n5356 ^ n5350 ^ 1'b0 ;
  assign n5358 = ( x30 & n453 ) | ( x30 & ~n4013 ) | ( n453 & ~n4013 ) ;
  assign n5359 = ( ~x185 & n593 ) | ( ~x185 & n3420 ) | ( n593 & n3420 ) ;
  assign n5360 = n4020 & n5359 ;
  assign n5361 = ( n4156 & ~n5358 ) | ( n4156 & n5360 ) | ( ~n5358 & n5360 ) ;
  assign n5363 = n1013 ^ n936 ^ n565 ;
  assign n5364 = x231 ^ x97 ^ x50 ;
  assign n5365 = ~n5363 & n5364 ;
  assign n5366 = n660 & ~n5365 ;
  assign n5362 = n3926 ^ n557 ^ 1'b0 ;
  assign n5367 = n5366 ^ n5362 ^ n4713 ;
  assign n5368 = ~x32 & n987 ;
  assign n5369 = n5368 ^ n1716 ^ 1'b0 ;
  assign n5370 = ~n2459 & n5369 ;
  assign n5371 = ( ~n344 & n2023 ) | ( ~n344 & n5370 ) | ( n2023 & n5370 ) ;
  assign n5372 = n1038 & n4039 ;
  assign n5373 = x44 & n2938 ;
  assign n5374 = n5372 & ~n5373 ;
  assign n5375 = n3516 ^ n1640 ^ 1'b0 ;
  assign n5376 = n2419 | n5375 ;
  assign n5377 = n3784 ^ n2070 ^ 1'b0 ;
  assign n5378 = n3264 & ~n5377 ;
  assign n5379 = n5378 ^ n3074 ^ 1'b0 ;
  assign n5380 = ~n810 & n4913 ;
  assign n5381 = n5379 & n5380 ;
  assign n5382 = x183 & ~n5381 ;
  assign n5383 = n5382 ^ n4046 ^ 1'b0 ;
  assign n5384 = n5376 | n5383 ;
  assign n5385 = n2159 & ~n5329 ;
  assign n5386 = n1985 ^ n652 ^ 1'b0 ;
  assign n5387 = n4552 ^ n2697 ^ n2471 ;
  assign n5388 = n4760 ^ n318 ^ x88 ;
  assign n5390 = n3494 | n4475 ;
  assign n5391 = n864 | n5390 ;
  assign n5392 = ~n2819 & n5391 ;
  assign n5393 = n5392 ^ n3845 ^ 1'b0 ;
  assign n5389 = n1950 | n2889 ;
  assign n5394 = n5393 ^ n5389 ^ 1'b0 ;
  assign n5395 = ( ~x245 & n4244 ) | ( ~x245 & n5394 ) | ( n4244 & n5394 ) ;
  assign n5396 = n4473 ^ n2642 ^ n1636 ;
  assign n5397 = ~n1203 & n1397 ;
  assign n5398 = n5397 ^ n3843 ^ n1813 ;
  assign n5401 = n3854 ^ n1354 ^ 1'b0 ;
  assign n5402 = n881 | n5401 ;
  assign n5399 = x224 & n3172 ;
  assign n5400 = n5399 ^ n1672 ^ 1'b0 ;
  assign n5403 = n5402 ^ n5400 ^ 1'b0 ;
  assign n5404 = ~n3615 & n5403 ;
  assign n5405 = ~n2315 & n3605 ;
  assign n5406 = ( n273 & n696 ) | ( n273 & ~n5405 ) | ( n696 & ~n5405 ) ;
  assign n5407 = ~n1468 & n2687 ;
  assign n5408 = n5407 ^ x250 ^ 1'b0 ;
  assign n5409 = ~n1555 & n2307 ;
  assign n5410 = n449 & n5409 ;
  assign n5411 = ( ~n2798 & n4457 ) | ( ~n2798 & n5410 ) | ( n4457 & n5410 ) ;
  assign n5412 = ~n286 & n1122 ;
  assign n5413 = n1016 & ~n5412 ;
  assign n5414 = n5413 ^ n3100 ^ 1'b0 ;
  assign n5415 = n5411 | n5414 ;
  assign n5416 = n3944 ^ n2463 ^ 1'b0 ;
  assign n5417 = ( n1343 & n1914 ) | ( n1343 & ~n3315 ) | ( n1914 & ~n3315 ) ;
  assign n5418 = n5417 ^ n3255 ^ 1'b0 ;
  assign n5419 = n4588 | n5418 ;
  assign n5420 = ~x113 & n4055 ;
  assign n5421 = n5308 ^ n738 ^ 1'b0 ;
  assign n5422 = ~n1144 & n5421 ;
  assign n5427 = n1249 ^ x182 ^ 1'b0 ;
  assign n5423 = n434 & ~n3758 ;
  assign n5424 = n2057 & n5423 ;
  assign n5425 = n1187 | n5424 ;
  assign n5426 = n5425 ^ n3492 ^ 1'b0 ;
  assign n5428 = n5427 ^ n5426 ^ n4471 ;
  assign n5429 = n4071 ^ n3744 ^ 1'b0 ;
  assign n5430 = n5428 | n5429 ;
  assign n5432 = n3455 & n5153 ;
  assign n5431 = n1343 & n2752 ;
  assign n5433 = n5432 ^ n5431 ^ 1'b0 ;
  assign n5434 = n2394 ^ n642 ^ 1'b0 ;
  assign n5435 = n5112 | n5434 ;
  assign n5436 = n5433 & ~n5435 ;
  assign n5437 = ( n1132 & n2936 ) | ( n1132 & n4517 ) | ( n2936 & n4517 ) ;
  assign n5444 = x76 & n2713 ;
  assign n5438 = n2061 ^ n1802 ^ n1201 ;
  assign n5439 = n4746 ^ n552 ^ 1'b0 ;
  assign n5440 = ( n2715 & n5438 ) | ( n2715 & ~n5439 ) | ( n5438 & ~n5439 ) ;
  assign n5441 = ~n1149 & n5440 ;
  assign n5442 = n3261 & n5441 ;
  assign n5443 = ~n4242 & n5442 ;
  assign n5445 = n5444 ^ n5443 ^ 1'b0 ;
  assign n5446 = n2425 ^ n2041 ^ 1'b0 ;
  assign n5447 = ~n3607 & n5446 ;
  assign n5448 = ~n895 & n3188 ;
  assign n5449 = ( n3339 & n3721 ) | ( n3339 & n5448 ) | ( n3721 & n5448 ) ;
  assign n5450 = n563 & n1249 ;
  assign n5451 = n5450 ^ n4421 ^ 1'b0 ;
  assign n5452 = x89 & ~n5451 ;
  assign n5453 = n5452 ^ x220 ^ 1'b0 ;
  assign n5454 = ~n1748 & n2443 ;
  assign n5455 = n4107 ^ n2740 ^ 1'b0 ;
  assign n5456 = n2145 & ~n5455 ;
  assign n5457 = n5456 ^ n2836 ^ 1'b0 ;
  assign n5458 = n1174 & ~n5457 ;
  assign n5459 = n3877 | n5458 ;
  assign n5460 = ( n2877 & ~n4026 ) | ( n2877 & n4148 ) | ( ~n4026 & n4148 ) ;
  assign n5461 = n4388 ^ n887 ^ 1'b0 ;
  assign n5462 = n3965 & n5461 ;
  assign n5463 = n5462 ^ n747 ^ 1'b0 ;
  assign n5464 = n2365 ^ n900 ^ x58 ;
  assign n5465 = n3242 & n5464 ;
  assign n5466 = n5465 ^ n1728 ^ 1'b0 ;
  assign n5467 = ( n1200 & ~n1201 ) | ( n1200 & n4053 ) | ( ~n1201 & n4053 ) ;
  assign n5468 = ( ~n1484 & n5466 ) | ( ~n1484 & n5467 ) | ( n5466 & n5467 ) ;
  assign n5470 = x93 & ~n823 ;
  assign n5469 = n1289 & n2983 ;
  assign n5471 = n5470 ^ n5469 ^ n4195 ;
  assign n5472 = n1454 ^ n505 ^ 1'b0 ;
  assign n5473 = ( n496 & n2295 ) | ( n496 & ~n3169 ) | ( n2295 & ~n3169 ) ;
  assign n5474 = n1781 & n2727 ;
  assign n5475 = n5474 ^ n1530 ^ 1'b0 ;
  assign n5476 = n3099 & ~n5475 ;
  assign n5477 = x41 & n1717 ;
  assign n5478 = ~n5476 & n5477 ;
  assign n5479 = ( n394 & ~n2038 ) | ( n394 & n5478 ) | ( ~n2038 & n5478 ) ;
  assign n5480 = ( n1665 & n1742 ) | ( n1665 & ~n2678 ) | ( n1742 & ~n2678 ) ;
  assign n5481 = ( x21 & ~n922 ) | ( x21 & n5480 ) | ( ~n922 & n5480 ) ;
  assign n5482 = n2238 ^ n2112 ^ 1'b0 ;
  assign n5483 = n1895 & n5482 ;
  assign n5484 = ( n2335 & n5481 ) | ( n2335 & ~n5483 ) | ( n5481 & ~n5483 ) ;
  assign n5485 = n3231 ^ n1203 ^ 1'b0 ;
  assign n5486 = n5485 ^ n3970 ^ n2976 ;
  assign n5490 = n1204 ^ x202 ^ 1'b0 ;
  assign n5491 = n4126 | n5490 ;
  assign n5489 = n1927 & n5193 ;
  assign n5492 = n5491 ^ n5489 ^ 1'b0 ;
  assign n5493 = n926 & n2189 ;
  assign n5494 = ~n5492 & n5493 ;
  assign n5487 = n2730 | n2964 ;
  assign n5488 = n5487 ^ n3105 ^ 1'b0 ;
  assign n5495 = n5494 ^ n5488 ^ 1'b0 ;
  assign n5497 = n3068 ^ n1951 ^ 1'b0 ;
  assign n5498 = n3097 & n5497 ;
  assign n5499 = n5498 ^ n3710 ^ 1'b0 ;
  assign n5500 = n5499 ^ n4693 ^ n804 ;
  assign n5496 = ( x245 & ~n2004 ) | ( x245 & n3979 ) | ( ~n2004 & n3979 ) ;
  assign n5501 = n5500 ^ n5496 ^ 1'b0 ;
  assign n5502 = n2157 ^ n1789 ^ n1352 ;
  assign n5503 = n5502 ^ n5274 ^ n509 ;
  assign n5504 = ( ~n3121 & n3361 ) | ( ~n3121 & n5503 ) | ( n3361 & n5503 ) ;
  assign n5505 = n4039 ^ n440 ^ 1'b0 ;
  assign n5506 = n2971 ^ n1720 ^ n1407 ;
  assign n5507 = n5506 ^ n3182 ^ x17 ;
  assign n5508 = n4695 & ~n5507 ;
  assign n5509 = n5508 ^ n1953 ^ 1'b0 ;
  assign n5510 = n1376 & ~n2118 ;
  assign n5511 = n5510 ^ n727 ^ 1'b0 ;
  assign n5512 = n1406 | n5511 ;
  assign n5513 = n297 & ~n5512 ;
  assign n5514 = n341 | n3305 ;
  assign n5515 = n259 & ~n5514 ;
  assign n5516 = n5513 & ~n5515 ;
  assign n5517 = n1361 | n2721 ;
  assign n5518 = n1058 | n5517 ;
  assign n5519 = n580 & n3656 ;
  assign n5520 = n5519 ^ n3037 ^ n1011 ;
  assign n5521 = ( x146 & ~n3130 ) | ( x146 & n3233 ) | ( ~n3130 & n3233 ) ;
  assign n5522 = ( n4776 & ~n5520 ) | ( n4776 & n5521 ) | ( ~n5520 & n5521 ) ;
  assign n5523 = ~n3821 & n5522 ;
  assign n5524 = ~n3568 & n5523 ;
  assign n5525 = n906 | n1497 ;
  assign n5526 = n3581 ^ n2619 ^ n1938 ;
  assign n5527 = n5526 ^ n4861 ^ 1'b0 ;
  assign n5528 = n3400 ^ n2921 ^ 1'b0 ;
  assign n5529 = n5528 ^ n2562 ^ 1'b0 ;
  assign n5530 = n5527 | n5529 ;
  assign n5531 = n5525 & ~n5530 ;
  assign n5532 = n1916 & n5531 ;
  assign n5533 = n3836 ^ n547 ^ 1'b0 ;
  assign n5534 = n911 | n5533 ;
  assign n5535 = n3454 ^ n2001 ^ 1'b0 ;
  assign n5537 = n1800 | n2802 ;
  assign n5538 = n5537 ^ n3795 ^ 1'b0 ;
  assign n5536 = n2046 ^ n275 ^ 1'b0 ;
  assign n5539 = n5538 ^ n5536 ^ 1'b0 ;
  assign n5540 = n565 | n2794 ;
  assign n5541 = n2227 & ~n5540 ;
  assign n5542 = n2019 & ~n5541 ;
  assign n5543 = n4421 ^ n1145 ^ 1'b0 ;
  assign n5544 = ( n807 & n5542 ) | ( n807 & ~n5543 ) | ( n5542 & ~n5543 ) ;
  assign n5545 = ( ~x169 & n1290 ) | ( ~x169 & n5069 ) | ( n1290 & n5069 ) ;
  assign n5546 = ( x201 & n1446 ) | ( x201 & ~n5545 ) | ( n1446 & ~n5545 ) ;
  assign n5547 = n516 & n874 ;
  assign n5548 = n4108 & n5547 ;
  assign n5549 = ( n1012 & n2403 ) | ( n1012 & n2852 ) | ( n2403 & n2852 ) ;
  assign n5550 = n843 & ~n5549 ;
  assign n5551 = n5550 ^ n4383 ^ 1'b0 ;
  assign n5552 = ~n5548 & n5551 ;
  assign n5553 = n2016 & n2204 ;
  assign n5554 = n970 & ~n1275 ;
  assign n5555 = n1280 & n2833 ;
  assign n5556 = n5554 & n5555 ;
  assign n5557 = ( n2245 & ~n2517 ) | ( n2245 & n3054 ) | ( ~n2517 & n3054 ) ;
  assign n5558 = n387 & n3067 ;
  assign n5559 = ~n3067 & n5558 ;
  assign n5560 = ~n633 & n5559 ;
  assign n5561 = x151 & ~n5560 ;
  assign n5562 = n5557 & n5561 ;
  assign n5563 = n1671 & n2106 ;
  assign n5564 = n5562 & n5563 ;
  assign n5565 = ( n1073 & ~n1480 ) | ( n1073 & n2680 ) | ( ~n1480 & n2680 ) ;
  assign n5566 = n1337 | n5565 ;
  assign n5567 = n1561 | n5566 ;
  assign n5568 = ~n3335 & n5567 ;
  assign n5569 = n3476 & n5568 ;
  assign n5573 = ~n1789 & n2924 ;
  assign n5574 = n2136 & n3299 ;
  assign n5575 = n5574 ^ n1558 ^ 1'b0 ;
  assign n5576 = ( x154 & ~n5573 ) | ( x154 & n5575 ) | ( ~n5573 & n5575 ) ;
  assign n5570 = ( x5 & ~x84 ) | ( x5 & n2205 ) | ( ~x84 & n2205 ) ;
  assign n5571 = n3169 | n5570 ;
  assign n5572 = n4592 & ~n5571 ;
  assign n5577 = n5576 ^ n5572 ^ n2341 ;
  assign n5578 = n5577 ^ n4084 ^ n2953 ;
  assign n5579 = n4009 & ~n4814 ;
  assign n5580 = n5579 ^ n3722 ^ n2204 ;
  assign n5581 = ~n499 & n2208 ;
  assign n5582 = n5581 ^ n2021 ^ 1'b0 ;
  assign n5585 = n459 ^ x191 ^ 1'b0 ;
  assign n5586 = n684 | n5585 ;
  assign n5587 = ~n722 & n1183 ;
  assign n5588 = n5586 & n5587 ;
  assign n5584 = n3526 ^ n1482 ^ 1'b0 ;
  assign n5583 = n2852 & ~n5185 ;
  assign n5589 = n5588 ^ n5584 ^ n5583 ;
  assign n5590 = ~n5582 & n5589 ;
  assign n5591 = ~n5580 & n5590 ;
  assign n5592 = n5376 ^ n2310 ^ n814 ;
  assign n5593 = n259 | n4932 ;
  assign n5594 = n1736 | n5593 ;
  assign n5595 = n2835 | n3533 ;
  assign n5596 = n4695 ^ n4121 ^ n1453 ;
  assign n5597 = ~n5595 & n5596 ;
  assign n5598 = ~n841 & n5597 ;
  assign n5599 = ( n559 & n5594 ) | ( n559 & ~n5598 ) | ( n5594 & ~n5598 ) ;
  assign n5601 = n5389 ^ n3544 ^ n642 ;
  assign n5600 = n1685 | n1707 ;
  assign n5602 = n5601 ^ n5600 ^ 1'b0 ;
  assign n5603 = n3074 ^ n2005 ^ n676 ;
  assign n5604 = ( n829 & n1276 ) | ( n829 & ~n1499 ) | ( n1276 & ~n1499 ) ;
  assign n5605 = n5604 ^ n3175 ^ 1'b0 ;
  assign n5606 = n1875 & n5605 ;
  assign n5607 = n3412 ^ n1499 ^ n1024 ;
  assign n5608 = ~n1108 & n5607 ;
  assign n5609 = n2706 ^ n2157 ^ x137 ;
  assign n5610 = n3072 & n5609 ;
  assign n5611 = n5610 ^ n4041 ^ 1'b0 ;
  assign n5612 = n3763 ^ n1590 ^ x11 ;
  assign n5613 = n5612 ^ n4236 ^ 1'b0 ;
  assign n5614 = n4456 ^ n3422 ^ 1'b0 ;
  assign n5615 = x114 & n5614 ;
  assign n5616 = n3819 ^ n1126 ^ 1'b0 ;
  assign n5617 = x250 & ~n515 ;
  assign n5618 = ~n983 & n5617 ;
  assign n5619 = n5618 ^ n4595 ^ n4060 ;
  assign n5620 = n4500 ^ n1702 ^ 1'b0 ;
  assign n5621 = ~n1133 & n5620 ;
  assign n5622 = ( n2279 & n5324 ) | ( n2279 & n5621 ) | ( n5324 & n5621 ) ;
  assign n5623 = n823 & ~n5613 ;
  assign n5624 = n4276 ^ n676 ^ 1'b0 ;
  assign n5625 = n5114 | n5624 ;
  assign n5626 = ( n1510 & ~n2844 ) | ( n1510 & n4587 ) | ( ~n2844 & n4587 ) ;
  assign n5628 = n1288 ^ x120 ^ 1'b0 ;
  assign n5627 = n363 | n3810 ;
  assign n5629 = n5628 ^ n5627 ^ n2284 ;
  assign n5630 = ~n4432 & n5629 ;
  assign n5631 = n4528 & n5630 ;
  assign n5632 = n5631 ^ n1103 ^ 1'b0 ;
  assign n5637 = n2462 ^ n741 ^ n535 ;
  assign n5633 = n1064 & n3242 ;
  assign n5634 = n5633 ^ n1243 ^ 1'b0 ;
  assign n5635 = n1031 & ~n5634 ;
  assign n5636 = ~n1923 & n5635 ;
  assign n5638 = n5637 ^ n5636 ^ 1'b0 ;
  assign n5639 = n1035 & n2667 ;
  assign n5640 = n5639 ^ n4153 ^ 1'b0 ;
  assign n5641 = ~n4645 & n5640 ;
  assign n5642 = ( x59 & ~n1232 ) | ( x59 & n2885 ) | ( ~n1232 & n2885 ) ;
  assign n5643 = n3519 ^ n1047 ^ 1'b0 ;
  assign n5645 = n2112 | n3349 ;
  assign n5644 = ~n1328 & n3528 ;
  assign n5646 = n5645 ^ n5644 ^ 1'b0 ;
  assign n5647 = x155 & ~n2451 ;
  assign n5648 = ~n922 & n5647 ;
  assign n5649 = ( n1492 & n2752 ) | ( n1492 & ~n5648 ) | ( n2752 & ~n5648 ) ;
  assign n5650 = ( ~n1399 & n3865 ) | ( ~n1399 & n4978 ) | ( n3865 & n4978 ) ;
  assign n5652 = x25 & x58 ;
  assign n5653 = ~n2242 & n5652 ;
  assign n5654 = n3317 | n5653 ;
  assign n5655 = n794 | n5654 ;
  assign n5656 = n5655 ^ n5373 ^ 1'b0 ;
  assign n5657 = n3710 & n5656 ;
  assign n5658 = n5657 ^ n1848 ^ 1'b0 ;
  assign n5651 = n5170 | n5621 ;
  assign n5659 = n5658 ^ n5651 ^ 1'b0 ;
  assign n5660 = ( n1588 & n2788 ) | ( n1588 & n4111 ) | ( n2788 & n4111 ) ;
  assign n5661 = n5660 ^ n3370 ^ 1'b0 ;
  assign n5662 = n4098 & ~n5661 ;
  assign n5664 = ( n703 & n1588 ) | ( n703 & n2270 ) | ( n1588 & n2270 ) ;
  assign n5663 = n1156 | n4829 ;
  assign n5665 = n5664 ^ n5663 ^ 1'b0 ;
  assign n5666 = n5665 ^ n4247 ^ n3885 ;
  assign n5667 = n1775 | n5358 ;
  assign n5668 = n2806 & ~n4618 ;
  assign n5669 = ~n5667 & n5668 ;
  assign n5670 = n5669 ^ n1755 ^ 1'b0 ;
  assign n5671 = n1527 | n1789 ;
  assign n5672 = x171 & n5671 ;
  assign n5673 = ~n3816 & n5672 ;
  assign n5674 = n5673 ^ n4791 ^ 1'b0 ;
  assign n5675 = n2919 ^ n1725 ^ 1'b0 ;
  assign n5676 = n4563 ^ n702 ^ 1'b0 ;
  assign n5677 = n2924 ^ n1197 ^ 1'b0 ;
  assign n5678 = n1715 & n4151 ;
  assign n5679 = n5677 & n5678 ;
  assign n5683 = n945 & n1455 ;
  assign n5684 = n5683 ^ n1040 ^ 1'b0 ;
  assign n5680 = n4475 ^ n1567 ^ 1'b0 ;
  assign n5681 = n1382 | n4107 ;
  assign n5682 = n5680 & n5681 ;
  assign n5685 = n5684 ^ n5682 ^ n4902 ;
  assign n5686 = ( ~n5088 & n5679 ) | ( ~n5088 & n5685 ) | ( n5679 & n5685 ) ;
  assign n5687 = n1613 | n1968 ;
  assign n5688 = n1258 ^ n1024 ^ 1'b0 ;
  assign n5689 = n5687 | n5688 ;
  assign n5690 = n3790 ^ n1107 ^ 1'b0 ;
  assign n5694 = ~n1365 & n3400 ;
  assign n5695 = n5694 ^ n3444 ^ 1'b0 ;
  assign n5691 = n838 ^ n711 ^ 1'b0 ;
  assign n5692 = n1943 & ~n5691 ;
  assign n5693 = n4457 & n5692 ;
  assign n5696 = n5695 ^ n5693 ^ 1'b0 ;
  assign n5697 = ( ~n1453 & n4411 ) | ( ~n1453 & n5696 ) | ( n4411 & n5696 ) ;
  assign n5698 = ( n1963 & n2445 ) | ( n1963 & ~n3755 ) | ( n2445 & ~n3755 ) ;
  assign n5699 = n2427 & n5698 ;
  assign n5700 = x182 & ~n2423 ;
  assign n5701 = n5700 ^ n2957 ^ 1'b0 ;
  assign n5702 = n5701 ^ n3990 ^ 1'b0 ;
  assign n5703 = n3091 & ~n4986 ;
  assign n5704 = n5703 ^ n434 ^ 1'b0 ;
  assign n5705 = ( n3128 & n3349 ) | ( n3128 & ~n4170 ) | ( n3349 & ~n4170 ) ;
  assign n5706 = ( x33 & n883 ) | ( x33 & n5705 ) | ( n883 & n5705 ) ;
  assign n5707 = n5706 ^ n3447 ^ n3039 ;
  assign n5708 = n3470 & n5707 ;
  assign n5709 = n5708 ^ n1133 ^ 1'b0 ;
  assign n5711 = x17 & n635 ;
  assign n5712 = n5711 ^ n2448 ^ 1'b0 ;
  assign n5710 = ~n1058 & n2306 ;
  assign n5713 = n5712 ^ n5710 ^ n3647 ;
  assign n5714 = n453 | n4781 ;
  assign n5715 = n1452 & ~n5714 ;
  assign n5716 = n838 & ~n5715 ;
  assign n5717 = ~n5713 & n5716 ;
  assign n5718 = ~n1635 & n3344 ;
  assign n5719 = n4346 ^ n2543 ^ 1'b0 ;
  assign n5720 = n5718 & ~n5719 ;
  assign n5721 = n5717 & n5720 ;
  assign n5722 = n587 ^ n479 ^ x158 ;
  assign n5723 = n2517 & n5722 ;
  assign n5724 = n973 & n2426 ;
  assign n5725 = ~n5723 & n5724 ;
  assign n5726 = n5725 ^ n3960 ^ 1'b0 ;
  assign n5727 = ~n2680 & n3178 ;
  assign n5728 = n1374 & n5727 ;
  assign n5729 = n3034 & ~n5728 ;
  assign n5730 = ~n297 & n1294 ;
  assign n5731 = n5730 ^ n3053 ^ 1'b0 ;
  assign n5732 = x104 | n815 ;
  assign n5733 = n5732 ^ n2994 ^ 1'b0 ;
  assign n5734 = n1094 & ~n5733 ;
  assign n5735 = n5731 & n5734 ;
  assign n5736 = ~n5729 & n5735 ;
  assign n5737 = n5736 ^ n5226 ^ n2907 ;
  assign n5738 = x242 & ~n5737 ;
  assign n5739 = n5738 ^ n957 ^ 1'b0 ;
  assign n5740 = n3047 ^ n1724 ^ n1213 ;
  assign n5741 = n5740 ^ n3304 ^ n2077 ;
  assign n5742 = n5741 ^ n4145 ^ n3185 ;
  assign n5743 = n5363 ^ n4027 ^ 1'b0 ;
  assign n5744 = n1890 | n5743 ;
  assign n5745 = n1324 & ~n1687 ;
  assign n5746 = ( n3181 & n5744 ) | ( n3181 & n5745 ) | ( n5744 & n5745 ) ;
  assign n5747 = n1671 & n3514 ;
  assign n5748 = n2478 & ~n5747 ;
  assign n5749 = n3771 ^ n1687 ^ 1'b0 ;
  assign n5750 = n3066 ^ x152 ^ 1'b0 ;
  assign n5751 = n2311 & ~n5750 ;
  assign n5752 = ( x115 & x163 ) | ( x115 & ~n771 ) | ( x163 & ~n771 ) ;
  assign n5753 = n2723 ^ n1040 ^ 1'b0 ;
  assign n5754 = ( x31 & n2945 ) | ( x31 & n5753 ) | ( n2945 & n5753 ) ;
  assign n5755 = ~n4554 & n5754 ;
  assign n5756 = n1206 & n1804 ;
  assign n5768 = n522 & ~n1671 ;
  assign n5757 = n2529 | n3532 ;
  assign n5758 = n2264 | n5757 ;
  assign n5759 = n1658 ^ n694 ^ 1'b0 ;
  assign n5760 = n5759 ^ n3573 ^ n360 ;
  assign n5763 = n1438 | n1647 ;
  assign n5761 = n1388 ^ n405 ^ 1'b0 ;
  assign n5762 = ( x8 & n2092 ) | ( x8 & ~n5761 ) | ( n2092 & ~n5761 ) ;
  assign n5764 = n5763 ^ n5762 ^ 1'b0 ;
  assign n5765 = n3474 & ~n5764 ;
  assign n5766 = n1372 & n5765 ;
  assign n5767 = ( n5758 & n5760 ) | ( n5758 & n5766 ) | ( n5760 & n5766 ) ;
  assign n5769 = n5768 ^ n5767 ^ 1'b0 ;
  assign n5770 = n1647 & ~n5769 ;
  assign n5771 = n1179 ^ n913 ^ x57 ;
  assign n5772 = ~n2605 & n5118 ;
  assign n5773 = ~n4756 & n5772 ;
  assign n5774 = n4113 & ~n5773 ;
  assign n5775 = ~n5771 & n5774 ;
  assign n5776 = n3223 ^ n2811 ^ 1'b0 ;
  assign n5780 = ~n3156 & n3920 ;
  assign n5781 = n987 & n5780 ;
  assign n5777 = n1731 ^ n1564 ^ n586 ;
  assign n5778 = n752 ^ n345 ^ 1'b0 ;
  assign n5779 = ( ~x8 & n5777 ) | ( ~x8 & n5778 ) | ( n5777 & n5778 ) ;
  assign n5782 = n5781 ^ n5779 ^ n5289 ;
  assign n5783 = ~n5776 & n5782 ;
  assign n5784 = ~n1155 & n5783 ;
  assign n5790 = n922 & n2222 ;
  assign n5791 = n5790 ^ n679 ^ 1'b0 ;
  assign n5785 = n1622 ^ n1506 ^ 1'b0 ;
  assign n5786 = x212 & ~n5785 ;
  assign n5787 = n5786 ^ n4661 ^ 1'b0 ;
  assign n5788 = n5787 ^ n2880 ^ 1'b0 ;
  assign n5789 = n4441 & ~n5788 ;
  assign n5792 = n5791 ^ n5789 ^ n539 ;
  assign n5793 = ( n4413 & n5055 ) | ( n4413 & ~n5285 ) | ( n5055 & ~n5285 ) ;
  assign n5794 = x159 & n4197 ;
  assign n5795 = n5794 ^ n1522 ^ 1'b0 ;
  assign n5796 = ( ~n2150 & n3761 ) | ( ~n2150 & n4825 ) | ( n3761 & n4825 ) ;
  assign n5797 = ~n1047 & n3087 ;
  assign n5798 = n5797 ^ n3097 ^ n493 ;
  assign n5805 = ( x83 & n1046 ) | ( x83 & ~n1494 ) | ( n1046 & ~n1494 ) ;
  assign n5799 = n1928 & n3402 ;
  assign n5800 = n5799 ^ n1079 ^ 1'b0 ;
  assign n5801 = ( x210 & n1120 ) | ( x210 & ~n5800 ) | ( n1120 & ~n5800 ) ;
  assign n5802 = n2035 & ~n2860 ;
  assign n5803 = n5802 ^ n604 ^ 1'b0 ;
  assign n5804 = ~n5801 & n5803 ;
  assign n5806 = n5805 ^ n5804 ^ n4635 ;
  assign n5807 = n2769 ^ n1598 ^ 1'b0 ;
  assign n5808 = n3831 ^ n795 ^ 1'b0 ;
  assign n5809 = n3184 & n5808 ;
  assign n5810 = ~n2875 & n5809 ;
  assign n5811 = n5807 & ~n5810 ;
  assign n5812 = n5811 ^ n4202 ^ 1'b0 ;
  assign n5813 = ( n4232 & n4735 ) | ( n4232 & ~n5812 ) | ( n4735 & ~n5812 ) ;
  assign n5814 = n3672 | n5813 ;
  assign n5815 = n1508 & n4747 ;
  assign n5816 = n5815 ^ n2942 ^ 1'b0 ;
  assign n5817 = ( n1252 & n5688 ) | ( n1252 & ~n5816 ) | ( n5688 & ~n5816 ) ;
  assign n5818 = n256 & n2279 ;
  assign n5819 = x243 | n1585 ;
  assign n5820 = n5819 ^ n3413 ^ 1'b0 ;
  assign n5821 = n5818 & ~n5820 ;
  assign n5822 = n4086 & n4614 ;
  assign n5823 = x169 & n5822 ;
  assign n5824 = n5632 ^ n1201 ^ 1'b0 ;
  assign n5825 = ~n1145 & n2396 ;
  assign n5826 = n3389 ^ n3117 ^ n1506 ;
  assign n5827 = n4783 ^ n1882 ^ n507 ;
  assign n5828 = ( n4862 & n5826 ) | ( n4862 & ~n5827 ) | ( n5826 & ~n5827 ) ;
  assign n5829 = x72 & n2558 ;
  assign n5830 = n2013 & n5829 ;
  assign n5831 = n5830 ^ n4815 ^ 1'b0 ;
  assign n5832 = n1707 | n5831 ;
  assign n5833 = n2520 ^ n1908 ^ 1'b0 ;
  assign n5834 = n2294 | n5833 ;
  assign n5835 = n3369 ^ n2509 ^ 1'b0 ;
  assign n5836 = x225 & n5835 ;
  assign n5837 = n1750 & n4118 ;
  assign n5838 = ( n5525 & ~n5768 ) | ( n5525 & n5837 ) | ( ~n5768 & n5837 ) ;
  assign n5839 = x4 | n913 ;
  assign n5840 = n4425 & n5839 ;
  assign n5841 = n5840 ^ n1322 ^ 1'b0 ;
  assign n5842 = n4935 ^ n4542 ^ x188 ;
  assign n5843 = ( ~n1226 & n3371 ) | ( ~n1226 & n5842 ) | ( n3371 & n5842 ) ;
  assign n5844 = n3781 | n5843 ;
  assign n5845 = n1044 | n2209 ;
  assign n5846 = n3839 | n5845 ;
  assign n5847 = ~n3675 & n5846 ;
  assign n5848 = n5847 ^ x247 ^ 1'b0 ;
  assign n5849 = n1074 & ~n3939 ;
  assign n5850 = n5849 ^ n3324 ^ 1'b0 ;
  assign n5855 = ( n2867 & n3915 ) | ( n2867 & ~n4001 ) | ( n3915 & ~n4001 ) ;
  assign n5851 = n5017 ^ n4080 ^ n3342 ;
  assign n5852 = ~n339 & n1628 ;
  assign n5853 = x164 & ~n5852 ;
  assign n5854 = ~n5851 & n5853 ;
  assign n5856 = n5855 ^ n5854 ^ 1'b0 ;
  assign n5857 = ( n264 & n1776 ) | ( n264 & ~n5108 ) | ( n1776 & ~n5108 ) ;
  assign n5858 = n5857 ^ n4927 ^ n4034 ;
  assign n5859 = ( n381 & ~n1537 ) | ( n381 & n4901 ) | ( ~n1537 & n4901 ) ;
  assign n5860 = x39 & ~n544 ;
  assign n5861 = n1334 | n1524 ;
  assign n5862 = n3545 | n5861 ;
  assign n5863 = n5862 ^ n3352 ^ 1'b0 ;
  assign n5864 = n5863 ^ n4400 ^ 1'b0 ;
  assign n5865 = n3762 | n5864 ;
  assign n5866 = n1978 | n5289 ;
  assign n5867 = x24 | n5866 ;
  assign n5868 = ( n897 & n2119 ) | ( n897 & ~n2884 ) | ( n2119 & ~n2884 ) ;
  assign n5869 = n5868 ^ n2827 ^ 1'b0 ;
  assign n5870 = n5345 ^ n2172 ^ n887 ;
  assign n5871 = n2582 & n3257 ;
  assign n5872 = n5871 ^ n3985 ^ 1'b0 ;
  assign n5873 = n5872 ^ n2287 ^ 1'b0 ;
  assign n5874 = n4510 ^ n4133 ^ n2105 ;
  assign n5875 = n1717 | n2292 ;
  assign n5876 = n2538 ^ n490 ^ 1'b0 ;
  assign n5877 = ~n5875 & n5876 ;
  assign n5878 = n3091 ^ n2329 ^ 1'b0 ;
  assign n5879 = n3002 | n5188 ;
  assign n5880 = n4132 & ~n5879 ;
  assign n5881 = ~n798 & n5880 ;
  assign n5882 = n5881 ^ n4443 ^ n3900 ;
  assign n5884 = n3196 ^ n1402 ^ n1389 ;
  assign n5885 = n5884 ^ n1553 ^ x173 ;
  assign n5883 = ( n632 & ~n733 ) | ( n632 & n4342 ) | ( ~n733 & n4342 ) ;
  assign n5886 = n5885 ^ n5883 ^ n3123 ;
  assign n5888 = n500 | n2355 ;
  assign n5889 = ( x113 & n3070 ) | ( x113 & n5888 ) | ( n3070 & n5888 ) ;
  assign n5890 = n2688 & n5889 ;
  assign n5891 = n464 & n5890 ;
  assign n5887 = ~n1772 & n3472 ;
  assign n5892 = n5891 ^ n5887 ^ 1'b0 ;
  assign n5893 = ~n4008 & n5892 ;
  assign n5894 = n5631 ^ n2039 ^ 1'b0 ;
  assign n5895 = ( n1291 & n4604 ) | ( n1291 & ~n4970 ) | ( n4604 & ~n4970 ) ;
  assign n5896 = n1301 & n2916 ;
  assign n5897 = ~n1455 & n5896 ;
  assign n5898 = ( n528 & ~n3712 ) | ( n528 & n5897 ) | ( ~n3712 & n5897 ) ;
  assign n5899 = n5159 | n5764 ;
  assign n5900 = n3910 ^ n3112 ^ 1'b0 ;
  assign n5901 = ~n1823 & n5900 ;
  assign n5903 = ( ~n672 & n1933 ) | ( ~n672 & n2414 ) | ( n1933 & n2414 ) ;
  assign n5902 = n3363 | n4424 ;
  assign n5904 = n5903 ^ n5902 ^ 1'b0 ;
  assign n5908 = n1985 ^ n1855 ^ 1'b0 ;
  assign n5909 = n1073 & n5908 ;
  assign n5905 = ( ~x114 & x231 ) | ( ~x114 & n575 ) | ( x231 & n575 ) ;
  assign n5906 = n3354 | n5905 ;
  assign n5907 = n4045 | n5906 ;
  assign n5910 = n5909 ^ n5907 ^ 1'b0 ;
  assign n5911 = n5904 & n5910 ;
  assign n5912 = ~n1224 & n2405 ;
  assign n5915 = n2416 ^ n1142 ^ 1'b0 ;
  assign n5916 = ( n2326 & n5139 ) | ( n2326 & n5915 ) | ( n5139 & n5915 ) ;
  assign n5913 = n5579 ^ n1094 ^ 1'b0 ;
  assign n5914 = n5913 ^ n4952 ^ 1'b0 ;
  assign n5917 = n5916 ^ n5914 ^ 1'b0 ;
  assign n5918 = ~n1602 & n5917 ;
  assign n5919 = n4535 ^ n4187 ^ 1'b0 ;
  assign n5920 = n5919 ^ n2526 ^ n839 ;
  assign n5921 = n1018 & n5920 ;
  assign n5922 = n5921 ^ n5762 ^ 1'b0 ;
  assign n5923 = n2299 ^ n2235 ^ n951 ;
  assign n5927 = n5114 ^ n1034 ^ 1'b0 ;
  assign n5924 = n294 & n764 ;
  assign n5925 = n1236 & n5924 ;
  assign n5926 = n5925 ^ n1200 ^ n925 ;
  assign n5928 = n5927 ^ n5926 ^ n2942 ;
  assign n5929 = ( ~x0 & x196 ) | ( ~x0 & n4601 ) | ( x196 & n4601 ) ;
  assign n5930 = n1484 & ~n5929 ;
  assign n5931 = n5928 & n5930 ;
  assign n5932 = n4975 | n5931 ;
  assign n5933 = n5923 | n5932 ;
  assign n5938 = n2794 & ~n3810 ;
  assign n5939 = n2957 & ~n3436 ;
  assign n5940 = ~n1549 & n5939 ;
  assign n5941 = n411 | n5940 ;
  assign n5942 = n5938 & ~n5941 ;
  assign n5934 = n3210 ^ n2651 ^ n1736 ;
  assign n5935 = n3410 & ~n5934 ;
  assign n5936 = n4940 ^ n2019 ^ 1'b0 ;
  assign n5937 = ( n4307 & n5935 ) | ( n4307 & n5936 ) | ( n5935 & n5936 ) ;
  assign n5943 = n5942 ^ n5937 ^ 1'b0 ;
  assign n5944 = n4745 & n5943 ;
  assign n5945 = n1116 & n3552 ;
  assign n5946 = ~n2549 & n3376 ;
  assign n5947 = n615 & n5946 ;
  assign n5948 = n5947 ^ n5573 ^ 1'b0 ;
  assign n5949 = n4257 | n5948 ;
  assign n5950 = ( n1051 & n1821 ) | ( n1051 & ~n5949 ) | ( n1821 & ~n5949 ) ;
  assign n5951 = n1275 & ~n3335 ;
  assign n5952 = n5951 ^ n1173 ^ 1'b0 ;
  assign n5953 = n1602 ^ n703 ^ 1'b0 ;
  assign n5954 = n4095 & ~n5953 ;
  assign n5955 = n2189 & ~n4128 ;
  assign n5956 = n1002 & n5955 ;
  assign n5957 = n5956 ^ n2971 ^ 1'b0 ;
  assign n5958 = n2141 & n5957 ;
  assign n5959 = ( n1516 & n3025 ) | ( n1516 & n3902 ) | ( n3025 & n3902 ) ;
  assign n5960 = n4689 ^ n288 ^ 1'b0 ;
  assign n5961 = x244 & n5960 ;
  assign n5962 = ~n4038 & n5961 ;
  assign n5963 = n1980 & n5962 ;
  assign n5965 = n3130 ^ n2861 ^ n1951 ;
  assign n5966 = n1203 | n5965 ;
  assign n5967 = n5966 ^ x251 ^ 1'b0 ;
  assign n5964 = ~n1334 & n2860 ;
  assign n5968 = n5967 ^ n5964 ^ 1'b0 ;
  assign n5969 = x170 & n5968 ;
  assign n5971 = n3615 ^ n913 ^ 1'b0 ;
  assign n5972 = n2221 & n5971 ;
  assign n5970 = n1633 & ~n2910 ;
  assign n5973 = n5972 ^ n5970 ^ 1'b0 ;
  assign n5974 = ~n818 & n1475 ;
  assign n5975 = n5974 ^ n2595 ^ 1'b0 ;
  assign n5976 = ( n1543 & n2860 ) | ( n1543 & n5975 ) | ( n2860 & n5975 ) ;
  assign n5977 = n3325 & ~n4162 ;
  assign n5978 = n5977 ^ n522 ^ 1'b0 ;
  assign n5979 = x57 & ~n4874 ;
  assign n5980 = n5979 ^ n676 ^ 1'b0 ;
  assign n5981 = ~n2315 & n5980 ;
  assign n5982 = x204 & n5981 ;
  assign n5983 = ~n2033 & n5903 ;
  assign n5984 = n5983 ^ n326 ^ 1'b0 ;
  assign n5985 = n2740 ^ n571 ^ 1'b0 ;
  assign n5986 = ( n1012 & n1302 ) | ( n1012 & ~n5985 ) | ( n1302 & ~n5985 ) ;
  assign n5987 = n3864 & n4237 ;
  assign n5988 = ( n5984 & ~n5986 ) | ( n5984 & n5987 ) | ( ~n5986 & n5987 ) ;
  assign n5989 = n5139 | n5988 ;
  assign n5990 = ( ~x76 & x116 ) | ( ~x76 & n1366 ) | ( x116 & n1366 ) ;
  assign n5991 = n756 ^ n460 ^ 1'b0 ;
  assign n5992 = ~x178 & n2589 ;
  assign n5993 = n5991 | n5992 ;
  assign n5994 = n1886 | n4760 ;
  assign n5995 = n5994 ^ n1115 ^ 1'b0 ;
  assign n5996 = n3361 & ~n5995 ;
  assign n5997 = n5996 ^ n1202 ^ 1'b0 ;
  assign n5998 = n1694 | n5997 ;
  assign n5999 = x48 & ~n3979 ;
  assign n6000 = n5620 ^ n2292 ^ n639 ;
  assign n6001 = ( n4049 & n4692 ) | ( n4049 & ~n6000 ) | ( n4692 & ~n6000 ) ;
  assign n6002 = n3853 & n6001 ;
  assign n6003 = n6002 ^ n4589 ^ 1'b0 ;
  assign n6006 = n259 | n3316 ;
  assign n6004 = x123 & n1388 ;
  assign n6005 = ~n4777 & n6004 ;
  assign n6007 = n6006 ^ n6005 ^ 1'b0 ;
  assign n6008 = n3532 | n6007 ;
  assign n6009 = x135 & n627 ;
  assign n6010 = n2661 & n6009 ;
  assign n6011 = n5786 ^ n3020 ^ 1'b0 ;
  assign n6012 = x86 & n715 ;
  assign n6013 = x239 & n5372 ;
  assign n6014 = n6013 ^ n1161 ^ 1'b0 ;
  assign n6015 = n2790 ^ n2204 ^ n740 ;
  assign n6016 = x197 & ~n1995 ;
  assign n6017 = n6016 ^ n4425 ^ 1'b0 ;
  assign n6018 = ~n6015 & n6017 ;
  assign n6019 = n6018 ^ n5584 ^ n2042 ;
  assign n6020 = n1236 ^ n876 ^ 1'b0 ;
  assign n6021 = ( n3583 & n4434 ) | ( n3583 & ~n5697 ) | ( n4434 & ~n5697 ) ;
  assign n6026 = n2098 & n2314 ;
  assign n6027 = ~n647 & n6026 ;
  assign n6022 = ~n1859 & n2462 ;
  assign n6023 = n6022 ^ x150 ^ 1'b0 ;
  assign n6024 = ( n559 & n740 ) | ( n559 & ~n6023 ) | ( n740 & ~n6023 ) ;
  assign n6025 = n6024 ^ n1583 ^ 1'b0 ;
  assign n6028 = n6027 ^ n6025 ^ n1580 ;
  assign n6029 = n1789 & n4767 ;
  assign n6030 = n1605 ^ x68 ^ 1'b0 ;
  assign n6031 = n6030 ^ n1500 ^ 1'b0 ;
  assign n6032 = n3240 | n6031 ;
  assign n6033 = x224 & ~n6032 ;
  assign n6034 = n6033 ^ n3561 ^ 1'b0 ;
  assign n6035 = n862 & n2105 ;
  assign n6036 = n6035 ^ n537 ^ 1'b0 ;
  assign n6037 = n4036 & n6036 ;
  assign n6038 = ( n4578 & n6034 ) | ( n4578 & n6037 ) | ( n6034 & n6037 ) ;
  assign n6039 = n1258 ^ n481 ^ 1'b0 ;
  assign n6040 = n5226 ^ n4882 ^ 1'b0 ;
  assign n6041 = n1434 & ~n6040 ;
  assign n6042 = n1451 & n3327 ;
  assign n6043 = n1115 & n6042 ;
  assign n6044 = n3160 | n6043 ;
  assign n6045 = n5429 & ~n6044 ;
  assign n6046 = ( ~n1653 & n2406 ) | ( ~n1653 & n4405 ) | ( n2406 & n4405 ) ;
  assign n6047 = n6046 ^ n4277 ^ n2654 ;
  assign n6048 = x170 | n6047 ;
  assign n6049 = n459 | n1189 ;
  assign n6050 = n471 | n6049 ;
  assign n6051 = ( ~x27 & n3826 ) | ( ~x27 & n6050 ) | ( n3826 & n6050 ) ;
  assign n6052 = n6051 ^ n557 ^ 1'b0 ;
  assign n6053 = n1270 & ~n3679 ;
  assign n6054 = ~n3188 & n5904 ;
  assign n6055 = n6054 ^ n343 ^ 1'b0 ;
  assign n6056 = n6053 & ~n6055 ;
  assign n6057 = n3843 & ~n5991 ;
  assign n6058 = ~n4149 & n6057 ;
  assign n6059 = n4432 ^ n2005 ^ 1'b0 ;
  assign n6060 = n3277 & ~n6059 ;
  assign n6063 = ( x91 & ~n2798 ) | ( x91 & n2821 ) | ( ~n2798 & n2821 ) ;
  assign n6061 = ~n1750 & n4777 ;
  assign n6062 = n6061 ^ n1597 ^ 1'b0 ;
  assign n6064 = n6063 ^ n6062 ^ 1'b0 ;
  assign n6065 = n6064 ^ n3963 ^ 1'b0 ;
  assign n6066 = n5745 & ~n6065 ;
  assign n6067 = n2752 & ~n4884 ;
  assign n6068 = ~n2004 & n6067 ;
  assign n6069 = ( x51 & n3275 ) | ( x51 & n6068 ) | ( n3275 & n6068 ) ;
  assign n6070 = ( n2449 & n3833 ) | ( n2449 & n6069 ) | ( n3833 & n6069 ) ;
  assign n6071 = ( ~n411 & n692 ) | ( ~n411 & n1080 ) | ( n692 & n1080 ) ;
  assign n6072 = n5291 & n6071 ;
  assign n6073 = n6072 ^ n1322 ^ 1'b0 ;
  assign n6074 = n6073 ^ n3097 ^ 1'b0 ;
  assign n6077 = n273 | n3409 ;
  assign n6075 = ( n862 & n1429 ) | ( n862 & n3593 ) | ( n1429 & n3593 ) ;
  assign n6076 = n4084 & n6075 ;
  assign n6078 = n6077 ^ n6076 ^ 1'b0 ;
  assign n6079 = n5058 ^ n4438 ^ 1'b0 ;
  assign n6080 = ~n1024 & n6079 ;
  assign n6081 = n5294 ^ n4865 ^ 1'b0 ;
  assign n6082 = ~n401 & n6081 ;
  assign n6083 = n6082 ^ x135 ^ 1'b0 ;
  assign n6084 = ~n381 & n6083 ;
  assign n6085 = ~n703 & n6084 ;
  assign n6086 = n1441 & ~n1870 ;
  assign n6087 = n4039 | n6086 ;
  assign n6088 = n1294 & ~n3185 ;
  assign n6089 = n4832 | n6088 ;
  assign n6090 = n4744 | n6089 ;
  assign n6091 = ( n2701 & n6087 ) | ( n2701 & ~n6090 ) | ( n6087 & ~n6090 ) ;
  assign n6092 = x218 | n861 ;
  assign n6093 = n6092 ^ n4298 ^ 1'b0 ;
  assign n6094 = n1418 ^ n1316 ^ 1'b0 ;
  assign n6095 = n3325 ^ n2335 ^ 1'b0 ;
  assign n6096 = n2903 & n6095 ;
  assign n6097 = n6096 ^ n4374 ^ n2824 ;
  assign n6098 = n6097 ^ n5298 ^ n4838 ;
  assign n6099 = x251 ^ x19 ^ 1'b0 ;
  assign n6100 = ( n1084 & n1602 ) | ( n1084 & ~n4034 ) | ( n1602 & ~n4034 ) ;
  assign n6104 = n326 | n3896 ;
  assign n6105 = n5118 | n6104 ;
  assign n6106 = ( ~n1723 & n5729 ) | ( ~n1723 & n6105 ) | ( n5729 & n6105 ) ;
  assign n6102 = n2259 ^ n415 ^ 1'b0 ;
  assign n6101 = n1939 & n4055 ;
  assign n6103 = n6102 ^ n6101 ^ 1'b0 ;
  assign n6107 = n6106 ^ n6103 ^ x134 ;
  assign n6108 = n371 & ~n4585 ;
  assign n6109 = n6108 ^ n4254 ^ 1'b0 ;
  assign n6110 = n1755 | n3426 ;
  assign n6111 = n4547 ^ x193 ^ 1'b0 ;
  assign n6116 = n1723 ^ n1179 ^ 1'b0 ;
  assign n6117 = n1666 & n6116 ;
  assign n6112 = n1240 & n1794 ;
  assign n6113 = n1760 | n4247 ;
  assign n6114 = n6112 | n6113 ;
  assign n6115 = n5057 & n6114 ;
  assign n6118 = n6117 ^ n6115 ^ 1'b0 ;
  assign n6119 = ~n2598 & n2737 ;
  assign n6120 = n5491 ^ n3363 ^ 1'b0 ;
  assign n6121 = n1666 & n6120 ;
  assign n6122 = n823 & n4812 ;
  assign n6123 = ~n6121 & n6122 ;
  assign n6124 = n1439 & n6123 ;
  assign n6125 = n2185 ^ n1423 ^ 1'b0 ;
  assign n6126 = n1958 ^ n631 ^ 1'b0 ;
  assign n6127 = n6125 | n6126 ;
  assign n6128 = n4029 ^ n1269 ^ 1'b0 ;
  assign n6129 = n3160 | n6128 ;
  assign n6130 = n4814 | n6129 ;
  assign n6131 = n6130 ^ n575 ^ 1'b0 ;
  assign n6132 = n6127 & n6131 ;
  assign n6133 = n4930 ^ n4350 ^ n2946 ;
  assign n6134 = n6133 ^ n4635 ^ n4514 ;
  assign n6135 = ( n5329 & n5922 ) | ( n5329 & n6134 ) | ( n5922 & n6134 ) ;
  assign n6136 = n2938 & ~n5914 ;
  assign n6137 = n6136 ^ n2429 ^ 1'b0 ;
  assign n6138 = n861 ^ n620 ^ 1'b0 ;
  assign n6139 = n6138 ^ n3027 ^ 1'b0 ;
  assign n6140 = n6137 & ~n6139 ;
  assign n6151 = ~n449 & n922 ;
  assign n6152 = n6151 ^ x245 ^ 1'b0 ;
  assign n6142 = x223 ^ x101 ^ 1'b0 ;
  assign n6143 = n914 & n6142 ;
  assign n6141 = n1727 ^ x148 ^ 1'b0 ;
  assign n6144 = n6143 ^ n6141 ^ 1'b0 ;
  assign n6145 = n2360 & ~n6144 ;
  assign n6146 = ~n3275 & n5593 ;
  assign n6147 = n6146 ^ n4176 ^ 1'b0 ;
  assign n6148 = n6147 ^ n5078 ^ 1'b0 ;
  assign n6149 = n6145 & n6148 ;
  assign n6150 = ~n1637 & n6149 ;
  assign n6153 = n6152 ^ n6150 ^ 1'b0 ;
  assign n6154 = n6001 ^ n2706 ^ 1'b0 ;
  assign n6155 = n1319 & ~n1533 ;
  assign n6156 = n6155 ^ n442 ^ 1'b0 ;
  assign n6157 = n1813 ^ n699 ^ 1'b0 ;
  assign n6158 = n6157 ^ n3157 ^ 1'b0 ;
  assign n6159 = n6156 | n6158 ;
  assign n6160 = ( n460 & n1593 ) | ( n460 & n3060 ) | ( n1593 & n3060 ) ;
  assign n6161 = n1616 | n6160 ;
  assign n6162 = n6161 ^ n3151 ^ 1'b0 ;
  assign n6163 = ~n1858 & n6162 ;
  assign n6164 = ~n1190 & n6163 ;
  assign n6169 = ~n1032 & n5089 ;
  assign n6170 = n6169 ^ n1307 ^ 1'b0 ;
  assign n6167 = n4944 ^ n1341 ^ 1'b0 ;
  assign n6165 = n3567 ^ n3222 ^ n2622 ;
  assign n6166 = x120 & ~n6165 ;
  assign n6168 = n6167 ^ n6166 ^ 1'b0 ;
  assign n6171 = n6170 ^ n6168 ^ 1'b0 ;
  assign n6172 = n3285 ^ n2055 ^ x216 ;
  assign n6173 = n2871 & n3315 ;
  assign n6174 = ~x61 & n6173 ;
  assign n6175 = ~n4995 & n6174 ;
  assign n6181 = n4029 ^ n1105 ^ 1'b0 ;
  assign n6182 = n4902 & ~n6181 ;
  assign n6180 = n4330 | n5298 ;
  assign n6183 = n6182 ^ n6180 ^ 1'b0 ;
  assign n6184 = ( ~n2233 & n4298 ) | ( ~n2233 & n6183 ) | ( n4298 & n6183 ) ;
  assign n6176 = ( ~n519 & n1727 ) | ( ~n519 & n3420 ) | ( n1727 & n3420 ) ;
  assign n6177 = n4957 ^ n3312 ^ n1249 ;
  assign n6178 = n6176 & n6177 ;
  assign n6179 = n6178 ^ n2888 ^ 1'b0 ;
  assign n6185 = n6184 ^ n6179 ^ x218 ;
  assign n6186 = x3 | n1851 ;
  assign n6187 = n382 ^ n341 ^ 1'b0 ;
  assign n6188 = n6186 & ~n6187 ;
  assign n6189 = n3002 ^ n2475 ^ 1'b0 ;
  assign n6190 = ( n256 & n6188 ) | ( n256 & n6189 ) | ( n6188 & n6189 ) ;
  assign n6194 = n2578 ^ n2311 ^ n1295 ;
  assign n6191 = x239 ^ x56 ^ 1'b0 ;
  assign n6192 = ( ~n713 & n2841 ) | ( ~n713 & n6191 ) | ( n2841 & n6191 ) ;
  assign n6193 = n1891 & ~n6192 ;
  assign n6195 = n6194 ^ n6193 ^ n3156 ;
  assign n6196 = n2619 ^ n1423 ^ n381 ;
  assign n6197 = n1173 & n6196 ;
  assign n6198 = ~n2644 & n6197 ;
  assign n6199 = n614 & ~n6198 ;
  assign n6200 = n6199 ^ n1350 ^ 1'b0 ;
  assign n6201 = n2329 | n6200 ;
  assign n6202 = n6201 ^ n2200 ^ 1'b0 ;
  assign n6203 = n4396 & n5999 ;
  assign n6204 = n6111 & n6203 ;
  assign n6205 = n5353 & ~n5775 ;
  assign n6206 = n3320 ^ n1965 ^ x250 ;
  assign n6207 = n5112 ^ n3729 ^ n3328 ;
  assign n6208 = n4101 ^ n1343 ^ 1'b0 ;
  assign n6209 = n6207 & n6208 ;
  assign n6210 = ~n6206 & n6209 ;
  assign n6211 = n6210 ^ n2155 ^ 1'b0 ;
  assign n6212 = n2574 | n6211 ;
  assign n6213 = n614 | n6212 ;
  assign n6214 = ~n268 & n1709 ;
  assign n6215 = n6214 ^ n3660 ^ 1'b0 ;
  assign n6216 = n3469 ^ n1285 ^ n1145 ;
  assign n6217 = ~n6215 & n6216 ;
  assign n6218 = n6217 ^ n4837 ^ 1'b0 ;
  assign n6219 = n4455 & ~n4550 ;
  assign n6220 = n6219 ^ n5265 ^ 1'b0 ;
  assign n6221 = n6066 | n6220 ;
  assign n6222 = n5123 ^ n4503 ^ 1'b0 ;
  assign n6223 = n3409 | n4311 ;
  assign n6224 = ~n829 & n4745 ;
  assign n6225 = ~n1838 & n6224 ;
  assign n6226 = n1629 & n2025 ;
  assign n6227 = n1772 & n6226 ;
  assign n6228 = n3935 ^ n3361 ^ 1'b0 ;
  assign n6229 = ( ~n829 & n2422 ) | ( ~n829 & n5318 ) | ( n2422 & n5318 ) ;
  assign n6230 = n6228 & ~n6229 ;
  assign n6231 = ~n2585 & n5593 ;
  assign n6232 = n3161 ^ n847 ^ 1'b0 ;
  assign n6233 = ~n3619 & n6232 ;
  assign n6234 = n3318 & n6233 ;
  assign n6235 = ~n1772 & n2236 ;
  assign n6236 = ~n1031 & n6235 ;
  assign n6237 = n6236 ^ n3517 ^ 1'b0 ;
  assign n6238 = n2968 | n6237 ;
  assign n6239 = n3502 & ~n6238 ;
  assign n6240 = n6075 ^ n2663 ^ 1'b0 ;
  assign n6241 = n5289 ^ n4502 ^ n3814 ;
  assign n6242 = ( n2760 & ~n6240 ) | ( n2760 & n6241 ) | ( ~n6240 & n6241 ) ;
  assign n6243 = n2957 ^ n2392 ^ n1789 ;
  assign n6244 = n6066 | n6243 ;
  assign n6245 = ( ~n428 & n704 ) | ( ~n428 & n2575 ) | ( n704 & n2575 ) ;
  assign n6246 = ~n5456 & n6245 ;
  assign n6247 = n2088 ^ x237 ^ 1'b0 ;
  assign n6248 = n5815 ^ n2397 ^ n1874 ;
  assign n6249 = n1820 | n6248 ;
  assign n6250 = n6249 ^ n4743 ^ n511 ;
  assign n6251 = n2447 ^ n603 ^ 1'b0 ;
  assign n6252 = n6250 & n6251 ;
  assign n6253 = ~n6247 & n6252 ;
  assign n6254 = n6246 & ~n6253 ;
  assign n6255 = n5388 ^ n2157 ^ n1716 ;
  assign n6256 = x179 | n775 ;
  assign n6257 = ( n3786 & n5042 ) | ( n3786 & n6256 ) | ( n5042 & n6256 ) ;
  assign n6258 = n1613 ^ n1361 ^ 1'b0 ;
  assign n6259 = n1316 | n6258 ;
  assign n6260 = n5368 ^ x74 ^ 1'b0 ;
  assign n6261 = ( n5812 & n6259 ) | ( n5812 & n6260 ) | ( n6259 & n6260 ) ;
  assign n6262 = n4132 & ~n4469 ;
  assign n6263 = n1435 ^ x121 ^ 1'b0 ;
  assign n6264 = x90 & ~n6263 ;
  assign n6265 = n3394 & n5119 ;
  assign n6266 = ~n6264 & n6265 ;
  assign n6267 = n6266 ^ n6133 ^ n3425 ;
  assign n6268 = n4768 ^ n3272 ^ 1'b0 ;
  assign n6269 = n6268 ^ n3619 ^ 1'b0 ;
  assign n6270 = n4619 ^ n2724 ^ 1'b0 ;
  assign n6271 = n1799 | n6270 ;
  assign n6272 = ~n6269 & n6271 ;
  assign n6274 = n2908 | n3373 ;
  assign n6275 = n6274 ^ n2045 ^ 1'b0 ;
  assign n6273 = n2397 & ~n3009 ;
  assign n6276 = n6275 ^ n6273 ^ 1'b0 ;
  assign n6277 = n2335 & ~n4805 ;
  assign n6278 = n6277 ^ n2995 ^ 1'b0 ;
  assign n6279 = n771 & ~n1024 ;
  assign n6280 = n3672 & n6279 ;
  assign n6281 = n6280 ^ n818 ^ 1'b0 ;
  assign n6282 = ~n6278 & n6281 ;
  assign n6283 = ~x185 & n3773 ;
  assign n6284 = n6283 ^ n5762 ^ 1'b0 ;
  assign n6286 = x28 & x99 ;
  assign n6287 = n6286 ^ n3317 ^ 1'b0 ;
  assign n6288 = n5761 ^ x9 ^ 1'b0 ;
  assign n6289 = n6287 & n6288 ;
  assign n6285 = n1401 | n6018 ;
  assign n6290 = n6289 ^ n6285 ^ 1'b0 ;
  assign n6291 = n5869 ^ x104 ^ 1'b0 ;
  assign n6292 = n4298 | n5865 ;
  assign n6293 = n2577 ^ n1994 ^ 1'b0 ;
  assign n6294 = n4020 ^ n1536 ^ 1'b0 ;
  assign n6295 = n6294 ^ x217 ^ 1'b0 ;
  assign n6296 = ( n4604 & n6293 ) | ( n4604 & ~n6295 ) | ( n6293 & ~n6295 ) ;
  assign n6297 = ( ~n2763 & n5486 ) | ( ~n2763 & n5618 ) | ( n5486 & n5618 ) ;
  assign n6298 = ~n1451 & n2105 ;
  assign n6299 = n4767 & n6298 ;
  assign n6300 = n6299 ^ x175 ^ 1'b0 ;
  assign n6306 = n5885 ^ n345 ^ 1'b0 ;
  assign n6301 = n1093 ^ n445 ^ 1'b0 ;
  assign n6302 = n1196 & ~n6301 ;
  assign n6303 = ~n966 & n6302 ;
  assign n6304 = n720 | n6303 ;
  assign n6305 = n4156 | n6304 ;
  assign n6307 = n6306 ^ n6305 ^ n4374 ;
  assign n6308 = n6228 ^ n5311 ^ 1'b0 ;
  assign n6309 = n1444 ^ n1103 ^ 1'b0 ;
  assign n6310 = n5577 | n6309 ;
  assign n6311 = n2847 | n3389 ;
  assign n6312 = n6310 & ~n6311 ;
  assign n6313 = n2255 | n6312 ;
  assign n6314 = n4240 & ~n4661 ;
  assign n6315 = n4004 & n5034 ;
  assign n6316 = n1739 | n3816 ;
  assign n6317 = n2572 ^ n2407 ^ 1'b0 ;
  assign n6318 = ~n6316 & n6317 ;
  assign n6319 = n1641 ^ n1457 ^ n883 ;
  assign n6320 = n5594 & ~n6319 ;
  assign n6321 = ~n1452 & n1978 ;
  assign n6322 = ~n808 & n6321 ;
  assign n6323 = n6322 ^ n4097 ^ 1'b0 ;
  assign n6324 = n6320 | n6323 ;
  assign n6325 = ( x121 & ~n847 ) | ( x121 & n3062 ) | ( ~n847 & n3062 ) ;
  assign n6326 = n759 & ~n1108 ;
  assign n6327 = x60 & ~n1189 ;
  assign n6328 = n6327 ^ n1802 ^ 1'b0 ;
  assign n6329 = n6328 ^ n2154 ^ n1115 ;
  assign n6330 = n6329 ^ n6170 ^ n3075 ;
  assign n6331 = n6326 & n6330 ;
  assign n6332 = n6331 ^ n841 ^ 1'b0 ;
  assign n6333 = n1234 & ~n6332 ;
  assign n6334 = ~n6325 & n6333 ;
  assign n6335 = n1048 ^ n678 ^ 1'b0 ;
  assign n6336 = n3093 ^ n2138 ^ 1'b0 ;
  assign n6337 = n3617 | n6336 ;
  assign n6338 = n4919 | n6337 ;
  assign n6344 = n3100 & n6086 ;
  assign n6339 = n5226 ^ n1420 ^ 1'b0 ;
  assign n6340 = ~n2154 & n6339 ;
  assign n6341 = n288 & n6340 ;
  assign n6342 = ( ~n535 & n1678 ) | ( ~n535 & n4327 ) | ( n1678 & n4327 ) ;
  assign n6343 = ~n6341 & n6342 ;
  assign n6345 = n6344 ^ n6343 ^ 1'b0 ;
  assign n6346 = n4569 & n5713 ;
  assign n6347 = n6345 & n6346 ;
  assign n6348 = x166 | n1733 ;
  assign n6349 = n4913 & ~n6348 ;
  assign n6350 = n4548 & n6349 ;
  assign n6351 = n2853 ^ x53 ^ 1'b0 ;
  assign n6352 = n2275 & n6351 ;
  assign n6353 = n6352 ^ n4492 ^ n1019 ;
  assign n6354 = n1951 ^ n1409 ^ 1'b0 ;
  assign n6355 = n2608 & ~n6354 ;
  assign n6356 = ~n1874 & n4697 ;
  assign n6357 = n2504 & n5606 ;
  assign n6358 = n4741 ^ n3219 ^ 1'b0 ;
  assign n6360 = n3169 ^ n1970 ^ 1'b0 ;
  assign n6361 = n5166 & ~n6360 ;
  assign n6359 = n2248 | n3052 ;
  assign n6362 = n6361 ^ n6359 ^ 1'b0 ;
  assign n6363 = ( n271 & n500 ) | ( n271 & n2164 ) | ( n500 & n2164 ) ;
  assign n6364 = n6363 ^ n1519 ^ n413 ;
  assign n6365 = n6364 ^ n2750 ^ 1'b0 ;
  assign n6366 = n1438 ^ n617 ^ 1'b0 ;
  assign n6367 = n6365 & ~n6366 ;
  assign n6371 = n1944 ^ n835 ^ 1'b0 ;
  assign n6372 = n6371 ^ n1018 ^ 1'b0 ;
  assign n6373 = ~n1912 & n6372 ;
  assign n6368 = n2340 ^ n1644 ^ n1554 ;
  assign n6369 = ~n3497 & n6368 ;
  assign n6370 = n6369 ^ n947 ^ 1'b0 ;
  assign n6374 = n6373 ^ n6370 ^ n5172 ;
  assign n6375 = n4639 ^ n2024 ^ 1'b0 ;
  assign n6376 = n6375 ^ n673 ^ x95 ;
  assign n6377 = n6376 ^ n1094 ^ 1'b0 ;
  assign n6378 = n4098 & ~n6377 ;
  assign n6379 = n6378 ^ n4499 ^ 1'b0 ;
  assign n6380 = n1569 & ~n1746 ;
  assign n6381 = ~n1496 & n6380 ;
  assign n6382 = n6257 ^ n1564 ^ 1'b0 ;
  assign n6383 = ~n1607 & n6382 ;
  assign n6384 = n6381 & n6383 ;
  assign n6385 = n1576 & n3494 ;
  assign n6386 = n6028 ^ n1888 ^ x29 ;
  assign n6388 = n573 & ~n2057 ;
  assign n6389 = n4369 & n6388 ;
  assign n6387 = n1579 ^ n775 ^ 1'b0 ;
  assign n6390 = n6389 ^ n6387 ^ 1'b0 ;
  assign n6391 = x213 & n5596 ;
  assign n6392 = n6123 & n6391 ;
  assign n6393 = ( x200 & n2523 ) | ( x200 & n6191 ) | ( n2523 & n6191 ) ;
  assign n6394 = n6393 ^ n3894 ^ 1'b0 ;
  assign n6395 = n1067 & n2993 ;
  assign n6400 = x59 & ~n405 ;
  assign n6396 = n2191 ^ n1552 ^ x177 ;
  assign n6397 = ~n1689 & n4088 ;
  assign n6398 = ~n6396 & n6397 ;
  assign n6399 = ( x82 & n3644 ) | ( x82 & ~n6398 ) | ( n3644 & ~n6398 ) ;
  assign n6401 = n6400 ^ n6399 ^ 1'b0 ;
  assign n6402 = ~n3070 & n6401 ;
  assign n6403 = n316 | n763 ;
  assign n6404 = n1713 & n6403 ;
  assign n6405 = ~n5275 & n6404 ;
  assign n6406 = n6405 ^ n5706 ^ 1'b0 ;
  assign n6407 = ( n1891 & n2570 ) | ( n1891 & ~n5103 ) | ( n2570 & ~n5103 ) ;
  assign n6408 = n6407 ^ x181 ^ 1'b0 ;
  assign n6409 = n6408 ^ n6312 ^ 1'b0 ;
  assign n6410 = n1425 | n6409 ;
  assign n6411 = n5636 ^ n1844 ^ 1'b0 ;
  assign n6412 = n6411 ^ n2338 ^ 1'b0 ;
  assign n6413 = x64 & n6412 ;
  assign n6414 = n368 & n6413 ;
  assign n6415 = n4296 ^ n3329 ^ 1'b0 ;
  assign n6416 = n5500 ^ n2299 ^ 1'b0 ;
  assign n6417 = ~n6415 & n6416 ;
  assign n6418 = n271 & n3502 ;
  assign n6419 = n738 ^ x62 ^ 1'b0 ;
  assign n6420 = x94 & n6419 ;
  assign n6421 = n1216 | n2137 ;
  assign n6422 = n561 & ~n6421 ;
  assign n6423 = n6420 & ~n6422 ;
  assign n6424 = ~n6418 & n6423 ;
  assign n6435 = ( n413 & n1650 ) | ( n413 & ~n2142 ) | ( n1650 & ~n2142 ) ;
  assign n6436 = n6435 ^ n3138 ^ 1'b0 ;
  assign n6433 = n2208 & ~n5275 ;
  assign n6434 = n6433 ^ n3147 ^ n1222 ;
  assign n6430 = n516 ^ x217 ^ 1'b0 ;
  assign n6431 = n6430 ^ n5344 ^ 1'b0 ;
  assign n6425 = x98 | n305 ;
  assign n6426 = n2804 ^ n343 ^ 1'b0 ;
  assign n6427 = ~n478 & n6426 ;
  assign n6428 = ( n2248 & n6425 ) | ( n2248 & n6427 ) | ( n6425 & n6427 ) ;
  assign n6429 = n2685 | n6428 ;
  assign n6432 = n6431 ^ n6429 ^ 1'b0 ;
  assign n6437 = n6436 ^ n6434 ^ n6432 ;
  assign n6438 = n5854 ^ n1351 ^ 1'b0 ;
  assign n6439 = n1829 & n1843 ;
  assign n6440 = n870 & ~n5275 ;
  assign n6441 = n850 & n6440 ;
  assign n6442 = n639 ^ n499 ^ n417 ;
  assign n6443 = n6441 | n6442 ;
  assign n6444 = n4557 | n6443 ;
  assign n6445 = ( n2636 & n6439 ) | ( n2636 & n6444 ) | ( n6439 & n6444 ) ;
  assign n6446 = n6109 ^ n773 ^ 1'b0 ;
  assign n6447 = n2548 & ~n5198 ;
  assign n6455 = n1270 & ~n2085 ;
  assign n6456 = n6455 ^ n1476 ^ 1'b0 ;
  assign n6450 = n3366 ^ n1773 ^ 1'b0 ;
  assign n6451 = n2991 ^ n1016 ^ 1'b0 ;
  assign n6452 = n6450 & n6451 ;
  assign n6453 = ( ~n1880 & n2824 ) | ( ~n1880 & n4906 ) | ( n2824 & n4906 ) ;
  assign n6454 = n6452 & n6453 ;
  assign n6457 = n6456 ^ n6454 ^ 1'b0 ;
  assign n6448 = n6024 ^ n3659 ^ n823 ;
  assign n6449 = ~n576 & n6448 ;
  assign n6458 = n6457 ^ n6449 ^ n4944 ;
  assign n6459 = n1383 | n3931 ;
  assign n6460 = n3322 & n6096 ;
  assign n6461 = n4391 & n6460 ;
  assign n6462 = n1208 ^ n621 ^ x241 ;
  assign n6463 = n402 ^ x184 ^ 1'b0 ;
  assign n6464 = n1727 & ~n6463 ;
  assign n6465 = n6464 ^ n1932 ^ 1'b0 ;
  assign n6466 = n4004 & ~n6465 ;
  assign n6467 = n6462 & n6466 ;
  assign n6468 = ( n2261 & n6461 ) | ( n2261 & ~n6467 ) | ( n6461 & ~n6467 ) ;
  assign n6473 = n6030 ^ n5160 ^ n1043 ;
  assign n6469 = ( n1765 & n3439 ) | ( n1765 & ~n4132 ) | ( n3439 & ~n4132 ) ;
  assign n6470 = n4985 ^ n2275 ^ 1'b0 ;
  assign n6471 = n2358 & ~n6470 ;
  assign n6472 = n6469 | n6471 ;
  assign n6474 = n6473 ^ n6472 ^ n1405 ;
  assign n6475 = n4879 | n5875 ;
  assign n6476 = n1341 | n6475 ;
  assign n6477 = ( n2680 & n3172 ) | ( n2680 & ~n3488 ) | ( n3172 & ~n3488 ) ;
  assign n6478 = ~x117 & n5361 ;
  assign n6479 = ( ~n4170 & n5325 ) | ( ~n4170 & n6478 ) | ( n5325 & n6478 ) ;
  assign n6480 = n4485 | n6479 ;
  assign n6482 = n4874 ^ n3080 ^ 1'b0 ;
  assign n6483 = n752 & ~n6482 ;
  assign n6484 = n6483 ^ n5088 ^ n1494 ;
  assign n6481 = n2922 & n5486 ;
  assign n6485 = n6484 ^ n6481 ^ 1'b0 ;
  assign n6486 = ( x192 & ~n514 ) | ( x192 & n4249 ) | ( ~n514 & n4249 ) ;
  assign n6487 = n661 & n888 ;
  assign n6488 = n5298 & n6487 ;
  assign n6489 = ( n3264 & n4223 ) | ( n3264 & n6488 ) | ( n4223 & n6488 ) ;
  assign n6490 = n1312 & ~n1869 ;
  assign n6491 = n6490 ^ n3107 ^ 1'b0 ;
  assign n6492 = n866 & n2676 ;
  assign n6493 = n6492 ^ n6368 ^ 1'b0 ;
  assign n6494 = n926 & ~n3704 ;
  assign n6495 = n6493 | n6494 ;
  assign n6496 = n6495 ^ n876 ^ 1'b0 ;
  assign n6497 = n6496 ^ n4149 ^ 1'b0 ;
  assign n6498 = x150 ^ x92 ^ 1'b0 ;
  assign n6499 = ( n387 & ~n1729 ) | ( n387 & n4371 ) | ( ~n1729 & n4371 ) ;
  assign n6500 = n2275 | n6499 ;
  assign n6501 = n6498 & ~n6500 ;
  assign n6502 = ( n2409 & n4617 ) | ( n2409 & ~n6501 ) | ( n4617 & ~n6501 ) ;
  assign n6503 = ~n3289 & n4902 ;
  assign n6504 = n1107 & n6503 ;
  assign n6505 = n3335 ^ n3237 ^ 1'b0 ;
  assign n6506 = n4630 ^ n2026 ^ 1'b0 ;
  assign n6507 = ( n3146 & ~n6505 ) | ( n3146 & n6506 ) | ( ~n6505 & n6506 ) ;
  assign n6508 = n3961 | n6036 ;
  assign n6509 = n2015 | n6508 ;
  assign n6510 = n4559 ^ n2155 ^ x43 ;
  assign n6511 = ( n3510 & n5928 ) | ( n3510 & n6510 ) | ( n5928 & n6510 ) ;
  assign n6512 = n6511 ^ n5722 ^ n5681 ;
  assign n6513 = n1524 & ~n1527 ;
  assign n6514 = n6513 ^ n405 ^ 1'b0 ;
  assign n6515 = n6514 ^ n2178 ^ n1462 ;
  assign n6516 = n6515 ^ n2929 ^ 1'b0 ;
  assign n6517 = n1410 ^ x52 ^ x12 ;
  assign n6518 = n2280 ^ n1308 ^ 1'b0 ;
  assign n6519 = n2577 | n6518 ;
  assign n6520 = ( ~n2172 & n6517 ) | ( ~n2172 & n6519 ) | ( n6517 & n6519 ) ;
  assign n6521 = n3898 & n5143 ;
  assign n6522 = n6521 ^ n2878 ^ 1'b0 ;
  assign n6523 = ( ~x109 & n273 ) | ( ~x109 & n2824 ) | ( n273 & n2824 ) ;
  assign n6524 = n6523 ^ n5723 ^ n4532 ;
  assign n6525 = n6522 | n6524 ;
  assign n6526 = n4202 & ~n6525 ;
  assign n6527 = ( n1871 & ~n5006 ) | ( n1871 & n5761 ) | ( ~n5006 & n5761 ) ;
  assign n6528 = ( n1211 & n1496 ) | ( n1211 & n2290 ) | ( n1496 & n2290 ) ;
  assign n6529 = n3967 | n6528 ;
  assign n6530 = n5464 | n6529 ;
  assign n6531 = ~x4 & n6530 ;
  assign n6532 = n5748 ^ n3409 ^ n3093 ;
  assign n6533 = ( n3345 & n3604 ) | ( n3345 & ~n6532 ) | ( n3604 & ~n6532 ) ;
  assign n6534 = n3585 ^ n1084 ^ 1'b0 ;
  assign n6535 = n1129 | n6534 ;
  assign n6536 = n6535 ^ n5445 ^ 1'b0 ;
  assign n6537 = n631 & n877 ;
  assign n6538 = ( n316 & n5992 ) | ( n316 & ~n6537 ) | ( n5992 & ~n6537 ) ;
  assign n6545 = ( n1630 & n1846 ) | ( n1630 & n4777 ) | ( n1846 & n4777 ) ;
  assign n6546 = n6545 ^ n5057 ^ n3717 ;
  assign n6540 = n3909 ^ n1168 ^ 1'b0 ;
  assign n6541 = n659 & ~n6540 ;
  assign n6542 = n6541 ^ n6396 ^ 1'b0 ;
  assign n6539 = ~n2214 & n2915 ;
  assign n6543 = n6542 ^ n6539 ^ 1'b0 ;
  assign n6544 = n3408 & n6543 ;
  assign n6547 = n6546 ^ n6544 ^ 1'b0 ;
  assign n6548 = n5223 & n5819 ;
  assign n6549 = n6548 ^ n2711 ^ 1'b0 ;
  assign n6550 = n4751 ^ n2669 ^ 1'b0 ;
  assign n6551 = n1847 & ~n6550 ;
  assign n6552 = ( ~n259 & n769 ) | ( ~n259 & n1108 ) | ( n769 & n1108 ) ;
  assign n6553 = x88 & ~n750 ;
  assign n6554 = n644 & n6553 ;
  assign n6555 = ( x196 & n322 ) | ( x196 & ~n2429 ) | ( n322 & ~n2429 ) ;
  assign n6556 = n6555 ^ n1126 ^ 1'b0 ;
  assign n6557 = n4604 ^ n1671 ^ x236 ;
  assign n6558 = ~n6556 & n6557 ;
  assign n6559 = ( n332 & ~n5148 ) | ( n332 & n6558 ) | ( ~n5148 & n6558 ) ;
  assign n6560 = ( n2128 & n4154 ) | ( n2128 & n6559 ) | ( n4154 & n6559 ) ;
  assign n6561 = ~n943 & n6560 ;
  assign n6562 = n6554 & n6561 ;
  assign n6563 = n6552 & n6562 ;
  assign n6564 = ~n5842 & n6563 ;
  assign n6565 = n6564 ^ n4815 ^ 1'b0 ;
  assign n6566 = n1584 & n3389 ;
  assign n6567 = n6566 ^ n6400 ^ 1'b0 ;
  assign n6568 = n4398 ^ n1343 ^ 1'b0 ;
  assign n6569 = n6135 ^ n5259 ^ n1727 ;
  assign n6578 = n2437 ^ x211 ^ 1'b0 ;
  assign n6579 = n4575 & ~n6578 ;
  assign n6580 = n4543 & n6579 ;
  assign n6570 = ~n2280 & n3065 ;
  assign n6571 = n6570 ^ n338 ^ 1'b0 ;
  assign n6572 = n6571 ^ n2078 ^ 1'b0 ;
  assign n6573 = n3268 | n6572 ;
  assign n6574 = n679 ^ n476 ^ 1'b0 ;
  assign n6575 = n2088 ^ n887 ^ 1'b0 ;
  assign n6576 = ~n6574 & n6575 ;
  assign n6577 = ~n6573 & n6576 ;
  assign n6581 = n6580 ^ n6577 ^ 1'b0 ;
  assign n6582 = n505 & ~n2409 ;
  assign n6583 = n2538 & n6582 ;
  assign n6584 = n3433 & ~n6583 ;
  assign n6585 = n6584 ^ n4330 ^ 1'b0 ;
  assign n6586 = n2208 & n6585 ;
  assign n6587 = n1980 & n6586 ;
  assign n6588 = ~n2780 & n3991 ;
  assign n6589 = n4592 ^ n3147 ^ n2907 ;
  assign n6590 = n4333 ^ n2920 ^ 1'b0 ;
  assign n6591 = ~n3125 & n6590 ;
  assign n6592 = n5942 ^ n4427 ^ n1979 ;
  assign n6593 = n5751 ^ n5646 ^ 1'b0 ;
  assign n6594 = ~n4227 & n6593 ;
  assign n6595 = n1037 | n2437 ;
  assign n6596 = n4029 & ~n6595 ;
  assign n6597 = n5357 ^ n718 ^ 1'b0 ;
  assign n6598 = n6596 | n6597 ;
  assign n6599 = n6598 ^ n2106 ^ 1'b0 ;
  assign n6601 = n3418 ^ n2974 ^ n520 ;
  assign n6600 = n2904 & ~n4692 ;
  assign n6602 = n6601 ^ n6600 ^ 1'b0 ;
  assign n6603 = x26 & n2842 ;
  assign n6604 = n3786 & n6603 ;
  assign n6605 = ~x2 & n6604 ;
  assign n6606 = x73 & n6605 ;
  assign n6607 = n5660 ^ n5567 ^ 1'b0 ;
  assign n6608 = ( ~n872 & n3802 ) | ( ~n872 & n4878 ) | ( n3802 & n4878 ) ;
  assign n6609 = ~n1000 & n4251 ;
  assign n6610 = n4678 ^ x222 ^ 1'b0 ;
  assign n6611 = n4100 ^ n3277 ^ n303 ;
  assign n6612 = n2690 ^ n365 ^ x69 ;
  assign n6613 = ( n2157 & n4197 ) | ( n2157 & n6612 ) | ( n4197 & n6612 ) ;
  assign n6614 = x107 & n6050 ;
  assign n6615 = ~n6613 & n6614 ;
  assign n6616 = ( ~n982 & n6611 ) | ( ~n982 & n6615 ) | ( n6611 & n6615 ) ;
  assign n6617 = n6610 | n6616 ;
  assign n6618 = n789 | n6617 ;
  assign n6619 = n2582 ^ n1024 ^ 1'b0 ;
  assign n6620 = ( ~n567 & n1158 ) | ( ~n567 & n6619 ) | ( n1158 & n6619 ) ;
  assign n6621 = n6620 ^ n3075 ^ n1521 ;
  assign n6623 = n2196 ^ n358 ^ 1'b0 ;
  assign n6622 = n957 & ~n4114 ;
  assign n6624 = n6623 ^ n6622 ^ 1'b0 ;
  assign n6626 = n5439 ^ n263 ^ 1'b0 ;
  assign n6627 = n6626 ^ n6075 ^ 1'b0 ;
  assign n6625 = x24 & n868 ;
  assign n6628 = n6627 ^ n6625 ^ 1'b0 ;
  assign n6629 = ~n3677 & n3786 ;
  assign n6630 = ~n684 & n5085 ;
  assign n6631 = ~n1270 & n6630 ;
  assign n6632 = n6631 ^ x117 ^ 1'b0 ;
  assign n6641 = x190 & ~n268 ;
  assign n6642 = n6641 ^ n3030 ^ 1'b0 ;
  assign n6633 = n449 ^ x173 ^ 1'b0 ;
  assign n6634 = n2310 & ~n6633 ;
  assign n6635 = x162 & ~n4729 ;
  assign n6636 = n6635 ^ n1713 ^ 1'b0 ;
  assign n6637 = n6328 | n6636 ;
  assign n6638 = n3896 & ~n6637 ;
  assign n6639 = n6634 & ~n6638 ;
  assign n6640 = n6639 ^ n2152 ^ 1'b0 ;
  assign n6643 = n6642 ^ n6640 ^ n2722 ;
  assign n6644 = n3456 | n6462 ;
  assign n6645 = ( ~n2116 & n4954 ) | ( ~n2116 & n6644 ) | ( n4954 & n6644 ) ;
  assign n6646 = n3928 ^ n3069 ^ n2524 ;
  assign n6647 = n1529 ^ n853 ^ 1'b0 ;
  assign n6648 = n4730 & ~n6647 ;
  assign n6649 = ~n6646 & n6648 ;
  assign n6650 = ~x46 & n2875 ;
  assign n6651 = n360 & n4995 ;
  assign n6652 = n6650 & n6651 ;
  assign n6653 = n6652 ^ n922 ^ 1'b0 ;
  assign n6654 = n6653 ^ n5544 ^ n4039 ;
  assign n6655 = n6649 | n6654 ;
  assign n6656 = n4367 | n6655 ;
  assign n6659 = n1244 ^ x150 ^ 1'b0 ;
  assign n6660 = n1999 & n6659 ;
  assign n6657 = ~n820 & n6105 ;
  assign n6658 = n6657 ^ n5513 ^ 1'b0 ;
  assign n6661 = n6660 ^ n6658 ^ n6501 ;
  assign n6662 = n3610 ^ n1012 ^ 1'b0 ;
  assign n6667 = ( ~n1975 & n2991 ) | ( ~n1975 & n4207 ) | ( n2991 & n4207 ) ;
  assign n6668 = n6667 ^ n4941 ^ 1'b0 ;
  assign n6663 = n3394 & n5221 ;
  assign n6664 = n1069 | n2178 ;
  assign n6665 = n459 | n6664 ;
  assign n6666 = n6663 & n6665 ;
  assign n6669 = n6668 ^ n6666 ^ 1'b0 ;
  assign n6670 = ( x86 & ~x178 ) | ( x86 & n1765 ) | ( ~x178 & n1765 ) ;
  assign n6671 = n2893 | n4282 ;
  assign n6672 = n6671 ^ n4588 ^ 1'b0 ;
  assign n6673 = n6672 ^ n468 ^ 1'b0 ;
  assign n6674 = n1324 & n6634 ;
  assign n6675 = ~n3721 & n6674 ;
  assign n6676 = n2889 & ~n4068 ;
  assign n6677 = ~n5303 & n6676 ;
  assign n6678 = n5880 & ~n6677 ;
  assign n6679 = n1806 ^ x105 ^ 1'b0 ;
  assign n6680 = n6679 ^ n1002 ^ 1'b0 ;
  assign n6681 = n4559 & n6680 ;
  assign n6682 = n3755 ^ n2200 ^ n2183 ;
  assign n6683 = n4945 & ~n6682 ;
  assign n6684 = n5042 ^ n2335 ^ x229 ;
  assign n6691 = ( n323 & n853 ) | ( n323 & n1252 ) | ( n853 & n1252 ) ;
  assign n6685 = n1802 ^ x76 ^ x7 ;
  assign n6686 = n2557 | n6152 ;
  assign n6687 = n6686 ^ n2355 ^ 1'b0 ;
  assign n6688 = n3370 & n6687 ;
  assign n6689 = n6688 ^ n3662 ^ n2595 ;
  assign n6690 = n6685 | n6689 ;
  assign n6692 = n6691 ^ n6690 ^ 1'b0 ;
  assign n6693 = n3049 & n6325 ;
  assign n6694 = ~x217 & n2378 ;
  assign n6695 = n3724 & n6694 ;
  assign n6696 = n6693 & n6695 ;
  assign n6697 = n6696 ^ n1452 ^ 1'b0 ;
  assign n6698 = n1220 ^ n943 ^ 1'b0 ;
  assign n6699 = n3075 ^ n424 ^ 1'b0 ;
  assign n6700 = n6699 ^ n2636 ^ 1'b0 ;
  assign n6701 = ~n4921 & n6700 ;
  assign n6702 = ~n6073 & n6660 ;
  assign n6703 = n6702 ^ n4254 ^ 1'b0 ;
  assign n6704 = n1970 & n3099 ;
  assign n6705 = n6704 ^ x198 ^ 1'b0 ;
  assign n6706 = ~n2165 & n6705 ;
  assign n6707 = n6706 ^ n1080 ^ 1'b0 ;
  assign n6708 = ~n5094 & n6707 ;
  assign n6709 = n1821 & n2146 ;
  assign n6710 = n6709 ^ n6031 ^ 1'b0 ;
  assign n6711 = ( n574 & n741 ) | ( n574 & ~n3369 ) | ( n741 & ~n3369 ) ;
  assign n6712 = n6711 ^ n4292 ^ 1'b0 ;
  assign n6713 = ~n3255 & n6712 ;
  assign n6714 = n6713 ^ n2251 ^ 1'b0 ;
  assign n6715 = n4269 & ~n6714 ;
  assign n6716 = n1538 & ~n1906 ;
  assign n6717 = n3724 ^ n2032 ^ x170 ;
  assign n6718 = x87 & ~n6717 ;
  assign n6719 = n1773 ^ n1107 ^ 1'b0 ;
  assign n6720 = ~n1514 & n3081 ;
  assign n6721 = n4084 & n6720 ;
  assign n6722 = n2113 & n2426 ;
  assign n6723 = n3943 ^ n2680 ^ n1155 ;
  assign n6724 = n6723 ^ n3158 ^ 1'b0 ;
  assign n6725 = n1497 ^ n1479 ^ x151 ;
  assign n6726 = ~n4861 & n6725 ;
  assign n6727 = n6726 ^ n1597 ^ 1'b0 ;
  assign n6728 = ( n1258 & ~n5193 ) | ( n1258 & n6727 ) | ( ~n5193 & n6727 ) ;
  assign n6729 = n6728 ^ x70 ^ 1'b0 ;
  assign n6730 = n6724 & ~n6729 ;
  assign n6731 = n425 & n6444 ;
  assign n6732 = n6731 ^ n1063 ^ 1'b0 ;
  assign n6733 = n3409 ^ n1496 ^ 1'b0 ;
  assign n6734 = n3553 | n6733 ;
  assign n6735 = n6734 ^ n5444 ^ n1586 ;
  assign n6736 = n3683 | n6735 ;
  assign n6737 = n3596 & ~n6736 ;
  assign n6738 = ~n1804 & n3373 ;
  assign n6739 = n6738 ^ x178 ^ 1'b0 ;
  assign n6740 = n6739 ^ n2120 ^ n1691 ;
  assign n6741 = n5760 ^ n3260 ^ 1'b0 ;
  assign n6742 = ~n5952 & n6741 ;
  assign n6743 = n3036 ^ n692 ^ 1'b0 ;
  assign n6744 = n968 & ~n6743 ;
  assign n6745 = n3510 ^ n1162 ^ n703 ;
  assign n6746 = n1133 ^ n973 ^ 1'b0 ;
  assign n6747 = ~n6018 & n6746 ;
  assign n6748 = ( n4754 & ~n6745 ) | ( n4754 & n6747 ) | ( ~n6745 & n6747 ) ;
  assign n6749 = n5800 ^ n1545 ^ 1'b0 ;
  assign n6750 = n6749 ^ n4857 ^ n4046 ;
  assign n6751 = n4653 & n6430 ;
  assign n6752 = n6751 ^ x24 ^ 1'b0 ;
  assign n6753 = n3049 & n6752 ;
  assign n6758 = ~n454 & n2734 ;
  assign n6754 = ( n887 & n2555 ) | ( n887 & ~n3078 ) | ( n2555 & ~n3078 ) ;
  assign n6755 = ~n6652 & n6754 ;
  assign n6756 = ~n2496 & n6755 ;
  assign n6757 = n6756 ^ n5878 ^ n1698 ;
  assign n6759 = n6758 ^ n6757 ^ 1'b0 ;
  assign n6760 = n2264 & n5394 ;
  assign n6761 = n3007 & n6760 ;
  assign n6762 = n2703 | n4662 ;
  assign n6763 = n6762 ^ n3516 ^ 1'b0 ;
  assign n6770 = n462 & n2257 ;
  assign n6764 = n2744 ^ n951 ^ x20 ;
  assign n6765 = n1194 ^ x28 ^ 1'b0 ;
  assign n6766 = n6545 ^ n3629 ^ 1'b0 ;
  assign n6767 = n6765 & n6766 ;
  assign n6768 = ~n6764 & n6767 ;
  assign n6769 = n6768 ^ n1079 ^ 1'b0 ;
  assign n6771 = n6770 ^ n6769 ^ n3349 ;
  assign n6772 = ( ~x66 & n3398 ) | ( ~x66 & n6771 ) | ( n3398 & n6771 ) ;
  assign n6773 = ~x129 & n6308 ;
  assign n6774 = n745 ^ x208 ^ 1'b0 ;
  assign n6775 = n371 & ~n2159 ;
  assign n6776 = ~n1632 & n6775 ;
  assign n6777 = ( n307 & n1657 ) | ( n307 & ~n1750 ) | ( n1657 & ~n1750 ) ;
  assign n6778 = n6777 ^ n3945 ^ n845 ;
  assign n6779 = ~n3288 & n6778 ;
  assign n6780 = n4797 & ~n6779 ;
  assign n6781 = ~n6776 & n6780 ;
  assign n6782 = ~n3432 & n5667 ;
  assign n6787 = n1349 & n3316 ;
  assign n6788 = ~x223 & n6787 ;
  assign n6783 = x242 | n1562 ;
  assign n6784 = ~n1251 & n6783 ;
  assign n6785 = n5274 & n6784 ;
  assign n6786 = n6785 ^ n1019 ^ 1'b0 ;
  assign n6789 = n6788 ^ n6786 ^ n895 ;
  assign n6790 = n715 & n1472 ;
  assign n6791 = ~x153 & n6790 ;
  assign n6792 = n5386 ^ n4528 ^ n748 ;
  assign n6793 = n6792 ^ n1076 ^ n519 ;
  assign n6794 = n6791 & n6793 ;
  assign n6795 = n2970 | n6032 ;
  assign n6796 = n6795 ^ n2728 ^ 1'b0 ;
  assign n6797 = n6796 ^ n5967 ^ x248 ;
  assign n6798 = ~n4499 & n6797 ;
  assign n6799 = ~n3039 & n6798 ;
  assign n6800 = n5667 & ~n5865 ;
  assign n6801 = ~n264 & n3488 ;
  assign n6802 = ~n6800 & n6801 ;
  assign n6804 = n2247 | n3309 ;
  assign n6803 = ~n1068 & n1322 ;
  assign n6805 = n6804 ^ n6803 ^ 1'b0 ;
  assign n6806 = n6783 ^ n1453 ^ 1'b0 ;
  assign n6807 = ~n4675 & n6806 ;
  assign n6810 = n1067 & n3100 ;
  assign n6808 = n1647 ^ x215 ^ 1'b0 ;
  assign n6809 = ~n2592 & n6808 ;
  assign n6811 = n6810 ^ n6809 ^ 1'b0 ;
  assign n6812 = ( x118 & n1593 ) | ( x118 & n1607 ) | ( n1593 & n1607 ) ;
  assign n6813 = n557 ^ x108 ^ 1'b0 ;
  assign n6814 = n2563 & ~n6813 ;
  assign n6815 = n6812 | n6814 ;
  assign n6816 = n3986 ^ n3273 ^ 1'b0 ;
  assign n6819 = n4120 & n4789 ;
  assign n6820 = n6819 ^ n2507 ^ 1'b0 ;
  assign n6817 = n1995 & n4173 ;
  assign n6818 = ~n2553 & n6817 ;
  assign n6821 = n6820 ^ n6818 ^ 1'b0 ;
  assign n6826 = n1944 ^ n1906 ^ n1828 ;
  assign n6823 = n1209 ^ n1138 ^ 1'b0 ;
  assign n6824 = ~n900 & n6823 ;
  assign n6825 = ~n2504 & n6824 ;
  assign n6827 = n6826 ^ n6825 ^ 1'b0 ;
  assign n6822 = n3369 ^ n702 ^ 1'b0 ;
  assign n6828 = n6827 ^ n6822 ^ n6677 ;
  assign n6829 = ( n1067 & ~n5761 ) | ( n1067 & n6828 ) | ( ~n5761 & n6828 ) ;
  assign n6830 = n1100 ^ n442 ^ 1'b0 ;
  assign n6831 = x243 & ~n6830 ;
  assign n6832 = n6831 ^ n637 ^ 1'b0 ;
  assign n6841 = n5837 ^ n2506 ^ 1'b0 ;
  assign n6833 = n499 | n1523 ;
  assign n6836 = n6727 ^ n5341 ^ 1'b0 ;
  assign n6834 = n2475 & n6560 ;
  assign n6835 = n6834 ^ n3557 ^ 1'b0 ;
  assign n6837 = n6836 ^ n6835 ^ 1'b0 ;
  assign n6838 = n5993 | n6837 ;
  assign n6839 = n6838 ^ x222 ^ 1'b0 ;
  assign n6840 = n6833 & n6839 ;
  assign n6842 = n6841 ^ n6840 ^ 1'b0 ;
  assign n6843 = n5522 ^ n5021 ^ n4052 ;
  assign n6844 = n347 & ~n1401 ;
  assign n6845 = n6844 ^ n1955 ^ 1'b0 ;
  assign n6846 = n6845 ^ n4768 ^ n854 ;
  assign n6847 = ~n5810 & n6846 ;
  assign n6848 = ~x24 & n475 ;
  assign n6849 = n3708 ^ n853 ^ 1'b0 ;
  assign n6850 = ~n5417 & n6849 ;
  assign n6851 = ( ~x83 & n6848 ) | ( ~x83 & n6850 ) | ( n6848 & n6850 ) ;
  assign n6852 = n6851 ^ n3389 ^ 1'b0 ;
  assign n6853 = n3247 & ~n6852 ;
  assign n6854 = ( n2968 & ~n3123 ) | ( n2968 & n6853 ) | ( ~n3123 & n6853 ) ;
  assign n6855 = ( n816 & n6847 ) | ( n816 & ~n6854 ) | ( n6847 & ~n6854 ) ;
  assign n6856 = n6452 ^ n4790 ^ n1164 ;
  assign n6857 = n3042 | n3949 ;
  assign n6858 = ( n1079 & ~n3654 ) | ( n1079 & n6857 ) | ( ~n3654 & n6857 ) ;
  assign n6859 = n4788 ^ n1236 ^ 1'b0 ;
  assign n6860 = n4991 | n6859 ;
  assign n6863 = n1881 ^ n363 ^ x147 ;
  assign n6864 = n3690 ^ n2154 ^ 1'b0 ;
  assign n6865 = n1495 & ~n6864 ;
  assign n6866 = ( n1128 & ~n6863 ) | ( n1128 & n6865 ) | ( ~n6863 & n6865 ) ;
  assign n6867 = n6866 ^ n4242 ^ n3406 ;
  assign n6861 = ( ~n735 & n1633 ) | ( ~n735 & n6688 ) | ( n1633 & n6688 ) ;
  assign n6862 = n1511 & ~n6861 ;
  assign n6868 = n6867 ^ n6862 ^ 1'b0 ;
  assign n6869 = n844 & ~n6868 ;
  assign n6870 = ( n716 & n2131 ) | ( n716 & ~n6869 ) | ( n2131 & ~n6869 ) ;
  assign n6871 = x73 & ~n3248 ;
  assign n6872 = n6871 ^ n3268 ^ 1'b0 ;
  assign n6873 = n737 | n1944 ;
  assign n6874 = n6872 | n6873 ;
  assign n6875 = n2462 | n5112 ;
  assign n6876 = n5582 ^ n1060 ^ 1'b0 ;
  assign n6877 = n5317 ^ n1120 ^ 1'b0 ;
  assign n6878 = ~n1327 & n6877 ;
  assign n6879 = n6878 ^ n1707 ^ 1'b0 ;
  assign n6884 = n633 | n4166 ;
  assign n6885 = n6884 ^ n1860 ^ 1'b0 ;
  assign n6880 = n1301 & ~n1707 ;
  assign n6881 = n672 & n6880 ;
  assign n6882 = n6881 ^ n729 ^ 1'b0 ;
  assign n6883 = n3542 & ~n6882 ;
  assign n6886 = n6885 ^ n6883 ^ 1'b0 ;
  assign n6887 = ~n1879 & n5526 ;
  assign n6888 = n6887 ^ n2491 ^ 1'b0 ;
  assign n6889 = ( x152 & ~n1995 ) | ( x152 & n3104 ) | ( ~n1995 & n3104 ) ;
  assign n6890 = n4286 | n6889 ;
  assign n6891 = n6888 | n6890 ;
  assign n6892 = n6846 ^ n6739 ^ 1'b0 ;
  assign n6893 = n6892 ^ n5335 ^ n1939 ;
  assign n6895 = n4027 ^ n3027 ^ 1'b0 ;
  assign n6896 = n2942 & ~n6895 ;
  assign n6897 = n6896 ^ n3854 ^ n877 ;
  assign n6894 = n2025 ^ n1647 ^ n1495 ;
  assign n6898 = n6897 ^ n6894 ^ 1'b0 ;
  assign n6899 = ( n1145 & n6893 ) | ( n1145 & n6898 ) | ( n6893 & n6898 ) ;
  assign n6900 = n922 & ~n2504 ;
  assign n6901 = n6900 ^ n1961 ^ 1'b0 ;
  assign n6902 = n6901 ^ n3000 ^ 1'b0 ;
  assign n6903 = ~n1918 & n6902 ;
  assign n6904 = n2459 ^ n1260 ^ 1'b0 ;
  assign n6908 = n4930 & ~n6193 ;
  assign n6905 = n4143 ^ n2589 ^ n1012 ;
  assign n6906 = n6905 ^ n2669 ^ 1'b0 ;
  assign n6907 = n3381 & ~n6906 ;
  assign n6909 = n6908 ^ n6907 ^ 1'b0 ;
  assign n6910 = n6904 | n6909 ;
  assign n6915 = n2534 ^ n1836 ^ 1'b0 ;
  assign n6916 = ~n4958 & n6915 ;
  assign n6913 = n6796 ^ x103 ^ 1'b0 ;
  assign n6911 = ~n4164 & n6050 ;
  assign n6912 = ~n3500 & n6911 ;
  assign n6914 = n6913 ^ n6912 ^ 1'b0 ;
  assign n6917 = n6916 ^ n6914 ^ n2016 ;
  assign n6918 = n1022 | n2700 ;
  assign n6919 = n890 | n6918 ;
  assign n6920 = n6919 ^ n3357 ^ 1'b0 ;
  assign n6921 = n1893 | n6920 ;
  assign n6922 = n6921 ^ n5203 ^ 1'b0 ;
  assign n6928 = n621 ^ n539 ^ 1'b0 ;
  assign n6929 = ~n273 & n6928 ;
  assign n6923 = n5386 ^ n1724 ^ 1'b0 ;
  assign n6924 = ~n1113 & n6923 ;
  assign n6925 = ~n1693 & n2416 ;
  assign n6926 = n6925 ^ n1204 ^ 1'b0 ;
  assign n6927 = ( n6425 & ~n6924 ) | ( n6425 & n6926 ) | ( ~n6924 & n6926 ) ;
  assign n6930 = n6929 ^ n6927 ^ n5688 ;
  assign n6931 = n990 & n5979 ;
  assign n6933 = ( n964 & n1899 ) | ( n964 & ~n3087 ) | ( n1899 & ~n3087 ) ;
  assign n6932 = n1011 | n6519 ;
  assign n6934 = n6933 ^ n6932 ^ 1'b0 ;
  assign n6935 = n4979 ^ n1928 ^ 1'b0 ;
  assign n6936 = x159 & n6935 ;
  assign n6937 = ~n6345 & n6936 ;
  assign n6938 = n6937 ^ n2277 ^ 1'b0 ;
  assign n6939 = n802 & n2524 ;
  assign n6940 = n5744 & n6939 ;
  assign n6943 = n4203 ^ n2583 ^ 1'b0 ;
  assign n6944 = n318 & ~n6943 ;
  assign n6945 = n3504 ^ n1328 ^ 1'b0 ;
  assign n6946 = ( n290 & ~n1403 ) | ( n290 & n6945 ) | ( ~n1403 & n6945 ) ;
  assign n6947 = n6946 ^ n3240 ^ 1'b0 ;
  assign n6948 = n6944 & n6947 ;
  assign n6941 = n3866 ^ n2412 ^ 1'b0 ;
  assign n6942 = ( x82 & n4091 ) | ( x82 & ~n6941 ) | ( n4091 & ~n6941 ) ;
  assign n6949 = n6948 ^ n6942 ^ 1'b0 ;
  assign n6950 = n2403 & n6949 ;
  assign n6951 = n3758 ^ n2373 ^ 1'b0 ;
  assign n6952 = n4657 | n6951 ;
  assign n6953 = n6952 ^ n1129 ^ 1'b0 ;
  assign n6954 = ~n2624 & n6953 ;
  assign n6960 = x131 & ~n1076 ;
  assign n6961 = n6960 ^ n3061 ^ n1429 ;
  assign n6955 = ~n970 & n3934 ;
  assign n6956 = n4296 & n6955 ;
  assign n6957 = n1570 | n6956 ;
  assign n6958 = n1943 | n6957 ;
  assign n6959 = ~n6047 & n6958 ;
  assign n6962 = n6961 ^ n6959 ^ 1'b0 ;
  assign n6966 = ~n2590 & n3592 ;
  assign n6967 = n6966 ^ x135 ^ 1'b0 ;
  assign n6963 = ( n455 & n511 ) | ( n455 & ~n6030 ) | ( n511 & ~n6030 ) ;
  assign n6964 = n5472 ^ n2307 ^ 1'b0 ;
  assign n6965 = n6963 | n6964 ;
  assign n6968 = n6967 ^ n6965 ^ n6295 ;
  assign n6972 = ( ~n1129 & n1448 ) | ( ~n1129 & n4045 ) | ( n1448 & n4045 ) ;
  assign n6970 = n980 | n1636 ;
  assign n6971 = n4179 & ~n6970 ;
  assign n6969 = n5410 ^ n3825 ^ n3268 ;
  assign n6973 = n6972 ^ n6971 ^ n6969 ;
  assign n6974 = x67 & ~n2450 ;
  assign n6975 = n6974 ^ n810 ^ 1'b0 ;
  assign n6976 = n3347 ^ x160 ^ 1'b0 ;
  assign n6977 = x40 & ~n3106 ;
  assign n6978 = ~n6976 & n6977 ;
  assign n6979 = n6975 | n6978 ;
  assign n6980 = ( ~n1763 & n2374 ) | ( ~n1763 & n3999 ) | ( n2374 & n3999 ) ;
  assign n6981 = ( x62 & ~n738 ) | ( x62 & n2957 ) | ( ~n738 & n2957 ) ;
  assign n6982 = n606 | n1552 ;
  assign n6983 = ( ~n3481 & n6345 ) | ( ~n3481 & n6982 ) | ( n6345 & n6982 ) ;
  assign n6984 = n499 | n6983 ;
  assign n6985 = n6984 ^ n2916 ^ 1'b0 ;
  assign n6986 = ( n1420 & ~n6981 ) | ( n1420 & n6985 ) | ( ~n6981 & n6985 ) ;
  assign n6987 = n3813 ^ n3531 ^ 1'b0 ;
  assign n6988 = ( x103 & n6863 ) | ( x103 & n6987 ) | ( n6863 & n6987 ) ;
  assign n6989 = ( x90 & n1081 ) | ( x90 & ~n1675 ) | ( n1081 & ~n1675 ) ;
  assign n6990 = n6989 ^ n6415 ^ n3984 ;
  assign n6991 = n5265 ^ n3892 ^ n3341 ;
  assign n6992 = n5065 ^ n4113 ^ n1182 ;
  assign n6993 = ( ~n4496 & n5160 ) | ( ~n4496 & n6992 ) | ( n5160 & n6992 ) ;
  assign n6994 = n3949 ^ n2554 ^ 1'b0 ;
  assign n6995 = n6994 ^ n6549 ^ n2188 ;
  assign n6996 = x196 | n4200 ;
  assign n6997 = n4767 | n6996 ;
  assign n6998 = n5094 ^ n2843 ^ n599 ;
  assign n6999 = n1093 | n4260 ;
  assign n7000 = n3126 ^ n3039 ^ 1'b0 ;
  assign n7001 = n1542 & n7000 ;
  assign n7002 = n7001 ^ n717 ^ 1'b0 ;
  assign n7003 = n1549 | n1836 ;
  assign n7004 = ( n1145 & n4933 ) | ( n1145 & ~n7003 ) | ( n4933 & ~n7003 ) ;
  assign n7005 = ( x183 & ~n7002 ) | ( x183 & n7004 ) | ( ~n7002 & n7004 ) ;
  assign n7006 = n1842 | n7005 ;
  assign n7007 = n6999 & ~n7006 ;
  assign n7008 = n7007 ^ n1759 ^ 1'b0 ;
  assign n7009 = n2005 & n6411 ;
  assign n7013 = ~n1066 & n1818 ;
  assign n7014 = n1774 & n7013 ;
  assign n7011 = n4018 ^ n2972 ^ n2191 ;
  assign n7010 = ( n2296 & n3305 ) | ( n2296 & ~n3555 ) | ( n3305 & ~n3555 ) ;
  assign n7012 = n7011 ^ n7010 ^ 1'b0 ;
  assign n7015 = n7014 ^ n7012 ^ 1'b0 ;
  assign n7016 = ( ~n2046 & n6484 ) | ( ~n2046 & n7015 ) | ( n6484 & n7015 ) ;
  assign n7025 = ~n1042 & n2306 ;
  assign n7026 = ~n3329 & n7025 ;
  assign n7021 = n4417 & ~n5033 ;
  assign n7022 = ~n2375 & n7021 ;
  assign n7017 = n3400 ^ n883 ^ 1'b0 ;
  assign n7018 = n2984 & ~n7017 ;
  assign n7019 = n7018 ^ n1935 ^ 1'b0 ;
  assign n7020 = ~n4351 & n7019 ;
  assign n7023 = n7022 ^ n7020 ^ 1'b0 ;
  assign n7024 = n7023 ^ n5926 ^ 1'b0 ;
  assign n7027 = n7026 ^ n7024 ^ 1'b0 ;
  assign n7028 = n5087 ^ n1910 ^ n1742 ;
  assign n7029 = n7028 ^ n6664 ^ n1709 ;
  assign n7030 = n4487 ^ n4448 ^ n1185 ;
  assign n7031 = n2967 ^ n926 ^ 1'b0 ;
  assign n7032 = n5437 | n7031 ;
  assign n7033 = n1423 & ~n6652 ;
  assign n7034 = n7033 ^ n5801 ^ 1'b0 ;
  assign n7035 = ( n1910 & n2311 ) | ( n1910 & n3390 ) | ( n2311 & n3390 ) ;
  assign n7036 = ~n378 & n2216 ;
  assign n7037 = n7036 ^ n1197 ^ 1'b0 ;
  assign n7038 = n295 & ~n1576 ;
  assign n7039 = ~n7037 & n7038 ;
  assign n7040 = n1927 ^ n1562 ^ n639 ;
  assign n7041 = ~n268 & n2351 ;
  assign n7042 = n7041 ^ n3962 ^ 1'b0 ;
  assign n7043 = n7040 & n7042 ;
  assign n7044 = n7043 ^ n5627 ^ n4026 ;
  assign n7045 = ( ~n7035 & n7039 ) | ( ~n7035 & n7044 ) | ( n7039 & n7044 ) ;
  assign n7046 = n5170 ^ n2557 ^ n1266 ;
  assign n7047 = n1943 ^ n1289 ^ 1'b0 ;
  assign n7048 = ~n7046 & n7047 ;
  assign n7049 = n1955 & n7048 ;
  assign n7050 = n678 & ~n4447 ;
  assign n7051 = n7050 ^ n3022 ^ 1'b0 ;
  assign n7052 = n325 | n1700 ;
  assign n7053 = n7052 ^ n3343 ^ 1'b0 ;
  assign n7056 = n1025 ^ x89 ^ 1'b0 ;
  assign n7057 = n6612 | n7056 ;
  assign n7058 = n7057 ^ n5433 ^ n1579 ;
  assign n7054 = ~n345 & n2885 ;
  assign n7055 = ~x24 & n7054 ;
  assign n7059 = n7058 ^ n7055 ^ 1'b0 ;
  assign n7060 = n7053 & n7059 ;
  assign n7061 = n1725 & n5006 ;
  assign n7062 = n7061 ^ n3795 ^ 1'b0 ;
  assign n7063 = n7060 & n7062 ;
  assign n7064 = n4955 | n6008 ;
  assign n7065 = ( n1378 & n1757 ) | ( n1378 & ~n1869 ) | ( n1757 & ~n1869 ) ;
  assign n7066 = ( n1519 & n5425 ) | ( n1519 & ~n7065 ) | ( n5425 & ~n7065 ) ;
  assign n7067 = n7066 ^ n5732 ^ n1678 ;
  assign n7068 = n2427 & ~n2539 ;
  assign n7069 = ( x159 & ~n3739 ) | ( x159 & n7068 ) | ( ~n3739 & n7068 ) ;
  assign n7070 = n7069 ^ n2958 ^ n936 ;
  assign n7071 = n7067 | n7070 ;
  assign n7072 = n5541 ^ n1733 ^ 1'b0 ;
  assign n7073 = n5609 & ~n7001 ;
  assign n7075 = n1452 ^ n560 ^ x86 ;
  assign n7074 = n1236 | n4340 ;
  assign n7076 = n7075 ^ n7074 ^ 1'b0 ;
  assign n7077 = ( n702 & n808 ) | ( n702 & n3902 ) | ( n808 & n3902 ) ;
  assign n7078 = n1219 & n7077 ;
  assign n7079 = n2915 & ~n4639 ;
  assign n7080 = ~n2648 & n6031 ;
  assign n7081 = n7080 ^ n816 ^ x51 ;
  assign n7082 = n3070 | n7081 ;
  assign n7083 = n3725 & ~n7082 ;
  assign n7084 = ( n6045 & n7079 ) | ( n6045 & n7083 ) | ( n7079 & n7083 ) ;
  assign n7085 = n7078 | n7084 ;
  assign n7086 = n5538 ^ n2577 ^ n864 ;
  assign n7087 = ~n6289 & n6608 ;
  assign n7092 = ~n4845 & n6483 ;
  assign n7088 = ~n1021 & n1427 ;
  assign n7089 = n7088 ^ n3091 ^ n2427 ;
  assign n7090 = n7089 ^ n5456 ^ 1'b0 ;
  assign n7091 = ( n1720 & ~n2100 ) | ( n1720 & n7090 ) | ( ~n2100 & n7090 ) ;
  assign n7093 = n7092 ^ n7091 ^ 1'b0 ;
  assign n7094 = n3200 & ~n7093 ;
  assign n7100 = n2215 | n3475 ;
  assign n7097 = n1326 ^ n1312 ^ n981 ;
  assign n7098 = n7097 ^ n3318 ^ x202 ;
  assign n7099 = n7098 ^ n2226 ^ 1'b0 ;
  assign n7095 = n1220 ^ x79 ^ 1'b0 ;
  assign n7096 = ~n7062 & n7095 ;
  assign n7101 = n7100 ^ n7099 ^ n7096 ;
  assign n7102 = x73 & n6484 ;
  assign n7103 = n5810 ^ n4154 ^ 1'b0 ;
  assign n7104 = n1814 & ~n7103 ;
  assign n7105 = n2022 | n4982 ;
  assign n7106 = x15 | n7105 ;
  assign n7107 = n6390 ^ x37 ^ 1'b0 ;
  assign n7108 = ~n4372 & n7107 ;
  assign n7109 = ~n4195 & n5275 ;
  assign n7110 = n7109 ^ n2899 ^ n1187 ;
  assign n7111 = n1884 ^ n1831 ^ n1787 ;
  assign n7112 = n402 & ~n1636 ;
  assign n7113 = n7112 ^ n6626 ^ 1'b0 ;
  assign n7114 = n2976 & n7113 ;
  assign n7115 = ~n7111 & n7114 ;
  assign n7116 = ( x51 & ~n5756 ) | ( x51 & n7115 ) | ( ~n5756 & n7115 ) ;
  assign n7117 = ( n1326 & n5406 ) | ( n1326 & ~n7116 ) | ( n5406 & ~n7116 ) ;
  assign n7118 = n3010 ^ n652 ^ 1'b0 ;
  assign n7119 = n1106 | n7118 ;
  assign n7120 = n4759 ^ n3317 ^ n816 ;
  assign n7121 = n7120 ^ n2780 ^ 1'b0 ;
  assign n7122 = n7119 | n7121 ;
  assign n7124 = ~n2643 & n3229 ;
  assign n7123 = n5078 & ~n5524 ;
  assign n7125 = n7124 ^ n7123 ^ 1'b0 ;
  assign n7126 = n528 ^ n318 ^ 1'b0 ;
  assign n7127 = ~n1032 & n7126 ;
  assign n7128 = n7127 ^ n3291 ^ n2019 ;
  assign n7129 = n6893 | n7128 ;
  assign n7130 = n7129 ^ n4327 ^ 1'b0 ;
  assign n7131 = n1320 & n2155 ;
  assign n7132 = ~n4980 & n7131 ;
  assign n7133 = n1012 | n1693 ;
  assign n7134 = n7132 & ~n7133 ;
  assign n7135 = ( n754 & n892 ) | ( n754 & ~n5448 ) | ( n892 & ~n5448 ) ;
  assign n7136 = n2990 | n3875 ;
  assign n7137 = n520 & ~n1011 ;
  assign n7138 = n2691 & n7137 ;
  assign n7139 = n2062 | n4364 ;
  assign n7140 = n3021 | n7139 ;
  assign n7141 = n920 ^ n850 ^ n442 ;
  assign n7142 = n868 & n3731 ;
  assign n7143 = n7142 ^ n4233 ^ 1'b0 ;
  assign n7144 = n7141 | n7143 ;
  assign n7145 = ( ~n6133 & n7140 ) | ( ~n6133 & n7144 ) | ( n7140 & n7144 ) ;
  assign n7146 = n4699 ^ n4282 ^ 1'b0 ;
  assign n7147 = n1209 | n7146 ;
  assign n7148 = n7147 ^ n1248 ^ 1'b0 ;
  assign n7149 = n4940 | n7148 ;
  assign n7151 = n3516 ^ n1107 ^ 1'b0 ;
  assign n7150 = ~n3862 & n4291 ;
  assign n7152 = n7151 ^ n7150 ^ 1'b0 ;
  assign n7153 = n3887 | n4689 ;
  assign n7154 = x74 | n7153 ;
  assign n7155 = x183 | n545 ;
  assign n7156 = n7155 ^ n2734 ^ 1'b0 ;
  assign n7157 = n2270 & n7156 ;
  assign n7158 = n7157 ^ x17 ^ 1'b0 ;
  assign n7159 = n2046 & n7158 ;
  assign n7160 = n4461 ^ n1861 ^ 1'b0 ;
  assign n7161 = n6514 ^ n2937 ^ x146 ;
  assign n7162 = n586 & ~n1037 ;
  assign n7163 = ~n2822 & n7162 ;
  assign n7164 = n2616 | n7163 ;
  assign n7165 = n7161 | n7164 ;
  assign n7166 = n1550 & n4228 ;
  assign n7167 = n5253 & n7166 ;
  assign n7168 = n3526 ^ n1382 ^ 1'b0 ;
  assign n7169 = n6647 ^ n4518 ^ 1'b0 ;
  assign n7170 = n7168 & ~n7169 ;
  assign n7171 = n7170 ^ n2256 ^ 1'b0 ;
  assign n7172 = ( x72 & ~n3642 ) | ( x72 & n4314 ) | ( ~n3642 & n4314 ) ;
  assign n7173 = ~n1680 & n7172 ;
  assign n7174 = n7173 ^ n4812 ^ n1999 ;
  assign n7175 = n3242 & n5327 ;
  assign n7176 = n7175 ^ n4319 ^ 1'b0 ;
  assign n7177 = n3994 ^ n1178 ^ 1'b0 ;
  assign n7178 = n2236 & ~n6376 ;
  assign n7179 = ~n3830 & n7178 ;
  assign n7180 = n7177 & ~n7179 ;
  assign n7181 = ~n5039 & n7180 ;
  assign n7182 = ( ~n675 & n1852 ) | ( ~n675 & n3086 ) | ( n1852 & n3086 ) ;
  assign n7183 = ~n1415 & n1999 ;
  assign n7184 = n7183 ^ n4541 ^ 1'b0 ;
  assign n7185 = n5034 & n7184 ;
  assign n7186 = n7185 ^ n2570 ^ 1'b0 ;
  assign n7187 = n7182 & n7186 ;
  assign n7188 = n3875 ^ n3789 ^ 1'b0 ;
  assign n7189 = ~n4357 & n7188 ;
  assign n7190 = n5426 | n7189 ;
  assign n7191 = n6462 ^ n3156 ^ 1'b0 ;
  assign n7192 = x1 & ~n7191 ;
  assign n7193 = n7192 ^ n2674 ^ n1870 ;
  assign n7194 = n1256 | n7193 ;
  assign n7195 = n1229 & ~n7194 ;
  assign n7196 = n6688 ^ n5472 ^ 1'b0 ;
  assign n7197 = ( n4502 & n7195 ) | ( n4502 & ~n7196 ) | ( n7195 & ~n7196 ) ;
  assign n7198 = n490 | n7197 ;
  assign n7199 = n2462 | n7198 ;
  assign n7200 = ( x210 & n3165 ) | ( x210 & ~n7128 ) | ( n3165 & ~n7128 ) ;
  assign n7201 = n3222 & n7200 ;
  assign n7202 = ~n7199 & n7201 ;
  assign n7203 = ~n2841 & n4063 ;
  assign n7204 = ~n3874 & n7203 ;
  assign n7205 = n7204 ^ n3158 ^ 1'b0 ;
  assign n7206 = n1261 & ~n7205 ;
  assign n7207 = ~n6387 & n7206 ;
  assign n7208 = n7207 ^ n939 ^ 1'b0 ;
  assign n7209 = n7208 ^ n7055 ^ 1'b0 ;
  assign n7210 = n2954 ^ n1523 ^ 1'b0 ;
  assign n7211 = n6866 ^ x138 ^ 1'b0 ;
  assign n7212 = n3640 & n7211 ;
  assign n7213 = ( ~n658 & n3370 ) | ( ~n658 & n4963 ) | ( n3370 & n4963 ) ;
  assign n7214 = n7213 ^ n2859 ^ n1744 ;
  assign n7215 = n1447 ^ n848 ^ x194 ;
  assign n7216 = ~n2116 & n7215 ;
  assign n7217 = n3692 | n7216 ;
  assign n7218 = n2215 | n7217 ;
  assign n7219 = n2714 & ~n4200 ;
  assign n7220 = ~n7218 & n7219 ;
  assign n7221 = n2346 ^ n1079 ^ 1'b0 ;
  assign n7222 = ~n7220 & n7221 ;
  assign n7223 = ( ~n5915 & n6624 ) | ( ~n5915 & n7222 ) | ( n6624 & n7222 ) ;
  assign n7226 = n3854 ^ n256 ^ 1'b0 ;
  assign n7224 = n690 & ~n3078 ;
  assign n7225 = n3535 & n7224 ;
  assign n7227 = n7226 ^ n7225 ^ n861 ;
  assign n7228 = ( n1671 & n4395 ) | ( n1671 & n7227 ) | ( n4395 & n7227 ) ;
  assign n7229 = ~n2302 & n7228 ;
  assign n7230 = n7229 ^ n2762 ^ 1'b0 ;
  assign n7231 = x24 | n936 ;
  assign n7232 = n7231 ^ n2348 ^ 1'b0 ;
  assign n7233 = ~n3797 & n7232 ;
  assign n7234 = n7233 ^ n6597 ^ 1'b0 ;
  assign n7235 = n5729 ^ n5261 ^ 1'b0 ;
  assign n7236 = ( n5413 & n5589 ) | ( n5413 & n7235 ) | ( n5589 & n7235 ) ;
  assign n7237 = x226 & n864 ;
  assign n7238 = n6881 ^ n5747 ^ 1'b0 ;
  assign n7239 = n3180 ^ n1016 ^ 1'b0 ;
  assign n7240 = n4383 & ~n7239 ;
  assign n7241 = ~n2126 & n7240 ;
  assign n7242 = n4265 & n7241 ;
  assign n7243 = ~n3967 & n7242 ;
  assign n7244 = ( n5717 & n7238 ) | ( n5717 & ~n7243 ) | ( n7238 & ~n7243 ) ;
  assign n7245 = n1209 & n1749 ;
  assign n7246 = n7245 ^ n1851 ^ 1'b0 ;
  assign n7247 = n7246 ^ n1204 ^ 1'b0 ;
  assign n7248 = n3099 & n7247 ;
  assign n7249 = n7248 ^ n6976 ^ 1'b0 ;
  assign n7250 = ~n7244 & n7249 ;
  assign n7251 = n4314 | n5732 ;
  assign n7252 = n7251 ^ n2822 ^ 1'b0 ;
  assign n7253 = n5815 ^ n850 ^ 1'b0 ;
  assign n7254 = ~n1987 & n7253 ;
  assign n7255 = n4845 ^ n3631 ^ 1'b0 ;
  assign n7256 = n7254 & n7255 ;
  assign n7257 = ( ~n3378 & n7252 ) | ( ~n3378 & n7256 ) | ( n7252 & n7256 ) ;
  assign n7258 = n1828 | n7257 ;
  assign n7259 = x223 | n7258 ;
  assign n7265 = n4239 ^ n3700 ^ 1'b0 ;
  assign n7260 = n4618 ^ n1665 ^ x227 ;
  assign n7261 = n7260 ^ n2823 ^ 1'b0 ;
  assign n7262 = n3263 | n7261 ;
  assign n7263 = n7262 ^ n2367 ^ n941 ;
  assign n7264 = n2837 & n7263 ;
  assign n7266 = n7265 ^ n7264 ^ 1'b0 ;
  assign n7267 = ( n356 & ~n4999 ) | ( n356 & n7266 ) | ( ~n4999 & n7266 ) ;
  assign n7268 = n1647 & n7267 ;
  assign n7269 = n369 & n7268 ;
  assign n7272 = n391 | n3575 ;
  assign n7273 = n7272 ^ n2820 ^ 1'b0 ;
  assign n7274 = n6352 & n7273 ;
  assign n7275 = n1452 & n7274 ;
  assign n7270 = ( ~n3227 & n5572 ) | ( ~n3227 & n6259 ) | ( n5572 & n6259 ) ;
  assign n7271 = ( n378 & n6513 ) | ( n378 & ~n7270 ) | ( n6513 & ~n7270 ) ;
  assign n7276 = n7275 ^ n7271 ^ n3956 ;
  assign n7277 = n6364 ^ n3835 ^ 1'b0 ;
  assign n7278 = n415 & ~n1759 ;
  assign n7279 = n7278 ^ n3791 ^ 1'b0 ;
  assign n7280 = n7279 ^ n3898 ^ n2577 ;
  assign n7281 = ~n1145 & n2358 ;
  assign n7282 = n7281 ^ x170 ^ 1'b0 ;
  assign n7283 = n7282 ^ n4458 ^ 1'b0 ;
  assign n7284 = ~n3620 & n7283 ;
  assign n7285 = n7284 ^ n535 ^ 1'b0 ;
  assign n7288 = ( ~n453 & n464 ) | ( ~n453 & n2658 ) | ( n464 & n2658 ) ;
  assign n7287 = n563 & ~n4591 ;
  assign n7289 = n7288 ^ n7287 ^ 1'b0 ;
  assign n7286 = n563 & ~n2022 ;
  assign n7290 = n7289 ^ n7286 ^ 1'b0 ;
  assign n7291 = n7285 | n7290 ;
  assign n7292 = n2443 ^ x156 ^ 1'b0 ;
  assign n7293 = n1133 & ~n7292 ;
  assign n7294 = n468 & n7293 ;
  assign n7295 = n7294 ^ n3066 ^ 1'b0 ;
  assign n7296 = n1028 & ~n2513 ;
  assign n7297 = n971 & n7296 ;
  assign n7298 = n1222 & n7297 ;
  assign n7299 = n4522 ^ n4314 ^ 1'b0 ;
  assign n7300 = n595 & ~n6698 ;
  assign n7301 = n565 | n1755 ;
  assign n7302 = n7301 ^ x138 ^ 1'b0 ;
  assign n7303 = n6519 & n7302 ;
  assign n7304 = n7259 ^ n3694 ^ 1'b0 ;
  assign n7305 = n4454 ^ n4095 ^ n3596 ;
  assign n7306 = n3343 & n7305 ;
  assign n7307 = n7306 ^ n4804 ^ 1'b0 ;
  assign n7308 = n4374 | n7125 ;
  assign n7309 = n4944 ^ n4787 ^ 1'b0 ;
  assign n7310 = n4614 & n5413 ;
  assign n7311 = n7310 ^ n853 ^ 1'b0 ;
  assign n7312 = n4050 ^ n3957 ^ 1'b0 ;
  assign n7313 = n5162 & ~n7312 ;
  assign n7314 = ~n3732 & n7313 ;
  assign n7315 = n7314 ^ n5305 ^ 1'b0 ;
  assign n7316 = n7315 ^ n3729 ^ 1'b0 ;
  assign n7317 = n2504 ^ n1657 ^ 1'b0 ;
  assign n7318 = ~n6024 & n7317 ;
  assign n7319 = n5053 & n7318 ;
  assign n7320 = n3093 | n6619 ;
  assign n7321 = n1211 & n7320 ;
  assign n7322 = n4046 ^ n3578 ^ 1'b0 ;
  assign n7323 = ~n7321 & n7322 ;
  assign n7324 = n4264 & n7323 ;
  assign n7326 = n2339 ^ n1850 ^ 1'b0 ;
  assign n7325 = x210 & ~n1863 ;
  assign n7327 = n7326 ^ n7325 ^ 1'b0 ;
  assign n7328 = n4500 ^ n3366 ^ 1'b0 ;
  assign n7329 = n7327 & n7328 ;
  assign n7330 = ~n3364 & n7329 ;
  assign n7331 = n7330 ^ n3456 ^ 1'b0 ;
  assign n7332 = n503 ^ n375 ^ 1'b0 ;
  assign n7333 = n2722 | n7332 ;
  assign n7334 = ~n3110 & n7333 ;
  assign n7335 = n3739 & n4318 ;
  assign n7336 = n7335 ^ n5470 ^ n1572 ;
  assign n7338 = x157 | n2248 ;
  assign n7337 = ( n1757 & n3178 ) | ( n1757 & n3440 ) | ( n3178 & n3440 ) ;
  assign n7339 = n7338 ^ n7337 ^ n4046 ;
  assign n7340 = n7339 ^ n2264 ^ n1187 ;
  assign n7341 = n3634 ^ n1182 ^ 1'b0 ;
  assign n7342 = ~n903 & n7341 ;
  assign n7343 = n3239 & n7342 ;
  assign n7344 = n7343 ^ n5459 ^ 1'b0 ;
  assign n7345 = ( ~n2835 & n4609 ) | ( ~n2835 & n4751 ) | ( n4609 & n4751 ) ;
  assign n7346 = n7345 ^ n578 ^ 1'b0 ;
  assign n7347 = n7337 ^ n3080 ^ n1928 ;
  assign n7348 = n7347 ^ n5638 ^ 1'b0 ;
  assign n7349 = ( n1482 & n2401 ) | ( n1482 & ~n2577 ) | ( n2401 & ~n2577 ) ;
  assign n7350 = ~n3449 & n7349 ;
  assign n7351 = n7350 ^ n1107 ^ 1'b0 ;
  assign n7352 = n860 | n5017 ;
  assign n7353 = n7352 ^ n3100 ^ 1'b0 ;
  assign n7354 = n3455 ^ n3429 ^ n1457 ;
  assign n7355 = ( ~n449 & n7353 ) | ( ~n449 & n7354 ) | ( n7353 & n7354 ) ;
  assign n7356 = ~n4469 & n7355 ;
  assign n7359 = x41 & ~n1851 ;
  assign n7360 = ~n6068 & n7359 ;
  assign n7357 = x173 & ~n2422 ;
  assign n7358 = n3891 & n7357 ;
  assign n7361 = n7360 ^ n7358 ^ n266 ;
  assign n7362 = ( n535 & ~n600 ) | ( n535 & n827 ) | ( ~n600 & n827 ) ;
  assign n7363 = n6717 & ~n7362 ;
  assign n7364 = n3939 & n7363 ;
  assign n7365 = n4230 ^ n715 ^ 1'b0 ;
  assign n7366 = x119 & n7365 ;
  assign n7367 = n5458 & n7366 ;
  assign n7368 = n7367 ^ n3091 ^ 1'b0 ;
  assign n7369 = n2573 | n4237 ;
  assign n7370 = n4945 ^ n2159 ^ 1'b0 ;
  assign n7371 = n7370 ^ n3839 ^ x178 ;
  assign n7372 = n6725 & n7371 ;
  assign n7373 = n7369 & n7372 ;
  assign n7374 = n1486 & ~n4458 ;
  assign n7375 = n4264 & n7374 ;
  assign n7376 = n1201 ^ n1185 ^ x137 ;
  assign n7377 = n6646 & ~n7376 ;
  assign n7378 = n7377 ^ n3133 ^ 1'b0 ;
  assign n7379 = x132 & n738 ;
  assign n7380 = n7379 ^ n1337 ^ n873 ;
  assign n7381 = n3286 & n4778 ;
  assign n7382 = n861 & n1080 ;
  assign n7383 = n7382 ^ n2282 ^ 1'b0 ;
  assign n7384 = n883 & ~n7383 ;
  assign n7385 = ~n1993 & n3563 ;
  assign n7392 = ( ~n2097 & n2394 ) | ( ~n2097 & n4895 ) | ( n2394 & n4895 ) ;
  assign n7390 = ~n1732 & n3845 ;
  assign n7386 = n2244 ^ n1088 ^ x249 ;
  assign n7387 = x215 & n7386 ;
  assign n7388 = n1435 & n7387 ;
  assign n7389 = n7388 ^ n2061 ^ n286 ;
  assign n7391 = n7390 ^ n7389 ^ n5235 ;
  assign n7393 = n7392 ^ n7391 ^ 1'b0 ;
  assign n7394 = ~n2023 & n2756 ;
  assign n7398 = n621 & ~n1275 ;
  assign n7399 = n7398 ^ n1763 ^ 1'b0 ;
  assign n7396 = n1943 ^ n1055 ^ x40 ;
  assign n7397 = ( ~n560 & n2931 ) | ( ~n560 & n7396 ) | ( n2931 & n7396 ) ;
  assign n7395 = n2679 | n6644 ;
  assign n7400 = n7399 ^ n7397 ^ n7395 ;
  assign n7401 = ~n5992 & n7400 ;
  assign n7402 = ~n6188 & n7401 ;
  assign n7406 = n1784 | n3550 ;
  assign n7407 = n7406 ^ n5373 ^ 1'b0 ;
  assign n7403 = n1406 & n6826 ;
  assign n7404 = n609 | n7403 ;
  assign n7405 = ~n4602 & n7404 ;
  assign n7408 = n7407 ^ n7405 ^ 1'b0 ;
  assign n7409 = x100 & n6562 ;
  assign n7410 = n7409 ^ n6027 ^ 1'b0 ;
  assign n7411 = n4933 | n6897 ;
  assign n7412 = n7411 ^ n6498 ^ n2145 ;
  assign n7413 = ( n1666 & n4170 ) | ( n1666 & n4421 ) | ( n4170 & n4421 ) ;
  assign n7414 = n7148 & n7413 ;
  assign n7415 = n7412 & n7414 ;
  assign n7416 = n5188 ^ n3545 ^ n1861 ;
  assign n7417 = n4482 ^ n2882 ^ n1161 ;
  assign n7418 = n2889 & ~n7417 ;
  assign n7419 = n7418 ^ n879 ^ 1'b0 ;
  assign n7420 = n4101 & n7419 ;
  assign n7421 = n1420 | n7245 ;
  assign n7422 = n7421 ^ n1615 ^ 1'b0 ;
  assign n7424 = n619 | n3806 ;
  assign n7425 = n3585 & ~n7424 ;
  assign n7426 = ( n2972 & n3631 ) | ( n2972 & n7425 ) | ( n3631 & n7425 ) ;
  assign n7423 = ~n4532 & n6770 ;
  assign n7427 = n7426 ^ n7423 ^ 1'b0 ;
  assign n7429 = n3636 | n5830 ;
  assign n7430 = n2323 & ~n7429 ;
  assign n7428 = n3385 | n5916 ;
  assign n7431 = n7430 ^ n7428 ^ 1'b0 ;
  assign n7434 = ~n2915 & n4456 ;
  assign n7432 = n756 | n5648 ;
  assign n7433 = n3318 & ~n7432 ;
  assign n7435 = n7434 ^ n7433 ^ n1980 ;
  assign n7436 = n7435 ^ n4654 ^ n1583 ;
  assign n7437 = n2479 & ~n6557 ;
  assign n7438 = n7437 ^ n6675 ^ 1'b0 ;
  assign n7439 = n2663 & n7438 ;
  assign n7440 = ~x57 & n7366 ;
  assign n7441 = n6505 ^ n292 ^ 1'b0 ;
  assign n7442 = n6627 & ~n7441 ;
  assign n7443 = ~n6307 & n7442 ;
  assign n7444 = n2651 & n7443 ;
  assign n7445 = n4203 & ~n6783 ;
  assign n7446 = n7445 ^ n1269 ^ 1'b0 ;
  assign n7448 = n673 & ~n2992 ;
  assign n7447 = ( n5264 & ~n5758 ) | ( n5264 & n6826 ) | ( ~n5758 & n6826 ) ;
  assign n7449 = n7448 ^ n7447 ^ 1'b0 ;
  assign n7450 = n1054 & ~n7449 ;
  assign n7451 = ~n2204 & n6147 ;
  assign n7452 = ( n1529 & n6581 ) | ( n1529 & n7451 ) | ( n6581 & n7451 ) ;
  assign n7453 = n1693 | n3521 ;
  assign n7454 = n5879 | n7453 ;
  assign n7455 = n2995 & n3814 ;
  assign n7456 = n7455 ^ n4631 ^ 1'b0 ;
  assign n7457 = n1770 ^ n1438 ^ 1'b0 ;
  assign n7458 = x251 & ~n5134 ;
  assign n7459 = n4855 & n7458 ;
  assign n7460 = n7457 & n7459 ;
  assign n7461 = n4305 ^ x159 ^ 1'b0 ;
  assign n7462 = n878 | n7461 ;
  assign n7463 = n4150 ^ n2908 ^ 1'b0 ;
  assign n7464 = n1630 & n7463 ;
  assign n7465 = ~n1080 & n2516 ;
  assign n7466 = n3592 & n6292 ;
  assign n7467 = n883 ^ x82 ^ 1'b0 ;
  assign n7468 = ~n6542 & n7467 ;
  assign n7469 = ( n3139 & ~n5485 ) | ( n3139 & n7468 ) | ( ~n5485 & n7468 ) ;
  assign n7470 = n7469 ^ n6140 ^ 1'b0 ;
  assign n7471 = ~n351 & n4975 ;
  assign n7472 = n7471 ^ n4120 ^ 1'b0 ;
  assign n7473 = n5419 | n5782 ;
  assign n7474 = n2026 & ~n5345 ;
  assign n7475 = n7474 ^ n6001 ^ 1'b0 ;
  assign n7476 = n2223 | n4327 ;
  assign n7477 = n4043 ^ n571 ^ 1'b0 ;
  assign n7478 = ~n2992 & n7477 ;
  assign n7479 = n7478 ^ n848 ^ 1'b0 ;
  assign n7480 = x176 & ~n7479 ;
  assign n7481 = n7480 ^ n6074 ^ x229 ;
  assign n7483 = n623 | n3475 ;
  assign n7482 = n3139 ^ n2352 ^ 1'b0 ;
  assign n7484 = n7483 ^ n7482 ^ n7245 ;
  assign n7485 = n7484 ^ n6685 ^ 1'b0 ;
  assign n7486 = n1401 ^ n1232 ^ n652 ;
  assign n7487 = n7486 ^ n3376 ^ 1'b0 ;
  assign n7488 = n3185 & n7487 ;
  assign n7489 = n970 ^ x1 ^ 1'b0 ;
  assign n7490 = n3390 | n7489 ;
  assign n7491 = n7490 ^ n1635 ^ 1'b0 ;
  assign n7492 = n7488 & n7491 ;
  assign n7493 = ( n619 & ~n623 ) | ( n619 & n2238 ) | ( ~n623 & n2238 ) ;
  assign n7494 = n6824 ^ n3854 ^ 1'b0 ;
  assign n7495 = n6411 ^ n2726 ^ 1'b0 ;
  assign n7496 = ~n7065 & n7495 ;
  assign n7497 = n5552 ^ n3421 ^ n3401 ;
  assign n7498 = n2307 & n3853 ;
  assign n7499 = ~n5456 & n7498 ;
  assign n7500 = n7499 ^ n4260 ^ 1'b0 ;
  assign n7501 = ~n7497 & n7500 ;
  assign n7502 = ~n7496 & n7501 ;
  assign n7503 = ( n519 & n1063 ) | ( n519 & ~n2352 ) | ( n1063 & ~n2352 ) ;
  assign n7504 = n7503 ^ n7358 ^ n2509 ;
  assign n7505 = ~n1172 & n1884 ;
  assign n7506 = n7505 ^ n468 ^ 1'b0 ;
  assign n7507 = n7506 ^ n4345 ^ 1'b0 ;
  assign n7508 = ( ~n1103 & n4229 ) | ( ~n1103 & n7507 ) | ( n4229 & n7507 ) ;
  assign n7509 = n7448 ^ n2964 ^ 1'b0 ;
  assign n7511 = n407 & ~n1492 ;
  assign n7512 = n286 & n7511 ;
  assign n7510 = n679 & ~n6638 ;
  assign n7513 = n7512 ^ n7510 ^ 1'b0 ;
  assign n7514 = n7513 ^ n4278 ^ 1'b0 ;
  assign n7515 = ~n4781 & n7514 ;
  assign n7516 = n4777 & ~n6963 ;
  assign n7517 = ~n6688 & n7516 ;
  assign n7518 = n3656 ^ n2136 ^ 1'b0 ;
  assign n7519 = n7517 | n7518 ;
  assign n7521 = ~x99 & x195 ;
  assign n7520 = x18 & ~n3810 ;
  assign n7522 = n7521 ^ n7520 ^ 1'b0 ;
  assign n7523 = n2720 | n4630 ;
  assign n7524 = n2245 ^ n609 ^ 1'b0 ;
  assign n7525 = n4079 & ~n7524 ;
  assign n7526 = n7525 ^ n2262 ^ n1492 ;
  assign n7528 = ( n327 & n1298 ) | ( n327 & n6086 ) | ( n1298 & n6086 ) ;
  assign n7527 = n560 | n1463 ;
  assign n7529 = n7528 ^ n7527 ^ n3094 ;
  assign n7530 = n6232 ^ n3328 ^ n1322 ;
  assign n7531 = ~n1863 & n5199 ;
  assign n7532 = ~n5163 & n7531 ;
  assign n7533 = n2454 | n7532 ;
  assign n7534 = n7530 | n7533 ;
  assign n7535 = n1713 & ~n1789 ;
  assign n7536 = n7535 ^ n6351 ^ n4142 ;
  assign n7537 = n2889 ^ n2017 ^ 1'b0 ;
  assign n7538 = n6112 & ~n7537 ;
  assign n7539 = n879 | n5717 ;
  assign n7540 = n7539 ^ n2948 ^ 1'b0 ;
  assign n7541 = n7540 ^ n533 ^ 1'b0 ;
  assign n7542 = n2425 & n7541 ;
  assign n7543 = n1022 & ~n6523 ;
  assign n7544 = n4154 & ~n4578 ;
  assign n7545 = n7543 & n7544 ;
  assign n7546 = n302 & n4554 ;
  assign n7547 = n5386 ^ n4019 ^ 1'b0 ;
  assign n7548 = ( n890 & ~n3231 ) | ( n890 & n3430 ) | ( ~n3231 & n3430 ) ;
  assign n7549 = x191 & ~n447 ;
  assign n7550 = ( n381 & n7184 ) | ( n381 & ~n7549 ) | ( n7184 & ~n7549 ) ;
  assign n7551 = ~n3803 & n7550 ;
  assign n7552 = ( n7547 & n7548 ) | ( n7547 & ~n7551 ) | ( n7548 & ~n7551 ) ;
  assign n7553 = n1076 ^ n790 ^ 1'b0 ;
  assign n7554 = n7553 ^ n1617 ^ 1'b0 ;
  assign n7555 = n5356 ^ n574 ^ 1'b0 ;
  assign n7556 = n6188 & ~n7555 ;
  assign n7557 = ~n2513 & n7556 ;
  assign n7558 = n7557 ^ n4291 ^ 1'b0 ;
  assign n7559 = ~n7554 & n7558 ;
  assign n7560 = n1549 ^ n970 ^ n577 ;
  assign n7561 = n7560 ^ n2826 ^ n2538 ;
  assign n7562 = ( x113 & n1038 ) | ( x113 & n5570 ) | ( n1038 & n5570 ) ;
  assign n7563 = n6046 & ~n7562 ;
  assign n7564 = ~n7561 & n7563 ;
  assign n7567 = x103 & ~n6846 ;
  assign n7568 = ~x239 & n7567 ;
  assign n7569 = n6620 & ~n7568 ;
  assign n7565 = ~n2486 & n5143 ;
  assign n7566 = n7565 ^ n305 ^ 1'b0 ;
  assign n7570 = n7569 ^ n7566 ^ n1571 ;
  assign n7571 = ( ~n410 & n7564 ) | ( ~n410 & n7570 ) | ( n7564 & n7570 ) ;
  assign n7572 = ~n1724 & n4220 ;
  assign n7573 = n7572 ^ n1094 ^ 1'b0 ;
  assign n7574 = x251 & ~n2472 ;
  assign n7575 = n7573 & n7574 ;
  assign n7576 = n6269 ^ n2006 ^ 1'b0 ;
  assign n7577 = n6278 ^ n4837 ^ n925 ;
  assign n7578 = n5345 ^ n2258 ^ n1543 ;
  assign n7580 = ( n1088 & n2200 ) | ( n1088 & ~n7417 ) | ( n2200 & ~n7417 ) ;
  assign n7579 = ~n2373 & n3093 ;
  assign n7581 = n7580 ^ n7579 ^ n3389 ;
  assign n7582 = n5441 ^ n3148 ^ 1'b0 ;
  assign n7583 = n3681 & n7582 ;
  assign n7584 = n7583 ^ n2677 ^ 1'b0 ;
  assign n7585 = n3604 & n7584 ;
  assign n7588 = ~n4904 & n5592 ;
  assign n7589 = n7588 ^ n4052 ^ 1'b0 ;
  assign n7586 = n3755 ^ n1205 ^ 1'b0 ;
  assign n7587 = n3034 & n7586 ;
  assign n7590 = n7589 ^ n7587 ^ 1'b0 ;
  assign n7591 = n5337 ^ n2331 ^ x61 ;
  assign n7592 = ~n4214 & n7591 ;
  assign n7593 = n6065 & n7592 ;
  assign n7594 = ~n4603 & n7593 ;
  assign n7595 = n5544 & n6903 ;
  assign n7597 = n906 & ~n7011 ;
  assign n7598 = n7597 ^ n5889 ^ 1'b0 ;
  assign n7596 = n2782 & n2798 ;
  assign n7599 = n7598 ^ n7596 ^ 1'b0 ;
  assign n7600 = n545 & n4143 ;
  assign n7601 = ~n5199 & n7600 ;
  assign n7602 = n5956 ^ n5740 ^ n914 ;
  assign n7605 = n595 & n1907 ;
  assign n7606 = ~n5351 & n7605 ;
  assign n7604 = x37 | n7115 ;
  assign n7607 = n7606 ^ n7604 ^ n2321 ;
  assign n7603 = n1550 & n6706 ;
  assign n7608 = n7607 ^ n7603 ^ 1'b0 ;
  assign n7615 = n430 & ~n1307 ;
  assign n7616 = n1021 & n7615 ;
  assign n7609 = ~n3307 & n6513 ;
  assign n7610 = n7609 ^ x173 ^ 1'b0 ;
  assign n7611 = n1696 ^ n1241 ^ 1'b0 ;
  assign n7612 = n2473 ^ n1438 ^ 1'b0 ;
  assign n7613 = n7611 & n7612 ;
  assign n7614 = ~n7610 & n7613 ;
  assign n7617 = n7616 ^ n7614 ^ 1'b0 ;
  assign n7618 = n7617 ^ n1144 ^ 1'b0 ;
  assign n7619 = ( n1152 & n4369 ) | ( n1152 & n4928 ) | ( n4369 & n4928 ) ;
  assign n7620 = n7001 | n7619 ;
  assign n7621 = n6545 & ~n7620 ;
  assign n7622 = ( n3305 & ~n3947 ) | ( n3305 & n7621 ) | ( ~n3947 & n7621 ) ;
  assign n7627 = x220 | n5579 ;
  assign n7624 = n3494 ^ n2637 ^ 1'b0 ;
  assign n7625 = n7624 ^ n925 ^ 1'b0 ;
  assign n7623 = n575 | n4351 ;
  assign n7626 = n7625 ^ n7623 ^ 1'b0 ;
  assign n7628 = n7627 ^ n7626 ^ n1067 ;
  assign n7629 = ( n347 & n2733 ) | ( n347 & ~n5258 ) | ( n2733 & ~n5258 ) ;
  assign n7630 = n5133 & n7629 ;
  assign n7631 = ~n795 & n7195 ;
  assign n7632 = n7631 ^ n1910 ^ 1'b0 ;
  assign n7633 = n7632 ^ n862 ^ 1'b0 ;
  assign n7634 = n7630 & n7633 ;
  assign n7635 = ( n704 & n1874 ) | ( n704 & n7488 ) | ( n1874 & n7488 ) ;
  assign n7636 = n621 & n690 ;
  assign n7637 = n7636 ^ n1164 ^ 1'b0 ;
  assign n7638 = ( n493 & ~n1980 ) | ( n493 & n7155 ) | ( ~n1980 & n7155 ) ;
  assign n7639 = n4391 ^ n1987 ^ n578 ;
  assign n7640 = x232 & ~n7639 ;
  assign n7641 = n7638 & n7640 ;
  assign n7642 = n1873 & ~n2486 ;
  assign n7643 = n7642 ^ x24 ^ 1'b0 ;
  assign n7644 = ( ~n933 & n1572 ) | ( ~n933 & n7643 ) | ( n1572 & n7643 ) ;
  assign n7645 = ~n7641 & n7644 ;
  assign n7646 = n7645 ^ n3959 ^ 1'b0 ;
  assign n7647 = n7637 & ~n7646 ;
  assign n7648 = n3394 ^ n2708 ^ 1'b0 ;
  assign n7649 = n927 & ~n7648 ;
  assign n7650 = ( n824 & ~n3714 ) | ( n824 & n4163 ) | ( ~n3714 & n4163 ) ;
  assign n7651 = n7649 & ~n7650 ;
  assign n7652 = n7651 ^ n3097 ^ 1'b0 ;
  assign n7657 = ( n718 & n843 ) | ( n718 & ~n4446 ) | ( n843 & ~n4446 ) ;
  assign n7653 = ( ~n697 & n1993 ) | ( ~n697 & n2970 ) | ( n1993 & n2970 ) ;
  assign n7654 = n4514 & n7653 ;
  assign n7655 = n2680 & n7654 ;
  assign n7656 = n1938 & ~n7655 ;
  assign n7658 = n7657 ^ n7656 ^ 1'b0 ;
  assign n7659 = n1934 | n7658 ;
  assign n7660 = n7652 | n7659 ;
  assign n7661 = ( n3122 & ~n3722 ) | ( n3122 & n3737 ) | ( ~n3722 & n3737 ) ;
  assign n7662 = ~n6752 & n7506 ;
  assign n7663 = ~x24 & n7662 ;
  assign n7664 = ( n7550 & ~n7661 ) | ( n7550 & n7663 ) | ( ~n7661 & n7663 ) ;
  assign n7665 = n718 & ~n769 ;
  assign n7666 = n4084 & ~n5967 ;
  assign n7667 = n7665 & n7666 ;
  assign n7668 = n1605 | n4137 ;
  assign n7669 = n489 & n1853 ;
  assign n7670 = n7669 ^ n6114 ^ 1'b0 ;
  assign n7672 = n902 ^ x192 ^ 1'b0 ;
  assign n7673 = n6793 ^ x205 ^ 1'b0 ;
  assign n7674 = ~n7672 & n7673 ;
  assign n7671 = n2852 & ~n6425 ;
  assign n7675 = n7674 ^ n7671 ^ 1'b0 ;
  assign n7676 = ( n686 & ~n2790 ) | ( n686 & n7675 ) | ( ~n2790 & n7675 ) ;
  assign n7679 = n2692 ^ n1047 ^ 1'b0 ;
  assign n7680 = n445 | n7679 ;
  assign n7681 = n3716 & ~n7680 ;
  assign n7682 = n7681 ^ n6287 ^ 1'b0 ;
  assign n7683 = n1083 & ~n7682 ;
  assign n7684 = n7683 ^ n2692 ^ 1'b0 ;
  assign n7677 = n3621 & n3687 ;
  assign n7678 = n7677 ^ n7184 ^ 1'b0 ;
  assign n7685 = n7684 ^ n7678 ^ 1'b0 ;
  assign n7686 = n507 & n7685 ;
  assign n7687 = ( ~n5710 & n7676 ) | ( ~n5710 & n7686 ) | ( n7676 & n7686 ) ;
  assign n7688 = n1247 & ~n5255 ;
  assign n7689 = n7688 ^ n2491 ^ 1'b0 ;
  assign n7690 = n7689 ^ n3945 ^ n3213 ;
  assign n7691 = ( n2214 & n7051 ) | ( n2214 & ~n7690 ) | ( n7051 & ~n7690 ) ;
  assign n7692 = ( n1486 & n6438 ) | ( n1486 & n7691 ) | ( n6438 & n7691 ) ;
  assign n7693 = ( n645 & n2752 ) | ( n645 & ~n3414 ) | ( n2752 & ~n3414 ) ;
  assign n7694 = n4174 & ~n6123 ;
  assign n7695 = n3188 & n7142 ;
  assign n7696 = n1804 | n4731 ;
  assign n7697 = n7359 ^ n4569 ^ n3042 ;
  assign n7698 = n5956 & n7697 ;
  assign n7699 = n7698 ^ n6981 ^ 1'b0 ;
  assign n7700 = n801 & n4496 ;
  assign n7701 = n7700 ^ x179 ^ 1'b0 ;
  assign n7702 = ( ~n2058 & n5248 ) | ( ~n2058 & n6846 ) | ( n5248 & n6846 ) ;
  assign n7703 = n2538 | n4170 ;
  assign n7704 = ~x150 & n2244 ;
  assign n7705 = n7704 ^ n1499 ^ 1'b0 ;
  assign n7706 = n4587 ^ n736 ^ 1'b0 ;
  assign n7707 = x164 & n7706 ;
  assign n7708 = n2615 & n7707 ;
  assign n7709 = n3381 ^ n3152 ^ 1'b0 ;
  assign n7710 = ~n629 & n7709 ;
  assign n7711 = n5376 & n7710 ;
  assign n7714 = n1602 ^ n1236 ^ 1'b0 ;
  assign n7715 = n2230 & n7714 ;
  assign n7716 = ~n1861 & n7715 ;
  assign n7717 = n1328 & n7716 ;
  assign n7718 = n7717 ^ n5169 ^ 1'b0 ;
  assign n7719 = n4679 | n7718 ;
  assign n7712 = n2900 ^ n2399 ^ 1'b0 ;
  assign n7713 = x59 & n7712 ;
  assign n7720 = n7719 ^ n7713 ^ 1'b0 ;
  assign n7721 = ( n2106 & n2651 ) | ( n2106 & ~n3072 ) | ( n2651 & ~n3072 ) ;
  assign n7722 = n1742 | n7721 ;
  assign n7723 = n7722 ^ n3263 ^ 1'b0 ;
  assign n7724 = ~n1229 & n2678 ;
  assign n7725 = ~n1999 & n7724 ;
  assign n7726 = n2251 ^ n1407 ^ n824 ;
  assign n7727 = n7726 ^ n5424 ^ n4725 ;
  assign n7728 = n7727 ^ n6808 ^ n3178 ;
  assign n7729 = ( n5505 & ~n5935 ) | ( n5505 & n7728 ) | ( ~n5935 & n7728 ) ;
  assign n7730 = ( ~n2658 & n7725 ) | ( ~n2658 & n7729 ) | ( n7725 & n7729 ) ;
  assign n7731 = n7730 ^ n5368 ^ 1'b0 ;
  assign n7732 = n3798 & n4679 ;
  assign n7733 = ( ~n2447 & n3062 ) | ( ~n2447 & n7732 ) | ( n3062 & n7732 ) ;
  assign n7734 = n7733 ^ n1989 ^ 1'b0 ;
  assign n7735 = n1058 & ~n7734 ;
  assign n7736 = ~n1861 & n7735 ;
  assign n7737 = n7462 & ~n7736 ;
  assign n7741 = n1302 & n4932 ;
  assign n7742 = n7741 ^ n2907 ^ 1'b0 ;
  assign n7743 = x111 & n7742 ;
  assign n7738 = n3994 ^ n3147 ^ 1'b0 ;
  assign n7739 = n3540 & ~n7738 ;
  assign n7740 = n3624 & ~n7739 ;
  assign n7744 = n7743 ^ n7740 ^ n3669 ;
  assign n7745 = n4611 ^ n4214 ^ 1'b0 ;
  assign n7746 = n7745 ^ n6510 ^ 1'b0 ;
  assign n7749 = n4263 ^ n1257 ^ 1'b0 ;
  assign n7747 = ( n866 & n2488 ) | ( n866 & ~n5883 ) | ( n2488 & ~n5883 ) ;
  assign n7748 = n5903 & n7747 ;
  assign n7750 = n7749 ^ n7748 ^ 1'b0 ;
  assign n7751 = n5351 & ~n7750 ;
  assign n7752 = n7751 ^ n2713 ^ 1'b0 ;
  assign n7753 = n2326 & ~n4427 ;
  assign n7754 = n7752 & n7753 ;
  assign n7755 = n1379 ^ n1365 ^ 1'b0 ;
  assign n7756 = n7755 ^ n6848 ^ 1'b0 ;
  assign n7757 = n4210 & n7756 ;
  assign n7758 = n3147 | n4552 ;
  assign n7759 = n5351 ^ n5177 ^ 1'b0 ;
  assign n7760 = n7759 ^ n5441 ^ n1592 ;
  assign n7761 = ( n4600 & ~n6463 ) | ( n4600 & n7760 ) | ( ~n6463 & n7760 ) ;
  assign n7762 = n6851 ^ n2800 ^ 1'b0 ;
  assign n7763 = n1080 & ~n7762 ;
  assign n7764 = n7763 ^ n2117 ^ 1'b0 ;
  assign n7765 = n7764 ^ n4561 ^ n1860 ;
  assign n7766 = n4741 & ~n7595 ;
  assign n7768 = x171 & n2304 ;
  assign n7769 = n7768 ^ n341 ^ 1'b0 ;
  assign n7767 = ( n857 & ~n3019 ) | ( n857 & n3551 ) | ( ~n3019 & n3551 ) ;
  assign n7770 = n7769 ^ n7767 ^ 1'b0 ;
  assign n7771 = n2052 ^ n639 ^ 1'b0 ;
  assign n7772 = n1816 | n7771 ;
  assign n7773 = ( ~n4469 & n7452 ) | ( ~n4469 & n7772 ) | ( n7452 & n7772 ) ;
  assign n7774 = ( n3704 & ~n3781 ) | ( n3704 & n5232 ) | ( ~n3781 & n5232 ) ;
  assign n7775 = n4542 & n7774 ;
  assign n7776 = ~n3263 & n7393 ;
  assign n7777 = n7650 ^ n841 ^ 1'b0 ;
  assign n7778 = ~n1908 & n5109 ;
  assign n7779 = n7778 ^ n5609 ^ 1'b0 ;
  assign n7780 = n5037 ^ n2292 ^ 1'b0 ;
  assign n7781 = n7779 | n7780 ;
  assign n7782 = n7777 & ~n7781 ;
  assign n7783 = x182 & n6062 ;
  assign n7784 = n7783 ^ n2995 ^ 1'b0 ;
  assign n7785 = ( n547 & ~n2378 ) | ( n547 & n7784 ) | ( ~n2378 & n7784 ) ;
  assign n7788 = n3014 ^ n2504 ^ 1'b0 ;
  assign n7786 = n1154 ^ n955 ^ 1'b0 ;
  assign n7787 = n2799 | n7786 ;
  assign n7789 = n7788 ^ n7787 ^ 1'b0 ;
  assign n7790 = ~n5255 & n7789 ;
  assign n7791 = n3040 ^ n2280 ^ 1'b0 ;
  assign n7792 = n5236 & ~n7791 ;
  assign n7793 = n1650 & ~n6818 ;
  assign n7794 = n7793 ^ n588 ^ 1'b0 ;
  assign n7795 = n879 & n3157 ;
  assign n7796 = n2357 ^ n2274 ^ n1640 ;
  assign n7797 = ~n5417 & n7796 ;
  assign n7798 = n7797 ^ n4402 ^ 1'b0 ;
  assign n7799 = n2914 | n7798 ;
  assign n7800 = n7795 | n7799 ;
  assign n7801 = ~n2283 & n5613 ;
  assign n7802 = n3873 & ~n7801 ;
  assign n7806 = n3360 & n3975 ;
  assign n7807 = n7806 ^ n5199 ^ n2326 ;
  assign n7804 = n2461 & n5028 ;
  assign n7805 = n7804 ^ n1867 ^ n1285 ;
  assign n7803 = n6991 ^ n2779 ^ 1'b0 ;
  assign n7808 = n7807 ^ n7805 ^ n7803 ;
  assign n7809 = n5412 | n5620 ;
  assign n7810 = n7809 ^ n2185 ^ 1'b0 ;
  assign n7811 = n2290 & ~n7810 ;
  assign n7812 = n2488 ^ n1494 ^ 1'b0 ;
  assign n7813 = n987 & ~n6316 ;
  assign n7814 = n7200 & ~n7813 ;
  assign n7815 = ( ~n6110 & n7812 ) | ( ~n6110 & n7814 ) | ( n7812 & n7814 ) ;
  assign n7818 = n7065 & n7649 ;
  assign n7816 = n1438 ^ x189 ^ 1'b0 ;
  assign n7817 = n6114 & ~n7816 ;
  assign n7819 = n7818 ^ n7817 ^ 1'b0 ;
  assign n7820 = n982 & n2852 ;
  assign n7821 = n7820 ^ n1131 ^ 1'b0 ;
  assign n7822 = n7821 ^ n931 ^ 1'b0 ;
  assign n7823 = ( n5771 & n7296 ) | ( n5771 & n7822 ) | ( n7296 & n7822 ) ;
  assign n7824 = ~n2150 & n3909 ;
  assign n7825 = n7824 ^ n609 ^ 1'b0 ;
  assign n7826 = n7825 ^ n1425 ^ 1'b0 ;
  assign n7827 = n6384 | n7826 ;
  assign n7828 = n4473 & ~n7827 ;
  assign n7829 = ~n7823 & n7828 ;
  assign n7830 = n3523 ^ n1750 ^ 1'b0 ;
  assign n7831 = n2522 | n4373 ;
  assign n7832 = n7665 & ~n7831 ;
  assign n7833 = n7832 ^ n6903 ^ 1'b0 ;
  assign n7835 = n1100 | n1778 ;
  assign n7834 = x53 & ~n1026 ;
  assign n7836 = n7835 ^ n7834 ^ 1'b0 ;
  assign n7837 = n7836 ^ n4995 ^ 1'b0 ;
  assign n7838 = n7837 ^ n1657 ^ 1'b0 ;
  assign n7839 = n1359 & ~n4501 ;
  assign n7840 = n7839 ^ n835 ^ 1'b0 ;
  assign n7841 = ( ~n1258 & n3458 ) | ( ~n1258 & n7840 ) | ( n3458 & n7840 ) ;
  assign n7842 = n7841 ^ n6228 ^ 1'b0 ;
  assign n7843 = n1506 & ~n3646 ;
  assign n7844 = n1253 | n6047 ;
  assign n7845 = n7844 ^ n3320 ^ n3033 ;
  assign n7846 = n4644 ^ n1422 ^ n1133 ;
  assign n7850 = n1690 & n2548 ;
  assign n7847 = n3931 ^ x16 ^ 1'b0 ;
  assign n7848 = ( n2674 & ~n6174 ) | ( n2674 & n7847 ) | ( ~n6174 & n7847 ) ;
  assign n7849 = n1463 | n7848 ;
  assign n7851 = n7850 ^ n7849 ^ 1'b0 ;
  assign n7852 = n4056 & n7851 ;
  assign n7853 = n4378 ^ n2735 ^ 1'b0 ;
  assign n7854 = n3617 | n7853 ;
  assign n7855 = n7854 ^ n7637 ^ 1'b0 ;
  assign n7856 = n1501 | n1860 ;
  assign n7857 = x205 & n7856 ;
  assign n7858 = n7196 ^ n4981 ^ n1161 ;
  assign n7859 = n2957 & n3500 ;
  assign n7860 = n7859 ^ n1257 ^ n951 ;
  assign n7861 = n7860 ^ n7818 ^ 1'b0 ;
  assign n7862 = ~n3961 & n7861 ;
  assign n7863 = n2976 ^ n2861 ^ n2798 ;
  assign n7864 = n2329 & n7863 ;
  assign n7865 = ( ~n589 & n2255 ) | ( ~n589 & n7864 ) | ( n2255 & n7864 ) ;
  assign n7866 = n6345 ^ x213 ^ 1'b0 ;
  assign n7867 = n7865 | n7866 ;
  assign n7868 = x143 & n5274 ;
  assign n7869 = n7868 ^ n808 ^ 1'b0 ;
  assign n7870 = n1884 ^ n335 ^ 1'b0 ;
  assign n7871 = n5706 & ~n7870 ;
  assign n7872 = n7871 ^ n7610 ^ n2919 ;
  assign n7873 = ~n552 & n6445 ;
  assign n7874 = n2827 & n7873 ;
  assign n7875 = n7872 | n7874 ;
  assign n7876 = n6450 ^ n5525 ^ 1'b0 ;
  assign n7877 = n7876 ^ n6730 ^ 1'b0 ;
  assign n7878 = n4616 ^ n3015 ^ n914 ;
  assign n7879 = n1838 & ~n4896 ;
  assign n7880 = n5565 ^ n2770 ^ 1'b0 ;
  assign n7881 = ( n4303 & n7879 ) | ( n4303 & ~n7880 ) | ( n7879 & ~n7880 ) ;
  assign n7882 = n7320 & n7804 ;
  assign n7883 = n7882 ^ n298 ^ 1'b0 ;
  assign n7884 = n5609 ^ n1336 ^ 1'b0 ;
  assign n7885 = n5518 & n7884 ;
  assign n7886 = ( ~n4528 & n7883 ) | ( ~n4528 & n7885 ) | ( n7883 & n7885 ) ;
  assign n7887 = x167 & ~n2259 ;
  assign n7888 = x40 | n7887 ;
  assign n7890 = ~n1603 & n2728 ;
  assign n7891 = n2169 & n7890 ;
  assign n7889 = x226 & n4868 ;
  assign n7892 = n7891 ^ n7889 ^ 1'b0 ;
  assign n7893 = n7892 ^ n5124 ^ 1'b0 ;
  assign n7894 = n1886 & ~n3896 ;
  assign n7895 = n1701 ^ x51 ^ 1'b0 ;
  assign n7896 = x80 & ~n7895 ;
  assign n7897 = n7896 ^ n4837 ^ 1'b0 ;
  assign n7898 = n1989 | n4108 ;
  assign n7899 = n7898 ^ n3429 ^ 1'b0 ;
  assign n7900 = n7899 ^ n3604 ^ 1'b0 ;
  assign n7901 = ~n2838 & n7900 ;
  assign n7902 = n390 & n1634 ;
  assign n7903 = n7902 ^ n3788 ^ 1'b0 ;
  assign n7904 = n7901 & n7903 ;
  assign n7905 = ( n7894 & n7897 ) | ( n7894 & n7904 ) | ( n7897 & n7904 ) ;
  assign n7906 = n3922 ^ n3779 ^ 1'b0 ;
  assign n7908 = n696 & ~n6063 ;
  assign n7907 = n2771 | n7891 ;
  assign n7909 = n7908 ^ n7907 ^ 1'b0 ;
  assign n7910 = x227 & ~n7909 ;
  assign n7911 = x229 & ~n7910 ;
  assign n7912 = n4659 & n7911 ;
  assign n7920 = n2207 & n4063 ;
  assign n7921 = n1966 & n7920 ;
  assign n7922 = n6326 & n7921 ;
  assign n7915 = n7726 ^ n2221 ^ 1'b0 ;
  assign n7916 = ~n3107 & n3691 ;
  assign n7917 = n7915 & n7916 ;
  assign n7918 = n6893 & n7917 ;
  assign n7913 = n2222 & n7899 ;
  assign n7914 = n4626 | n7913 ;
  assign n7919 = n7918 ^ n7914 ^ 1'b0 ;
  assign n7923 = n7922 ^ n7919 ^ 1'b0 ;
  assign n7924 = ~n2507 & n2769 ;
  assign n7925 = ~x155 & n7924 ;
  assign n7926 = n2794 ^ x214 ^ 1'b0 ;
  assign n7927 = n2626 | n7926 ;
  assign n7928 = n2052 | n5056 ;
  assign n7929 = n7928 ^ n7026 ^ 1'b0 ;
  assign n7930 = n7929 ^ n7634 ^ n5929 ;
  assign n7931 = n2582 & n3375 ;
  assign n7932 = n7931 ^ x197 ^ 1'b0 ;
  assign n7933 = n5619 | n7932 ;
  assign n7934 = n2287 & ~n7933 ;
  assign n7935 = ~n2486 & n6867 ;
  assign n7936 = ~n1047 & n7935 ;
  assign n7937 = n7934 | n7936 ;
  assign n7938 = n7937 ^ n6170 ^ 1'b0 ;
  assign n7941 = n1543 & ~n5237 ;
  assign n7942 = n825 & n7941 ;
  assign n7939 = n597 | n3549 ;
  assign n7940 = n482 | n7939 ;
  assign n7943 = n7942 ^ n7940 ^ 1'b0 ;
  assign n7944 = n6011 & ~n7943 ;
  assign n7945 = n2986 & ~n3473 ;
  assign n7946 = n7945 ^ n1024 ^ 1'b0 ;
  assign n7947 = x241 & ~n4155 ;
  assign n7948 = n7947 ^ n6023 ^ 1'b0 ;
  assign n7949 = ~n1672 & n7948 ;
  assign n7950 = n7949 ^ n832 ^ 1'b0 ;
  assign n7951 = n3000 & n7950 ;
  assign n7952 = ~n2820 & n7951 ;
  assign n7953 = n7952 ^ n1690 ^ 1'b0 ;
  assign n7954 = n7946 & n7953 ;
  assign n7955 = n7954 ^ n5006 ^ 1'b0 ;
  assign n7956 = n4474 & n7955 ;
  assign n7957 = ~n3304 & n7956 ;
  assign n7958 = n3283 ^ n2350 ^ 1'b0 ;
  assign n7959 = n7765 ^ n5221 ^ 1'b0 ;
  assign n7969 = n667 | n5134 ;
  assign n7970 = n961 | n7969 ;
  assign n7971 = n7970 ^ n531 ^ 1'b0 ;
  assign n7960 = ~n665 & n759 ;
  assign n7961 = n7960 ^ n3739 ^ 1'b0 ;
  assign n7962 = n2529 ^ n1145 ^ 1'b0 ;
  assign n7963 = ~n7961 & n7962 ;
  assign n7966 = n863 | n2047 ;
  assign n7964 = n635 & n1675 ;
  assign n7965 = n7964 ^ n5428 ^ 1'b0 ;
  assign n7967 = n7966 ^ n7965 ^ 1'b0 ;
  assign n7968 = n7963 & ~n7967 ;
  assign n7972 = n7971 ^ n7968 ^ 1'b0 ;
  assign n7973 = ~n7690 & n7972 ;
  assign n7974 = n341 & ~n6003 ;
  assign n7975 = n2769 ^ x44 ^ 1'b0 ;
  assign n7976 = n5469 | n7975 ;
  assign n7977 = n7976 ^ n6691 ^ 1'b0 ;
  assign n7978 = ~n3567 & n7977 ;
  assign n7979 = ( n2433 & n5613 ) | ( n2433 & n7978 ) | ( n5613 & n7978 ) ;
  assign n7980 = n6919 ^ n6207 ^ 1'b0 ;
  assign n7981 = n4713 & ~n7980 ;
  assign n7982 = ~n6973 & n7981 ;
  assign n7985 = n1588 ^ x97 ^ 1'b0 ;
  assign n7983 = n1452 & n6373 ;
  assign n7984 = ~n2919 & n7983 ;
  assign n7986 = n7985 ^ n7984 ^ 1'b0 ;
  assign n7987 = n2798 ^ n2009 ^ 1'b0 ;
  assign n7988 = n7987 ^ n5206 ^ 1'b0 ;
  assign n7989 = n5904 ^ n2502 ^ 1'b0 ;
  assign n7990 = n4707 | n7989 ;
  assign n7991 = n6711 ^ n3991 ^ n3527 ;
  assign n7992 = ( ~n1415 & n4424 ) | ( ~n1415 & n7991 ) | ( n4424 & n7991 ) ;
  assign n7993 = n2940 ^ n2354 ^ 1'b0 ;
  assign n7994 = ~n6554 & n7993 ;
  assign n7995 = n3813 ^ n3722 ^ n2138 ;
  assign n7996 = n1691 ^ n659 ^ 1'b0 ;
  assign n7997 = n7284 ^ n4340 ^ 1'b0 ;
  assign n7998 = n7996 | n7997 ;
  assign n7999 = n1043 | n7998 ;
  assign n8000 = n7995 & ~n7999 ;
  assign n8001 = n7994 | n8000 ;
  assign n8002 = n7968 ^ n390 ^ 1'b0 ;
  assign n8003 = n3507 & ~n8002 ;
  assign n8004 = n4097 ^ n1847 ^ x161 ;
  assign n8005 = ~n1574 & n8004 ;
  assign n8006 = n1958 & ~n8005 ;
  assign n8007 = ~n5072 & n8006 ;
  assign n8008 = n8007 ^ n421 ^ 1'b0 ;
  assign n8009 = n3689 ^ n1742 ^ 1'b0 ;
  assign n8011 = n1310 & ~n1438 ;
  assign n8012 = n8011 ^ n6462 ^ 1'b0 ;
  assign n8010 = n4008 & ~n7769 ;
  assign n8013 = n8012 ^ n8010 ^ 1'b0 ;
  assign n8014 = x169 & n5006 ;
  assign n8015 = n8014 ^ n2854 ^ 1'b0 ;
  assign n8016 = n8013 | n8015 ;
  assign n8017 = n8016 ^ x121 ^ 1'b0 ;
  assign n8018 = x96 & ~n8017 ;
  assign n8021 = n6165 ^ n655 ^ n559 ;
  assign n8022 = ( ~n462 & n5283 ) | ( ~n462 & n8021 ) | ( n5283 & n8021 ) ;
  assign n8019 = n3905 & n5674 ;
  assign n8020 = n3424 & n8019 ;
  assign n8023 = n8022 ^ n8020 ^ 1'b0 ;
  assign n8026 = ( x81 & n1707 ) | ( x81 & n2718 ) | ( n1707 & n2718 ) ;
  assign n8024 = n3069 ^ n891 ^ 1'b0 ;
  assign n8025 = ( n1372 & n5586 ) | ( n1372 & ~n8024 ) | ( n5586 & ~n8024 ) ;
  assign n8027 = n8026 ^ n8025 ^ 1'b0 ;
  assign n8028 = n3329 ^ n2155 ^ 1'b0 ;
  assign n8029 = ( ~n591 & n4446 ) | ( ~n591 & n8028 ) | ( n4446 & n8028 ) ;
  assign n8030 = x128 | n740 ;
  assign n8031 = n2379 | n8030 ;
  assign n8032 = n8029 | n8031 ;
  assign n8033 = n1160 ^ x211 ^ 1'b0 ;
  assign n8034 = n1285 & n8033 ;
  assign n8035 = n1399 & ~n4667 ;
  assign n8036 = n8035 ^ n518 ^ 1'b0 ;
  assign n8037 = ~n7606 & n8036 ;
  assign n8038 = n8037 ^ n2590 ^ 1'b0 ;
  assign n8039 = n5317 & n8038 ;
  assign n8040 = n8039 ^ n273 ^ 1'b0 ;
  assign n8041 = n6448 | n8040 ;
  assign n8042 = ( x229 & n5219 ) | ( x229 & ~n8041 ) | ( n5219 & ~n8041 ) ;
  assign n8043 = n444 & n1965 ;
  assign n8044 = n8043 ^ n3166 ^ 1'b0 ;
  assign n8045 = n5905 & n8044 ;
  assign n8047 = n1484 & n5106 ;
  assign n8046 = ( n921 & ~n2711 ) | ( n921 & n7836 ) | ( ~n2711 & n7836 ) ;
  assign n8048 = n8047 ^ n8046 ^ n515 ;
  assign n8049 = ( n2319 & n5609 ) | ( n2319 & ~n7582 ) | ( n5609 & ~n7582 ) ;
  assign n8050 = n6032 ^ n1374 ^ x14 ;
  assign n8051 = n6960 & n7232 ;
  assign n8052 = ( n961 & n4847 ) | ( n961 & ~n8051 ) | ( n4847 & ~n8051 ) ;
  assign n8053 = n8050 | n8052 ;
  assign n8054 = n8053 ^ n7548 ^ 1'b0 ;
  assign n8055 = n824 & ~n3215 ;
  assign n8056 = n8055 ^ n2665 ^ 1'b0 ;
  assign n8057 = ~n1349 & n6725 ;
  assign n8058 = n3213 ^ n1394 ^ 1'b0 ;
  assign n8059 = ~n8057 & n8058 ;
  assign n8060 = ~n8056 & n8059 ;
  assign n8061 = ~n7069 & n8060 ;
  assign n8062 = ( n2874 & n3613 ) | ( n2874 & n7284 ) | ( n3613 & n7284 ) ;
  assign n8063 = n8062 ^ n6123 ^ 1'b0 ;
  assign n8064 = n3507 & ~n5063 ;
  assign n8065 = n8064 ^ n2280 ^ 1'b0 ;
  assign n8066 = ~n6441 & n7006 ;
  assign n8067 = n4493 ^ n4347 ^ 1'b0 ;
  assign n8068 = ( n542 & n7978 ) | ( n542 & n8067 ) | ( n7978 & n8067 ) ;
  assign n8069 = ~n1091 & n3015 ;
  assign n8070 = n2852 & n8069 ;
  assign n8071 = n8070 ^ n3570 ^ 1'b0 ;
  assign n8072 = n1534 & n1536 ;
  assign n8073 = n8072 ^ n4378 ^ 1'b0 ;
  assign n8074 = n6442 ^ n1094 ^ 1'b0 ;
  assign n8075 = n8074 ^ n4891 ^ n2403 ;
  assign n8076 = n8075 ^ n4237 ^ 1'b0 ;
  assign n8077 = ( n861 & n8073 ) | ( n861 & n8076 ) | ( n8073 & n8076 ) ;
  assign n8078 = n5931 ^ n1189 ^ n1156 ;
  assign n8079 = ( n1937 & n4009 ) | ( n1937 & ~n7943 ) | ( n4009 & ~n7943 ) ;
  assign n8083 = n3519 ^ n3410 ^ n2295 ;
  assign n8080 = n1126 ^ n1086 ^ 1'b0 ;
  assign n8081 = n5676 & ~n8080 ;
  assign n8082 = n3342 | n8081 ;
  assign n8084 = n8083 ^ n8082 ^ 1'b0 ;
  assign n8085 = n3762 & n8084 ;
  assign n8086 = ~n4280 & n8072 ;
  assign n8087 = n943 | n2802 ;
  assign n8088 = n3196 | n8087 ;
  assign n8089 = ( ~n3932 & n5233 ) | ( ~n3932 & n8088 ) | ( n5233 & n8088 ) ;
  assign n8090 = n4630 ^ n903 ^ 1'b0 ;
  assign n8091 = ~n6389 & n8090 ;
  assign n8092 = n2321 & ~n2370 ;
  assign n8093 = n7419 ^ n3375 ^ n1447 ;
  assign n8094 = n3980 ^ n2842 ^ 1'b0 ;
  assign n8095 = ~n3694 & n7885 ;
  assign n8096 = n741 & n8095 ;
  assign n8097 = n516 & ~n4190 ;
  assign n8098 = ~n4760 & n8097 ;
  assign n8099 = n8098 ^ n5382 ^ 1'b0 ;
  assign n8100 = ( x206 & ~n1696 ) | ( x206 & n3344 ) | ( ~n1696 & n3344 ) ;
  assign n8101 = ~n3237 & n8100 ;
  assign n8102 = n1968 ^ n1435 ^ n785 ;
  assign n8103 = n1200 & n7088 ;
  assign n8104 = ~n7397 & n8103 ;
  assign n8105 = ( n3990 & n4378 ) | ( n3990 & n4458 ) | ( n4378 & n4458 ) ;
  assign n8106 = n4604 & ~n8105 ;
  assign n8107 = ( ~n2680 & n8104 ) | ( ~n2680 & n8106 ) | ( n8104 & n8106 ) ;
  assign n8108 = n8102 | n8107 ;
  assign n8109 = n6663 ^ n5588 ^ 1'b0 ;
  assign n8110 = n4644 | n8109 ;
  assign n8111 = n8110 ^ n741 ^ 1'b0 ;
  assign n8114 = n891 ^ n706 ^ 1'b0 ;
  assign n8115 = n3553 & ~n8114 ;
  assign n8116 = n8115 ^ n8036 ^ 1'b0 ;
  assign n8112 = n2735 ^ n2676 ^ n277 ;
  assign n8113 = n7739 & ~n8112 ;
  assign n8117 = n8116 ^ n8113 ^ 1'b0 ;
  assign n8118 = ~n1541 & n6054 ;
  assign n8119 = n8118 ^ n1174 ^ 1'b0 ;
  assign n8120 = n7108 ^ n5746 ^ n2509 ;
  assign n8121 = n2458 ^ n1113 ^ 1'b0 ;
  assign n8122 = n1615 | n2301 ;
  assign n8123 = ~n4369 & n8122 ;
  assign n8124 = n8123 ^ n2491 ^ 1'b0 ;
  assign n8125 = n2078 | n8124 ;
  assign n8126 = n412 & ~n2893 ;
  assign n8127 = ~n4631 & n8126 ;
  assign n8128 = n1860 ^ n1805 ^ n989 ;
  assign n8129 = ( ~n2538 & n8127 ) | ( ~n2538 & n8128 ) | ( n8127 & n8128 ) ;
  assign n8130 = ( ~x138 & n1281 ) | ( ~x138 & n4438 ) | ( n1281 & n4438 ) ;
  assign n8131 = n8129 | n8130 ;
  assign n8132 = n8131 ^ n6298 ^ 1'b0 ;
  assign n8133 = n8132 ^ n4755 ^ 1'b0 ;
  assign n8134 = n8125 | n8133 ;
  assign n8135 = n6337 ^ n3237 ^ n2494 ;
  assign n8136 = n8135 ^ n717 ^ 1'b0 ;
  assign n8137 = n2465 | n8136 ;
  assign n8140 = n2433 ^ n2025 ^ 1'b0 ;
  assign n8138 = ~n1593 & n4029 ;
  assign n8139 = ( ~n2429 & n3763 ) | ( ~n2429 & n8138 ) | ( n3763 & n8138 ) ;
  assign n8141 = n8140 ^ n8139 ^ 1'b0 ;
  assign n8142 = ~n8137 & n8141 ;
  assign n8143 = n5021 ^ n4589 ^ n3428 ;
  assign n8144 = n704 & ~n8143 ;
  assign n8145 = x91 | n4364 ;
  assign n8146 = n5328 & ~n8145 ;
  assign n8147 = x48 & ~n3931 ;
  assign n8148 = n8147 ^ n5694 ^ 1'b0 ;
  assign n8152 = x234 & ~n3385 ;
  assign n8153 = n8152 ^ n5264 ^ 1'b0 ;
  assign n8154 = n2671 & n8153 ;
  assign n8155 = ~n1718 & n8154 ;
  assign n8156 = n2407 & ~n8155 ;
  assign n8157 = n2255 & n8156 ;
  assign n8149 = ( ~x26 & n2121 ) | ( ~x26 & n2523 ) | ( n2121 & n2523 ) ;
  assign n8150 = n8149 ^ n3305 ^ n1081 ;
  assign n8151 = x230 | n8150 ;
  assign n8158 = n8157 ^ n8151 ^ n6102 ;
  assign n8159 = n3239 | n8158 ;
  assign n8160 = n4464 ^ n3585 ^ n1326 ;
  assign n8161 = n3404 & n8160 ;
  assign n8167 = n3234 | n5323 ;
  assign n8168 = ( ~x58 & n2003 ) | ( ~x58 & n8167 ) | ( n2003 & n8167 ) ;
  assign n8162 = x186 & ~n410 ;
  assign n8163 = n8162 ^ n363 ^ 1'b0 ;
  assign n8164 = x148 & ~n2615 ;
  assign n8165 = ( ~n2927 & n8163 ) | ( ~n2927 & n8164 ) | ( n8163 & n8164 ) ;
  assign n8166 = ~n4104 & n8165 ;
  assign n8169 = n8168 ^ n8166 ^ 1'b0 ;
  assign n8170 = n584 ^ x121 ^ 1'b0 ;
  assign n8171 = n5684 ^ n3774 ^ 1'b0 ;
  assign n8172 = n8171 ^ n3160 ^ 1'b0 ;
  assign n8173 = ( n2594 & n7665 ) | ( n2594 & ~n8172 ) | ( n7665 & ~n8172 ) ;
  assign n8174 = ~n1881 & n4080 ;
  assign n8175 = n3866 & n8174 ;
  assign n8176 = ~n1128 & n7664 ;
  assign n8177 = n8175 & n8176 ;
  assign n8178 = ~n325 & n1553 ;
  assign n8179 = ~x253 & n8178 ;
  assign n8180 = n8179 ^ x110 ^ 1'b0 ;
  assign n8181 = n3649 & ~n4105 ;
  assign n8182 = n3508 & ~n8181 ;
  assign n8183 = n2333 | n8182 ;
  assign n8184 = n8183 ^ n4784 ^ 1'b0 ;
  assign n8185 = n1104 & n8184 ;
  assign n8186 = ~n8180 & n8185 ;
  assign n8188 = n3868 ^ n3404 ^ n567 ;
  assign n8187 = n5436 ^ n3934 ^ n3316 ;
  assign n8189 = n8188 ^ n8187 ^ n7040 ;
  assign n8190 = n1895 & ~n7425 ;
  assign n8191 = ~x81 & n8190 ;
  assign n8193 = n3826 & ~n8073 ;
  assign n8192 = n7560 ^ n4089 ^ n2695 ;
  assign n8194 = n8193 ^ n8192 ^ 1'b0 ;
  assign n8195 = n8194 ^ n7333 ^ 1'b0 ;
  assign n8196 = ~n8191 & n8195 ;
  assign n8197 = ( ~n1026 & n3100 ) | ( ~n1026 & n6123 ) | ( n3100 & n6123 ) ;
  assign n8198 = ( n2058 & ~n2118 ) | ( n2058 & n3387 ) | ( ~n2118 & n3387 ) ;
  assign n8199 = n6082 ^ n1951 ^ 1'b0 ;
  assign n8200 = n8198 & n8199 ;
  assign n8201 = n2306 ^ n1068 ^ 1'b0 ;
  assign n8202 = n909 & n3321 ;
  assign n8203 = n5276 ^ n1432 ^ 1'b0 ;
  assign n8204 = n913 | n8203 ;
  assign n8205 = n8202 | n8204 ;
  assign n8206 = n8205 ^ x194 ^ 1'b0 ;
  assign n8207 = n3133 & n8206 ;
  assign n8208 = n7172 ^ n1103 ^ 1'b0 ;
  assign n8209 = n1567 | n8208 ;
  assign n8210 = ~n275 & n907 ;
  assign n8211 = n8210 ^ n4469 ^ 1'b0 ;
  assign n8212 = ( n4370 & ~n4381 ) | ( n4370 & n8211 ) | ( ~n4381 & n8211 ) ;
  assign n8213 = n476 ^ x97 ^ 1'b0 ;
  assign n8214 = ~n3046 & n8213 ;
  assign n8215 = n464 | n8214 ;
  assign n8216 = n1571 & ~n8215 ;
  assign n8217 = n8216 ^ n7389 ^ 1'b0 ;
  assign n8218 = n1527 & ~n8217 ;
  assign n8219 = n8218 ^ n691 ^ 1'b0 ;
  assign n8220 = n3199 ^ n974 ^ 1'b0 ;
  assign n8221 = n5681 & n8220 ;
  assign n8222 = ( n863 & n8219 ) | ( n863 & n8221 ) | ( n8219 & n8221 ) ;
  assign n8223 = ( n8209 & ~n8212 ) | ( n8209 & n8222 ) | ( ~n8212 & n8222 ) ;
  assign n8224 = ~n667 & n8223 ;
  assign n8225 = n6990 & n8224 ;
  assign n8226 = n8207 & ~n8225 ;
  assign n8227 = n8201 & n8226 ;
  assign n8228 = ( ~x224 & n2504 ) | ( ~x224 & n2531 ) | ( n2504 & n2531 ) ;
  assign n8229 = n2523 | n8228 ;
  assign n8230 = n8229 ^ n2186 ^ 1'b0 ;
  assign n8231 = n5115 & n8230 ;
  assign n8232 = n8231 ^ n2611 ^ 1'b0 ;
  assign n8233 = ~n4652 & n8232 ;
  assign n8234 = n2286 | n8233 ;
  assign n8235 = n1039 ^ n856 ^ 1'b0 ;
  assign n8236 = n1617 & ~n4067 ;
  assign n8237 = n8098 & n8236 ;
  assign n8241 = n3676 ^ n3155 ^ 1'b0 ;
  assign n8242 = n8175 | n8241 ;
  assign n8238 = n5705 ^ x206 ^ 1'b0 ;
  assign n8239 = x238 & ~n8238 ;
  assign n8240 = n5752 & ~n8239 ;
  assign n8243 = n8242 ^ n8240 ^ 1'b0 ;
  assign n8244 = x184 ^ x169 ^ 1'b0 ;
  assign n8245 = n8244 ^ n986 ^ 1'b0 ;
  assign n8246 = n5692 & ~n8245 ;
  assign n8247 = n3759 ^ n3516 ^ n2315 ;
  assign n8248 = n3736 | n7417 ;
  assign n8249 = n8248 ^ n6865 ^ n5408 ;
  assign n8250 = n2708 | n3172 ;
  assign n8251 = n1814 | n3053 ;
  assign n8252 = n1378 | n8251 ;
  assign n8254 = n3883 | n6693 ;
  assign n8253 = n2670 & n3464 ;
  assign n8255 = n8254 ^ n8253 ^ 1'b0 ;
  assign n8256 = n1329 ^ x182 ^ 1'b0 ;
  assign n8257 = n5646 ^ n4698 ^ n673 ;
  assign n8258 = n3066 ^ n375 ^ 1'b0 ;
  assign n8259 = n8258 ^ n2174 ^ 1'b0 ;
  assign n8271 = n1950 ^ n1495 ^ n1482 ;
  assign n8263 = n861 & n2405 ;
  assign n8260 = n3605 | n6848 ;
  assign n8261 = ~x77 & n3955 ;
  assign n8262 = n8260 | n8261 ;
  assign n8264 = n8263 ^ n8262 ^ 1'b0 ;
  assign n8265 = n4007 | n5429 ;
  assign n8266 = n8264 & ~n8265 ;
  assign n8267 = n1624 | n2879 ;
  assign n8268 = n8267 ^ n2406 ^ 1'b0 ;
  assign n8269 = n8268 ^ n1412 ^ 1'b0 ;
  assign n8270 = ~n8266 & n8269 ;
  assign n8272 = n8271 ^ n8270 ^ 1'b0 ;
  assign n8273 = n3944 ^ n3776 ^ n3578 ;
  assign n8274 = n1862 & ~n5627 ;
  assign n8275 = n5569 & n8274 ;
  assign n8276 = n8167 ^ x21 ^ 1'b0 ;
  assign n8277 = n2889 ^ n2671 ^ 1'b0 ;
  assign n8278 = n8277 ^ n7317 ^ n2223 ;
  assign n8279 = ( n5875 & ~n7411 ) | ( n5875 & n8278 ) | ( ~n7411 & n8278 ) ;
  assign n8280 = n8279 ^ n3568 ^ n1322 ;
  assign n8281 = n8012 ^ n4274 ^ n426 ;
  assign n8282 = n4144 & ~n8281 ;
  assign n8283 = n7496 ^ n3541 ^ 1'b0 ;
  assign n8284 = n1928 & n8283 ;
  assign n8285 = n1126 | n2518 ;
  assign n8286 = n682 | n8285 ;
  assign n8287 = n2325 & ~n8286 ;
  assign n8288 = n4961 ^ x124 ^ 1'b0 ;
  assign n8289 = n2250 | n5636 ;
  assign n8290 = n8289 ^ n3631 ^ 1'b0 ;
  assign n8291 = n2884 & ~n4510 ;
  assign n8292 = n2284 & n8291 ;
  assign n8293 = ~n500 & n8292 ;
  assign n8294 = n8293 ^ n2293 ^ 1'b0 ;
  assign n8295 = ~n1545 & n6678 ;
  assign n8300 = n1339 | n7053 ;
  assign n8296 = n4020 ^ n2889 ^ 1'b0 ;
  assign n8297 = n1487 | n8296 ;
  assign n8298 = n5732 & ~n8297 ;
  assign n8299 = n8298 ^ n3639 ^ n3567 ;
  assign n8301 = n8300 ^ n8299 ^ n512 ;
  assign n8302 = ( n515 & n953 ) | ( n515 & n8036 ) | ( n953 & n8036 ) ;
  assign n8303 = n6629 ^ n3639 ^ 1'b0 ;
  assign n8304 = ~n368 & n8303 ;
  assign n8305 = ~n8302 & n8304 ;
  assign n8306 = n7805 ^ n4958 ^ 1'b0 ;
  assign n8307 = n2048 ^ n1760 ^ 1'b0 ;
  assign n8308 = n8307 ^ n1684 ^ 1'b0 ;
  assign n8309 = ~n5436 & n8308 ;
  assign n8310 = ( n2447 & n7934 ) | ( n2447 & n8309 ) | ( n7934 & n8309 ) ;
  assign n8311 = n423 | n651 ;
  assign n8312 = n8311 ^ n2827 ^ 1'b0 ;
  assign n8317 = ( x24 & n2106 ) | ( x24 & n3110 ) | ( n2106 & n3110 ) ;
  assign n8313 = n3105 ^ x179 ^ 1'b0 ;
  assign n8314 = n6514 | n8313 ;
  assign n8315 = n8314 ^ n3227 ^ n1054 ;
  assign n8316 = n8315 ^ n6363 ^ 1'b0 ;
  assign n8318 = n8317 ^ n8316 ^ n3049 ;
  assign n8319 = ( n351 & n3418 ) | ( n351 & n3936 ) | ( n3418 & n3936 ) ;
  assign n8320 = ~n2790 & n8319 ;
  assign n8321 = n7046 & n8320 ;
  assign n8322 = n8138 ^ n5882 ^ 1'b0 ;
  assign n8323 = n8165 & ~n8322 ;
  assign n8324 = n4595 & ~n4824 ;
  assign n8325 = n8324 ^ n6546 ^ 1'b0 ;
  assign n8326 = n7182 ^ n7047 ^ 1'b0 ;
  assign n8327 = n382 & n8326 ;
  assign n8328 = n6068 ^ n3165 ^ 1'b0 ;
  assign n8329 = n8328 ^ n4210 ^ 1'b0 ;
  assign n8330 = n8329 ^ n2229 ^ 1'b0 ;
  assign n8331 = n8327 & ~n8330 ;
  assign n8338 = n2150 & n3804 ;
  assign n8333 = n3803 ^ x8 ^ 1'b0 ;
  assign n8334 = n5066 ^ n2435 ^ 1'b0 ;
  assign n8335 = n1912 | n8334 ;
  assign n8336 = n8333 & ~n8335 ;
  assign n8337 = n8336 ^ n6643 ^ 1'b0 ;
  assign n8332 = ~n2842 & n6031 ;
  assign n8339 = n8338 ^ n8337 ^ n8332 ;
  assign n8340 = n2441 & ~n5191 ;
  assign n8341 = ( n904 & ~n5002 ) | ( n904 & n8340 ) | ( ~n5002 & n8340 ) ;
  assign n8342 = n3758 ^ n958 ^ 1'b0 ;
  assign n8343 = ~n6385 & n8342 ;
  assign n8344 = n559 & ~n2185 ;
  assign n8345 = n1971 & n8344 ;
  assign n8346 = ~n282 & n8345 ;
  assign n8347 = ~n4520 & n8346 ;
  assign n8348 = n8347 ^ n4480 ^ 1'b0 ;
  assign n8349 = x215 & n8199 ;
  assign n8350 = ~n7190 & n8349 ;
  assign n8351 = n4060 ^ n3547 ^ n2317 ;
  assign n8352 = ~n1144 & n7741 ;
  assign n8356 = n7127 ^ n3892 ^ n619 ;
  assign n8353 = n3364 | n4282 ;
  assign n8354 = n405 | n8353 ;
  assign n8355 = n8354 ^ n3853 ^ n1749 ;
  assign n8357 = n8356 ^ n8355 ^ n2411 ;
  assign n8358 = ( n5388 & n8352 ) | ( n5388 & ~n8357 ) | ( n8352 & ~n8357 ) ;
  assign n8359 = n5104 | n7456 ;
  assign n8360 = n8359 ^ n1741 ^ 1'b0 ;
  assign n8361 = n4334 ^ n2589 ^ 1'b0 ;
  assign n8362 = n5078 ^ n4197 ^ n2106 ;
  assign n8363 = n4668 ^ n2390 ^ n2216 ;
  assign n8364 = ( ~n2179 & n5926 ) | ( ~n2179 & n8363 ) | ( n5926 & n8363 ) ;
  assign n8365 = ( n1622 & n5424 ) | ( n1622 & n6777 ) | ( n5424 & n6777 ) ;
  assign n8366 = n1671 | n8365 ;
  assign n8367 = n8366 ^ n8253 ^ 1'b0 ;
  assign n8368 = n1010 & n3507 ;
  assign n8369 = n3009 & ~n4635 ;
  assign n8370 = n8368 & n8369 ;
  assign n8371 = ~n2338 & n2367 ;
  assign n8372 = n5732 & n8371 ;
  assign n8373 = n5775 | n8372 ;
  assign n8374 = n2603 | n8373 ;
  assign n8375 = n2105 ^ n1821 ^ n1262 ;
  assign n8376 = n754 | n8375 ;
  assign n8377 = n2396 | n4293 ;
  assign n8378 = ( n3069 & n8376 ) | ( n3069 & n8377 ) | ( n8376 & n8377 ) ;
  assign n8379 = n4773 & n8378 ;
  assign n8380 = ~n8374 & n8379 ;
  assign n8385 = n5586 ^ n457 ^ 1'b0 ;
  assign n8386 = n587 | n8385 ;
  assign n8387 = n8386 ^ n991 ^ 1'b0 ;
  assign n8388 = n3260 | n8387 ;
  assign n8381 = n4766 & ~n7562 ;
  assign n8382 = n2172 ^ n1923 ^ 1'b0 ;
  assign n8383 = n8382 ^ n2764 ^ 1'b0 ;
  assign n8384 = n8381 & n8383 ;
  assign n8389 = n8388 ^ n8384 ^ n3024 ;
  assign n8390 = n368 | n8114 ;
  assign n8391 = x109 & ~n3113 ;
  assign n8392 = n2317 & n8391 ;
  assign n8393 = n341 & n8392 ;
  assign n8394 = ( n1715 & n3007 ) | ( n1715 & n3640 ) | ( n3007 & n3640 ) ;
  assign n8395 = n3412 & n5308 ;
  assign n8396 = n8395 ^ n2888 ^ 1'b0 ;
  assign n8397 = n426 | n1370 ;
  assign n8398 = n8397 ^ n854 ^ 1'b0 ;
  assign n8399 = ( n1111 & n2964 ) | ( n1111 & n8398 ) | ( n2964 & n8398 ) ;
  assign n8400 = n1893 | n8399 ;
  assign n8401 = n8400 ^ n2130 ^ 1'b0 ;
  assign n8402 = ~n4388 & n7243 ;
  assign n8403 = ~n4083 & n8402 ;
  assign n8404 = n5586 ^ n1820 ^ n747 ;
  assign n8405 = n3267 & ~n8404 ;
  assign n8406 = n8405 ^ n3632 ^ 1'b0 ;
  assign n8407 = n8406 ^ n1718 ^ 1'b0 ;
  assign n8408 = n4151 & n8251 ;
  assign n8409 = n2191 & n8408 ;
  assign n8410 = n4041 | n8409 ;
  assign n8411 = n8407 & ~n8410 ;
  assign n8412 = ( n6436 & n8403 ) | ( n6436 & n8411 ) | ( n8403 & n8411 ) ;
  assign n8428 = n3581 ^ n2734 ^ 1'b0 ;
  assign n8429 = n8428 ^ n5648 ^ n4447 ;
  assign n8414 = n810 | n3231 ;
  assign n8415 = x96 | n8414 ;
  assign n8413 = n720 | n6032 ;
  assign n8416 = n8415 ^ n8413 ^ 1'b0 ;
  assign n8417 = n8416 ^ n5883 ^ 1'b0 ;
  assign n8418 = n3368 | n8417 ;
  assign n8419 = n8418 ^ n3440 ^ 1'b0 ;
  assign n8420 = ( n4045 & n5859 ) | ( n4045 & n8419 ) | ( n5859 & n8419 ) ;
  assign n8421 = n1149 & ~n2489 ;
  assign n8422 = n8421 ^ n2466 ^ 1'b0 ;
  assign n8423 = n6480 ^ n5031 ^ 1'b0 ;
  assign n8424 = n8422 & ~n8423 ;
  assign n8425 = ~n8420 & n8424 ;
  assign n8426 = n3436 & n8425 ;
  assign n8427 = n1500 & ~n8426 ;
  assign n8430 = n8429 ^ n8427 ^ 1'b0 ;
  assign n8431 = n515 ^ n344 ^ 1'b0 ;
  assign n8432 = ( ~n2706 & n3406 ) | ( ~n2706 & n6018 ) | ( n3406 & n6018 ) ;
  assign n8433 = ( n3113 & ~n3645 ) | ( n3113 & n8432 ) | ( ~n3645 & n8432 ) ;
  assign n8434 = n8431 & ~n8433 ;
  assign n8435 = n8434 ^ n4965 ^ 1'b0 ;
  assign n8436 = n1108 | n1151 ;
  assign n8437 = n8436 ^ n1046 ^ 1'b0 ;
  assign n8438 = ( n5049 & n7653 ) | ( n5049 & ~n8437 ) | ( n7653 & ~n8437 ) ;
  assign n8439 = ( n2901 & ~n4305 ) | ( n2901 & n8438 ) | ( ~n4305 & n8438 ) ;
  assign n8440 = n2468 ^ n1521 ^ 1'b0 ;
  assign n8441 = n5327 ^ n2887 ^ 1'b0 ;
  assign n8442 = n5456 & ~n8441 ;
  assign n8443 = x49 ^ x10 ^ 1'b0 ;
  assign n8444 = ~n2085 & n8443 ;
  assign n8445 = n8442 & n8444 ;
  assign n8446 = ~n8440 & n8445 ;
  assign n8447 = x30 & n8446 ;
  assign n8448 = n1803 & ~n8447 ;
  assign n8449 = n5914 ^ n2734 ^ 1'b0 ;
  assign n8450 = n356 & n4703 ;
  assign n8451 = n8450 ^ n3168 ^ 1'b0 ;
  assign n8452 = ~n1124 & n4428 ;
  assign n8453 = ~n4367 & n8452 ;
  assign n8454 = n8453 ^ n4749 ^ 1'b0 ;
  assign n8455 = n3416 & n8454 ;
  assign n8456 = n8455 ^ n4519 ^ 1'b0 ;
  assign n8457 = n6430 ^ n1294 ^ n1161 ;
  assign n8458 = n4852 | n8457 ;
  assign n8459 = n8006 ^ x147 ^ 1'b0 ;
  assign n8460 = ( n5950 & ~n8458 ) | ( n5950 & n8459 ) | ( ~n8458 & n8459 ) ;
  assign n8461 = n6084 ^ x218 ^ 1'b0 ;
  assign n8463 = n2342 ^ n307 ^ 1'b0 ;
  assign n8464 = n1327 & ~n4583 ;
  assign n8465 = n8463 & n8464 ;
  assign n8466 = n1044 | n8465 ;
  assign n8462 = n686 | n8299 ;
  assign n8467 = n8466 ^ n8462 ^ 1'b0 ;
  assign n8468 = n935 | n1007 ;
  assign n8469 = n7437 ^ n6703 ^ n569 ;
  assign n8470 = n1711 ^ n1118 ^ 1'b0 ;
  assign n8471 = ~n780 & n8470 ;
  assign n8472 = x71 & n1664 ;
  assign n8473 = n2793 & n8472 ;
  assign n8474 = ( n7910 & n8471 ) | ( n7910 & ~n8473 ) | ( n8471 & ~n8473 ) ;
  assign n8475 = ~n1594 & n4904 ;
  assign n8476 = n2938 & n4872 ;
  assign n8477 = ~n5764 & n8476 ;
  assign n8478 = ( ~n493 & n4301 ) | ( ~n493 & n5798 ) | ( n4301 & n5798 ) ;
  assign n8479 = n8478 ^ n7494 ^ 1'b0 ;
  assign n8480 = n8177 | n8479 ;
  assign n8481 = ( n358 & n4441 ) | ( n358 & ~n4528 ) | ( n4441 & ~n4528 ) ;
  assign n8482 = n3576 & n8163 ;
  assign n8483 = ~n7168 & n8482 ;
  assign n8484 = ( n5615 & n8375 ) | ( n5615 & n8483 ) | ( n8375 & n8483 ) ;
  assign n8485 = ~n7499 & n8384 ;
  assign n8486 = ~n6444 & n8485 ;
  assign n8487 = n1264 & n5990 ;
  assign n8488 = n8487 ^ n3662 ^ 1'b0 ;
  assign n8489 = n1324 ^ x63 ^ 1'b0 ;
  assign n8490 = ~n8488 & n8489 ;
  assign n8491 = n8490 ^ n6111 ^ n4670 ;
  assign n8495 = n2534 ^ n809 ^ 1'b0 ;
  assign n8496 = n2966 & n8495 ;
  assign n8497 = ( n415 & n5318 ) | ( n415 & ~n8496 ) | ( n5318 & ~n8496 ) ;
  assign n8492 = n3974 | n5637 ;
  assign n8493 = n4247 | n8492 ;
  assign n8494 = n8493 ^ n2125 ^ 1'b0 ;
  assign n8498 = n8497 ^ n8494 ^ n1557 ;
  assign n8499 = n1558 | n3318 ;
  assign n8500 = n8499 ^ n565 ^ 1'b0 ;
  assign n8501 = n2151 | n8500 ;
  assign n8502 = n8501 ^ n4217 ^ 1'b0 ;
  assign n8503 = ~n8046 & n8502 ;
  assign n8504 = n413 & n8503 ;
  assign n8505 = x224 ^ x15 ^ 1'b0 ;
  assign n8506 = n615 | n8505 ;
  assign n8507 = n1247 | n8506 ;
  assign n8508 = n3732 ^ n3723 ^ n747 ;
  assign n8509 = n8508 ^ n1734 ^ 1'b0 ;
  assign n8510 = x190 & ~n8509 ;
  assign n8511 = n8510 ^ n5872 ^ 1'b0 ;
  assign n8516 = n1680 & n5438 ;
  assign n8517 = ~n4430 & n8516 ;
  assign n8514 = n2929 | n3125 ;
  assign n8515 = n8514 ^ n820 ^ 1'b0 ;
  assign n8518 = n8517 ^ n8515 ^ 1'b0 ;
  assign n8519 = ~n4996 & n8518 ;
  assign n8512 = ( x239 & n2169 ) | ( x239 & n4228 ) | ( n2169 & n4228 ) ;
  assign n8513 = ~n7376 & n8512 ;
  assign n8520 = n8519 ^ n8513 ^ 1'b0 ;
  assign n8521 = n6574 ^ n4855 ^ 1'b0 ;
  assign n8522 = n4792 ^ n3566 ^ 1'b0 ;
  assign n8523 = n7078 | n8522 ;
  assign n8524 = ~n3979 & n8523 ;
  assign n8525 = n1893 & ~n2487 ;
  assign n8526 = n3403 ^ n2209 ^ 1'b0 ;
  assign n8527 = n8526 ^ n3580 ^ 1'b0 ;
  assign n8530 = n668 ^ x76 ^ 1'b0 ;
  assign n8531 = n1613 & ~n8530 ;
  assign n8528 = ( n461 & n885 ) | ( n461 & n1851 ) | ( n885 & n1851 ) ;
  assign n8529 = ( n1791 & n5382 ) | ( n1791 & ~n8528 ) | ( n5382 & ~n8528 ) ;
  assign n8532 = n8531 ^ n8529 ^ n3658 ;
  assign n8533 = ( n1140 & n1786 ) | ( n1140 & ~n3763 ) | ( n1786 & ~n3763 ) ;
  assign n8534 = n8533 ^ n8362 ^ 1'b0 ;
  assign n8539 = n5473 ^ n5246 ^ n586 ;
  assign n8535 = n920 | n2032 ;
  assign n8536 = n6316 & ~n8535 ;
  assign n8537 = n8536 ^ n1231 ^ x86 ;
  assign n8538 = n3881 & n8537 ;
  assign n8540 = n8539 ^ n8538 ^ 1'b0 ;
  assign n8541 = n829 | n7520 ;
  assign n8542 = ( n4693 & n4988 ) | ( n4693 & ~n6228 ) | ( n4988 & ~n6228 ) ;
  assign n8543 = n8541 & n8542 ;
  assign n8544 = n5848 ^ x243 ^ 1'b0 ;
  assign n8545 = n3088 & ~n7629 ;
  assign n8547 = ~n377 & n3086 ;
  assign n8548 = ~n4249 & n8547 ;
  assign n8549 = n8548 ^ n6627 ^ 1'b0 ;
  assign n8550 = n2401 & ~n8549 ;
  assign n8546 = n4791 ^ n4385 ^ 1'b0 ;
  assign n8551 = n8550 ^ n8546 ^ 1'b0 ;
  assign n8552 = n8551 ^ n2808 ^ n1650 ;
  assign n8558 = ( n5648 & n6661 ) | ( n5648 & n8260 ) | ( n6661 & n8260 ) ;
  assign n8554 = ~n525 & n1916 ;
  assign n8553 = ~n287 & n5009 ;
  assign n8555 = n8554 ^ n8553 ^ 1'b0 ;
  assign n8556 = n6496 & n8555 ;
  assign n8557 = x114 & n8556 ;
  assign n8559 = n8558 ^ n8557 ^ 1'b0 ;
  assign n8560 = n1831 ^ x203 ^ 1'b0 ;
  assign n8561 = n1209 | n8560 ;
  assign n8562 = n6856 & ~n8155 ;
  assign n8563 = n8561 & n8562 ;
  assign n8564 = n310 | n576 ;
  assign n8565 = n363 & ~n8564 ;
  assign n8566 = n4305 ^ n2481 ^ 1'b0 ;
  assign n8567 = ~n8565 & n8566 ;
  assign n8568 = n591 & ~n3125 ;
  assign n8569 = n8568 ^ n703 ^ 1'b0 ;
  assign n8570 = n7549 ^ n4807 ^ 1'b0 ;
  assign n8571 = n8569 & n8570 ;
  assign n8572 = ( n337 & n1583 ) | ( n337 & n8311 ) | ( n1583 & n8311 ) ;
  assign n8573 = n990 & ~n8572 ;
  assign n8574 = n5475 ^ n2511 ^ 1'b0 ;
  assign n8575 = n903 | n8574 ;
  assign n8576 = n3283 ^ n2406 ^ n1541 ;
  assign n8577 = n8576 ^ n927 ^ 1'b0 ;
  assign n8578 = ~n8575 & n8577 ;
  assign n8579 = n7741 ^ n1944 ^ 1'b0 ;
  assign n8580 = n6399 & n8579 ;
  assign n8581 = n8580 ^ n3599 ^ 1'b0 ;
  assign n8582 = n7917 & n8581 ;
  assign n8583 = n3156 & n8582 ;
  assign n8584 = n7805 & n8583 ;
  assign n8585 = n2986 & n4985 ;
  assign n8586 = n7186 ^ n5207 ^ 1'b0 ;
  assign n8587 = ~n4048 & n8586 ;
  assign n8588 = n8587 ^ n5078 ^ n3361 ;
  assign n8589 = n3982 ^ n874 ^ 1'b0 ;
  assign n8590 = ~n4475 & n8589 ;
  assign n8591 = n8588 & n8590 ;
  assign n8592 = x106 & n1584 ;
  assign n8593 = n8592 ^ n2167 ^ 1'b0 ;
  assign n8594 = n5964 ^ n4027 ^ 1'b0 ;
  assign n8595 = n8593 | n8594 ;
  assign n8596 = n1392 | n4720 ;
  assign n8597 = n4592 & ~n8596 ;
  assign n8598 = ( n4180 & ~n8595 ) | ( n4180 & n8597 ) | ( ~n8595 & n8597 ) ;
  assign n8599 = n7403 & ~n8598 ;
  assign n8600 = ~n5918 & n8599 ;
  assign n8601 = n3698 & n8600 ;
  assign n8610 = ~n2889 & n4804 ;
  assign n8611 = n8610 ^ n7586 ^ 1'b0 ;
  assign n8612 = n8611 ^ n1168 ^ 1'b0 ;
  assign n8607 = n7099 ^ n4982 ^ 1'b0 ;
  assign n8608 = n6841 & ~n8607 ;
  assign n8606 = n6316 ^ n6062 ^ n663 ;
  assign n8609 = n8608 ^ n8606 ^ n4343 ;
  assign n8604 = n6777 & n7393 ;
  assign n8602 = ~n4114 & n7548 ;
  assign n8603 = n8602 ^ n5262 ^ 1'b0 ;
  assign n8605 = n8604 ^ n8603 ^ 1'b0 ;
  assign n8613 = n8612 ^ n8609 ^ n8605 ;
  assign n8615 = n2425 | n2546 ;
  assign n8616 = n509 & ~n8615 ;
  assign n8614 = ( n789 & n1817 ) | ( n789 & n5264 ) | ( n1817 & n5264 ) ;
  assign n8617 = n8616 ^ n8614 ^ 1'b0 ;
  assign n8618 = ~n1258 & n8617 ;
  assign n8619 = n4258 & n8618 ;
  assign n8620 = n8619 ^ n841 ^ 1'b0 ;
  assign n8622 = n519 | n7058 ;
  assign n8621 = n2006 & n4242 ;
  assign n8623 = n8622 ^ n8621 ^ 1'b0 ;
  assign n8624 = n8623 ^ n584 ^ 1'b0 ;
  assign n8625 = n6783 ^ n5694 ^ 1'b0 ;
  assign n8626 = n1312 & ~n8625 ;
  assign n8627 = ( n1741 & n3854 ) | ( n1741 & ~n8626 ) | ( n3854 & ~n8626 ) ;
  assign n8628 = n5298 & ~n8627 ;
  assign n8629 = n8628 ^ n8231 ^ 1'b0 ;
  assign n8630 = ( n2236 & ~n4561 ) | ( n2236 & n6494 ) | ( ~n4561 & n6494 ) ;
  assign n8631 = n5439 | n8630 ;
  assign n8632 = n3403 ^ x218 ^ 1'b0 ;
  assign n8633 = n8632 ^ n4229 ^ n4162 ;
  assign n8634 = ~n401 & n8633 ;
  assign n8636 = x190 & ~n3638 ;
  assign n8637 = n8636 ^ n4761 ^ 1'b0 ;
  assign n8638 = n4395 & n8637 ;
  assign n8635 = n2836 | n3945 ;
  assign n8639 = n8638 ^ n8635 ^ 1'b0 ;
  assign n8640 = n7046 ^ n4363 ^ n1527 ;
  assign n8641 = n3400 ^ n3091 ^ 1'b0 ;
  assign n8642 = n8641 ^ n6406 ^ 1'b0 ;
  assign n8643 = n5230 ^ n3557 ^ x207 ;
  assign n8644 = ( n4809 & n6084 ) | ( n4809 & ~n8643 ) | ( n6084 & ~n8643 ) ;
  assign n8645 = n7965 & n7990 ;
  assign n8646 = ~n8644 & n8645 ;
  assign n8649 = ~n1365 & n3590 ;
  assign n8650 = n8649 ^ n547 ^ 1'b0 ;
  assign n8647 = ( x200 & ~n4457 ) | ( x200 & n5580 ) | ( ~n4457 & n5580 ) ;
  assign n8648 = ~n7936 & n8647 ;
  assign n8651 = n8650 ^ n8648 ^ 1'b0 ;
  assign n8652 = ( n1214 & n7176 ) | ( n1214 & ~n8481 ) | ( n7176 & ~n8481 ) ;
  assign n8653 = ~n2102 & n5779 ;
  assign n8657 = ( ~n3432 & n3804 ) | ( ~n3432 & n3819 ) | ( n3804 & n3819 ) ;
  assign n8654 = n3972 ^ n1307 ^ 1'b0 ;
  assign n8655 = ( x182 & n795 ) | ( x182 & ~n8654 ) | ( n795 & ~n8654 ) ;
  assign n8656 = ~n8529 & n8655 ;
  assign n8658 = n8657 ^ n8656 ^ 1'b0 ;
  assign n8659 = n6669 ^ n5083 ^ n1276 ;
  assign n8660 = n1106 ^ n300 ^ 1'b0 ;
  assign n8661 = n837 & ~n8660 ;
  assign n8662 = n8661 ^ n4729 ^ 1'b0 ;
  assign n8663 = x168 & n8662 ;
  assign n8664 = n8663 ^ n3196 ^ 1'b0 ;
  assign n8665 = n578 ^ x121 ^ 1'b0 ;
  assign n8666 = n2993 ^ n1655 ^ 1'b0 ;
  assign n8667 = n1919 | n8666 ;
  assign n8668 = n8665 & ~n8667 ;
  assign n8669 = ( n3786 & n5576 ) | ( n3786 & ~n8668 ) | ( n5576 & ~n8668 ) ;
  assign n8672 = n8328 ^ n5294 ^ 1'b0 ;
  assign n8673 = n8672 ^ n1141 ^ 1'b0 ;
  assign n8670 = n3922 ^ n1024 ^ n360 ;
  assign n8671 = n8670 ^ n5275 ^ n378 ;
  assign n8674 = n8673 ^ n8671 ^ 1'b0 ;
  assign n8675 = x156 & n3934 ;
  assign n8676 = ( n3934 & ~n6552 ) | ( n3934 & n8675 ) | ( ~n6552 & n8675 ) ;
  assign n8677 = n5725 | n6799 ;
  assign n8678 = n8676 | n8677 ;
  assign n8679 = ( ~n1870 & n4801 ) | ( ~n1870 & n6351 ) | ( n4801 & n6351 ) ;
  assign n8680 = n1684 | n8321 ;
  assign n8681 = n8679 | n8680 ;
  assign n8682 = n8500 ^ n2614 ^ 1'b0 ;
  assign n8683 = n8682 ^ n6778 ^ 1'b0 ;
  assign n8684 = n5411 ^ n5123 ^ x73 ;
  assign n8685 = ~n2385 & n7497 ;
  assign n8686 = ~n5557 & n7916 ;
  assign n8687 = ~n7486 & n8686 ;
  assign n8688 = n2310 & ~n3105 ;
  assign n8689 = n1678 & n7520 ;
  assign n8690 = n8689 ^ n2386 ^ n1116 ;
  assign n8691 = n8690 ^ x166 ^ 1'b0 ;
  assign n8692 = x19 & ~n8691 ;
  assign n8693 = n8692 ^ n5937 ^ 1'b0 ;
  assign n8694 = n6699 | n8693 ;
  assign n8695 = n6774 | n8694 ;
  assign n8696 = n8129 ^ n5128 ^ n1669 ;
  assign n8697 = ( n1069 & n8695 ) | ( n1069 & ~n8696 ) | ( n8695 & ~n8696 ) ;
  assign n8698 = n584 | n1328 ;
  assign n8699 = n3257 & ~n8698 ;
  assign n8700 = n1831 & n8699 ;
  assign n8701 = n8700 ^ n5190 ^ 1'b0 ;
  assign n8702 = n7289 & ~n8701 ;
  assign n8703 = n8702 ^ n6223 ^ n4139 ;
  assign n8704 = ( ~n3806 & n4308 ) | ( ~n3806 & n8703 ) | ( n4308 & n8703 ) ;
  assign n8705 = n8704 ^ n2427 ^ 1'b0 ;
  assign n8712 = x102 & ~n7680 ;
  assign n8713 = ~x159 & n8712 ;
  assign n8706 = n3521 ^ n659 ^ 1'b0 ;
  assign n8707 = n3234 & ~n8706 ;
  assign n8708 = n8707 ^ n578 ^ 1'b0 ;
  assign n8709 = n3590 & n8708 ;
  assign n8710 = n5107 | n5991 ;
  assign n8711 = n8709 | n8710 ;
  assign n8714 = n8713 ^ n8711 ^ 1'b0 ;
  assign n8715 = n4024 & ~n8714 ;
  assign n8718 = n2233 ^ n1548 ^ x104 ;
  assign n8716 = ( ~x230 & n703 ) | ( ~x230 & n1261 ) | ( n703 & n1261 ) ;
  assign n8717 = ( n1254 & n2157 ) | ( n1254 & n8716 ) | ( n2157 & n8716 ) ;
  assign n8719 = n8718 ^ n8717 ^ 1'b0 ;
  assign n8720 = n8715 & ~n8719 ;
  assign n8721 = ~n4008 & n8720 ;
  assign n8722 = ( n2852 & ~n3343 ) | ( n2852 & n4559 ) | ( ~n3343 & n4559 ) ;
  assign n8723 = n1969 ^ n1543 ^ 1'b0 ;
  assign n8724 = n8722 & n8723 ;
  assign n8725 = n2884 ^ n303 ^ 1'b0 ;
  assign n8726 = n8725 ^ n2642 ^ n911 ;
  assign n8727 = n1175 ^ n697 ^ 1'b0 ;
  assign n8728 = n1791 & ~n3266 ;
  assign n8729 = n8728 ^ n5582 ^ 1'b0 ;
  assign n8730 = ~n4451 & n8729 ;
  assign n8731 = ~n2167 & n8730 ;
  assign n8732 = ( x209 & n1562 ) | ( x209 & n1596 ) | ( n1562 & n1596 ) ;
  assign n8733 = ~n3591 & n3773 ;
  assign n8734 = ~n5447 & n7317 ;
  assign n8735 = n4200 | n7100 ;
  assign n8736 = n8735 ^ n694 ^ 1'b0 ;
  assign n8741 = n7726 ^ n2718 ^ 1'b0 ;
  assign n8742 = x68 & ~n8741 ;
  assign n8737 = n2229 & ~n2865 ;
  assign n8738 = n2554 & n8737 ;
  assign n8739 = n8738 ^ n474 ^ 1'b0 ;
  assign n8740 = ~n1971 & n8739 ;
  assign n8743 = n8742 ^ n8740 ^ x9 ;
  assign n8744 = ~n4803 & n5471 ;
  assign n8745 = n8744 ^ n2562 ^ 1'b0 ;
  assign n8746 = ( n1885 & n5576 ) | ( n1885 & ~n5713 ) | ( n5576 & ~n5713 ) ;
  assign n8747 = n3948 & ~n8746 ;
  assign n8748 = ~n8745 & n8747 ;
  assign n8749 = n7155 ^ n2769 ^ 1'b0 ;
  assign n8750 = ~n8286 & n8384 ;
  assign n8751 = n8094 ^ n7517 ^ n6252 ;
  assign n8752 = n4386 & n7686 ;
  assign n8753 = n1564 & ~n8752 ;
  assign n8754 = n6448 | n6753 ;
  assign n8755 = n1867 ^ n1724 ^ 1'b0 ;
  assign n8756 = n8755 ^ n4413 ^ 1'b0 ;
  assign n8757 = n4666 ^ n2861 ^ n1852 ;
  assign n8758 = ~n1088 & n3113 ;
  assign n8761 = ( ~n4244 & n6303 ) | ( ~n4244 & n7769 ) | ( n6303 & n7769 ) ;
  assign n8762 = n8761 ^ n5265 ^ n2658 ;
  assign n8760 = n4876 ^ n1739 ^ n591 ;
  assign n8763 = n8762 ^ n8760 ^ n4141 ;
  assign n8759 = n377 | n7929 ;
  assign n8764 = n8763 ^ n8759 ^ 1'b0 ;
  assign n8765 = n4228 & n5786 ;
  assign n8766 = n3073 & n8765 ;
  assign n8767 = n8766 ^ n334 ^ 1'b0 ;
  assign n8768 = n5353 | n6679 ;
  assign n8769 = n8768 ^ n2841 ^ 1'b0 ;
  assign n8770 = n8767 & ~n8769 ;
  assign n8771 = n8770 ^ x9 ^ 1'b0 ;
  assign n8772 = n2767 & ~n6499 ;
  assign n8773 = n8772 ^ n4947 ^ n2447 ;
  assign n8774 = ( n1750 & ~n7106 ) | ( n1750 & n8773 ) | ( ~n7106 & n8773 ) ;
  assign n8775 = ~n1639 & n3067 ;
  assign n8776 = n4628 | n8775 ;
  assign n8777 = ~n1799 & n5436 ;
  assign n8778 = n3717 | n6236 ;
  assign n8779 = n7155 ^ n1258 ^ 1'b0 ;
  assign n8780 = n8778 & n8779 ;
  assign n8781 = x181 & n8780 ;
  assign n8782 = ( n4137 & ~n8777 ) | ( n4137 & n8781 ) | ( ~n8777 & n8781 ) ;
  assign n8783 = n1755 & n8469 ;
  assign n8784 = n4884 ^ n1385 ^ n745 ;
  assign n8785 = n8784 ^ n6921 ^ 1'b0 ;
  assign n8786 = ~n898 & n8785 ;
  assign n8787 = n1933 ^ x218 ^ 1'b0 ;
  assign n8788 = n2137 & n8787 ;
  assign n8789 = n5681 & ~n7801 ;
  assign n8790 = ~n6085 & n8789 ;
  assign n8791 = n8790 ^ x70 ^ 1'b0 ;
  assign n8792 = n1761 ^ n1569 ^ 1'b0 ;
  assign n8804 = n3040 ^ n2622 ^ 1'b0 ;
  assign n8805 = ~n363 & n8804 ;
  assign n8799 = n256 | n2469 ;
  assign n8800 = n7916 ^ n4874 ^ 1'b0 ;
  assign n8801 = n8800 ^ n6389 ^ 1'b0 ;
  assign n8802 = n8801 ^ n7639 ^ n4303 ;
  assign n8803 = n8799 & n8802 ;
  assign n8806 = n8805 ^ n8803 ^ 1'b0 ;
  assign n8793 = x13 & ~n5586 ;
  assign n8794 = n8793 ^ n1283 ^ 1'b0 ;
  assign n8795 = n675 & ~n1701 ;
  assign n8796 = n8794 & n8795 ;
  assign n8797 = n8078 ^ n8041 ^ 1'b0 ;
  assign n8798 = n8796 | n8797 ;
  assign n8807 = n8806 ^ n8798 ^ n7088 ;
  assign n8808 = n4462 ^ n2416 ^ 1'b0 ;
  assign n8809 = n5679 ^ n5044 ^ 1'b0 ;
  assign n8810 = n8808 & ~n8809 ;
  assign n8811 = n2680 & n8810 ;
  assign n8812 = ~x77 & n8811 ;
  assign n8813 = n6528 ^ n4219 ^ n2162 ;
  assign n8814 = ~n7811 & n8813 ;
  assign n8815 = n1695 & n8814 ;
  assign n8816 = ( n5532 & n6078 ) | ( n5532 & ~n8815 ) | ( n6078 & ~n8815 ) ;
  assign n8817 = n3680 & n5339 ;
  assign n8818 = ~n4278 & n8817 ;
  assign n8819 = ~n5214 & n8818 ;
  assign n8824 = n913 | n6845 ;
  assign n8820 = n2023 | n2577 ;
  assign n8821 = n7769 & ~n8820 ;
  assign n8822 = n3909 & n6563 ;
  assign n8823 = n8821 & n8822 ;
  assign n8825 = n8824 ^ n8823 ^ 1'b0 ;
  assign n8826 = ~n8819 & n8825 ;
  assign n8827 = n341 & n979 ;
  assign n8828 = n1813 & ~n3992 ;
  assign n8829 = n8828 ^ n7515 ^ 1'b0 ;
  assign n8830 = n4496 ^ n3566 ^ 1'b0 ;
  assign n8831 = n6914 ^ n4364 ^ 1'b0 ;
  assign n8832 = n7925 ^ n2095 ^ 1'b0 ;
  assign n8833 = n8824 | n8832 ;
  assign n8834 = x139 & n5545 ;
  assign n8835 = n5548 ^ n2147 ^ 1'b0 ;
  assign n8836 = n8835 ^ n7610 ^ 1'b0 ;
  assign n8837 = n6425 ^ n4543 ^ n3636 ;
  assign n8838 = n2121 & n8837 ;
  assign n8839 = n8836 & n8838 ;
  assign n8840 = n8834 & ~n8839 ;
  assign n8841 = ~n7773 & n8840 ;
  assign n8842 = n6262 ^ n3021 ^ 1'b0 ;
  assign n8843 = n8502 | n8842 ;
  assign n8844 = n2770 & n6143 ;
  assign n8845 = n8844 ^ n5553 ^ 1'b0 ;
  assign n8846 = n4915 & n7024 ;
  assign n8847 = ( ~n2573 & n8845 ) | ( ~n2573 & n8846 ) | ( n8845 & n8846 ) ;
  assign n8848 = n8847 ^ n6125 ^ 1'b0 ;
  assign n8849 = ~n2058 & n5689 ;
  assign n8850 = n6649 & n8849 ;
  assign n8851 = n8850 ^ n6543 ^ 1'b0 ;
  assign n8852 = n1664 & ~n2718 ;
  assign n8853 = ~n8851 & n8852 ;
  assign n8854 = n2718 ^ n1585 ^ 1'b0 ;
  assign n8855 = n3315 & n8854 ;
  assign n8856 = n2619 & n4148 ;
  assign n8857 = n8856 ^ n6717 ^ 1'b0 ;
  assign n8858 = n8855 & n8857 ;
  assign n8859 = n7777 & n8858 ;
  assign n8860 = n4203 & n5800 ;
  assign n8861 = ~n1459 & n8860 ;
  assign n8862 = n3341 ^ n522 ^ 1'b0 ;
  assign n8863 = ( n3471 & n8861 ) | ( n3471 & ~n8862 ) | ( n8861 & ~n8862 ) ;
  assign n8864 = n7762 ^ n4633 ^ 1'b0 ;
  assign n8865 = n3383 & n8864 ;
  assign n8866 = n1185 & n3507 ;
  assign n8867 = ~n6914 & n8866 ;
  assign n8868 = n1895 & n6015 ;
  assign n8869 = n8868 ^ n7674 ^ 1'b0 ;
  assign n8870 = n3429 & n7830 ;
  assign n8872 = n459 & ~n3636 ;
  assign n8871 = n4398 | n8218 ;
  assign n8873 = n8872 ^ n8871 ^ 1'b0 ;
  assign n8874 = ~n1487 & n3570 ;
  assign n8875 = n8874 ^ n8181 ^ 1'b0 ;
  assign n8876 = n8875 ^ n6193 ^ 1'b0 ;
  assign n8877 = n2539 & ~n6164 ;
  assign n8878 = n8877 ^ n6930 ^ 1'b0 ;
  assign n8879 = n5323 ^ n2488 ^ 1'b0 ;
  assign n8880 = n4631 & n8879 ;
  assign n8881 = ~n2794 & n8880 ;
  assign n8882 = n8881 ^ n877 ^ 1'b0 ;
  assign n8883 = ( x82 & n861 ) | ( x82 & ~n2147 ) | ( n861 & ~n2147 ) ;
  assign n8884 = n3457 & ~n8883 ;
  assign n8885 = n8884 ^ n1345 ^ 1'b0 ;
  assign n8886 = n3549 & n8885 ;
  assign n8887 = n8886 ^ n5840 ^ 1'b0 ;
  assign n8888 = n5187 ^ n1000 ^ 1'b0 ;
  assign n8889 = n557 & ~n929 ;
  assign n8890 = n1278 & n8889 ;
  assign n8891 = ( n752 & ~n3423 ) | ( n752 & n5055 ) | ( ~n3423 & n5055 ) ;
  assign n8892 = n8891 ^ n1768 ^ 1'b0 ;
  assign n8893 = n4053 & n8892 ;
  assign n8894 = n7157 ^ n3336 ^ 1'b0 ;
  assign n8895 = n8894 ^ n5043 ^ n2253 ;
  assign n8896 = n8317 ^ n7592 ^ 1'b0 ;
  assign n8897 = ( x140 & n8426 ) | ( x140 & ~n8896 ) | ( n8426 & ~n8896 ) ;
  assign n8898 = n911 ^ n834 ^ 1'b0 ;
  assign n8899 = n8898 ^ n1247 ^ n511 ;
  assign n8903 = n7243 ^ n4230 ^ 1'b0 ;
  assign n8900 = n2827 & n4197 ;
  assign n8901 = ~n2847 & n8900 ;
  assign n8902 = ~n8662 & n8901 ;
  assign n8904 = n8903 ^ n8902 ^ x176 ;
  assign n8907 = ~x137 & n1996 ;
  assign n8908 = ( ~n2977 & n4078 ) | ( ~n2977 & n7017 ) | ( n4078 & n7017 ) ;
  assign n8909 = n2278 & ~n8908 ;
  assign n8910 = n1754 & ~n8909 ;
  assign n8911 = n7989 & n8910 ;
  assign n8912 = n1260 & ~n8911 ;
  assign n8913 = ~n8907 & n8912 ;
  assign n8905 = n5003 ^ n4569 ^ 1'b0 ;
  assign n8906 = ~n3802 & n8905 ;
  assign n8914 = n8913 ^ n8906 ^ 1'b0 ;
  assign n8915 = n5926 ^ n3920 ^ 1'b0 ;
  assign n8916 = n3941 & n8915 ;
  assign n8917 = n8916 ^ n3872 ^ 1'b0 ;
  assign n8918 = n8835 | n8917 ;
  assign n8919 = n8657 ^ n3979 ^ 1'b0 ;
  assign n8920 = n4303 | n8919 ;
  assign n8921 = n7186 ^ n3361 ^ 1'b0 ;
  assign n8922 = ~n2911 & n8921 ;
  assign n8923 = n2720 & ~n8922 ;
  assign n8924 = n6147 ^ n5947 ^ 1'b0 ;
  assign n8925 = n4304 | n8924 ;
  assign n8926 = n8201 ^ n2116 ^ n349 ;
  assign n8927 = ( n4113 & ~n8925 ) | ( n4113 & n8926 ) | ( ~n8925 & n8926 ) ;
  assign n8928 = ( ~x31 & n3774 ) | ( ~x31 & n7726 ) | ( n3774 & n7726 ) ;
  assign n8929 = n5797 ^ n3923 ^ n1891 ;
  assign n8930 = ( n6717 & n8928 ) | ( n6717 & ~n8929 ) | ( n8928 & ~n8929 ) ;
  assign n8931 = n4027 ^ n450 ^ 1'b0 ;
  assign n8932 = n5344 | n8931 ;
  assign n8933 = n4664 ^ n2517 ^ 1'b0 ;
  assign n8934 = ~n8932 & n8933 ;
  assign n8935 = ( ~n5541 & n6685 ) | ( ~n5541 & n8934 ) | ( n6685 & n8934 ) ;
  assign n8936 = n8935 ^ n5316 ^ n4091 ;
  assign n8937 = n7880 ^ n6710 ^ n5135 ;
  assign n8938 = n8936 & n8937 ;
  assign n8939 = n8938 ^ x137 ^ 1'b0 ;
  assign n8940 = n1596 ^ n1090 ^ n382 ;
  assign n8941 = ~n3160 & n8940 ;
  assign n8942 = n8165 ^ n4069 ^ 1'b0 ;
  assign n8943 = n8942 ^ n6504 ^ 1'b0 ;
  assign n8944 = n8186 & ~n8943 ;
  assign n8945 = ( n3037 & n3106 ) | ( n3037 & ~n7718 ) | ( n3106 & ~n7718 ) ;
  assign n8946 = n341 & ~n4950 ;
  assign n8947 = ( x101 & ~n2942 ) | ( x101 & n3857 ) | ( ~n2942 & n3857 ) ;
  assign n8948 = ~n3219 & n8947 ;
  assign n8949 = ( x162 & n1895 ) | ( x162 & n2523 ) | ( n1895 & n2523 ) ;
  assign n8950 = n5207 & n8949 ;
  assign n8951 = n8950 ^ n5479 ^ 1'b0 ;
  assign n8952 = ( n415 & n2019 ) | ( n415 & ~n2936 ) | ( n2019 & ~n2936 ) ;
  assign n8964 = n8689 ^ n1886 ^ 1'b0 ;
  assign n8965 = n8964 ^ n6414 ^ 1'b0 ;
  assign n8962 = ~n625 & n774 ;
  assign n8955 = n6797 ^ n3596 ^ n2541 ;
  assign n8956 = n4031 | n8955 ;
  assign n8957 = n957 & n8956 ;
  assign n8958 = n7326 ^ n6487 ^ n3504 ;
  assign n8959 = n5033 | n8958 ;
  assign n8960 = n8957 | n8959 ;
  assign n8953 = ~n2009 & n8722 ;
  assign n8954 = ~n3680 & n8953 ;
  assign n8961 = n8960 ^ n8954 ^ 1'b0 ;
  assign n8963 = n8962 ^ n8961 ^ 1'b0 ;
  assign n8966 = n8965 ^ n8963 ^ 1'b0 ;
  assign n8967 = ( n8951 & n8952 ) | ( n8951 & ~n8966 ) | ( n8952 & ~n8966 ) ;
  assign n8968 = n2171 ^ n659 ^ 1'b0 ;
  assign n8969 = x17 & ~n8968 ;
  assign n8970 = n8969 ^ n5039 ^ 1'b0 ;
  assign n8971 = ( ~n756 & n2835 ) | ( ~n756 & n4510 ) | ( n2835 & n4510 ) ;
  assign n8972 = n8971 ^ n3525 ^ 1'b0 ;
  assign n8973 = ~n3481 & n8972 ;
  assign n8974 = n7806 ^ n6540 ^ 1'b0 ;
  assign n8975 = n4948 & n8974 ;
  assign n8976 = n8975 ^ n6711 ^ 1'b0 ;
  assign n8977 = n1809 & ~n8193 ;
  assign n8978 = ~x124 & n8977 ;
  assign n8979 = n8978 ^ n365 ^ 1'b0 ;
  assign n8981 = ( n980 & ~n1951 ) | ( n980 & n4703 ) | ( ~n1951 & n4703 ) ;
  assign n8980 = n606 & n2769 ;
  assign n8982 = n8981 ^ n8980 ^ 1'b0 ;
  assign n8983 = ~n7867 & n8982 ;
  assign n8984 = n3069 | n3140 ;
  assign n8985 = n1564 | n8984 ;
  assign n8986 = ~n7665 & n8985 ;
  assign n8987 = n6064 ^ n5189 ^ 1'b0 ;
  assign n8988 = n7995 | n8987 ;
  assign n8989 = n8986 | n8988 ;
  assign n8990 = n1580 ^ n1266 ^ 1'b0 ;
  assign n8991 = x191 & n8990 ;
  assign n8992 = n4751 & n8991 ;
  assign n8993 = ~n8391 & n8992 ;
  assign n8994 = n3624 & ~n8437 ;
  assign n8995 = n8994 ^ n6558 ^ 1'b0 ;
  assign n8996 = ( n1853 & ~n2006 ) | ( n1853 & n5625 ) | ( ~n2006 & n5625 ) ;
  assign n9000 = ~n606 & n4471 ;
  assign n9001 = n9000 ^ n1842 ^ 1'b0 ;
  assign n9002 = ~n8657 & n9001 ;
  assign n8997 = n2411 ^ n826 ^ 1'b0 ;
  assign n8998 = n3596 & ~n8997 ;
  assign n8999 = n2804 & n8998 ;
  assign n9003 = n9002 ^ n8999 ^ 1'b0 ;
  assign n9004 = n8996 | n9003 ;
  assign n9007 = n868 & ~n4200 ;
  assign n9008 = ~n4811 & n9007 ;
  assign n9009 = n9008 ^ n5669 ^ 1'b0 ;
  assign n9010 = n4245 & n9009 ;
  assign n9006 = n2786 | n3656 ;
  assign n9011 = n9010 ^ n9006 ^ 1'b0 ;
  assign n9005 = n4258 ^ n576 ^ 1'b0 ;
  assign n9012 = n9011 ^ n9005 ^ 1'b0 ;
  assign n9015 = n5480 ^ n806 ^ 1'b0 ;
  assign n9016 = n9015 ^ n4899 ^ 1'b0 ;
  assign n9017 = n2560 | n9016 ;
  assign n9013 = ~n478 & n3358 ;
  assign n9014 = n9013 ^ n7774 ^ 1'b0 ;
  assign n9018 = n9017 ^ n9014 ^ 1'b0 ;
  assign n9019 = n3049 ^ n1045 ^ 1'b0 ;
  assign n9020 = n9019 ^ n8124 ^ 1'b0 ;
  assign n9021 = n2875 ^ n824 ^ 1'b0 ;
  assign n9022 = ( n277 & n652 ) | ( n277 & n1440 ) | ( n652 & n1440 ) ;
  assign n9023 = n9022 ^ n7348 ^ 1'b0 ;
  assign n9024 = n9021 & n9023 ;
  assign n9025 = ( n798 & n863 ) | ( n798 & ~n1032 ) | ( n863 & ~n1032 ) ;
  assign n9026 = ( n2045 & n4338 ) | ( n2045 & ~n9025 ) | ( n4338 & ~n9025 ) ;
  assign n9027 = n6562 | n9026 ;
  assign n9028 = n5814 & ~n9027 ;
  assign n9029 = ~n2588 & n4288 ;
  assign n9030 = n9029 ^ n1795 ^ 1'b0 ;
  assign n9031 = n3000 & ~n9030 ;
  assign n9032 = n1554 & n9031 ;
  assign n9033 = n3302 ^ n915 ^ x1 ;
  assign n9034 = ~n9032 & n9033 ;
  assign n9035 = n9034 ^ n723 ^ 1'b0 ;
  assign n9036 = n4851 ^ n3279 ^ 1'b0 ;
  assign n9037 = ~n5337 & n9036 ;
  assign n9038 = n9037 ^ n5595 ^ n2697 ;
  assign n9039 = ~n4048 & n9038 ;
  assign n9040 = ~n6390 & n9039 ;
  assign n9041 = ( x88 & n3140 ) | ( x88 & ~n8900 ) | ( n3140 & ~n8900 ) ;
  assign n9042 = n3237 & n7435 ;
  assign n9043 = ~n5287 & n9042 ;
  assign n9044 = n5857 | n9043 ;
  assign n9045 = n1390 & n1602 ;
  assign n9046 = ( n4958 & n6856 ) | ( n4958 & n8119 ) | ( n6856 & n8119 ) ;
  assign n9047 = ~n3192 & n9046 ;
  assign n9050 = ( n2634 & n3835 ) | ( n2634 & n8155 ) | ( n3835 & n8155 ) ;
  assign n9051 = ~n887 & n9050 ;
  assign n9048 = n8311 ^ n545 ^ 1'b0 ;
  assign n9049 = n9048 ^ n5713 ^ n1203 ;
  assign n9052 = n9051 ^ n9049 ^ 1'b0 ;
  assign n9053 = n1283 & n2954 ;
  assign n9054 = n9053 ^ n3657 ^ 1'b0 ;
  assign n9055 = n3403 & ~n9054 ;
  assign n9056 = ~n3731 & n9055 ;
  assign n9057 = n8684 ^ n3728 ^ 1'b0 ;
  assign n9058 = n2308 & n9057 ;
  assign n9059 = n9041 ^ n3184 ^ n472 ;
  assign n9060 = n3637 | n4007 ;
  assign n9061 = n9060 ^ n2598 ^ 1'b0 ;
  assign n9062 = n9061 ^ n6087 ^ n2737 ;
  assign n9063 = n1677 | n8658 ;
  assign n9064 = ( ~n1515 & n3332 ) | ( ~n1515 & n4024 ) | ( n3332 & n4024 ) ;
  assign n9065 = n1547 | n1719 ;
  assign n9066 = n9065 ^ n5658 ^ 1'b0 ;
  assign n9067 = n9064 | n9066 ;
  assign n9069 = ( n968 & ~n6514 ) | ( n968 & n8157 ) | ( ~n6514 & n8157 ) ;
  assign n9068 = n4039 | n4138 ;
  assign n9070 = n9069 ^ n9068 ^ 1'b0 ;
  assign n9071 = n7639 | n8717 ;
  assign n9072 = n2260 & ~n2487 ;
  assign n9073 = n3217 & n9072 ;
  assign n9074 = ( ~n4141 & n6831 ) | ( ~n4141 & n9073 ) | ( n6831 & n9073 ) ;
  assign n9075 = n3196 ^ n3064 ^ 1'b0 ;
  assign n9076 = ~n780 & n3695 ;
  assign n9077 = n5731 & ~n9076 ;
  assign n9078 = n6620 ^ n2837 ^ 1'b0 ;
  assign n9079 = n5436 ^ n5255 ^ n843 ;
  assign n9080 = n9079 ^ n1769 ^ n1462 ;
  assign n9081 = n5134 ^ x209 ^ 1'b0 ;
  assign n9083 = ~n5863 & n5869 ;
  assign n9082 = ( x171 & n1038 ) | ( x171 & ~n4744 ) | ( n1038 & ~n4744 ) ;
  assign n9084 = n9083 ^ n9082 ^ n1613 ;
  assign n9089 = ~x108 & n6758 ;
  assign n9085 = n1362 & ~n1442 ;
  assign n9086 = n9085 ^ n7525 ^ 1'b0 ;
  assign n9087 = n2230 & n9086 ;
  assign n9088 = n9087 ^ n953 ^ 1'b0 ;
  assign n9090 = n9089 ^ n9088 ^ n7784 ;
  assign n9091 = n9090 ^ n1154 ^ 1'b0 ;
  assign n9092 = n1138 | n9091 ;
  assign n9093 = n292 & n4975 ;
  assign n9094 = n9093 ^ n3914 ^ 1'b0 ;
  assign n9095 = ( n1774 & n2517 ) | ( n1774 & ~n5153 ) | ( n2517 & ~n5153 ) ;
  assign n9096 = n9094 & n9095 ;
  assign n9097 = n5139 ^ n2242 ^ 1'b0 ;
  assign n9098 = n9097 ^ n5413 ^ 1'b0 ;
  assign n9099 = ( n1199 & ~n3429 ) | ( n1199 & n8193 ) | ( ~n3429 & n8193 ) ;
  assign n9100 = ~n9098 & n9099 ;
  assign n9101 = n2047 & n8145 ;
  assign n9102 = n394 & n3935 ;
  assign n9103 = ( x105 & n1572 ) | ( x105 & ~n6106 ) | ( n1572 & ~n6106 ) ;
  assign n9104 = ( n2906 & ~n9102 ) | ( n2906 & n9103 ) | ( ~n9102 & n9103 ) ;
  assign n9105 = ~n9101 & n9104 ;
  assign n9106 = n9105 ^ n5091 ^ 1'b0 ;
  assign n9107 = n273 | n2772 ;
  assign n9108 = n9107 ^ x65 ^ 1'b0 ;
  assign n9109 = n8428 ^ n4342 ^ 1'b0 ;
  assign n9110 = n8049 ^ n627 ^ 1'b0 ;
  assign n9112 = n5382 ^ n1851 ^ 1'b0 ;
  assign n9111 = n1843 & n2314 ;
  assign n9113 = n9112 ^ n9111 ^ n2645 ;
  assign n9114 = x27 & x193 ;
  assign n9115 = n9114 ^ n3599 ^ 1'b0 ;
  assign n9116 = n2575 & ~n9115 ;
  assign n9117 = ~n6938 & n9116 ;
  assign n9118 = n2663 & n3600 ;
  assign n9119 = n8260 ^ n6936 ^ 1'b0 ;
  assign n9120 = n1877 | n9119 ;
  assign n9121 = ~n1482 & n8496 ;
  assign n9122 = n7366 ^ n5374 ^ n1541 ;
  assign n9123 = n4174 ^ n2526 ^ 1'b0 ;
  assign n9126 = n633 & ~n2194 ;
  assign n9127 = n297 | n9126 ;
  assign n9128 = n2216 | n9127 ;
  assign n9129 = ~n4299 & n9128 ;
  assign n9124 = n4462 ^ n3235 ^ 1'b0 ;
  assign n9125 = n9088 & ~n9124 ;
  assign n9130 = n9129 ^ n9125 ^ 1'b0 ;
  assign n9131 = n3568 & n9130 ;
  assign n9132 = n503 | n3948 ;
  assign n9133 = n973 & ~n2024 ;
  assign n9134 = n9133 ^ n4268 ^ 1'b0 ;
  assign n9135 = n7863 ^ n2329 ^ 1'b0 ;
  assign n9136 = n9134 & ~n9135 ;
  assign n9140 = x31 & ~n1063 ;
  assign n9141 = n9140 ^ n2660 ^ 1'b0 ;
  assign n9142 = n9141 ^ n7840 ^ n5342 ;
  assign n9137 = n7637 ^ n1368 ^ 1'b0 ;
  assign n9138 = n595 & n9137 ;
  assign n9139 = n5109 & ~n9138 ;
  assign n9143 = n9142 ^ n9139 ^ n428 ;
  assign n9144 = n4994 ^ n433 ^ 1'b0 ;
  assign n9145 = ~n512 & n9144 ;
  assign n9146 = ( ~x116 & n1532 ) | ( ~x116 & n9145 ) | ( n1532 & n9145 ) ;
  assign n9147 = n6034 & ~n8718 ;
  assign n9148 = n1266 & n9147 ;
  assign n9151 = n545 & ~n7621 ;
  assign n9152 = n9151 ^ n5157 ^ 1'b0 ;
  assign n9153 = n5819 & ~n9152 ;
  assign n9154 = n4239 & ~n9153 ;
  assign n9149 = ( x81 & n3875 ) | ( x81 & n4448 ) | ( n3875 & n4448 ) ;
  assign n9150 = n2216 & ~n9149 ;
  assign n9155 = n9154 ^ n9150 ^ 1'b0 ;
  assign n9156 = ( n4107 & n4372 ) | ( n4107 & ~n4579 ) | ( n4372 & ~n4579 ) ;
  assign n9157 = ~n387 & n9156 ;
  assign n9158 = n9157 ^ n4999 ^ 1'b0 ;
  assign n9159 = ( n2280 & n6581 ) | ( n2280 & n7348 ) | ( n6581 & n7348 ) ;
  assign n9160 = n4045 & ~n4690 ;
  assign n9163 = ( x164 & n866 ) | ( x164 & n5148 ) | ( n866 & n5148 ) ;
  assign n9161 = n2636 | n2794 ;
  assign n9162 = n5599 & ~n9161 ;
  assign n9164 = n9163 ^ n9162 ^ 1'b0 ;
  assign n9165 = n8737 & n9164 ;
  assign n9166 = n6364 | n9165 ;
  assign n9167 = n9166 ^ n2341 ^ 1'b0 ;
  assign n9168 = ( x0 & n335 ) | ( x0 & ~n2551 ) | ( n335 & ~n2551 ) ;
  assign n9169 = n9168 ^ n7521 ^ 1'b0 ;
  assign n9170 = n1413 & n9169 ;
  assign n9174 = n2399 ^ n1852 ^ 1'b0 ;
  assign n9171 = ~n449 & n990 ;
  assign n9172 = ~n4365 & n9171 ;
  assign n9173 = ( n493 & n3147 ) | ( n493 & ~n9172 ) | ( n3147 & ~n9172 ) ;
  assign n9175 = n9174 ^ n9173 ^ 1'b0 ;
  assign n9176 = n6086 & ~n9175 ;
  assign n9177 = ( x43 & ~n3670 ) | ( x43 & n5628 ) | ( ~n3670 & n5628 ) ;
  assign n9178 = n9177 ^ n2590 ^ 1'b0 ;
  assign n9179 = ( n4855 & n7218 ) | ( n4855 & n9178 ) | ( n7218 & n9178 ) ;
  assign n9180 = ( n1744 & ~n3651 ) | ( n1744 & n9179 ) | ( ~n3651 & n9179 ) ;
  assign n9181 = n3531 ^ n2708 ^ 1'b0 ;
  assign n9182 = n3959 ^ n2121 ^ 1'b0 ;
  assign n9183 = n358 | n1138 ;
  assign n9184 = n9183 ^ n3629 ^ 1'b0 ;
  assign n9185 = n9182 & n9184 ;
  assign n9186 = n1653 | n6710 ;
  assign n9187 = n3275 | n5476 ;
  assign n9188 = n3328 & ~n9187 ;
  assign n9189 = n9188 ^ n8932 ^ n4961 ;
  assign n9190 = ~n980 & n9189 ;
  assign n9191 = n9190 ^ n2092 ^ 1'b0 ;
  assign n9192 = n9186 & ~n9191 ;
  assign n9193 = ( n955 & n3982 ) | ( n955 & ~n7520 ) | ( n3982 & ~n7520 ) ;
  assign n9194 = n4187 & ~n7961 ;
  assign n9195 = n2208 & n9194 ;
  assign n9196 = n9193 & n9195 ;
  assign n9197 = n944 & n6149 ;
  assign n9198 = n1487 ^ n1022 ^ n629 ;
  assign n9199 = n496 & n9198 ;
  assign n9200 = ~n4895 & n9199 ;
  assign n9201 = n7841 & ~n9200 ;
  assign n9202 = n528 & n9201 ;
  assign n9203 = n9202 ^ n7416 ^ 1'b0 ;
  assign n9205 = ~n1506 & n2231 ;
  assign n9206 = n2302 & n9205 ;
  assign n9204 = n1350 | n1497 ;
  assign n9207 = n9206 ^ n9204 ^ 1'b0 ;
  assign n9208 = n8067 | n9207 ;
  assign n9209 = n9203 & ~n9208 ;
  assign n9210 = n6402 | n9209 ;
  assign n9211 = n2985 ^ n1542 ^ 1'b0 ;
  assign n9212 = n752 & ~n9211 ;
  assign n9213 = ~x134 & n9212 ;
  assign n9214 = n8964 ^ n358 ^ 1'b0 ;
  assign n9215 = ~n4922 & n9214 ;
  assign n9216 = n4383 & ~n4394 ;
  assign n9217 = n9216 ^ n3059 ^ 1'b0 ;
  assign n9218 = n4814 & n8363 ;
  assign n9219 = n9218 ^ n1709 ^ 1'b0 ;
  assign n9220 = ~n2338 & n9219 ;
  assign n9221 = n9217 & n9220 ;
  assign n9222 = n5575 ^ n3958 ^ n2070 ;
  assign n9223 = n6973 & ~n9222 ;
  assign n9224 = ~n5579 & n9223 ;
  assign n9232 = n5815 ^ n2719 ^ 1'b0 ;
  assign n9229 = n6863 ^ n6770 ^ 1'b0 ;
  assign n9230 = n2957 & ~n9229 ;
  assign n9231 = ~n3689 & n9230 ;
  assign n9225 = ~n2165 & n6319 ;
  assign n9226 = ~n5203 & n9225 ;
  assign n9227 = n1260 & n5895 ;
  assign n9228 = n9226 & n9227 ;
  assign n9233 = n9232 ^ n9231 ^ n9228 ;
  assign n9235 = n2376 & n7887 ;
  assign n9234 = x25 & ~n3067 ;
  assign n9236 = n9235 ^ n9234 ^ n8893 ;
  assign n9240 = ( ~n752 & n1613 ) | ( ~n752 & n3033 ) | ( n1613 & n3033 ) ;
  assign n9237 = n7148 & ~n7252 ;
  assign n9238 = n9237 ^ n4630 ^ 1'b0 ;
  assign n9239 = n8744 | n9238 ;
  assign n9241 = n9240 ^ n9239 ^ 1'b0 ;
  assign n9242 = n449 & ~n3239 ;
  assign n9243 = ~x202 & n4365 ;
  assign n9244 = n9242 & n9243 ;
  assign n9245 = n9244 ^ n6795 ^ 1'b0 ;
  assign n9246 = n6631 ^ n3873 ^ 1'b0 ;
  assign n9247 = n6603 ^ n4278 ^ n3316 ;
  assign n9248 = x76 & ~n9247 ;
  assign n9249 = ~n2772 & n7691 ;
  assign n9255 = x72 & ~n903 ;
  assign n9256 = n9201 & n9255 ;
  assign n9257 = n9256 ^ n823 ^ 1'b0 ;
  assign n9250 = n1057 ^ x203 ^ 1'b0 ;
  assign n9251 = n1573 & ~n9250 ;
  assign n9252 = n844 | n5974 ;
  assign n9253 = n9251 | n9252 ;
  assign n9254 = n6496 & n9253 ;
  assign n9258 = n9257 ^ n9254 ^ 1'b0 ;
  assign n9259 = ( ~n302 & n3504 ) | ( ~n302 & n7134 ) | ( n3504 & n7134 ) ;
  assign n9260 = n2333 | n9259 ;
  assign n9261 = ~n3940 & n7897 ;
  assign n9262 = ~n5095 & n5710 ;
  assign n9263 = n1655 & n9262 ;
  assign n9264 = n7747 | n9263 ;
  assign n9265 = n7760 ^ n1179 ^ 1'b0 ;
  assign n9266 = n6259 ^ n3481 ^ 1'b0 ;
  assign n9267 = n9266 ^ n1579 ^ 1'b0 ;
  assign n9268 = n2121 & ~n9267 ;
  assign n9269 = n3432 & ~n4729 ;
  assign n9270 = n2355 | n3314 ;
  assign n9271 = n9270 ^ x210 ^ 1'b0 ;
  assign n9272 = n5055 & ~n8381 ;
  assign n9273 = ~n4390 & n5528 ;
  assign n9274 = n9273 ^ n4646 ^ 1'b0 ;
  assign n9275 = n2304 & n5317 ;
  assign n9276 = ~n1422 & n9275 ;
  assign n9277 = n9276 ^ n8206 ^ 1'b0 ;
  assign n9278 = n3268 ^ n2942 ^ n1847 ;
  assign n9279 = n6293 | n7006 ;
  assign n9280 = n1452 & ~n8911 ;
  assign n9281 = n5306 ^ n992 ^ 1'b0 ;
  assign n9284 = n7568 ^ n2270 ^ 1'b0 ;
  assign n9285 = n6172 & ~n9284 ;
  assign n9282 = n4398 ^ n2562 ^ n1278 ;
  assign n9283 = n9282 ^ n6462 ^ n3051 ;
  assign n9286 = n9285 ^ n9283 ^ n8967 ;
  assign n9287 = ( ~n3857 & n9212 ) | ( ~n3857 & n9233 ) | ( n9212 & n9233 ) ;
  assign n9288 = n4725 ^ n4193 ^ 1'b0 ;
  assign n9289 = x151 & n9288 ;
  assign n9290 = n8018 & n9289 ;
  assign n9291 = n2128 ^ n1805 ^ 1'b0 ;
  assign n9292 = n3690 & ~n9291 ;
  assign n9293 = n7835 & n9292 ;
  assign n9294 = n9293 ^ n6264 ^ 1'b0 ;
  assign n9296 = x251 & n545 ;
  assign n9297 = n9296 ^ n4411 ^ 1'b0 ;
  assign n9298 = n5269 & ~n9297 ;
  assign n9299 = n9298 ^ n5575 ^ 1'b0 ;
  assign n9295 = n978 ^ x17 ^ 1'b0 ;
  assign n9300 = n9299 ^ n9295 ^ 1'b0 ;
  assign n9301 = ( ~n1258 & n7895 ) | ( ~n1258 & n8660 ) | ( n7895 & n8660 ) ;
  assign n9302 = n9301 ^ n4539 ^ 1'b0 ;
  assign n9303 = n1938 | n9302 ;
  assign n9304 = n8067 | n9303 ;
  assign n9305 = n9304 ^ n8065 ^ 1'b0 ;
  assign n9306 = n6310 & n9305 ;
  assign n9307 = n308 & ~n2487 ;
  assign n9308 = n9307 ^ n6868 ^ 1'b0 ;
  assign n9309 = ~n396 & n4612 ;
  assign n9310 = n883 & ~n1427 ;
  assign n9311 = n9310 ^ n703 ^ 1'b0 ;
  assign n9312 = ( ~n266 & n1310 ) | ( ~n266 & n9311 ) | ( n1310 & n9311 ) ;
  assign n9313 = n5763 ^ x188 ^ 1'b0 ;
  assign n9314 = ~n3957 & n9313 ;
  assign n9315 = n9314 ^ n938 ^ 1'b0 ;
  assign n9316 = n9312 & ~n9315 ;
  assign n9317 = n986 ^ n539 ^ 1'b0 ;
  assign n9318 = n2909 & n9317 ;
  assign n9319 = n9318 ^ n6936 ^ 1'b0 ;
  assign n9320 = n9319 ^ n402 ^ 1'b0 ;
  assign n9321 = n6194 ^ n1197 ^ 1'b0 ;
  assign n9322 = ~n929 & n9321 ;
  assign n9323 = n1038 & n9322 ;
  assign n9324 = n5370 & ~n9323 ;
  assign n9325 = n9324 ^ n1057 ^ 1'b0 ;
  assign n9326 = ( n451 & ~n5545 ) | ( n451 & n9198 ) | ( ~n5545 & n9198 ) ;
  assign n9327 = n3945 & n9326 ;
  assign n9328 = n4619 ^ n1720 ^ 1'b0 ;
  assign n9329 = x34 & ~n9328 ;
  assign n9330 = n9329 ^ n7100 ^ 1'b0 ;
  assign n9331 = n2389 ^ n1047 ^ 1'b0 ;
  assign n9332 = n9276 ^ n4061 ^ n2788 ;
  assign n9333 = n335 & n9332 ;
  assign n9334 = n9331 & ~n9333 ;
  assign n9335 = ~n3944 & n9334 ;
  assign n9337 = n3936 ^ n1133 ^ 1'b0 ;
  assign n9336 = n2644 ^ x249 ^ 1'b0 ;
  assign n9338 = n9337 ^ n9336 ^ n1203 ;
  assign n9339 = n2257 & n3049 ;
  assign n9340 = ~n6694 & n9339 ;
  assign n9341 = ( n1200 & ~n2313 ) | ( n1200 & n5513 ) | ( ~n2313 & n5513 ) ;
  assign n9342 = n1629 & n9341 ;
  assign n9343 = ( n8315 & n9340 ) | ( n8315 & ~n9342 ) | ( n9340 & ~n9342 ) ;
  assign n9344 = n5342 ^ n5323 ^ n368 ;
  assign n9345 = n6822 ^ n4198 ^ n2837 ;
  assign n9346 = n3002 & ~n3312 ;
  assign n9347 = n2846 | n5913 ;
  assign n9348 = n9347 ^ n9273 ^ 1'b0 ;
  assign n9349 = n9346 & n9348 ;
  assign n9350 = n8354 ^ n3894 ^ n520 ;
  assign n9351 = n978 & ~n9350 ;
  assign n9352 = n5584 ^ n1962 ^ n580 ;
  assign n9353 = n9352 ^ x6 ^ 1'b0 ;
  assign n9354 = n9353 ^ x28 ^ 1'b0 ;
  assign n9355 = n4301 & n8955 ;
  assign n9356 = n9355 ^ n6459 ^ 1'b0 ;
  assign n9357 = ( n1476 & n7535 ) | ( n1476 & ~n9356 ) | ( n7535 & ~n9356 ) ;
  assign n9358 = n4306 ^ n2192 ^ n1448 ;
  assign n9359 = n8762 & ~n9358 ;
  assign n9360 = n3546 ^ n3135 ^ 1'b0 ;
  assign n9361 = ( n3633 & n6783 ) | ( n3633 & ~n9360 ) | ( n6783 & ~n9360 ) ;
  assign n9364 = n1294 ^ n500 ^ x99 ;
  assign n9365 = ( n326 & ~n723 ) | ( n326 & n9364 ) | ( ~n723 & n9364 ) ;
  assign n9366 = ~n2892 & n9365 ;
  assign n9362 = n2779 & n2831 ;
  assign n9363 = ~n2705 & n9362 ;
  assign n9367 = n9366 ^ n9363 ^ n3604 ;
  assign n9368 = n6271 & n9367 ;
  assign n9369 = ~n6833 & n9368 ;
  assign n9370 = n9369 ^ n6816 ^ n1755 ;
  assign n9371 = n933 | n9370 ;
  assign n9372 = n6326 & ~n6438 ;
  assign n9373 = ~n3100 & n9372 ;
  assign n9374 = n2482 & n4370 ;
  assign n9375 = n9374 ^ n7037 ^ 1'b0 ;
  assign n9376 = n3570 ^ n2701 ^ n549 ;
  assign n9377 = n606 & ~n6881 ;
  assign n9378 = n1635 & n2733 ;
  assign n9379 = n9378 ^ n6253 ^ n4978 ;
  assign n9380 = n7568 ^ n7336 ^ 1'b0 ;
  assign n9381 = ~n9379 & n9380 ;
  assign n9382 = n1688 | n9381 ;
  assign n9383 = ~n1166 & n1472 ;
  assign n9384 = n7733 ^ n3680 ^ 1'b0 ;
  assign n9385 = n9383 | n9384 ;
  assign n9386 = n2603 & n9385 ;
  assign n9387 = n4927 ^ x172 ^ 1'b0 ;
  assign n9388 = n5823 | n9387 ;
  assign n9389 = n9388 ^ x201 ^ 1'b0 ;
  assign n9390 = n5464 & ~n9389 ;
  assign n9391 = n1999 & n9032 ;
  assign n9392 = n9390 & n9391 ;
  assign n9393 = n6052 ^ n5135 ^ x200 ;
  assign n9394 = n9393 ^ n8435 ^ n2067 ;
  assign n9395 = n7277 | n7546 ;
  assign n9396 = n9395 ^ n2033 ^ 1'b0 ;
  assign n9404 = n1395 ^ n951 ^ n787 ;
  assign n9397 = n1110 | n3060 ;
  assign n9398 = n9397 ^ x86 ^ 1'b0 ;
  assign n9399 = ( n1262 & n3182 ) | ( n1262 & n3732 ) | ( n3182 & n3732 ) ;
  assign n9400 = ( n287 & n1206 ) | ( n287 & n6749 ) | ( n1206 & n6749 ) ;
  assign n9401 = n9399 & n9400 ;
  assign n9402 = n9401 ^ n6134 ^ 1'b0 ;
  assign n9403 = n9398 & n9402 ;
  assign n9405 = n9404 ^ n9403 ^ 1'b0 ;
  assign n9406 = n3692 ^ n966 ^ 1'b0 ;
  assign n9407 = n1378 ^ n1106 ^ 1'b0 ;
  assign n9408 = ~n3664 & n9407 ;
  assign n9409 = ~n5556 & n9408 ;
  assign n9410 = n5556 & n9409 ;
  assign n9411 = ~n1336 & n5334 ;
  assign n9412 = ( n9406 & n9410 ) | ( n9406 & n9411 ) | ( n9410 & n9411 ) ;
  assign n9413 = n1206 ^ n900 ^ 1'b0 ;
  assign n9414 = x112 & n6211 ;
  assign n9417 = n656 & n1622 ;
  assign n9416 = n6758 ^ n4396 ^ n3528 ;
  assign n9418 = n9417 ^ n9416 ^ n3275 ;
  assign n9415 = n3563 & ~n7394 ;
  assign n9419 = n9418 ^ n9415 ^ 1'b0 ;
  assign n9420 = n9228 ^ n9153 ^ 1'b0 ;
  assign n9422 = n3439 ^ n1248 ^ n966 ;
  assign n9421 = ~x146 & n1090 ;
  assign n9423 = n9422 ^ n9421 ^ n330 ;
  assign n9424 = n1705 & ~n3702 ;
  assign n9425 = n4789 ^ n1155 ^ 1'b0 ;
  assign n9426 = n3056 & n9425 ;
  assign n9427 = n7726 ^ n4242 ^ 1'b0 ;
  assign n9428 = n3402 & n9427 ;
  assign n9429 = n9428 ^ n8528 ^ 1'b0 ;
  assign n9430 = n9426 & n9429 ;
  assign n9431 = n9424 & ~n9430 ;
  assign n9432 = n2114 & n3723 ;
  assign n9433 = ~n3728 & n9432 ;
  assign n9434 = ( n1492 & ~n3797 ) | ( n1492 & n9433 ) | ( ~n3797 & n9433 ) ;
  assign n9435 = n9431 & ~n9434 ;
  assign n9436 = n9435 ^ n7791 ^ 1'b0 ;
  assign n9437 = ( ~n1716 & n3327 ) | ( ~n1716 & n8230 ) | ( n3327 & n8230 ) ;
  assign n9438 = n300 & ~n2159 ;
  assign n9439 = n9438 ^ n6016 ^ n5203 ;
  assign n9440 = n2818 & ~n9439 ;
  assign n9441 = ~n9437 & n9440 ;
  assign n9442 = n9441 ^ n1079 ^ 1'b0 ;
  assign n9443 = n1523 & n9442 ;
  assign n9444 = n4550 ^ n3561 ^ 1'b0 ;
  assign n9445 = n4655 ^ n2899 ^ 1'b0 ;
  assign n9446 = ~n3425 & n4987 ;
  assign n9447 = n9446 ^ n7115 ^ 1'b0 ;
  assign n9448 = ( n1248 & n7821 ) | ( n1248 & ~n9447 ) | ( n7821 & ~n9447 ) ;
  assign n9449 = n9448 ^ n5586 ^ n1607 ;
  assign n9450 = n1937 | n9449 ;
  assign n9451 = n3119 & ~n9450 ;
  assign n9452 = n4314 ^ n2976 ^ n1296 ;
  assign n9453 = n9452 ^ n6088 ^ n1550 ;
  assign n9454 = n2315 & n2770 ;
  assign n9457 = n256 & n1286 ;
  assign n9455 = x183 & ~n2936 ;
  assign n9456 = n9455 ^ n1849 ^ 1'b0 ;
  assign n9458 = n9457 ^ n9456 ^ n2085 ;
  assign n9459 = ( n522 & n9454 ) | ( n522 & ~n9458 ) | ( n9454 & ~n9458 ) ;
  assign n9460 = n7489 & ~n9327 ;
  assign n9461 = n1522 | n8523 ;
  assign n9462 = n4126 | n9386 ;
  assign n9463 = n9461 | n9462 ;
  assign n9464 = n4999 & ~n6374 ;
  assign n9465 = n4083 & ~n5744 ;
  assign n9466 = n9465 ^ x166 ^ 1'b0 ;
  assign n9467 = n840 ^ x74 ^ 1'b0 ;
  assign n9468 = n4236 | n8891 ;
  assign n9469 = n9422 | n9468 ;
  assign n9470 = n9467 | n9469 ;
  assign n9471 = n3549 & n9470 ;
  assign n9472 = n9466 & n9471 ;
  assign n9473 = n2903 & n4086 ;
  assign n9474 = n844 & n1586 ;
  assign n9475 = n3934 ^ n1208 ^ 1'b0 ;
  assign n9476 = n9327 ^ n7576 ^ 1'b0 ;
  assign n9477 = n9475 & n9476 ;
  assign n9478 = ( n302 & ~n4056 ) | ( n302 & n7787 ) | ( ~n4056 & n7787 ) ;
  assign n9483 = n2723 ^ n1932 ^ n794 ;
  assign n9484 = n9483 ^ n8058 ^ n2731 ;
  assign n9480 = n7070 & ~n8689 ;
  assign n9481 = n9480 ^ n1011 ^ 1'b0 ;
  assign n9482 = n6402 & ~n9481 ;
  assign n9485 = n9484 ^ n9482 ^ 1'b0 ;
  assign n9479 = ~n4323 & n9113 ;
  assign n9486 = n9485 ^ n9479 ^ 1'b0 ;
  assign n9487 = ~n9478 & n9486 ;
  assign n9488 = n9487 ^ n4793 ^ 1'b0 ;
  assign n9489 = n3093 ^ n2861 ^ 1'b0 ;
  assign n9490 = n6027 | n9489 ;
  assign n9491 = ( n4039 & n5107 ) | ( n4039 & ~n9490 ) | ( n5107 & ~n9490 ) ;
  assign n9492 = n5451 ^ n3200 ^ 1'b0 ;
  assign n9493 = n2682 ^ x213 ^ 1'b0 ;
  assign n9494 = n6027 & ~n9493 ;
  assign n9495 = n1604 & ~n9494 ;
  assign n9496 = n8466 & n9495 ;
  assign n9497 = n4767 ^ n862 ^ 1'b0 ;
  assign n9498 = ( ~n3878 & n3969 ) | ( ~n3878 & n9497 ) | ( n3969 & n9497 ) ;
  assign n9499 = n1067 & ~n5379 ;
  assign n9500 = ~n9498 & n9499 ;
  assign n9501 = n9319 ^ n9139 ^ n5437 ;
  assign n9502 = n3831 | n7252 ;
  assign n9503 = n9502 ^ x12 ^ 1'b0 ;
  assign n9504 = n9503 ^ n7378 ^ n4484 ;
  assign n9505 = ~n4767 & n8554 ;
  assign n9506 = n9505 ^ n1760 ^ 1'b0 ;
  assign n9507 = n5376 & n7404 ;
  assign n9508 = n5949 ^ n1828 ^ 1'b0 ;
  assign n9509 = ~n820 & n9508 ;
  assign n9510 = n4678 & ~n9509 ;
  assign n9511 = ( n2553 & ~n4471 ) | ( n2553 & n5686 ) | ( ~n4471 & n5686 ) ;
  assign n9512 = ( n1981 & ~n3581 ) | ( n1981 & n9240 ) | ( ~n3581 & n9240 ) ;
  assign n9513 = n5033 ^ n3312 ^ 1'b0 ;
  assign n9514 = n4013 ^ n1935 ^ n1291 ;
  assign n9515 = n3504 & ~n9514 ;
  assign n9516 = n4055 ^ n4004 ^ n1249 ;
  assign n9517 = ( n4788 & ~n9515 ) | ( n4788 & n9516 ) | ( ~n9515 & n9516 ) ;
  assign n9518 = n6392 ^ n1258 ^ 1'b0 ;
  assign n9519 = n9518 ^ n6528 ^ 1'b0 ;
  assign n9520 = n9519 ^ n8237 ^ n7613 ;
  assign n9521 = ~n603 & n7856 ;
  assign n9522 = n7970 | n9521 ;
  assign n9523 = ( ~n2275 & n4112 ) | ( ~n2275 & n5643 ) | ( n4112 & n5643 ) ;
  assign n9524 = n9523 ^ n284 ^ 1'b0 ;
  assign n9525 = x139 & n9524 ;
  assign n9526 = n827 & ~n2971 ;
  assign n9527 = n9526 ^ n9018 ^ 1'b0 ;
  assign n9529 = ( n3105 & ~n6328 ) | ( n3105 & n6846 ) | ( ~n6328 & n6846 ) ;
  assign n9528 = n2897 | n9014 ;
  assign n9530 = n9529 ^ n9528 ^ 1'b0 ;
  assign n9531 = n1940 ^ n275 ^ 1'b0 ;
  assign n9532 = n2775 & ~n9531 ;
  assign n9533 = ( ~n3696 & n6574 ) | ( ~n3696 & n9532 ) | ( n6574 & n9532 ) ;
  assign n9534 = n9533 ^ n6175 ^ n1769 ;
  assign n9538 = n6861 ^ n5805 ^ x53 ;
  assign n9539 = n9538 ^ n263 ^ 1'b0 ;
  assign n9540 = n1016 & ~n1720 ;
  assign n9541 = n6793 ^ n891 ^ 1'b0 ;
  assign n9542 = ~n409 & n9541 ;
  assign n9543 = ~n9540 & n9542 ;
  assign n9544 = n9543 ^ n5183 ^ 1'b0 ;
  assign n9545 = n9539 & n9544 ;
  assign n9546 = ( n6160 & n7749 ) | ( n6160 & n9545 ) | ( n7749 & n9545 ) ;
  assign n9535 = ~n2411 & n5904 ;
  assign n9536 = n9535 ^ n6127 ^ 1'b0 ;
  assign n9537 = n843 & ~n9536 ;
  assign n9547 = n9546 ^ n9537 ^ 1'b0 ;
  assign n9548 = ( ~n2541 & n2598 ) | ( ~n2541 & n3216 ) | ( n2598 & n3216 ) ;
  assign n9549 = n9548 ^ n2449 ^ 1'b0 ;
  assign n9550 = n2075 | n9549 ;
  assign n9551 = n932 | n9550 ;
  assign n9552 = n9551 ^ n6472 ^ n3016 ;
  assign n9553 = n5361 ^ n1709 ^ 1'b0 ;
  assign n9554 = ( n905 & ~n9552 ) | ( n905 & n9553 ) | ( ~n9552 & n9553 ) ;
  assign n9555 = n970 & n3170 ;
  assign n9556 = n6436 ^ n2092 ^ 1'b0 ;
  assign n9557 = n5721 | n9556 ;
  assign n9558 = n9557 ^ n325 ^ 1'b0 ;
  assign n9559 = ( x107 & n1335 ) | ( x107 & ~n2078 ) | ( n1335 & ~n2078 ) ;
  assign n9560 = n9559 ^ n4689 ^ x49 ;
  assign n9561 = n9560 ^ x213 ^ 1'b0 ;
  assign n9562 = ( n723 & n8406 ) | ( n723 & ~n9561 ) | ( n8406 & ~n9561 ) ;
  assign n9563 = n967 | n6750 ;
  assign n9564 = n5075 ^ n1713 ^ x197 ;
  assign n9565 = n5778 & n8778 ;
  assign n9566 = n9564 & n9565 ;
  assign n9567 = n5927 ^ n1603 ^ n1580 ;
  assign n9568 = ( n1927 & ~n4273 ) | ( n1927 & n5925 ) | ( ~n4273 & n5925 ) ;
  assign n9569 = ( n2940 & ~n3156 ) | ( n2940 & n8363 ) | ( ~n3156 & n8363 ) ;
  assign n9570 = n6764 | n9569 ;
  assign n9571 = n435 | n9570 ;
  assign n9572 = n5112 ^ n2822 ^ 1'b0 ;
  assign n9573 = n9572 ^ n8924 ^ 1'b0 ;
  assign n9574 = n4668 | n9573 ;
  assign n9575 = ~n2459 & n9574 ;
  assign n9576 = n9575 ^ n8356 ^ 1'b0 ;
  assign n9577 = n706 & n7062 ;
  assign n9578 = n4600 ^ n3097 ^ 1'b0 ;
  assign n9579 = ( n1013 & n3842 ) | ( n1013 & ~n6133 ) | ( n3842 & ~n6133 ) ;
  assign n9580 = ~n1503 & n9579 ;
  assign n9585 = n4221 & n5567 ;
  assign n9586 = n9585 ^ n7282 ^ 1'b0 ;
  assign n9587 = ( n3439 & n4342 ) | ( n3439 & n9586 ) | ( n4342 & n9586 ) ;
  assign n9581 = n3187 & ~n5276 ;
  assign n9582 = n9581 ^ n5698 ^ x134 ;
  assign n9583 = ~n4913 & n9582 ;
  assign n9584 = n7227 | n9583 ;
  assign n9588 = n9587 ^ n9584 ^ 1'b0 ;
  assign n9589 = n9588 ^ n5281 ^ 1'b0 ;
  assign n9590 = n9580 | n9589 ;
  assign n9591 = ( x189 & n7176 ) | ( x189 & n9014 ) | ( n7176 & n9014 ) ;
  assign n9592 = n4448 | n9591 ;
  assign n9593 = n6592 & n8228 ;
  assign n9594 = n1975 ^ n1617 ^ 1'b0 ;
  assign n9595 = n6824 ^ n1835 ^ 1'b0 ;
  assign n9596 = n3086 & ~n9595 ;
  assign n9597 = ( ~n5201 & n7894 ) | ( ~n5201 & n9596 ) | ( n7894 & n9596 ) ;
  assign n9598 = ~n7142 & n9597 ;
  assign n9599 = n6754 & n9598 ;
  assign n9604 = ( ~n2059 & n3659 ) | ( ~n2059 & n3880 ) | ( n3659 & n3880 ) ;
  assign n9600 = ( n2589 & n5353 ) | ( n2589 & n7715 ) | ( n5353 & n7715 ) ;
  assign n9601 = n2469 & n4434 ;
  assign n9602 = n9601 ^ n9230 ^ 1'b0 ;
  assign n9603 = n9600 & n9602 ;
  assign n9605 = n9604 ^ n9603 ^ 1'b0 ;
  assign n9606 = n9605 ^ n8303 ^ 1'b0 ;
  assign n9607 = n3571 ^ n3531 ^ n1740 ;
  assign n9608 = x112 & n949 ;
  assign n9609 = n2106 & n3962 ;
  assign n9610 = n9609 ^ n4686 ^ 1'b0 ;
  assign n9611 = ( ~n2167 & n2567 ) | ( ~n2167 & n7613 ) | ( n2567 & n7613 ) ;
  assign n9612 = ( n6448 & n9610 ) | ( n6448 & n9611 ) | ( n9610 & n9611 ) ;
  assign n9613 = n2566 | n3755 ;
  assign n9614 = n2520 & ~n9613 ;
  assign n9615 = ( n4332 & ~n7304 ) | ( n4332 & n9614 ) | ( ~n7304 & n9614 ) ;
  assign n9616 = n4308 ^ n1781 ^ 1'b0 ;
  assign n9617 = ~n2429 & n9616 ;
  assign n9623 = n3820 | n3869 ;
  assign n9619 = n2003 | n2897 ;
  assign n9620 = n3797 & ~n9619 ;
  assign n9621 = n2100 | n9620 ;
  assign n9622 = n9621 ^ n5659 ^ 1'b0 ;
  assign n9624 = n9623 ^ n9622 ^ n2984 ;
  assign n9618 = ( n1635 & ~n2478 ) | ( n1635 & n7488 ) | ( ~n2478 & n7488 ) ;
  assign n9625 = n9624 ^ n9618 ^ 1'b0 ;
  assign n9626 = n3226 | n9625 ;
  assign n9628 = n2838 ^ n433 ^ 1'b0 ;
  assign n9627 = ( n440 & ~n3426 ) | ( n440 & n6054 ) | ( ~n3426 & n6054 ) ;
  assign n9629 = n9628 ^ n9627 ^ 1'b0 ;
  assign n9630 = n7646 | n9629 ;
  assign n9631 = n3206 ^ n567 ^ n513 ;
  assign n9634 = n2769 & ~n8114 ;
  assign n9632 = n7362 ^ n1505 ^ 1'b0 ;
  assign n9633 = ~n4628 & n9632 ;
  assign n9635 = n9634 ^ n9633 ^ 1'b0 ;
  assign n9636 = n2510 & ~n4263 ;
  assign n9637 = n2032 & n9636 ;
  assign n9638 = n9637 ^ n1296 ^ 1'b0 ;
  assign n9639 = n3104 | n9638 ;
  assign n9640 = n9635 | n9639 ;
  assign n9641 = n3404 & n4369 ;
  assign n9642 = n2718 ^ n661 ^ 1'b0 ;
  assign n9643 = n9642 ^ n8004 ^ n752 ;
  assign n9644 = n7745 & ~n9643 ;
  assign n9645 = ( ~n2953 & n3187 ) | ( ~n2953 & n9644 ) | ( n3187 & n9644 ) ;
  assign n9646 = ~n9641 & n9645 ;
  assign n9647 = n9646 ^ n5297 ^ 1'b0 ;
  assign n9648 = n1463 & n9647 ;
  assign n9649 = n2742 & n9648 ;
  assign n9650 = n3222 & ~n8222 ;
  assign n9651 = n3800 & ~n5265 ;
  assign n9652 = n9651 ^ n2817 ^ 1'b0 ;
  assign n9653 = ~n1166 & n9652 ;
  assign n9654 = n4638 | n9516 ;
  assign n9655 = n5770 ^ n2793 ^ 1'b0 ;
  assign n9656 = n3731 & ~n9655 ;
  assign n9657 = ~n5165 & n9656 ;
  assign n9658 = n4109 & n9657 ;
  assign n9659 = ~n1306 & n4999 ;
  assign n9660 = ( n4913 & ~n7893 ) | ( n4913 & n9659 ) | ( ~n7893 & n9659 ) ;
  assign n9661 = n1763 ^ n816 ^ 1'b0 ;
  assign n9662 = n1696 & n9661 ;
  assign n9667 = n8404 | n9000 ;
  assign n9668 = n9667 ^ n1597 ^ 1'b0 ;
  assign n9664 = n2675 ^ n1516 ^ n922 ;
  assign n9665 = ~n2157 & n9664 ;
  assign n9663 = n4929 & n5763 ;
  assign n9666 = n9665 ^ n9663 ^ 1'b0 ;
  assign n9669 = n9668 ^ n9666 ^ 1'b0 ;
  assign n9670 = x209 & ~n9669 ;
  assign n9671 = n9662 & n9670 ;
  assign n9672 = ~n3378 & n9671 ;
  assign n9673 = n6330 ^ n904 ^ 1'b0 ;
  assign n9674 = ~n1145 & n7236 ;
  assign n9675 = n9674 ^ n2256 ^ 1'b0 ;
  assign n9676 = n4203 ^ n2005 ^ n1266 ;
  assign n9677 = n9676 ^ n4346 ^ n1239 ;
  assign n9681 = n2217 & n2506 ;
  assign n9680 = n2723 & ~n3439 ;
  assign n9682 = n9681 ^ n9680 ^ 1'b0 ;
  assign n9678 = n862 & ~n2095 ;
  assign n9679 = n415 & ~n9678 ;
  assign n9683 = n9682 ^ n9679 ^ 1'b0 ;
  assign n9684 = x2 & n1849 ;
  assign n9685 = n9684 ^ x103 ^ 1'b0 ;
  assign n9686 = n9685 ^ n2389 ^ 1'b0 ;
  assign n9687 = n5039 & ~n9686 ;
  assign n9688 = n9687 ^ n9250 ^ 1'b0 ;
  assign n9689 = n1320 | n9688 ;
  assign n9690 = n9689 ^ n5689 ^ 1'b0 ;
  assign n9691 = ~n9683 & n9690 ;
  assign n9692 = n904 & n9691 ;
  assign n9693 = n4528 | n6018 ;
  assign n9694 = n9693 ^ n3519 ^ 1'b0 ;
  assign n9695 = n9694 ^ n6551 ^ 1'b0 ;
  assign n9696 = n6436 ^ n3924 ^ n2828 ;
  assign n9697 = ~n6952 & n9696 ;
  assign n9698 = ~n3233 & n9697 ;
  assign n9699 = ~n4027 & n7337 ;
  assign n9700 = n9699 ^ n4690 ^ 1'b0 ;
  assign n9701 = n6491 | n9700 ;
  assign n9702 = n7788 ^ n3550 ^ 1'b0 ;
  assign n9703 = n9702 ^ n325 ^ 1'b0 ;
  assign n9704 = ~n9701 & n9703 ;
  assign n9705 = n9704 ^ n6274 ^ 1'b0 ;
  assign n9708 = n7824 ^ n980 ^ n715 ;
  assign n9706 = n4840 ^ n4314 ^ 1'b0 ;
  assign n9707 = n4997 | n9706 ;
  assign n9709 = n9708 ^ n9707 ^ 1'b0 ;
  assign n9710 = n6465 ^ n1448 ^ 1'b0 ;
  assign n9711 = n9710 ^ n2294 ^ 1'b0 ;
  assign n9712 = ~n9709 & n9711 ;
  assign n9713 = x182 & n6942 ;
  assign n9714 = n9713 ^ n4294 ^ 1'b0 ;
  assign n9715 = n6322 & ~n9714 ;
  assign n9716 = n9715 ^ x156 ^ 1'b0 ;
  assign n9717 = n9611 ^ n5818 ^ 1'b0 ;
  assign n9720 = x163 & n4740 ;
  assign n9721 = n4022 & n9720 ;
  assign n9722 = n9721 ^ n3674 ^ 1'b0 ;
  assign n9723 = n763 | n9722 ;
  assign n9719 = n2660 ^ n2238 ^ n1042 ;
  assign n9718 = n7466 ^ n5993 ^ 1'b0 ;
  assign n9724 = n9723 ^ n9719 ^ n9718 ;
  assign n9728 = n669 & ~n3060 ;
  assign n9729 = n9728 ^ x39 ^ 1'b0 ;
  assign n9726 = ( n2092 & n4053 ) | ( n2092 & ~n6913 ) | ( n4053 & ~n6913 ) ;
  assign n9727 = n2179 | n9726 ;
  assign n9730 = n9729 ^ n9727 ^ 1'b0 ;
  assign n9725 = ~n1203 & n7990 ;
  assign n9731 = n9730 ^ n9725 ^ 1'b0 ;
  assign n9732 = n5072 ^ n1800 ^ 1'b0 ;
  assign n9733 = n6781 | n9732 ;
  assign n9734 = n8412 & ~n9733 ;
  assign n9735 = n6094 & ~n7837 ;
  assign n9737 = ( n1362 & n1479 ) | ( n1362 & ~n2006 ) | ( n1479 & ~n2006 ) ;
  assign n9736 = n998 | n3819 ;
  assign n9738 = n9737 ^ n9736 ^ 1'b0 ;
  assign n9739 = n913 & ~n3408 ;
  assign n9740 = x121 & n957 ;
  assign n9741 = ~n9739 & n9740 ;
  assign n9742 = n9431 ^ n9155 ^ n7190 ;
  assign n9743 = n5612 ^ n1108 ^ n1032 ;
  assign n9744 = n1995 & ~n4254 ;
  assign n9745 = n9744 ^ n2036 ^ 1'b0 ;
  assign n9746 = ( n4437 & ~n9743 ) | ( n4437 & n9745 ) | ( ~n9743 & n9745 ) ;
  assign n9747 = ~n5513 & n9605 ;
  assign n9748 = n8192 ^ n3915 ^ 1'b0 ;
  assign n9749 = n801 & ~n9748 ;
  assign n9750 = ~n4319 & n6783 ;
  assign n9751 = n9750 ^ n9578 ^ n6330 ;
  assign n9752 = n1353 & ~n1450 ;
  assign n9753 = n8375 ^ n2473 ^ 1'b0 ;
  assign n9754 = n2461 & n9753 ;
  assign n9755 = ( ~n550 & n5598 ) | ( ~n550 & n9754 ) | ( n5598 & n9754 ) ;
  assign n9756 = ( n2332 & n9752 ) | ( n2332 & ~n9755 ) | ( n9752 & ~n9755 ) ;
  assign n9757 = n7220 ^ n6945 ^ 1'b0 ;
  assign n9758 = n514 & n2833 ;
  assign n9759 = n9758 ^ n3977 ^ 1'b0 ;
  assign n9760 = ~n9064 & n9759 ;
  assign n9761 = n9757 & n9760 ;
  assign n9762 = ~n6227 & n9761 ;
  assign n9763 = n3100 & n9037 ;
  assign n9764 = n9763 ^ x226 ^ 1'b0 ;
  assign n9765 = n2207 & n9764 ;
  assign n9766 = n9765 ^ n5319 ^ 1'b0 ;
  assign n9767 = n5123 & n9766 ;
  assign n9768 = n4303 ^ n2703 ^ n453 ;
  assign n9769 = n2640 ^ n1468 ^ 1'b0 ;
  assign n9770 = ~n3649 & n9769 ;
  assign n9771 = n3383 ^ n877 ^ 1'b0 ;
  assign n9772 = n1780 & n9771 ;
  assign n9773 = n2443 & n9772 ;
  assign n9774 = n300 & ~n1916 ;
  assign n9775 = ~n1657 & n9774 ;
  assign n9776 = ( ~n1856 & n4915 ) | ( ~n1856 & n9775 ) | ( n4915 & n9775 ) ;
  assign n9777 = n4838 ^ n1940 ^ n257 ;
  assign n9778 = ( ~n4090 & n9776 ) | ( ~n4090 & n9777 ) | ( n9776 & n9777 ) ;
  assign n9779 = ( n9770 & ~n9773 ) | ( n9770 & n9778 ) | ( ~n9773 & n9778 ) ;
  assign n9780 = ~n1418 & n5671 ;
  assign n9781 = n9780 ^ n1267 ^ 1'b0 ;
  assign n9782 = n4398 & n9781 ;
  assign n9783 = n7966 ^ n2117 ^ 1'b0 ;
  assign n9784 = n5999 ^ n3770 ^ 1'b0 ;
  assign n9785 = ~n3848 & n9784 ;
  assign n9786 = n1618 | n9707 ;
  assign n9787 = n4245 | n9786 ;
  assign n9788 = n1853 & n5408 ;
  assign n9789 = ( n1022 & n4212 ) | ( n1022 & n8214 ) | ( n4212 & n8214 ) ;
  assign n9790 = ~n4018 & n9789 ;
  assign n9791 = n9790 ^ n1010 ^ 1'b0 ;
  assign n9792 = n4661 & ~n9791 ;
  assign n9793 = x205 & n8508 ;
  assign n9794 = n9793 ^ n8017 ^ n2783 ;
  assign n9795 = n1739 & n9794 ;
  assign n9796 = n621 & ~n9795 ;
  assign n9797 = n9527 & n9796 ;
  assign n9798 = n6560 & ~n7758 ;
  assign n9799 = n7163 & n9798 ;
  assign n9800 = n6043 ^ n6031 ^ 1'b0 ;
  assign n9801 = n4392 | n9800 ;
  assign n9802 = ( n3424 & ~n9799 ) | ( n3424 & n9801 ) | ( ~n9799 & n9801 ) ;
  assign n9805 = n1493 ^ n1397 ^ 1'b0 ;
  assign n9806 = n4379 & n9805 ;
  assign n9803 = n4806 | n9301 ;
  assign n9804 = n5998 | n9803 ;
  assign n9807 = n9806 ^ n9804 ^ 1'b0 ;
  assign n9808 = n4705 & n9807 ;
  assign n9809 = n9802 & n9808 ;
  assign n9810 = x160 & ~n949 ;
  assign n9811 = n1684 & n9810 ;
  assign n9812 = n9811 ^ n6289 ^ n4065 ;
  assign n9813 = n5078 & n5801 ;
  assign n9814 = n1037 & n9813 ;
  assign n9815 = ( x66 & ~n2319 ) | ( x66 & n2408 ) | ( ~n2319 & n2408 ) ;
  assign n9816 = ( n1534 & ~n2425 ) | ( n1534 & n9815 ) | ( ~n2425 & n9815 ) ;
  assign n9817 = ~n9814 & n9816 ;
  assign n9818 = ~n4322 & n9817 ;
  assign n9819 = n5736 | n7370 ;
  assign n9820 = n2897 & ~n9819 ;
  assign n9821 = n5070 ^ n447 ^ 1'b0 ;
  assign n9822 = n9820 | n9821 ;
  assign n9823 = n9822 ^ n1051 ^ 1'b0 ;
  assign n9824 = ( n3483 & n9818 ) | ( n3483 & ~n9823 ) | ( n9818 & ~n9823 ) ;
  assign n9825 = n9812 & ~n9824 ;
  assign n9826 = ~n6170 & n9825 ;
  assign n9827 = n9025 ^ n6408 ^ 1'b0 ;
  assign n9828 = n5020 & ~n6677 ;
  assign n9829 = ( ~n7747 & n9198 ) | ( ~n7747 & n9297 ) | ( n9198 & n9297 ) ;
  assign n9830 = n7132 ^ n3521 ^ n2035 ;
  assign n9831 = ( n2174 & n3030 ) | ( n2174 & ~n9230 ) | ( n3030 & ~n9230 ) ;
  assign n9832 = n4703 ^ n2534 ^ n950 ;
  assign n9833 = ~n9831 & n9832 ;
  assign n9834 = ~n2098 & n9833 ;
  assign n9835 = ~n277 & n1257 ;
  assign n9836 = n5588 & ~n6306 ;
  assign n9837 = ( n7125 & n7568 ) | ( n7125 & n9836 ) | ( n7568 & n9836 ) ;
  assign n9838 = ( n1172 & n9835 ) | ( n1172 & ~n9837 ) | ( n9835 & ~n9837 ) ;
  assign n9839 = n9838 ^ n2766 ^ n2538 ;
  assign n9840 = n5583 ^ n4039 ^ n2543 ;
  assign n9841 = n8985 ^ n2595 ^ n1644 ;
  assign n9842 = ( n3859 & ~n9840 ) | ( n3859 & n9841 ) | ( ~n9840 & n9841 ) ;
  assign n9843 = n7840 ^ n2125 ^ 1'b0 ;
  assign n9844 = n6711 ^ n3990 ^ 1'b0 ;
  assign n9845 = ( n1732 & ~n7971 ) | ( n1732 & n9417 ) | ( ~n7971 & n9417 ) ;
  assign n9846 = n8084 ^ n2885 ^ 1'b0 ;
  assign n9847 = n1933 & n2496 ;
  assign n9848 = n9847 ^ n8930 ^ 1'b0 ;
  assign n9849 = ~n2780 & n9848 ;
  assign n9850 = n2651 & ~n3037 ;
  assign n9851 = n5472 ^ n4303 ^ n1554 ;
  assign n9852 = n5793 & n9851 ;
  assign n9853 = n382 & n993 ;
  assign n9854 = ~n8365 & n9853 ;
  assign n9855 = n9854 ^ n4026 ^ 1'b0 ;
  assign n9856 = ~n6846 & n9099 ;
  assign n9857 = n9856 ^ n3583 ^ 1'b0 ;
  assign n9858 = n7686 & ~n9857 ;
  assign n9859 = ( x87 & n1873 ) | ( x87 & n7055 ) | ( n1873 & n7055 ) ;
  assign n9860 = n9859 ^ n5739 ^ 1'b0 ;
  assign n9861 = n292 & ~n6745 ;
  assign n9862 = n5001 | n9861 ;
  assign n9863 = n3223 & ~n9862 ;
  assign n9864 = n5153 & ~n9863 ;
  assign n9865 = n2874 ^ n428 ^ 1'b0 ;
  assign n9866 = n2339 & ~n9865 ;
  assign n9867 = n2951 ^ n1810 ^ 1'b0 ;
  assign n9868 = n5339 & n9867 ;
  assign n9869 = n4815 & ~n9868 ;
  assign n9870 = n9869 ^ n958 ^ 1'b0 ;
  assign n9871 = n9866 & ~n9870 ;
  assign n9872 = n9732 ^ n8188 ^ n3181 ;
  assign n9873 = n1530 | n5852 ;
  assign n9874 = n9873 ^ n6337 ^ n2381 ;
  assign n9875 = n7987 ^ n5579 ^ n1239 ;
  assign n9876 = n2496 & ~n3279 ;
  assign n9877 = n2023 & n9876 ;
  assign n9878 = n9877 ^ n8725 ^ n8722 ;
  assign n9879 = n9878 ^ n7976 ^ n4214 ;
  assign n9880 = ( n9874 & ~n9875 ) | ( n9874 & n9879 ) | ( ~n9875 & n9879 ) ;
  assign n9883 = x231 & ~n1724 ;
  assign n9884 = ~n2396 & n9883 ;
  assign n9885 = n9884 ^ n1810 ^ 1'b0 ;
  assign n9881 = n9378 ^ n5631 ^ 1'b0 ;
  assign n9882 = n9881 ^ n5133 ^ n1766 ;
  assign n9886 = n9885 ^ n9882 ^ 1'b0 ;
  assign n9887 = n9608 ^ n1616 ^ 1'b0 ;
  assign n9888 = n2656 ^ n489 ^ 1'b0 ;
  assign n9889 = n7716 & ~n9888 ;
  assign n9890 = n8398 ^ n7047 ^ n482 ;
  assign n9891 = n920 | n1308 ;
  assign n9892 = n8181 ^ n6016 ^ n2845 ;
  assign n9893 = n9892 ^ n464 ^ 1'b0 ;
  assign n9894 = n763 | n9893 ;
  assign n9895 = n2643 & ~n7777 ;
  assign n9896 = n9895 ^ n7509 ^ 1'b0 ;
  assign n9897 = n5397 ^ n4889 ^ 1'b0 ;
  assign n9898 = n3597 & n7690 ;
  assign n9899 = n9897 | n9898 ;
  assign n9900 = n6851 ^ n4353 ^ 1'b0 ;
  assign n9901 = n2403 & ~n9900 ;
  assign n9902 = ( n3433 & n4089 ) | ( n3433 & n9901 ) | ( n4089 & n9901 ) ;
  assign n9903 = n5090 & ~n5737 ;
  assign n9904 = x27 | n9903 ;
  assign n9905 = n6086 ^ n3939 ^ 1'b0 ;
  assign n9906 = x12 & ~n9905 ;
  assign n9907 = n4128 | n9906 ;
  assign n9908 = n9907 ^ n7530 ^ n6001 ;
  assign n9909 = ~n7848 & n9908 ;
  assign n9910 = n9909 ^ n9358 ^ 1'b0 ;
  assign n9912 = n2672 & n5903 ;
  assign n9913 = n1105 & n9912 ;
  assign n9911 = n2173 & n4722 ;
  assign n9914 = n9913 ^ n9911 ^ 1'b0 ;
  assign n9917 = n4685 ^ n4115 ^ n518 ;
  assign n9915 = n7481 ^ n1487 ^ 1'b0 ;
  assign n9916 = x238 & ~n9915 ;
  assign n9918 = n9917 ^ n9916 ^ 1'b0 ;
  assign n9919 = n6160 ^ n3066 ^ n2414 ;
  assign n9920 = n7978 & ~n9919 ;
  assign n9921 = n9365 & n9920 ;
  assign n9922 = ( n792 & n6201 ) | ( n792 & ~n7216 ) | ( n6201 & ~n7216 ) ;
  assign n9923 = n2334 ^ n479 ^ 1'b0 ;
  assign n9924 = ~n817 & n9923 ;
  assign n9925 = ( n3390 & ~n9922 ) | ( n3390 & n9924 ) | ( ~n9922 & n9924 ) ;
  assign n9926 = n7902 ^ x21 ^ 1'b0 ;
  assign n9927 = n5725 | n9926 ;
  assign n9928 = n9925 & n9927 ;
  assign n9929 = n4013 ^ n2691 ^ n2437 ;
  assign n9930 = n4699 & ~n9929 ;
  assign n9931 = n5755 & n9930 ;
  assign n9932 = n9538 & ~n9931 ;
  assign n9933 = n5886 ^ n5874 ^ n2538 ;
  assign n9934 = n4388 ^ n3630 ^ n1734 ;
  assign n9935 = n9934 ^ n3978 ^ 1'b0 ;
  assign n9936 = ~n9933 & n9935 ;
  assign n9937 = n6448 ^ n986 ^ 1'b0 ;
  assign n9938 = n8183 | n9937 ;
  assign n9939 = n7416 | n9938 ;
  assign n9944 = n9561 ^ n545 ^ 1'b0 ;
  assign n9945 = n9944 ^ n6167 ^ n4901 ;
  assign n9940 = n6170 ^ n1035 ^ 1'b0 ;
  assign n9941 = n2740 | n9940 ;
  assign n9942 = n9941 ^ n6048 ^ 1'b0 ;
  assign n9943 = ~n7011 & n9942 ;
  assign n9946 = n9945 ^ n9943 ^ 1'b0 ;
  assign n9947 = n9464 & n9946 ;
  assign n9951 = n2247 & ~n7638 ;
  assign n9952 = ~n436 & n9951 ;
  assign n9953 = ( n682 & ~n4029 ) | ( n682 & n9952 ) | ( ~n4029 & n9952 ) ;
  assign n9948 = n6715 ^ n4437 ^ n3865 ;
  assign n9949 = n9948 ^ n7269 ^ n3702 ;
  assign n9950 = ~n9246 & n9949 ;
  assign n9954 = n9953 ^ n9950 ^ 1'b0 ;
  assign n9955 = n6418 & ~n9954 ;
  assign n9956 = n9318 ^ n4985 ^ 1'b0 ;
  assign n9957 = n2405 & n9956 ;
  assign n9958 = n748 & n2222 ;
  assign n9959 = n9958 ^ n9518 ^ 1'b0 ;
  assign n9960 = n9957 & n9959 ;
  assign n9961 = n1366 & ~n6242 ;
  assign n9962 = n9551 ^ n7296 ^ 1'b0 ;
  assign n9963 = ~n6783 & n9962 ;
  assign n9964 = n9963 ^ n6813 ^ 1'b0 ;
  assign n9965 = ~n2131 & n2640 ;
  assign n9966 = n9965 ^ n4005 ^ 1'b0 ;
  assign n9967 = n9966 ^ n7353 ^ 1'b0 ;
  assign n9968 = n3781 & n9967 ;
  assign n9969 = ~n8507 & n9968 ;
  assign n9970 = n1042 | n5430 ;
  assign n9971 = n7014 & ~n9970 ;
  assign n9972 = ( n1291 & n4127 ) | ( n1291 & n9971 ) | ( n4127 & n9971 ) ;
  assign n9973 = ~n9969 & n9972 ;
  assign n9974 = n9973 ^ n2312 ^ 1'b0 ;
  assign n9975 = n5110 & n5156 ;
  assign n9976 = n9975 ^ n5676 ^ 1'b0 ;
  assign n9977 = n2073 & n9976 ;
  assign n9978 = n9974 & n9977 ;
  assign n9979 = n2256 & ~n7008 ;
  assign n9980 = ~n6379 & n9979 ;
  assign n9981 = n9564 ^ n7265 ^ 1'b0 ;
  assign n9982 = n1877 ^ x195 ^ 1'b0 ;
  assign n9983 = n3872 ^ n2817 ^ 1'b0 ;
  assign n9986 = n1609 ^ n1126 ^ 1'b0 ;
  assign n9984 = n3961 ^ n2217 ^ 1'b0 ;
  assign n9985 = n9644 | n9984 ;
  assign n9987 = n9986 ^ n9985 ^ n8639 ;
  assign n9988 = n9688 ^ n3716 ^ n3457 ;
  assign n9989 = n1909 & n9988 ;
  assign n9990 = n9989 ^ n3027 ^ 1'b0 ;
  assign n9991 = n6758 ^ n2258 ^ 1'b0 ;
  assign n9992 = n5313 ^ n3641 ^ n1482 ;
  assign n9993 = n5626 & n9168 ;
  assign n9994 = n3796 | n9921 ;
  assign n9995 = n9994 ^ n4148 ^ 1'b0 ;
  assign n9996 = n7737 ^ n5075 ^ 1'b0 ;
  assign n9998 = n9659 ^ n2128 ^ x159 ;
  assign n9997 = ( n2296 & n5020 ) | ( n2296 & ~n9596 ) | ( n5020 & ~n9596 ) ;
  assign n9999 = n9998 ^ n9997 ^ 1'b0 ;
  assign n10000 = n7399 & n9999 ;
  assign n10001 = n1976 | n7358 ;
  assign n10002 = n5106 ^ n2278 ^ n998 ;
  assign n10003 = ( ~n3117 & n4287 ) | ( ~n3117 & n5325 ) | ( n4287 & n5325 ) ;
  assign n10004 = n9037 & n10003 ;
  assign n10005 = n10004 ^ n2825 ^ 1'b0 ;
  assign n10006 = n3185 & ~n5666 ;
  assign n10007 = n10006 ^ n3464 ^ 1'b0 ;
  assign n10008 = ~n2179 & n6555 ;
  assign n10009 = n10007 & n10008 ;
  assign n10010 = ( ~n469 & n884 ) | ( ~n469 & n3814 ) | ( n884 & n3814 ) ;
  assign n10011 = n1168 & n10010 ;
  assign n10012 = n7961 ^ n3766 ^ 1'b0 ;
  assign n10013 = n1022 | n10012 ;
  assign n10014 = n10013 ^ n2790 ^ 1'b0 ;
  assign n10015 = ~n10011 & n10014 ;
  assign n10016 = ~n955 & n10015 ;
  assign n10017 = ( n3064 & n4677 ) | ( n3064 & ~n10016 ) | ( n4677 & ~n10016 ) ;
  assign n10018 = ~n10009 & n10017 ;
  assign n10019 = n10005 & n10018 ;
  assign n10020 = ~n10002 & n10019 ;
  assign n10021 = n1352 & ~n3909 ;
  assign n10022 = x218 | n6043 ;
  assign n10023 = n10021 | n10022 ;
  assign n10024 = ( n1274 & n1345 ) | ( n1274 & ~n3924 ) | ( n1345 & ~n3924 ) ;
  assign n10025 = ~n2680 & n8238 ;
  assign n10026 = n10024 & ~n10025 ;
  assign n10027 = ~n2287 & n4132 ;
  assign n10028 = ~x1 & n10027 ;
  assign n10029 = n5128 | n9803 ;
  assign n10030 = n2130 & ~n10029 ;
  assign n10031 = ( n1628 & ~n1853 ) | ( n1628 & n2636 ) | ( ~n1853 & n2636 ) ;
  assign n10032 = x81 & n1199 ;
  assign n10033 = n10031 & n10032 ;
  assign n10034 = n10033 ^ n4039 ^ 1'b0 ;
  assign n10035 = n4045 & n4177 ;
  assign n10036 = n10034 & n10035 ;
  assign n10037 = n10030 | n10036 ;
  assign n10038 = n10037 ^ x64 ^ 1'b0 ;
  assign n10039 = ( n6070 & n10028 ) | ( n6070 & n10038 ) | ( n10028 & n10038 ) ;
  assign n10040 = n2028 ^ n500 ^ 1'b0 ;
  assign n10041 = n5850 & n10040 ;
  assign n10042 = ( n1457 & n4438 ) | ( n1457 & n10041 ) | ( n4438 & n10041 ) ;
  assign n10043 = n6627 ^ n1963 ^ 1'b0 ;
  assign n10044 = x189 & n10043 ;
  assign n10045 = n10044 ^ n3970 ^ n825 ;
  assign n10046 = x82 & n10045 ;
  assign n10047 = x182 & ~n604 ;
  assign n10048 = n10047 ^ n2819 ^ 1'b0 ;
  assign n10049 = n2055 & n10048 ;
  assign n10050 = n2968 & n10049 ;
  assign n10051 = n8924 | n10050 ;
  assign n10052 = n3248 & ~n10051 ;
  assign n10053 = n4946 ^ n1787 ^ n807 ;
  assign n10054 = ( n2878 & ~n7482 ) | ( n2878 & n10053 ) | ( ~n7482 & n10053 ) ;
  assign n10055 = ~n1160 & n3746 ;
  assign n10056 = n10055 ^ n6922 ^ n1442 ;
  assign n10057 = ~n10054 & n10056 ;
  assign n10058 = n10052 & n10057 ;
  assign n10059 = n5657 ^ n4577 ^ x0 ;
  assign n10060 = n821 ^ n771 ^ 1'b0 ;
  assign n10061 = n1770 & ~n10060 ;
  assign n10062 = n6518 ^ n3322 ^ 1'b0 ;
  assign n10063 = n10062 ^ n4685 ^ n2769 ;
  assign n10064 = n10063 ^ n3069 ^ n775 ;
  assign n10065 = n5805 ^ n3404 ^ n955 ;
  assign n10066 = n824 & ~n4162 ;
  assign n10067 = n10066 ^ n3905 ^ 1'b0 ;
  assign n10068 = n9783 | n10067 ;
  assign n10069 = n3261 & n3853 ;
  assign n10070 = n10069 ^ n9818 ^ 1'b0 ;
  assign n10071 = n5328 ^ n3540 ^ 1'b0 ;
  assign n10072 = n1604 & ~n3953 ;
  assign n10074 = n7788 ^ n1641 ^ 1'b0 ;
  assign n10075 = ~n8300 & n10074 ;
  assign n10073 = n6441 ^ n3042 ^ n2771 ;
  assign n10076 = n10075 ^ n10073 ^ 1'b0 ;
  assign n10077 = n2498 & ~n3145 ;
  assign n10078 = n10076 & n10077 ;
  assign n10080 = n5732 ^ n3240 ^ n1074 ;
  assign n10079 = n1237 & ~n9319 ;
  assign n10081 = n10080 ^ n10079 ^ 1'b0 ;
  assign n10082 = n10081 ^ n8913 ^ 1'b0 ;
  assign n10083 = n1602 ^ n1107 ^ 1'b0 ;
  assign n10084 = n3599 & n10083 ;
  assign n10085 = n3050 ^ n2806 ^ n2502 ;
  assign n10086 = ( x39 & x100 ) | ( x39 & n9247 ) | ( x100 & n9247 ) ;
  assign n10087 = n10085 & n10086 ;
  assign n10088 = ( n6858 & n10084 ) | ( n6858 & n10087 ) | ( n10084 & n10087 ) ;
  assign n10089 = n1907 | n2509 ;
  assign n10090 = n10089 ^ n5451 ^ n3233 ;
  assign n10091 = n6876 ^ n2831 ^ 1'b0 ;
  assign n10092 = n5453 ^ n2572 ^ 1'b0 ;
  assign n10093 = n10092 ^ n3379 ^ 1'b0 ;
  assign n10094 = n2522 ^ n1350 ^ 1'b0 ;
  assign n10095 = ( n2264 & n3110 ) | ( n2264 & ~n10094 ) | ( n3110 & ~n10094 ) ;
  assign n10096 = n10095 ^ n8149 ^ 1'b0 ;
  assign n10098 = x251 & ~n2650 ;
  assign n10099 = n10098 ^ n7289 ^ 1'b0 ;
  assign n10097 = n2174 & n7813 ;
  assign n10100 = n10099 ^ n10097 ^ 1'b0 ;
  assign n10101 = ( n1039 & ~n10096 ) | ( n1039 & n10100 ) | ( ~n10096 & n10100 ) ;
  assign n10102 = n5275 ^ n1578 ^ 1'b0 ;
  assign n10103 = n10102 ^ n3944 ^ 1'b0 ;
  assign n10104 = n1204 | n10103 ;
  assign n10108 = n3808 ^ n2043 ^ n1418 ;
  assign n10109 = n1495 ^ n264 ^ 1'b0 ;
  assign n10110 = n10109 ^ n5803 ^ 1'b0 ;
  assign n10111 = n10108 & ~n10110 ;
  assign n10112 = ( n877 & ~n8861 ) | ( n877 & n10111 ) | ( ~n8861 & n10111 ) ;
  assign n10105 = n3299 ^ n3056 ^ n1536 ;
  assign n10106 = n6361 ^ n3683 ^ n3100 ;
  assign n10107 = n10105 | n10106 ;
  assign n10113 = n10112 ^ n10107 ^ 1'b0 ;
  assign n10114 = n3146 ^ n2989 ^ n1151 ;
  assign n10115 = x218 & ~n1254 ;
  assign n10116 = n2883 & n10115 ;
  assign n10117 = n1182 & ~n10116 ;
  assign n10118 = ~n577 & n743 ;
  assign n10119 = n403 & n10118 ;
  assign n10120 = ( n10114 & ~n10117 ) | ( n10114 & n10119 ) | ( ~n10117 & n10119 ) ;
  assign n10121 = n10120 ^ n3621 ^ 1'b0 ;
  assign n10122 = n1362 & ~n2816 ;
  assign n10123 = ( ~n485 & n2662 ) | ( ~n485 & n10122 ) | ( n2662 & n10122 ) ;
  assign n10124 = ( n8294 & n9536 ) | ( n8294 & ~n10123 ) | ( n9536 & ~n10123 ) ;
  assign n10125 = n8504 ^ n6123 ^ 1'b0 ;
  assign n10126 = n3961 | n6573 ;
  assign n10127 = n1943 | n10126 ;
  assign n10128 = ~n5967 & n10127 ;
  assign n10129 = n3947 & n10128 ;
  assign n10130 = ( n7417 & n8278 ) | ( n7417 & ~n10129 ) | ( n8278 & ~n10129 ) ;
  assign n10131 = n1145 ^ n591 ^ 1'b0 ;
  assign n10132 = n8368 ^ n2733 ^ x21 ;
  assign n10133 = ~n10131 & n10132 ;
  assign n10134 = n2893 & n10133 ;
  assign n10135 = n10134 ^ n3248 ^ 1'b0 ;
  assign n10136 = n4515 ^ n580 ^ 1'b0 ;
  assign n10137 = x229 | n10136 ;
  assign n10138 = n6999 | n8155 ;
  assign n10139 = n10138 ^ n9824 ^ 1'b0 ;
  assign n10140 = n8298 ^ n1607 ^ n692 ;
  assign n10141 = n4448 ^ n3349 ^ 1'b0 ;
  assign n10142 = n10140 & n10141 ;
  assign n10143 = ~n4270 & n4378 ;
  assign n10144 = n3389 & n10143 ;
  assign n10145 = n9884 & ~n10144 ;
  assign n10146 = n10142 & ~n10145 ;
  assign n10147 = n10146 ^ n9547 ^ 1'b0 ;
  assign n10148 = n3386 & ~n8225 ;
  assign n10149 = n10148 ^ n2147 ^ 1'b0 ;
  assign n10150 = n9058 & ~n10149 ;
  assign n10151 = ( x209 & n4200 ) | ( x209 & ~n5840 ) | ( n4200 & ~n5840 ) ;
  assign n10152 = n9018 & ~n10151 ;
  assign n10153 = n8781 ^ n4703 ^ n2097 ;
  assign n10154 = n8300 ^ n4468 ^ n2708 ;
  assign n10155 = n2769 & n6177 ;
  assign n10156 = n308 | n2635 ;
  assign n10157 = n10156 ^ n2348 ^ 1'b0 ;
  assign n10161 = n2867 & ~n6032 ;
  assign n10162 = n10161 ^ n3487 ^ 1'b0 ;
  assign n10159 = n6904 ^ n3731 ^ 1'b0 ;
  assign n10160 = n740 | n10159 ;
  assign n10163 = n10162 ^ n10160 ^ 1'b0 ;
  assign n10158 = n293 | n4388 ;
  assign n10164 = n10163 ^ n10158 ^ 1'b0 ;
  assign n10165 = n1066 & ~n3670 ;
  assign n10166 = ~n6941 & n10165 ;
  assign n10167 = n10166 ^ x211 ^ 1'b0 ;
  assign n10168 = n8328 ^ n7836 ^ x155 ;
  assign n10169 = ( ~n1249 & n2448 ) | ( ~n1249 & n3507 ) | ( n2448 & n3507 ) ;
  assign n10170 = n10169 ^ n3773 ^ n3620 ;
  assign n10171 = ~n1037 & n3575 ;
  assign n10172 = n10171 ^ n7672 ^ 1'b0 ;
  assign n10173 = n10070 & n10172 ;
  assign n10174 = n6837 | n10173 ;
  assign n10175 = n6924 ^ n6198 ^ 1'b0 ;
  assign n10176 = n1689 | n10175 ;
  assign n10177 = n10176 ^ n2209 ^ 1'b0 ;
  assign n10178 = ~n1316 & n10177 ;
  assign n10179 = n2516 ^ n344 ^ 1'b0 ;
  assign n10180 = n1763 ^ n356 ^ 1'b0 ;
  assign n10181 = n4086 & n10180 ;
  assign n10182 = ( n4980 & n5569 ) | ( n4980 & n10181 ) | ( n5569 & n10181 ) ;
  assign n10183 = ( n3931 & n10179 ) | ( n3931 & n10182 ) | ( n10179 & n10182 ) ;
  assign n10184 = n2504 ^ n915 ^ 1'b0 ;
  assign n10185 = n2667 & n10184 ;
  assign n10186 = n6174 ^ n2759 ^ 1'b0 ;
  assign n10187 = n4950 & n10186 ;
  assign n10188 = n5004 & n10187 ;
  assign n10189 = n10188 ^ n5276 ^ 1'b0 ;
  assign n10190 = ( n9677 & n10185 ) | ( n9677 & ~n10189 ) | ( n10185 & ~n10189 ) ;
  assign n10191 = n8409 ^ n8012 ^ n2628 ;
  assign n10192 = n4529 & n7483 ;
  assign n10193 = ( n4870 & ~n10191 ) | ( n4870 & n10192 ) | ( ~n10191 & n10192 ) ;
  assign n10194 = n5439 ^ n3314 ^ 1'b0 ;
  assign n10195 = n10194 ^ n7799 ^ n6567 ;
  assign n10196 = ( n5698 & n9467 ) | ( n5698 & ~n10195 ) | ( n9467 & ~n10195 ) ;
  assign n10197 = n2547 ^ n264 ^ 1'b0 ;
  assign n10198 = ~n1908 & n3370 ;
  assign n10199 = ~n10197 & n10198 ;
  assign n10200 = n3067 & n3396 ;
  assign n10202 = ( n2496 & n6982 ) | ( n2496 & ~n7128 ) | ( n6982 & ~n7128 ) ;
  assign n10201 = n2030 ^ n539 ^ x231 ;
  assign n10203 = n10202 ^ n10201 ^ n6188 ;
  assign n10204 = ~n1919 & n8429 ;
  assign n10205 = n10204 ^ n5596 ^ 1'b0 ;
  assign n10206 = n1172 | n3071 ;
  assign n10210 = n3576 & ~n4726 ;
  assign n10211 = n6987 & n10210 ;
  assign n10209 = n7426 ^ n7028 ^ 1'b0 ;
  assign n10212 = n10211 ^ n10209 ^ n3519 ;
  assign n10213 = n4047 | n10212 ;
  assign n10214 = n10213 ^ n5752 ^ 1'b0 ;
  assign n10207 = n2945 & n6361 ;
  assign n10208 = ~n1664 & n10207 ;
  assign n10215 = n10214 ^ n10208 ^ 1'b0 ;
  assign n10216 = n10206 | n10215 ;
  assign n10217 = n10205 | n10216 ;
  assign n10218 = n10203 & ~n10217 ;
  assign n10219 = n5670 ^ n4971 ^ 1'b0 ;
  assign n10220 = n2207 & n10219 ;
  assign n10221 = n10220 ^ n4652 ^ 1'b0 ;
  assign n10222 = n10151 ^ n347 ^ 1'b0 ;
  assign n10223 = n522 & n10222 ;
  assign n10224 = n10223 ^ x149 ^ 1'b0 ;
  assign n10225 = ~n2580 & n3669 ;
  assign n10226 = n2472 & n10225 ;
  assign n10227 = n4450 | n10226 ;
  assign n10228 = n3194 | n10227 ;
  assign n10229 = n10228 ^ n8448 ^ n2812 ;
  assign n10230 = n4763 ^ n1657 ^ 1'b0 ;
  assign n10231 = n10230 ^ n9417 ^ 1'b0 ;
  assign n10232 = ( n4749 & ~n10229 ) | ( n4749 & n10231 ) | ( ~n10229 & n10231 ) ;
  assign n10233 = n7599 & ~n8077 ;
  assign n10234 = n10233 ^ n1004 ^ 1'b0 ;
  assign n10235 = n3381 ^ n1852 ^ 1'b0 ;
  assign n10236 = n4827 | n10235 ;
  assign n10237 = n1425 | n7850 ;
  assign n10238 = ~n1250 & n10237 ;
  assign n10239 = n10236 & n10238 ;
  assign n10240 = n6473 ^ n2106 ^ 1'b0 ;
  assign n10241 = n7886 & ~n10240 ;
  assign n10242 = ~n1659 & n10241 ;
  assign n10243 = ~n1817 & n6776 ;
  assign n10244 = n10243 ^ n3414 ^ n2598 ;
  assign n10245 = ( ~n447 & n3819 ) | ( ~n447 & n10244 ) | ( n3819 & n10244 ) ;
  assign n10246 = n7942 | n10180 ;
  assign n10247 = n3821 & ~n10246 ;
  assign n10248 = ( n920 & n3755 ) | ( n920 & ~n9030 ) | ( n3755 & ~n9030 ) ;
  assign n10249 = n5006 ^ n2397 ^ 1'b0 ;
  assign n10250 = n9467 & n10249 ;
  assign n10251 = n4228 & ~n6264 ;
  assign n10252 = ( n829 & ~n4521 ) | ( n829 & n6831 ) | ( ~n4521 & n6831 ) ;
  assign n10253 = ~n7833 & n10252 ;
  assign n10254 = n10251 & n10253 ;
  assign n10255 = n10254 ^ n6875 ^ 1'b0 ;
  assign n10256 = n3282 | n3442 ;
  assign n10257 = n10256 ^ n1908 ^ 1'b0 ;
  assign n10258 = n6915 ^ n5319 ^ 1'b0 ;
  assign n10259 = ~n6246 & n7624 ;
  assign n10260 = n10259 ^ n9945 ^ 1'b0 ;
  assign n10261 = ( n2794 & ~n9754 ) | ( n2794 & n9838 ) | ( ~n9754 & n9838 ) ;
  assign n10264 = n6328 ^ n2618 ^ 1'b0 ;
  assign n10262 = n2055 & n4269 ;
  assign n10263 = n10262 ^ n5405 ^ n3947 ;
  assign n10265 = n10264 ^ n10263 ^ 1'b0 ;
  assign n10266 = n10265 ^ n3252 ^ 1'b0 ;
  assign n10267 = n4227 ^ n1534 ^ 1'b0 ;
  assign n10268 = n10267 ^ n10171 ^ 1'b0 ;
  assign n10269 = n1543 & ~n10268 ;
  assign n10270 = n10269 ^ n3640 ^ 1'b0 ;
  assign n10271 = n1247 & ~n10270 ;
  assign n10272 = n1972 ^ n1562 ^ 1'b0 ;
  assign n10273 = n10271 & n10272 ;
  assign n10274 = n10273 ^ x24 ^ 1'b0 ;
  assign n10275 = n10274 ^ n5230 ^ n2317 ;
  assign n10276 = x51 & n873 ;
  assign n10277 = ~n677 & n10276 ;
  assign n10278 = n10080 ^ n1090 ^ 1'b0 ;
  assign n10279 = n10277 | n10278 ;
  assign n10280 = n10279 ^ n1635 ^ 1'b0 ;
  assign n10281 = ~n5363 & n10280 ;
  assign n10282 = n8821 ^ n1363 ^ 1'b0 ;
  assign n10283 = n1757 | n10282 ;
  assign n10284 = n10283 ^ n9552 ^ 1'b0 ;
  assign n10285 = n5203 & n10284 ;
  assign n10286 = n10281 & ~n10285 ;
  assign n10287 = n780 ^ n464 ^ 1'b0 ;
  assign n10288 = n1873 & ~n7658 ;
  assign n10289 = ( ~n487 & n10287 ) | ( ~n487 & n10288 ) | ( n10287 & n10288 ) ;
  assign n10290 = n4321 ^ n1958 ^ 1'b0 ;
  assign n10291 = n10290 ^ n2050 ^ 1'b0 ;
  assign n10292 = n8949 & n10291 ;
  assign n10293 = n10289 & n10292 ;
  assign n10294 = n10293 ^ n6428 ^ 1'b0 ;
  assign n10295 = x141 & n347 ;
  assign n10296 = n10028 & n10295 ;
  assign n10297 = n542 | n10296 ;
  assign n10298 = n10297 ^ n3789 ^ 1'b0 ;
  assign n10299 = n10298 ^ n4741 ^ 1'b0 ;
  assign n10300 = n4088 & n8317 ;
  assign n10301 = n10300 ^ n8288 ^ 1'b0 ;
  assign n10302 = n3086 & n3219 ;
  assign n10303 = n1204 & n10302 ;
  assign n10304 = n1510 & ~n10303 ;
  assign n10305 = x246 & n1781 ;
  assign n10306 = n10305 ^ n980 ^ 1'b0 ;
  assign n10307 = n10306 ^ n8278 ^ 1'b0 ;
  assign n10308 = ~n1582 & n10307 ;
  assign n10309 = n10308 ^ n5565 ^ 1'b0 ;
  assign n10310 = n5813 ^ n2771 ^ 1'b0 ;
  assign n10311 = n6056 ^ n3868 ^ 1'b0 ;
  assign n10312 = n6850 & n10311 ;
  assign n10313 = n9333 & n10312 ;
  assign n10314 = ( n639 & n659 ) | ( n639 & ~n8508 ) | ( n659 & ~n8508 ) ;
  assign n10315 = n2287 | n10314 ;
  assign n10316 = n2024 | n5926 ;
  assign n10317 = n10316 ^ n2387 ^ 1'b0 ;
  assign n10318 = n10317 ^ n3373 ^ 1'b0 ;
  assign n10319 = x149 & ~n8515 ;
  assign n10320 = n3012 & n10319 ;
  assign n10321 = n4517 ^ n4397 ^ 1'b0 ;
  assign n10322 = ( ~n2462 & n4013 ) | ( ~n2462 & n10321 ) | ( n4013 & n10321 ) ;
  assign n10323 = n6587 ^ n3237 ^ n1444 ;
  assign n10324 = n1178 ^ n891 ^ 1'b0 ;
  assign n10325 = n10324 ^ n6907 ^ 1'b0 ;
  assign n10326 = ( n6914 & ~n7883 ) | ( n6914 & n9321 ) | ( ~n7883 & n9321 ) ;
  assign n10327 = ( n2429 & ~n4219 ) | ( n2429 & n10326 ) | ( ~n4219 & n10326 ) ;
  assign n10328 = n10325 & n10327 ;
  assign n10329 = n10328 ^ n2642 ^ 1'b0 ;
  assign n10330 = n10323 & n10329 ;
  assign n10331 = ~n2804 & n6433 ;
  assign n10332 = n10331 ^ n4003 ^ n3368 ;
  assign n10333 = n7761 ^ n7665 ^ x17 ;
  assign n10334 = n9044 ^ n7741 ^ n3604 ;
  assign n10335 = n10334 ^ n10182 ^ 1'b0 ;
  assign n10336 = ~n10333 & n10335 ;
  assign n10337 = n10336 ^ n4572 ^ 1'b0 ;
  assign n10338 = n7537 ^ n861 ^ 1'b0 ;
  assign n10339 = n1689 | n10338 ;
  assign n10340 = ( n2592 & n6944 ) | ( n2592 & ~n10339 ) | ( n6944 & ~n10339 ) ;
  assign n10341 = n1024 | n2603 ;
  assign n10342 = ( n7358 & n10340 ) | ( n7358 & ~n10341 ) | ( n10340 & ~n10341 ) ;
  assign n10343 = n2118 ^ n1718 ^ 1'b0 ;
  assign n10344 = n1388 & ~n10343 ;
  assign n10345 = ~n5761 & n10344 ;
  assign n10346 = n2351 ^ n1206 ^ 1'b0 ;
  assign n10347 = n5671 ^ x24 ^ 1'b0 ;
  assign n10348 = n10346 | n10347 ;
  assign n10349 = n5091 ^ n2378 ^ n565 ;
  assign n10350 = ( n741 & n2912 ) | ( n741 & ~n10349 ) | ( n2912 & ~n10349 ) ;
  assign n10351 = ( n7740 & ~n10348 ) | ( n7740 & n10350 ) | ( ~n10348 & n10350 ) ;
  assign n10352 = ~n4925 & n10351 ;
  assign n10353 = n10352 ^ n4389 ^ 1'b0 ;
  assign n10354 = ~n632 & n3596 ;
  assign n10355 = n10354 ^ n2178 ^ 1'b0 ;
  assign n10356 = n4447 ^ n1343 ^ n528 ;
  assign n10357 = n10356 ^ n4367 ^ n1170 ;
  assign n10358 = n704 & n4080 ;
  assign n10359 = n5281 ^ n1359 ^ 1'b0 ;
  assign n10360 = n10358 & ~n10359 ;
  assign n10361 = n3059 ^ n2500 ^ 1'b0 ;
  assign n10362 = n2977 | n10361 ;
  assign n10363 = n6127 | n10362 ;
  assign n10364 = n2435 ^ n1258 ^ n310 ;
  assign n10365 = n10364 ^ n10025 ^ n7753 ;
  assign n10366 = ~n9463 & n10365 ;
  assign n10368 = n7996 ^ n4600 ^ 1'b0 ;
  assign n10369 = n10368 ^ n8618 ^ 1'b0 ;
  assign n10367 = n2838 ^ n2289 ^ x169 ;
  assign n10370 = n10369 ^ n10367 ^ 1'b0 ;
  assign n10371 = n10370 ^ n3416 ^ n990 ;
  assign n10373 = n6622 ^ x138 ^ 1'b0 ;
  assign n10374 = x210 & ~n10373 ;
  assign n10375 = n3821 & n10374 ;
  assign n10376 = n10375 ^ n3687 ^ n1895 ;
  assign n10372 = n560 & n8439 ;
  assign n10377 = n10376 ^ n10372 ^ 1'b0 ;
  assign n10378 = n5747 ^ n950 ^ n797 ;
  assign n10379 = n4929 ^ n4889 ^ 1'b0 ;
  assign n10380 = ( n5854 & n6646 ) | ( n5854 & n10379 ) | ( n6646 & n10379 ) ;
  assign n10381 = n10021 & ~n10380 ;
  assign n10382 = n3374 & n5246 ;
  assign n10383 = ~n8209 & n10382 ;
  assign n10384 = n2720 & ~n10383 ;
  assign n10385 = n10384 ^ n4625 ^ 1'b0 ;
  assign n10390 = n3779 & n6896 ;
  assign n10386 = n1366 & ~n3215 ;
  assign n10387 = n3961 & n10386 ;
  assign n10388 = n10387 ^ n3632 ^ n531 ;
  assign n10389 = n6000 & n10388 ;
  assign n10391 = n10390 ^ n10389 ^ 1'b0 ;
  assign n10392 = n2331 | n4392 ;
  assign n10393 = n1858 ^ n1711 ^ 1'b0 ;
  assign n10394 = n775 | n10393 ;
  assign n10395 = n10394 ^ n2759 ^ 1'b0 ;
  assign n10396 = n10010 & ~n10395 ;
  assign n10397 = n7892 & ~n8775 ;
  assign n10398 = ~n10396 & n10397 ;
  assign n10399 = n10392 & ~n10398 ;
  assign n10400 = n10399 ^ n4823 ^ 1'b0 ;
  assign n10401 = n971 & ~n9559 ;
  assign n10402 = n8324 & n10401 ;
  assign n10403 = n4858 ^ n3320 ^ 1'b0 ;
  assign n10404 = n10402 & n10403 ;
  assign n10405 = ~n8800 & n10404 ;
  assign n10406 = n10405 ^ n5056 ^ 1'b0 ;
  assign n10407 = ~n10400 & n10406 ;
  assign n10408 = n7245 | n10407 ;
  assign n10409 = n4983 ^ x38 ^ 1'b0 ;
  assign n10410 = n6596 ^ n3898 ^ 1'b0 ;
  assign n10411 = n10409 | n10410 ;
  assign n10413 = n632 | n2583 ;
  assign n10412 = n6056 ^ n1948 ^ 1'b0 ;
  assign n10414 = n10413 ^ n10412 ^ n8150 ;
  assign n10415 = n702 & ~n2754 ;
  assign n10416 = ~n2594 & n10415 ;
  assign n10417 = n2421 | n10416 ;
  assign n10418 = n3960 ^ n3070 ^ 1'b0 ;
  assign n10419 = n1494 | n10418 ;
  assign n10420 = n5731 & ~n10419 ;
  assign n10421 = n10420 ^ n1550 ^ 1'b0 ;
  assign n10422 = n926 & n981 ;
  assign n10423 = n399 & n2946 ;
  assign n10424 = ~n10422 & n10423 ;
  assign n10425 = ( n10020 & ~n10421 ) | ( n10020 & n10424 ) | ( ~n10421 & n10424 ) ;
  assign n10426 = n5759 & n8364 ;
  assign n10429 = x219 & ~n2994 ;
  assign n10428 = n6368 ^ n2117 ^ 1'b0 ;
  assign n10430 = n10429 ^ n10428 ^ 1'b0 ;
  assign n10427 = n3357 | n9064 ;
  assign n10431 = n10430 ^ n10427 ^ 1'b0 ;
  assign n10434 = n6328 ^ n356 ^ 1'b0 ;
  assign n10432 = n2727 ^ n1079 ^ x209 ;
  assign n10433 = n5497 & ~n10432 ;
  assign n10435 = n10434 ^ n10433 ^ 1'b0 ;
  assign n10436 = n6647 | n10435 ;
  assign n10437 = ( n1702 & n10431 ) | ( n1702 & ~n10436 ) | ( n10431 & ~n10436 ) ;
  assign n10440 = n5612 ^ n1427 ^ x130 ;
  assign n10438 = n381 | n6174 ;
  assign n10439 = n3519 | n10438 ;
  assign n10441 = n10440 ^ n10439 ^ 1'b0 ;
  assign n10442 = ~n4612 & n10441 ;
  assign n10456 = n9683 ^ n3797 ^ 1'b0 ;
  assign n10443 = n5193 ^ x169 ^ x165 ;
  assign n10444 = n5134 ^ x31 ^ 1'b0 ;
  assign n10445 = n5335 | n10444 ;
  assign n10446 = ( n1517 & ~n10443 ) | ( n1517 & n10445 ) | ( ~n10443 & n10445 ) ;
  assign n10447 = ~n7858 & n10446 ;
  assign n10448 = n1858 ^ n905 ^ x222 ;
  assign n10449 = n4911 & ~n10448 ;
  assign n10450 = n2032 & n10449 ;
  assign n10451 = ( n6930 & n10447 ) | ( n6930 & n10450 ) | ( n10447 & n10450 ) ;
  assign n10452 = n2106 & n3260 ;
  assign n10453 = n10452 ^ n6450 ^ 1'b0 ;
  assign n10454 = n10453 ^ n8729 ^ n3823 ;
  assign n10455 = n10451 | n10454 ;
  assign n10457 = n10456 ^ n10455 ^ 1'b0 ;
  assign n10460 = n2826 ^ n2640 ^ 1'b0 ;
  assign n10461 = n5696 | n10460 ;
  assign n10458 = ~n633 & n9853 ;
  assign n10459 = n2045 & n10458 ;
  assign n10462 = n10461 ^ n10459 ^ 1'b0 ;
  assign n10463 = ( n4588 & n5629 ) | ( n4588 & ~n10462 ) | ( n5629 & ~n10462 ) ;
  assign n10470 = ( ~x83 & n1702 ) | ( ~x83 & n7796 ) | ( n1702 & n7796 ) ;
  assign n10468 = n996 ^ x120 ^ 1'b0 ;
  assign n10467 = n2080 | n3782 ;
  assign n10469 = n10468 ^ n10467 ^ 1'b0 ;
  assign n10465 = n7069 ^ n3464 ^ x149 ;
  assign n10464 = ~n2426 & n7457 ;
  assign n10466 = n10465 ^ n10464 ^ n1368 ;
  assign n10471 = n10470 ^ n10469 ^ n10466 ;
  assign n10472 = n10471 ^ n7325 ^ n3488 ;
  assign n10473 = n5929 & ~n6908 ;
  assign n10474 = n6491 ^ n3585 ^ 1'b0 ;
  assign n10475 = ~n4598 & n10474 ;
  assign n10476 = n10475 ^ n8719 ^ 1'b0 ;
  assign n10477 = x184 & n344 ;
  assign n10478 = n3866 & ~n9588 ;
  assign n10479 = n7037 & n9477 ;
  assign n10480 = n10479 ^ n9630 ^ 1'b0 ;
  assign n10482 = n4243 ^ n1446 ^ 1'b0 ;
  assign n10483 = n5969 & ~n10482 ;
  assign n10481 = ~n4316 & n9457 ;
  assign n10484 = n10483 ^ n10481 ^ n8144 ;
  assign n10485 = ( n870 & n4465 ) | ( n870 & n5686 ) | ( n4465 & n5686 ) ;
  assign n10486 = ( ~n782 & n9597 ) | ( ~n782 & n10485 ) | ( n9597 & n10485 ) ;
  assign n10487 = n10486 ^ n5436 ^ n3545 ;
  assign n10488 = n3730 & n10487 ;
  assign n10489 = ~x17 & n6287 ;
  assign n10490 = n10489 ^ n7073 ^ 1'b0 ;
  assign n10491 = n10488 & n10490 ;
  assign n10492 = n10491 ^ n7355 ^ 1'b0 ;
  assign n10495 = x27 & n3406 ;
  assign n10496 = n10495 ^ n9350 ^ 1'b0 ;
  assign n10493 = ( ~n857 & n5215 ) | ( ~n857 & n5257 ) | ( n5215 & n5257 ) ;
  assign n10494 = n1675 & n10493 ;
  assign n10497 = n10496 ^ n10494 ^ 1'b0 ;
  assign n10498 = n3260 & n6218 ;
  assign n10501 = n7721 ^ n6919 ^ n2777 ;
  assign n10502 = n10501 ^ n1655 ^ 1'b0 ;
  assign n10503 = ~n3321 & n10502 ;
  assign n10499 = n2680 & ~n5524 ;
  assign n10500 = ~n4129 & n10499 ;
  assign n10504 = n10503 ^ n10500 ^ n1415 ;
  assign n10505 = ~n1702 & n4978 ;
  assign n10506 = n5269 & ~n6894 ;
  assign n10507 = n5359 & ~n7825 ;
  assign n10508 = n3620 ^ x75 ^ 1'b0 ;
  assign n10509 = n1746 | n10508 ;
  assign n10510 = n10509 ^ n7927 ^ 1'b0 ;
  assign n10511 = ( n3744 & n6717 ) | ( n3744 & ~n6719 ) | ( n6717 & ~n6719 ) ;
  assign n10512 = n10511 ^ n7858 ^ 1'b0 ;
  assign n10514 = n6243 ^ n411 ^ 1'b0 ;
  assign n10513 = n379 | n8878 ;
  assign n10515 = n10514 ^ n10513 ^ 1'b0 ;
  assign n10516 = n6717 ^ n3091 ^ 1'b0 ;
  assign n10517 = n5126 ^ n1145 ^ 1'b0 ;
  assign n10518 = n7661 | n10517 ;
  assign n10519 = n639 | n8473 ;
  assign n10522 = n4867 & n9559 ;
  assign n10523 = n10522 ^ n9587 ^ 1'b0 ;
  assign n10520 = n8381 ^ x45 ^ 1'b0 ;
  assign n10521 = n10520 ^ n5744 ^ 1'b0 ;
  assign n10524 = n10523 ^ n10521 ^ n2193 ;
  assign n10525 = ( n1948 & n9740 ) | ( n1948 & ~n10524 ) | ( n9740 & ~n10524 ) ;
  assign n10526 = n4447 | n8945 ;
  assign n10527 = n599 & ~n9814 ;
  assign n10528 = n10526 & n10527 ;
  assign n10529 = ~n3521 & n8183 ;
  assign n10530 = n4243 & ~n10529 ;
  assign n10531 = n5170 & n10530 ;
  assign n10532 = n9874 & ~n10531 ;
  assign n10533 = n2901 ^ n606 ^ 1'b0 ;
  assign n10534 = n2306 & ~n9299 ;
  assign n10535 = n10533 & n10534 ;
  assign n10543 = n10050 ^ n747 ^ 1'b0 ;
  assign n10536 = ~n7109 & n9729 ;
  assign n10537 = n3324 ^ n1512 ^ 1'b0 ;
  assign n10538 = n10537 ^ n2942 ^ 1'b0 ;
  assign n10539 = n9276 | n10538 ;
  assign n10540 = x85 & ~n10539 ;
  assign n10541 = n10540 ^ n7694 ^ 1'b0 ;
  assign n10542 = ( n6793 & n10536 ) | ( n6793 & ~n10541 ) | ( n10536 & ~n10541 ) ;
  assign n10544 = n10543 ^ n10542 ^ 1'b0 ;
  assign n10545 = n7812 ^ n5844 ^ 1'b0 ;
  assign n10551 = n6927 ^ n3654 ^ 1'b0 ;
  assign n10546 = n6571 ^ n5637 ^ 1'b0 ;
  assign n10547 = n1846 ^ n588 ^ 1'b0 ;
  assign n10548 = n10546 & n10547 ;
  assign n10549 = n10548 ^ n4626 ^ 1'b0 ;
  assign n10550 = n10549 ^ n2506 ^ 1'b0 ;
  assign n10552 = n10551 ^ n10550 ^ n10432 ;
  assign n10553 = n10552 ^ n7079 ^ 1'b0 ;
  assign n10554 = n654 & ~n6425 ;
  assign n10555 = n4254 & n10554 ;
  assign n10556 = n10555 ^ n4585 ^ 1'b0 ;
  assign n10557 = n5077 & n10556 ;
  assign n10558 = n4068 | n10557 ;
  assign n10559 = n656 & ~n885 ;
  assign n10560 = n10559 ^ n6573 ^ n4522 ;
  assign n10561 = n6314 & ~n10560 ;
  assign n10562 = n9685 ^ n7961 ^ 1'b0 ;
  assign n10563 = n979 ^ n415 ^ 1'b0 ;
  assign n10564 = n10563 ^ n402 ^ x196 ;
  assign n10565 = n8017 & ~n8382 ;
  assign n10566 = n7371 ^ n6064 ^ n2411 ;
  assign n10567 = n10566 ^ n4994 ^ 1'b0 ;
  assign n10568 = n2894 & ~n10567 ;
  assign n10569 = n7243 ^ n4198 ^ 1'b0 ;
  assign n10570 = n6985 & n10569 ;
  assign n10571 = ( n2429 & ~n8284 ) | ( n2429 & n8956 ) | ( ~n8284 & n8956 ) ;
  assign n10572 = n3040 | n3969 ;
  assign n10573 = n861 | n10572 ;
  assign n10574 = n9106 ^ n2026 ^ 1'b0 ;
  assign n10575 = n10573 & ~n10574 ;
  assign n10578 = n616 & n4223 ;
  assign n10579 = n10578 ^ n354 ^ 1'b0 ;
  assign n10580 = ~n4553 & n10579 ;
  assign n10581 = n10580 ^ n6603 ^ 1'b0 ;
  assign n10576 = ~n8449 & n10396 ;
  assign n10577 = n10576 ^ n472 ^ 1'b0 ;
  assign n10582 = n10581 ^ n10577 ^ n305 ;
  assign n10583 = n10582 ^ n3539 ^ n1701 ;
  assign n10584 = n5726 ^ n4913 ^ n4581 ;
  assign n10585 = n298 | n4583 ;
  assign n10586 = ~n9884 & n10585 ;
  assign n10587 = ~n9255 & n10586 ;
  assign n10593 = n3924 & ~n4199 ;
  assign n10588 = x250 & ~n890 ;
  assign n10589 = ~n6347 & n10588 ;
  assign n10590 = n10589 ^ n4230 ^ 1'b0 ;
  assign n10591 = n2314 & ~n10590 ;
  assign n10592 = n10591 ^ n7226 ^ 1'b0 ;
  assign n10594 = n10593 ^ n10592 ^ 1'b0 ;
  assign n10595 = n10587 | n10594 ;
  assign n10596 = ~n1874 & n4913 ;
  assign n10597 = ~n3194 & n10596 ;
  assign n10598 = n1322 | n10597 ;
  assign n10599 = n4144 & n10598 ;
  assign n10600 = x146 & ~n10599 ;
  assign n10601 = n8928 ^ n2293 ^ 1'b0 ;
  assign n10602 = n7417 ^ n2373 ^ n845 ;
  assign n10603 = n10602 ^ n6638 ^ n2951 ;
  assign n10604 = n7171 | n10603 ;
  assign n10605 = x47 & n1537 ;
  assign n10606 = ~n778 & n10605 ;
  assign n10607 = n7440 ^ x200 ^ 1'b0 ;
  assign n10608 = n5803 & n10607 ;
  assign n10609 = n10606 & n10608 ;
  assign n10610 = n8818 ^ n3239 ^ 1'b0 ;
  assign n10611 = n10609 | n10610 ;
  assign n10612 = n5556 ^ n1804 ^ 1'b0 ;
  assign n10613 = n3920 | n10612 ;
  assign n10614 = n892 | n6777 ;
  assign n10615 = ( ~n8372 & n10613 ) | ( ~n8372 & n10614 ) | ( n10613 & n10614 ) ;
  assign n10616 = n843 & n10615 ;
  assign n10617 = n2447 ^ n368 ^ x199 ;
  assign n10618 = n10617 ^ n4958 ^ n4591 ;
  assign n10619 = n10618 ^ n9157 ^ n3096 ;
  assign n10621 = n1362 & n10324 ;
  assign n10620 = ( n337 & n987 ) | ( n337 & ~n3182 ) | ( n987 & ~n3182 ) ;
  assign n10622 = n10621 ^ n10620 ^ 1'b0 ;
  assign n10623 = n4227 ^ n3086 ^ 1'b0 ;
  assign n10624 = n10623 ^ n10492 ^ 1'b0 ;
  assign n10628 = n6069 | n6229 ;
  assign n10629 = ~n3087 & n10628 ;
  assign n10625 = n1438 ^ n1298 ^ 1'b0 ;
  assign n10626 = n3374 & n10625 ;
  assign n10627 = n10626 ^ n1709 ^ n1593 ;
  assign n10630 = n10629 ^ n10627 ^ 1'b0 ;
  assign n10631 = ~n7848 & n10630 ;
  assign n10632 = n2633 ^ x16 ^ 1'b0 ;
  assign n10633 = ~n4947 & n10632 ;
  assign n10634 = n1479 & ~n10633 ;
  assign n10635 = x205 & ~n10634 ;
  assign n10636 = ~n10631 & n10635 ;
  assign n10637 = n9377 ^ n8043 ^ 1'b0 ;
  assign n10639 = n9255 ^ n1965 ^ 1'b0 ;
  assign n10640 = ( n559 & n1322 ) | ( n559 & n10639 ) | ( n1322 & n10639 ) ;
  assign n10641 = n10640 ^ n511 ^ 1'b0 ;
  assign n10642 = n10641 ^ n5094 ^ 1'b0 ;
  assign n10643 = n10642 ^ n6016 ^ 1'b0 ;
  assign n10638 = n4115 & n4891 ;
  assign n10644 = n10643 ^ n10638 ^ n9812 ;
  assign n10645 = n6400 ^ n495 ^ 1'b0 ;
  assign n10646 = ( n1270 & n2634 ) | ( n1270 & n3636 ) | ( n2634 & n3636 ) ;
  assign n10647 = ~n9685 & n10646 ;
  assign n10648 = n10647 ^ n5621 ^ 1'b0 ;
  assign n10649 = n2885 | n5947 ;
  assign n10650 = n10648 | n10649 ;
  assign n10651 = n1374 | n2968 ;
  assign n10652 = n10651 ^ n3494 ^ 1'b0 ;
  assign n10653 = n1424 & n7481 ;
  assign n10654 = n10653 ^ n7665 ^ 1'b0 ;
  assign n10655 = ( n6384 & ~n10652 ) | ( n6384 & n10654 ) | ( ~n10652 & n10654 ) ;
  assign n10656 = ( x167 & n257 ) | ( x167 & n718 ) | ( n257 & n718 ) ;
  assign n10657 = n10656 ^ n1694 ^ n716 ;
  assign n10658 = n10657 ^ n1105 ^ x18 ;
  assign n10659 = ( n405 & ~n4685 ) | ( n405 & n9025 ) | ( ~n4685 & n9025 ) ;
  assign n10660 = n10171 ^ n1042 ^ n270 ;
  assign n10661 = n6446 & ~n10660 ;
  assign n10663 = n7769 ^ n2386 ^ 1'b0 ;
  assign n10662 = n7486 ^ n3667 ^ 1'b0 ;
  assign n10664 = n10663 ^ n10662 ^ n298 ;
  assign n10665 = n8182 ^ n843 ^ 1'b0 ;
  assign n10666 = n6135 | n9861 ;
  assign n10667 = x78 | n10666 ;
  assign n10668 = ~n5301 & n10667 ;
  assign n10669 = n10665 & n10668 ;
  assign n10670 = ( n7686 & n10664 ) | ( n7686 & ~n10669 ) | ( n10664 & ~n10669 ) ;
  assign n10671 = n8361 ^ n6933 ^ n5518 ;
  assign n10672 = n2068 ^ n2013 ^ 1'b0 ;
  assign n10673 = n10626 ^ n430 ^ 1'b0 ;
  assign n10674 = n4107 & n10673 ;
  assign n10675 = ( n8548 & ~n10370 ) | ( n8548 & n10674 ) | ( ~n10370 & n10674 ) ;
  assign n10679 = n807 & n3892 ;
  assign n10680 = n10679 ^ n4397 ^ 1'b0 ;
  assign n10678 = x224 & n1260 ;
  assign n10681 = n10680 ^ n10678 ^ 1'b0 ;
  assign n10676 = n8360 & ~n9168 ;
  assign n10677 = n6211 & n10676 ;
  assign n10682 = n10681 ^ n10677 ^ n8630 ;
  assign n10683 = n3349 ^ n1254 ^ 1'b0 ;
  assign n10684 = n7486 & ~n8129 ;
  assign n10685 = n10684 ^ n638 ^ 1'b0 ;
  assign n10686 = n1611 & n2885 ;
  assign n10687 = n5818 ^ n4730 ^ n991 ;
  assign n10688 = ( n2605 & n5408 ) | ( n2605 & ~n10687 ) | ( n5408 & ~n10687 ) ;
  assign n10689 = n5580 ^ n559 ^ 1'b0 ;
  assign n10690 = n10688 & n10689 ;
  assign n10691 = ( n597 & ~n3390 ) | ( n597 & n10690 ) | ( ~n3390 & n10690 ) ;
  assign n10692 = n10691 ^ n2677 ^ 1'b0 ;
  assign n10693 = x2 | n9966 ;
  assign n10694 = n10693 ^ n7440 ^ 1'b0 ;
  assign n10695 = n5926 | n8821 ;
  assign n10696 = n5575 ^ n3749 ^ 1'b0 ;
  assign n10697 = n1004 ^ x60 ^ 1'b0 ;
  assign n10698 = n1140 | n10697 ;
  assign n10699 = n10696 & ~n10698 ;
  assign n10700 = n10699 ^ n2223 ^ 1'b0 ;
  assign n10701 = ~n6931 & n10700 ;
  assign n10702 = n10701 ^ n2647 ^ 1'b0 ;
  assign n10703 = n10695 | n10702 ;
  assign n10704 = n2763 & n3788 ;
  assign n10705 = n1339 & n3328 ;
  assign n10706 = n10705 ^ n6177 ^ 1'b0 ;
  assign n10707 = n2106 ^ n848 ^ 1'b0 ;
  assign n10708 = n10212 ^ n4219 ^ n1413 ;
  assign n10709 = n2636 ^ n2169 ^ 1'b0 ;
  assign n10710 = ( n5804 & n10708 ) | ( n5804 & n10709 ) | ( n10708 & n10709 ) ;
  assign n10711 = n3719 ^ n1807 ^ 1'b0 ;
  assign n10712 = ( ~n1667 & n6202 ) | ( ~n1667 & n10711 ) | ( n6202 & n10711 ) ;
  assign n10713 = n2085 & n7528 ;
  assign n10714 = n10713 ^ n3775 ^ n1705 ;
  assign n10715 = x172 & n1761 ;
  assign n10716 = ~n6870 & n10715 ;
  assign n10717 = n3949 | n8575 ;
  assign n10718 = n10717 ^ n9090 ^ 1'b0 ;
  assign n10721 = ( n3068 & n7226 ) | ( n3068 & ~n7333 ) | ( n7226 & ~n7333 ) ;
  assign n10719 = n356 & ~n10522 ;
  assign n10720 = ~n1913 & n10719 ;
  assign n10722 = n10721 ^ n10720 ^ n4357 ;
  assign n10723 = ( ~x1 & n841 ) | ( ~x1 & n2314 ) | ( n841 & n2314 ) ;
  assign n10724 = n3022 & ~n3654 ;
  assign n10725 = n3567 | n10724 ;
  assign n10726 = n10725 ^ n6958 ^ 1'b0 ;
  assign n10727 = n2099 & ~n5607 ;
  assign n10728 = n3995 ^ n1618 ^ 1'b0 ;
  assign n10729 = n10728 ^ n10606 ^ n6717 ;
  assign n10730 = n1304 | n3947 ;
  assign n10731 = n10730 ^ n2009 ^ 1'b0 ;
  assign n10732 = n769 & n5500 ;
  assign n10733 = n10732 ^ n3245 ^ 1'b0 ;
  assign n10734 = ~n1541 & n10733 ;
  assign n10735 = n10734 ^ n3514 ^ 1'b0 ;
  assign n10736 = n7932 ^ n5030 ^ n652 ;
  assign n10737 = ~n7860 & n9011 ;
  assign n10738 = ~n2182 & n9605 ;
  assign n10739 = ( ~n1460 & n8548 ) | ( ~n1460 & n10021 ) | ( n8548 & n10021 ) ;
  assign n10740 = n1665 & n10739 ;
  assign n10741 = n7992 ^ n7840 ^ 1'b0 ;
  assign n10742 = n7060 ^ n3851 ^ n1463 ;
  assign n10743 = ~n1728 & n5065 ;
  assign n10744 = n4879 ^ n2798 ^ n559 ;
  assign n10745 = ( n3791 & n6201 ) | ( n3791 & n10744 ) | ( n6201 & n10744 ) ;
  assign n10746 = n10745 ^ n7280 ^ 1'b0 ;
  assign n10747 = n5432 & n10746 ;
  assign n10750 = n5022 & ~n6724 ;
  assign n10751 = n10750 ^ n4637 ^ n1797 ;
  assign n10748 = n3775 ^ x146 ^ 1'b0 ;
  assign n10749 = n9288 & ~n10748 ;
  assign n10752 = n10751 ^ n10749 ^ 1'b0 ;
  assign n10753 = n4428 & n4628 ;
  assign n10754 = n4931 & n7001 ;
  assign n10755 = n10753 | n10754 ;
  assign n10756 = n8388 ^ n785 ^ 1'b0 ;
  assign n10757 = n10755 | n10756 ;
  assign n10758 = ( n9683 & ~n10464 ) | ( n9683 & n10757 ) | ( ~n10464 & n10757 ) ;
  assign n10759 = n10758 ^ n8739 ^ 1'b0 ;
  assign n10764 = n1832 ^ n894 ^ 1'b0 ;
  assign n10762 = ~n2341 & n6403 ;
  assign n10760 = n3434 & ~n4818 ;
  assign n10761 = n589 & ~n10760 ;
  assign n10763 = n10762 ^ n10761 ^ 1'b0 ;
  assign n10765 = n10764 ^ n10763 ^ n8006 ;
  assign n10766 = n6711 ^ n6574 ^ 1'b0 ;
  assign n10767 = ~n3160 & n10766 ;
  assign n10768 = ~n5582 & n10767 ;
  assign n10772 = n4884 ^ n4583 ^ 1'b0 ;
  assign n10773 = n3196 & n10772 ;
  assign n10769 = n4224 ^ n1908 ^ 1'b0 ;
  assign n10770 = n2654 & n10769 ;
  assign n10771 = ( n4937 & n5912 ) | ( n4937 & n10770 ) | ( n5912 & n10770 ) ;
  assign n10774 = n10773 ^ n10771 ^ 1'b0 ;
  assign n10775 = n3121 & n5248 ;
  assign n10776 = n10775 ^ n1296 ^ 1'b0 ;
  assign n10780 = ~n4563 & n7616 ;
  assign n10777 = n4899 ^ n2807 ^ 1'b0 ;
  assign n10778 = n10777 ^ n5436 ^ n2513 ;
  assign n10779 = n8898 | n10778 ;
  assign n10781 = n10780 ^ n10779 ^ 1'b0 ;
  assign n10782 = n5535 ^ n3356 ^ 1'b0 ;
  assign n10783 = n6241 ^ n1835 ^ 1'b0 ;
  assign n10784 = n10782 & n10783 ;
  assign n10785 = n10784 ^ n5376 ^ x145 ;
  assign n10786 = n10785 ^ n7832 ^ 1'b0 ;
  assign n10787 = n10781 | n10786 ;
  assign n10788 = n3361 & ~n8932 ;
  assign n10789 = n10788 ^ n1450 ^ 1'b0 ;
  assign n10790 = n4699 ^ n2912 ^ 1'b0 ;
  assign n10791 = n6452 & n10790 ;
  assign n10792 = n10789 & n10791 ;
  assign n10793 = n10792 ^ n2638 ^ 1'b0 ;
  assign n10794 = n1877 & ~n4523 ;
  assign n10795 = ~n542 & n1149 ;
  assign n10796 = n10794 & n10795 ;
  assign n10797 = n10793 | n10796 ;
  assign n10798 = n1867 | n10797 ;
  assign n10799 = ( n947 & ~n4974 ) | ( n947 & n10798 ) | ( ~n4974 & n10798 ) ;
  assign n10810 = n5430 | n6642 ;
  assign n10811 = n10810 ^ n9002 ^ 1'b0 ;
  assign n10801 = n7468 ^ n6319 ^ n923 ;
  assign n10802 = n3044 & n10801 ;
  assign n10803 = n10802 ^ n394 ^ 1'b0 ;
  assign n10800 = n2351 & n8985 ;
  assign n10804 = n10803 ^ n10800 ^ 1'b0 ;
  assign n10805 = n10804 ^ n6870 ^ 1'b0 ;
  assign n10806 = ( n715 & n8456 ) | ( n715 & ~n10805 ) | ( n8456 & ~n10805 ) ;
  assign n10807 = n8361 ^ n7808 ^ 1'b0 ;
  assign n10808 = n10806 | n10807 ;
  assign n10809 = n5471 | n10808 ;
  assign n10812 = n10811 ^ n10809 ^ 1'b0 ;
  assign n10813 = n5156 ^ n1285 ^ 1'b0 ;
  assign n10814 = ~n863 & n10813 ;
  assign n10815 = ~n1110 & n10814 ;
  assign n10816 = ~n5706 & n10815 ;
  assign n10817 = ~n2942 & n7719 ;
  assign n10818 = n10816 | n10817 ;
  assign n10820 = n8406 ^ n559 ^ 1'b0 ;
  assign n10819 = ~n7209 & n8715 ;
  assign n10821 = n10820 ^ n10819 ^ 1'b0 ;
  assign n10822 = ~n1755 & n6913 ;
  assign n10823 = n4443 | n9800 ;
  assign n10824 = n10823 ^ n5948 ^ 1'b0 ;
  assign n10825 = x42 | n10824 ;
  assign n10826 = n4498 & ~n5975 ;
  assign n10827 = ~n4637 & n5549 ;
  assign n10828 = n10728 & n10827 ;
  assign n10829 = n10122 ^ n4376 ^ n3433 ;
  assign n10830 = n10829 ^ n3211 ^ n1133 ;
  assign n10831 = n10830 ^ n4371 ^ 1'b0 ;
  assign n10832 = n10828 | n10831 ;
  assign n10833 = n9299 ^ n2230 ^ 1'b0 ;
  assign n10834 = n4498 & n7373 ;
  assign n10835 = n5801 & n10102 ;
  assign n10836 = n8315 ^ n5198 ^ 1'b0 ;
  assign n10837 = n5938 ^ n399 ^ 1'b0 ;
  assign n10838 = ~n10836 & n10837 ;
  assign n10839 = ( ~n1475 & n3406 ) | ( ~n1475 & n5058 ) | ( n3406 & n5058 ) ;
  assign n10840 = n10839 ^ n967 ^ 1'b0 ;
  assign n10841 = ( ~n2118 & n3607 ) | ( ~n2118 & n4388 ) | ( n3607 & n4388 ) ;
  assign n10842 = ( n3016 & n5288 ) | ( n3016 & ~n6615 ) | ( n5288 & ~n6615 ) ;
  assign n10843 = n10842 ^ n3196 ^ 1'b0 ;
  assign n10844 = n6232 & n10843 ;
  assign n10845 = n6661 | n9743 ;
  assign n10846 = ( ~n2697 & n3132 ) | ( ~n2697 & n9230 ) | ( n3132 & n9230 ) ;
  assign n10847 = n10846 ^ n2086 ^ 1'b0 ;
  assign n10848 = n563 & n10847 ;
  assign n10849 = n5789 ^ n2767 ^ 1'b0 ;
  assign n10850 = n10140 & ~n10849 ;
  assign n10851 = n10850 ^ n6958 ^ 1'b0 ;
  assign n10852 = ( n3160 & n10848 ) | ( n3160 & ~n10851 ) | ( n10848 & ~n10851 ) ;
  assign n10853 = n10058 ^ n2278 ^ 1'b0 ;
  assign n10854 = n4559 ^ n4209 ^ n2381 ;
  assign n10855 = n3547 & n10854 ;
  assign n10856 = n10855 ^ n7919 ^ 1'b0 ;
  assign n10857 = n10856 ^ n6093 ^ 1'b0 ;
  assign n10858 = ~n1825 & n10753 ;
  assign n10859 = n4977 & n10858 ;
  assign n10860 = n8403 ^ n2987 ^ 1'b0 ;
  assign n10861 = n10860 ^ n6910 ^ n6256 ;
  assign n10862 = n5027 | n6041 ;
  assign n10863 = n4743 & n4875 ;
  assign n10864 = n5770 & n10680 ;
  assign n10865 = n10863 & n10864 ;
  assign n10866 = ( ~n1254 & n10862 ) | ( ~n1254 & n10865 ) | ( n10862 & n10865 ) ;
  assign n10867 = ~n3866 & n4308 ;
  assign n10868 = ~n4308 & n10867 ;
  assign n10869 = n1923 & ~n10868 ;
  assign n10870 = n10868 & n10869 ;
  assign n10871 = n10870 ^ n10830 ^ n5712 ;
  assign n10872 = n1685 | n9025 ;
  assign n10873 = n10872 ^ n4988 ^ 1'b0 ;
  assign n10874 = n1284 & n8442 ;
  assign n10875 = n10874 ^ n576 ^ 1'b0 ;
  assign n10876 = ~n1298 & n10875 ;
  assign n10877 = ~n4301 & n10876 ;
  assign n10878 = n4493 & ~n10877 ;
  assign n10879 = n10878 ^ n10814 ^ 1'b0 ;
  assign n10880 = n10873 & ~n10879 ;
  assign n10881 = n10880 ^ n7559 ^ 1'b0 ;
  assign n10882 = n2009 & ~n9217 ;
  assign n10883 = ~n6456 & n10272 ;
  assign n10884 = n3836 & n10883 ;
  assign n10885 = ( n5032 & n9765 ) | ( n5032 & ~n10884 ) | ( n9765 & ~n10884 ) ;
  assign n10886 = n5761 ^ n4441 ^ n1361 ;
  assign n10891 = n2387 ^ n1523 ^ 1'b0 ;
  assign n10887 = n2055 & ~n2921 ;
  assign n10888 = n9729 & n10887 ;
  assign n10889 = ( n802 & ~n2236 ) | ( n802 & n5807 ) | ( ~n2236 & n5807 ) ;
  assign n10890 = ~n10888 & n10889 ;
  assign n10892 = n10891 ^ n10890 ^ 1'b0 ;
  assign n10893 = ~n5798 & n7125 ;
  assign n10894 = ~n10892 & n10893 ;
  assign n10895 = ~n3113 & n7101 ;
  assign n10896 = n3157 ^ n952 ^ x7 ;
  assign n10897 = n5093 & ~n10896 ;
  assign n10898 = ~n7948 & n10897 ;
  assign n10899 = n2259 | n10898 ;
  assign n10906 = ~n2819 & n3970 ;
  assign n10907 = ( n1953 & n8492 ) | ( n1953 & n10906 ) | ( n8492 & n10906 ) ;
  assign n10908 = n4228 & ~n10907 ;
  assign n10909 = ~n1495 & n10908 ;
  assign n10900 = n5759 ^ n1902 ^ 1'b0 ;
  assign n10901 = n1976 & n10900 ;
  assign n10902 = n10901 ^ n3658 ^ 1'b0 ;
  assign n10903 = n3928 & ~n10902 ;
  assign n10904 = n2488 & n10903 ;
  assign n10905 = n9147 | n10904 ;
  assign n10910 = n10909 ^ n10905 ^ 1'b0 ;
  assign n10911 = n1840 & ~n4723 ;
  assign n10912 = n10911 ^ n5923 ^ 1'b0 ;
  assign n10913 = ( n1895 & ~n9290 ) | ( n1895 & n10912 ) | ( ~n9290 & n10912 ) ;
  assign n10914 = n3849 ^ n2726 ^ n1128 ;
  assign n10915 = n10914 ^ n9567 ^ n5747 ;
  assign n10916 = n10264 ^ x197 ^ 1'b0 ;
  assign n10917 = n1201 & ~n10916 ;
  assign n10918 = ~n6861 & n10917 ;
  assign n10919 = n3022 ^ n771 ^ 1'b0 ;
  assign n10920 = n3624 & ~n4495 ;
  assign n10921 = ~n5311 & n10920 ;
  assign n10922 = ( n2389 & ~n2396 ) | ( n2389 & n8463 ) | ( ~n2396 & n8463 ) ;
  assign n10923 = ( n3219 & ~n3413 ) | ( n3219 & n10922 ) | ( ~n3413 & n10922 ) ;
  assign n10924 = n10923 ^ n8171 ^ n2356 ;
  assign n10925 = n5747 | n5976 ;
  assign n10926 = n10925 ^ n8009 ^ n5355 ;
  assign n10927 = n1310 ^ n1190 ^ 1'b0 ;
  assign n10928 = n10927 ^ n3919 ^ 1'b0 ;
  assign n10929 = n10928 ^ n2857 ^ 1'b0 ;
  assign n10930 = n5739 & ~n10929 ;
  assign n10931 = n263 ^ x176 ^ 1'b0 ;
  assign n10932 = ~n5219 & n7263 ;
  assign n10933 = ~n992 & n10932 ;
  assign n10934 = ~n1946 & n10933 ;
  assign n10935 = n10934 ^ n2261 ^ 1'b0 ;
  assign n10936 = ~n3007 & n10935 ;
  assign n10937 = n936 ^ x20 ^ 1'b0 ;
  assign n10938 = ( n1081 & ~n10416 ) | ( n1081 & n10937 ) | ( ~n10416 & n10937 ) ;
  assign n10939 = n3847 & n5052 ;
  assign n10941 = n3492 ^ n3100 ^ 1'b0 ;
  assign n10940 = n4059 ^ n3900 ^ 1'b0 ;
  assign n10942 = n10941 ^ n10940 ^ n6738 ;
  assign n10943 = n10942 ^ n4013 ^ n3432 ;
  assign n10944 = n4797 & ~n8520 ;
  assign n10945 = ~n4455 & n10944 ;
  assign n10946 = n3545 & ~n3821 ;
  assign n10947 = n3314 & n10946 ;
  assign n10948 = ~n2742 & n10947 ;
  assign n10949 = x202 & ~n2823 ;
  assign n10950 = ~n2719 & n10949 ;
  assign n10951 = n10950 ^ n3401 ^ 1'b0 ;
  assign n10952 = x180 & ~n10951 ;
  assign n10954 = ( n3504 & ~n6196 ) | ( n3504 & n6463 ) | ( ~n6196 & n6463 ) ;
  assign n10953 = n10777 ^ n7617 ^ n2095 ;
  assign n10955 = n10954 ^ n10953 ^ n3600 ;
  assign n10956 = x68 & n10955 ;
  assign n10957 = n10956 ^ n3153 ^ 1'b0 ;
  assign n10959 = n1399 ^ n1149 ^ x199 ;
  assign n10960 = n559 & n10959 ;
  assign n10961 = n10453 ^ n7390 ^ 1'b0 ;
  assign n10962 = n1433 & n10961 ;
  assign n10963 = n10960 & n10962 ;
  assign n10958 = n1937 & ~n2332 ;
  assign n10964 = n10963 ^ n10958 ^ n5928 ;
  assign n10965 = ~n6206 & n10964 ;
  assign n10966 = n10965 ^ n688 ^ 1'b0 ;
  assign n10967 = n3679 ^ n2703 ^ 1'b0 ;
  assign n10968 = ~n3212 & n10967 ;
  assign n10969 = n10968 ^ n3896 ^ n667 ;
  assign n10970 = n7789 ^ n2822 ^ 1'b0 ;
  assign n10971 = ( ~n5177 & n10969 ) | ( ~n5177 & n10970 ) | ( n10969 & n10970 ) ;
  assign n10972 = n3731 & ~n9882 ;
  assign n10973 = ~n6014 & n10972 ;
  assign n10974 = n7361 ^ n6993 ^ 1'b0 ;
  assign n10975 = ~n1113 & n9406 ;
  assign n10976 = ~n2990 & n10975 ;
  assign n10977 = ( ~n3755 & n5594 ) | ( ~n3755 & n10976 ) | ( n5594 & n10976 ) ;
  assign n10978 = ( n1440 & n2021 ) | ( n1440 & n10977 ) | ( n2021 & n10977 ) ;
  assign n10979 = n10041 & ~n10978 ;
  assign n10980 = ~n8029 & n10979 ;
  assign n10981 = n7573 ^ n6850 ^ n4500 ;
  assign n10982 = n7755 ^ n2182 ^ 1'b0 ;
  assign n10983 = n10982 ^ n4829 ^ 1'b0 ;
  assign n10984 = n10981 & ~n10983 ;
  assign n10985 = ~n6540 & n10984 ;
  assign n10986 = ~n4792 & n10985 ;
  assign n10987 = n1923 & n4888 ;
  assign n10988 = n10987 ^ n10751 ^ 1'b0 ;
  assign n10990 = n9586 ^ n3839 ^ 1'b0 ;
  assign n10991 = n1955 ^ n1672 ^ 1'b0 ;
  assign n10992 = ~n10990 & n10991 ;
  assign n10989 = n9864 ^ n5433 ^ 1'b0 ;
  assign n10993 = n10992 ^ n10989 ^ n9415 ;
  assign n10994 = n10993 ^ n4615 ^ 1'b0 ;
  assign n10995 = n2643 & ~n4016 ;
  assign n10996 = n10995 ^ n1909 ^ 1'b0 ;
  assign n10997 = n6597 ^ n4736 ^ 1'b0 ;
  assign n10998 = n4617 & ~n10997 ;
  assign n10999 = n9729 & n10998 ;
  assign n11000 = n10999 ^ n6384 ^ n2043 ;
  assign n11001 = n2102 ^ x227 ^ 1'b0 ;
  assign n11002 = n8422 ^ n1037 ^ 1'b0 ;
  assign n11003 = n5160 | n11002 ;
  assign n11004 = n2654 & ~n11003 ;
  assign n11005 = ~n2208 & n11004 ;
  assign n11006 = ~n8071 & n9306 ;
  assign n11007 = n11005 & n11006 ;
  assign n11008 = ( n9297 & n11001 ) | ( n9297 & ~n11007 ) | ( n11001 & ~n11007 ) ;
  assign n11010 = n3702 | n5710 ;
  assign n11009 = n3900 & ~n4713 ;
  assign n11011 = n11010 ^ n11009 ^ n6449 ;
  assign n11012 = ( n1943 & n4911 ) | ( n1943 & ~n11011 ) | ( n4911 & ~n11011 ) ;
  assign n11014 = n1850 | n4747 ;
  assign n11015 = n11014 ^ n9659 ^ 1'b0 ;
  assign n11013 = ( n574 & n1794 ) | ( n574 & n6653 ) | ( n1794 & n6653 ) ;
  assign n11016 = n11015 ^ n11013 ^ 1'b0 ;
  assign n11017 = ~n6159 & n11016 ;
  assign n11018 = n6688 & n10323 ;
  assign n11019 = n11018 ^ n3307 ^ 1'b0 ;
  assign n11021 = n4138 ^ n904 ^ 1'b0 ;
  assign n11022 = n1821 & ~n11021 ;
  assign n11020 = ( n256 & ~n2116 ) | ( n256 & n3475 ) | ( ~n2116 & n3475 ) ;
  assign n11023 = n11022 ^ n11020 ^ n7800 ;
  assign n11024 = n9101 | n9822 ;
  assign n11025 = n1194 | n11024 ;
  assign n11026 = n6222 ^ n1442 ^ 1'b0 ;
  assign n11027 = n8398 ^ n2513 ^ 1'b0 ;
  assign n11028 = ( n6538 & n11026 ) | ( n6538 & ~n11027 ) | ( n11026 & ~n11027 ) ;
  assign n11029 = n10555 ^ n7827 ^ n5376 ;
  assign n11030 = n4913 ^ n1332 ^ 1'b0 ;
  assign n11031 = n955 | n11030 ;
  assign n11032 = n11031 ^ n1821 ^ n1468 ;
  assign n11033 = n11032 ^ n3826 ^ n1977 ;
  assign n11035 = ( ~n5317 & n9198 ) | ( ~n5317 & n10522 ) | ( n9198 & n10522 ) ;
  assign n11034 = n8183 | n10116 ;
  assign n11036 = n11035 ^ n11034 ^ 1'b0 ;
  assign n11037 = ~n898 & n11036 ;
  assign n11038 = n3432 ^ n717 ^ 1'b0 ;
  assign n11039 = ~n6558 & n11038 ;
  assign n11040 = ~n1211 & n11039 ;
  assign n11041 = ~n6870 & n11040 ;
  assign n11042 = ~n1131 & n3795 ;
  assign n11043 = n11042 ^ n966 ^ 1'b0 ;
  assign n11047 = n8338 ^ n7887 ^ n1336 ;
  assign n11048 = ~n5931 & n11047 ;
  assign n11045 = n2737 ^ n1981 ^ 1'b0 ;
  assign n11044 = n1504 ^ n1174 ^ 1'b0 ;
  assign n11046 = n11045 ^ n11044 ^ n8969 ;
  assign n11049 = n11048 ^ n11046 ^ 1'b0 ;
  assign n11050 = n11043 & ~n11049 ;
  assign n11051 = n3978 & n6695 ;
  assign n11052 = n11051 ^ n6041 ^ n4496 ;
  assign n11053 = n303 | n2746 ;
  assign n11054 = ( n3776 & n7213 ) | ( n3776 & ~n11053 ) | ( n7213 & ~n11053 ) ;
  assign n11055 = n11054 ^ n6996 ^ 1'b0 ;
  assign n11056 = ~n1937 & n5554 ;
  assign n11057 = n3204 ^ n2937 ^ 1'b0 ;
  assign n11058 = ~n4977 & n11057 ;
  assign n11059 = n11058 ^ n6802 ^ 1'b0 ;
  assign n11060 = ~n5503 & n7442 ;
  assign n11061 = n11059 & n11060 ;
  assign n11062 = ~n11056 & n11061 ;
  assign n11063 = ~n1579 & n4760 ;
  assign n11064 = n11063 ^ n9381 ^ 1'b0 ;
  assign n11065 = n2567 & ~n2842 ;
  assign n11066 = n8372 & n11065 ;
  assign n11069 = n5744 ^ n810 ^ 1'b0 ;
  assign n11070 = ~n2185 & n11069 ;
  assign n11067 = n962 | n6024 ;
  assign n11068 = n591 | n11067 ;
  assign n11071 = n11070 ^ n11068 ^ 1'b0 ;
  assign n11072 = ~n11066 & n11071 ;
  assign n11073 = ( n8124 & n10378 ) | ( n8124 & ~n11072 ) | ( n10378 & ~n11072 ) ;
  assign n11074 = ( n1863 & n5752 ) | ( n1863 & n5817 ) | ( n5752 & n5817 ) ;
  assign n11076 = n5397 ^ n2157 ^ n1448 ;
  assign n11075 = n1138 | n5118 ;
  assign n11077 = n11076 ^ n11075 ^ 1'b0 ;
  assign n11079 = n3776 & n7404 ;
  assign n11080 = n11079 ^ n900 ^ 1'b0 ;
  assign n11078 = n10688 ^ n3907 ^ n706 ;
  assign n11081 = n11080 ^ n11078 ^ n6620 ;
  assign n11082 = ~n11077 & n11081 ;
  assign n11083 = ~n2085 & n9620 ;
  assign n11084 = n11083 ^ n4993 ^ 1'b0 ;
  assign n11085 = n8623 ^ n3296 ^ n1115 ;
  assign n11086 = n11085 ^ n1053 ^ 1'b0 ;
  assign n11087 = n3998 & ~n11086 ;
  assign n11088 = n10129 ^ n1182 ^ 1'b0 ;
  assign n11089 = ~n8449 & n11088 ;
  assign n11090 = ( n1506 & n3784 ) | ( n1506 & n6688 ) | ( n3784 & n6688 ) ;
  assign n11091 = n6914 & ~n11090 ;
  assign n11092 = n1639 & n2157 ;
  assign n11093 = ~n1187 & n11092 ;
  assign n11094 = ~n2205 & n10875 ;
  assign n11095 = n3113 & n11094 ;
  assign n11096 = n11093 | n11095 ;
  assign n11097 = n11096 ^ n9656 ^ 1'b0 ;
  assign n11098 = ~n1039 & n1354 ;
  assign n11099 = n11098 ^ n966 ^ 1'b0 ;
  assign n11100 = n11099 ^ n8153 ^ n6109 ;
  assign n11101 = n11100 ^ n6888 ^ n2183 ;
  assign n11102 = n2924 ^ n866 ^ 1'b0 ;
  assign n11103 = n11101 & n11102 ;
  assign n11107 = x90 & ~n2138 ;
  assign n11108 = n11107 ^ n3696 ^ 1'b0 ;
  assign n11106 = n7165 ^ n5584 ^ n3591 ;
  assign n11104 = n7180 ^ n573 ^ 1'b0 ;
  assign n11105 = n11104 ^ n8563 ^ n5492 ;
  assign n11109 = n11108 ^ n11106 ^ n11105 ;
  assign n11110 = ( n572 & n3835 ) | ( n572 & n6229 ) | ( n3835 & n6229 ) ;
  assign n11111 = n6667 & n11110 ;
  assign n11112 = n3231 & ~n7220 ;
  assign n11113 = n7104 | n11112 ;
  assign n11114 = n10130 & ~n11113 ;
  assign n11115 = n5859 & ~n6223 ;
  assign n11116 = n3437 ^ n3254 ^ n1201 ;
  assign n11117 = n11116 ^ n7752 ^ 1'b0 ;
  assign n11118 = n8971 | n11117 ;
  assign n11119 = n6624 ^ x98 ^ 1'b0 ;
  assign n11120 = ~n11118 & n11119 ;
  assign n11121 = n1476 & n11120 ;
  assign n11122 = ~n5935 & n9803 ;
  assign n11127 = n3304 ^ x214 ^ 1'b0 ;
  assign n11128 = n3049 & ~n11127 ;
  assign n11124 = ~n2133 & n10801 ;
  assign n11125 = n11124 ^ n3051 ^ 1'b0 ;
  assign n11123 = n1530 | n1701 ;
  assign n11126 = n11125 ^ n11123 ^ 1'b0 ;
  assign n11129 = n11128 ^ n11126 ^ 1'b0 ;
  assign n11130 = n7425 ^ n2615 ^ 1'b0 ;
  assign n11131 = n11129 & n11130 ;
  assign n11132 = n5699 & ~n7430 ;
  assign n11133 = n10333 & n11132 ;
  assign n11134 = ~n440 & n9332 ;
  assign n11135 = n11134 ^ n351 ^ 1'b0 ;
  assign n11136 = n1851 & n11135 ;
  assign n11137 = n11136 ^ n3277 ^ 1'b0 ;
  assign n11138 = n4162 ^ x233 ^ 1'b0 ;
  assign n11139 = n3423 & ~n11138 ;
  assign n11140 = n2621 ^ n1131 ^ n928 ;
  assign n11141 = n11140 ^ n7017 ^ 1'b0 ;
  assign n11142 = n3759 | n11141 ;
  assign n11143 = ( n6737 & n6767 ) | ( n6737 & ~n7708 ) | ( n6767 & ~n7708 ) ;
  assign n11144 = n8979 ^ n6373 ^ 1'b0 ;
  assign n11145 = n10804 & ~n11144 ;
  assign n11146 = n11145 ^ n7384 ^ n1480 ;
  assign n11152 = n7046 ^ n1550 ^ n390 ;
  assign n11153 = n6046 ^ x33 ^ 1'b0 ;
  assign n11154 = ~n11152 & n11153 ;
  assign n11151 = n7333 ^ n4318 ^ n1703 ;
  assign n11155 = n11154 ^ n11151 ^ 1'b0 ;
  assign n11156 = ~n958 & n11155 ;
  assign n11147 = n7715 ^ n6634 ^ 1'b0 ;
  assign n11148 = n11147 ^ n6875 ^ n2860 ;
  assign n11149 = n11148 ^ n10564 ^ 1'b0 ;
  assign n11150 = n3700 & ~n11149 ;
  assign n11157 = n11156 ^ n11150 ^ 1'b0 ;
  assign n11158 = n7047 ^ n973 ^ 1'b0 ;
  assign n11159 = ~n1042 & n11158 ;
  assign n11160 = n2015 & n2042 ;
  assign n11161 = n8831 & n11160 ;
  assign n11162 = n10301 ^ n8145 ^ n7305 ;
  assign n11163 = ( n6515 & n8926 ) | ( n6515 & n9775 ) | ( n8926 & n9775 ) ;
  assign n11164 = ~n500 & n4306 ;
  assign n11165 = n11164 ^ n5377 ^ 1'b0 ;
  assign n11166 = ~n11163 & n11165 ;
  assign n11167 = n7316 & n11166 ;
  assign n11168 = n2688 & n3637 ;
  assign n11169 = n7973 & ~n11168 ;
  assign n11170 = n1755 | n1795 ;
  assign n11171 = ~n2635 & n11170 ;
  assign n11173 = n7386 ^ n576 ^ 1'b0 ;
  assign n11172 = n3939 ^ n2406 ^ 1'b0 ;
  assign n11174 = n11173 ^ n11172 ^ n1050 ;
  assign n11175 = n8559 ^ n337 ^ 1'b0 ;
  assign n11176 = n1755 & n11175 ;
  assign n11177 = n9285 & ~n9561 ;
  assign n11178 = n11177 ^ n4258 ^ 1'b0 ;
  assign n11179 = ( ~n2344 & n3915 ) | ( ~n2344 & n4004 ) | ( n3915 & n4004 ) ;
  assign n11180 = n11178 & n11179 ;
  assign n11181 = ~n5119 & n5699 ;
  assign n11182 = ( ~n5345 & n9598 ) | ( ~n5345 & n11181 ) | ( n9598 & n11181 ) ;
  assign n11183 = n3236 ^ n2222 ^ 1'b0 ;
  assign n11184 = x74 & n11183 ;
  assign n11185 = n11184 ^ n11056 ^ n4747 ;
  assign n11187 = n3338 ^ n1666 ^ 1'b0 ;
  assign n11186 = ( n3730 & n3784 ) | ( n3730 & n6439 ) | ( n3784 & n6439 ) ;
  assign n11188 = n11187 ^ n11186 ^ n2967 ;
  assign n11189 = n11185 & ~n11188 ;
  assign n11190 = n10409 ^ n2386 ^ n266 ;
  assign n11191 = n3587 | n9986 ;
  assign n11192 = n7721 ^ n2174 ^ n335 ;
  assign n11193 = n3737 & n11192 ;
  assign n11194 = ~x79 & n11193 ;
  assign n11196 = n8172 ^ n639 ^ 1'b0 ;
  assign n11197 = n11196 ^ n831 ^ 1'b0 ;
  assign n11195 = ~n2451 & n7743 ;
  assign n11198 = n11197 ^ n11195 ^ 1'b0 ;
  assign n11199 = ( ~n6014 & n11194 ) | ( ~n6014 & n11198 ) | ( n11194 & n11198 ) ;
  assign n11200 = n11199 ^ n6914 ^ 1'b0 ;
  assign n11201 = n4689 ^ n2391 ^ 1'b0 ;
  assign n11202 = ~n7285 & n11201 ;
  assign n11203 = ( n1442 & n3169 ) | ( n1442 & ~n9818 ) | ( n3169 & ~n9818 ) ;
  assign n11204 = n11203 ^ n6046 ^ 1'b0 ;
  assign n11205 = n11202 | n11204 ;
  assign n11206 = n2699 & ~n11205 ;
  assign n11213 = n11135 ^ n500 ^ 1'b0 ;
  assign n11214 = n859 | n11213 ;
  assign n11207 = n7570 ^ n826 ^ 1'b0 ;
  assign n11208 = n4703 ^ n1725 ^ 1'b0 ;
  assign n11209 = ~n9794 & n11208 ;
  assign n11210 = ( n5213 & n10095 ) | ( n5213 & n11209 ) | ( n10095 & n11209 ) ;
  assign n11211 = n11210 ^ n4197 ^ n2259 ;
  assign n11212 = ~n11207 & n11211 ;
  assign n11215 = n11214 ^ n11212 ^ 1'b0 ;
  assign n11216 = n2476 & n7573 ;
  assign n11217 = ~n1435 & n9222 ;
  assign n11218 = n4256 & n11217 ;
  assign n11219 = n3985 & n11218 ;
  assign n11220 = n3723 & ~n11219 ;
  assign n11221 = n11220 ^ n5541 ^ 1'b0 ;
  assign n11222 = ~n10413 & n11221 ;
  assign n11223 = ~n11216 & n11222 ;
  assign n11224 = n9097 ^ n7338 ^ 1'b0 ;
  assign n11225 = n4256 & n11224 ;
  assign n11226 = n8104 ^ n7801 ^ 1'b0 ;
  assign n11227 = n11225 & n11226 ;
  assign n11228 = n4397 | n6779 ;
  assign n11229 = n11228 ^ n3842 ^ 1'b0 ;
  assign n11230 = ( n3919 & n9147 ) | ( n3919 & n11229 ) | ( n9147 & n11229 ) ;
  assign n11231 = n3638 & n9660 ;
  assign n11232 = n7077 ^ x79 ^ 1'b0 ;
  assign n11233 = n3394 & ~n7721 ;
  assign n11234 = ~n6929 & n11233 ;
  assign n11235 = n11234 ^ n2536 ^ x57 ;
  assign n11236 = ( n4529 & ~n11232 ) | ( n4529 & n11235 ) | ( ~n11232 & n11235 ) ;
  assign n11239 = n877 & n7238 ;
  assign n11240 = n4558 & n11239 ;
  assign n11237 = ~n489 & n1713 ;
  assign n11238 = n11237 ^ n7416 ^ 1'b0 ;
  assign n11241 = n11240 ^ n11238 ^ 1'b0 ;
  assign n11242 = x12 & n11241 ;
  assign n11243 = ( n5472 & n9332 ) | ( n5472 & ~n11242 ) | ( n9332 & ~n11242 ) ;
  assign n11244 = n3952 | n9391 ;
  assign n11245 = n11244 ^ n8102 ^ 1'b0 ;
  assign n11246 = n3204 ^ n1467 ^ 1'b0 ;
  assign n11247 = n11246 ^ n5126 ^ n269 ;
  assign n11248 = n11247 ^ n4013 ^ n939 ;
  assign n11249 = ( n5445 & ~n6606 ) | ( n5445 & n6847 ) | ( ~n6606 & n6847 ) ;
  assign n11250 = n6636 ^ n4817 ^ 1'b0 ;
  assign n11251 = n9845 & n11250 ;
  assign n11252 = ( n327 & n6990 ) | ( n327 & n11251 ) | ( n6990 & n11251 ) ;
  assign n11253 = n11252 ^ n8829 ^ 1'b0 ;
  assign n11254 = n10964 & ~n11253 ;
  assign n11255 = n1043 | n3539 ;
  assign n11256 = n11255 ^ n4060 ^ 1'b0 ;
  assign n11257 = n7240 ^ n3575 ^ n490 ;
  assign n11258 = n8043 & ~n11257 ;
  assign n11259 = n403 & ~n5294 ;
  assign n11260 = n5639 | n6892 ;
  assign n11261 = n3585 | n11260 ;
  assign n11262 = n11259 & ~n11261 ;
  assign n11263 = n7305 & ~n7532 ;
  assign n11264 = ~n2279 & n11263 ;
  assign n11265 = ~n4172 & n6430 ;
  assign n11266 = ~n1201 & n11265 ;
  assign n11267 = n3152 & ~n11266 ;
  assign n11268 = n11267 ^ n6264 ^ 1'b0 ;
  assign n11269 = n11268 ^ n7163 ^ 1'b0 ;
  assign n11270 = n6747 ^ n5287 ^ n2911 ;
  assign n11271 = n8404 ^ n3516 ^ 1'b0 ;
  assign n11272 = n1104 & ~n11271 ;
  assign n11273 = n11272 ^ n1273 ^ 1'b0 ;
  assign n11274 = n3487 | n11273 ;
  assign n11275 = n11270 & n11274 ;
  assign n11276 = ~n11269 & n11275 ;
  assign n11277 = n1350 | n5919 ;
  assign n11278 = n11277 ^ n1963 ^ 1'b0 ;
  assign n11279 = n9326 & ~n11278 ;
  assign n11280 = n11279 ^ n571 ^ 1'b0 ;
  assign n11281 = n11276 | n11280 ;
  assign n11282 = n4449 ^ n1994 ^ 1'b0 ;
  assign n11283 = n266 & ~n11282 ;
  assign n11284 = n11283 ^ n2006 ^ 1'b0 ;
  assign n11285 = ( ~n608 & n1593 ) | ( ~n608 & n2888 ) | ( n1593 & n2888 ) ;
  assign n11286 = n11285 ^ n4744 ^ n4449 ;
  assign n11288 = n10537 ^ n6182 ^ n410 ;
  assign n11287 = n6532 | n6773 ;
  assign n11289 = n11288 ^ n11287 ^ 1'b0 ;
  assign n11290 = ( n1403 & ~n10394 ) | ( n1403 & n11289 ) | ( ~n10394 & n11289 ) ;
  assign n11291 = n9954 ^ n468 ^ 1'b0 ;
  assign n11293 = n4827 ^ n1002 ^ 1'b0 ;
  assign n11294 = n7376 | n11293 ;
  assign n11295 = n11294 ^ n8017 ^ 1'b0 ;
  assign n11292 = ~n1047 & n8965 ;
  assign n11296 = n11295 ^ n11292 ^ 1'b0 ;
  assign n11297 = n6624 ^ n3242 ^ 1'b0 ;
  assign n11298 = n9582 & ~n11297 ;
  assign n11302 = n1549 & n9000 ;
  assign n11299 = n5353 ^ n1820 ^ n1522 ;
  assign n11300 = n2066 & ~n5642 ;
  assign n11301 = ( n8818 & n11299 ) | ( n8818 & ~n11300 ) | ( n11299 & ~n11300 ) ;
  assign n11303 = n11302 ^ n11301 ^ 1'b0 ;
  assign n11304 = n5213 | n8937 ;
  assign n11305 = n402 | n4048 ;
  assign n11306 = n11305 ^ n9658 ^ 1'b0 ;
  assign n11307 = n8909 ^ n6643 ^ 1'b0 ;
  assign n11308 = ~n11306 & n11307 ;
  assign n11309 = n6250 & n9677 ;
  assign n11310 = n11309 ^ n7384 ^ 1'b0 ;
  assign n11311 = n5952 ^ n2991 ^ 1'b0 ;
  assign n11312 = n9050 | n9627 ;
  assign n11314 = x9 & ~n5215 ;
  assign n11315 = n11314 ^ n7293 ^ 1'b0 ;
  assign n11313 = n6820 ^ n3100 ^ n654 ;
  assign n11316 = n11315 ^ n11313 ^ 1'b0 ;
  assign n11317 = n2083 & ~n11316 ;
  assign n11318 = n2078 & ~n2901 ;
  assign n11319 = n3674 & ~n11318 ;
  assign n11320 = n11319 ^ n5397 ^ 1'b0 ;
  assign n11321 = n10811 ^ n5843 ^ 1'b0 ;
  assign n11322 = ~n11320 & n11321 ;
  assign n11323 = n9812 & n11322 ;
  assign n11324 = ~n10463 & n11323 ;
  assign n11325 = ( ~n1620 & n2110 ) | ( ~n1620 & n9156 ) | ( n2110 & n9156 ) ;
  assign n11326 = n6274 & ~n10748 ;
  assign n11327 = n11326 ^ x140 ^ 1'b0 ;
  assign n11328 = n5973 ^ n4930 ^ 1'b0 ;
  assign n11329 = n5111 ^ n4751 ^ n4234 ;
  assign n11330 = n2867 ^ n405 ^ 1'b0 ;
  assign n11331 = n4202 ^ n986 ^ x6 ;
  assign n11332 = n11331 ^ n2791 ^ n1321 ;
  assign n11333 = n7919 | n11332 ;
  assign n11334 = n2806 | n11333 ;
  assign n11335 = n11330 & n11334 ;
  assign n11336 = ~x155 & n11335 ;
  assign n11337 = n4147 ^ n757 ^ 1'b0 ;
  assign n11338 = n4411 & ~n11337 ;
  assign n11340 = ( n518 & n717 ) | ( n518 & n5712 ) | ( n717 & n5712 ) ;
  assign n11341 = n11340 ^ n9161 ^ n3798 ;
  assign n11339 = n6571 & ~n6752 ;
  assign n11342 = n11341 ^ n11339 ^ 1'b0 ;
  assign n11343 = n11342 ^ n2401 ^ 1'b0 ;
  assign n11344 = n6783 & n11343 ;
  assign n11346 = x232 & ~n335 ;
  assign n11347 = n11346 ^ n4458 ^ 1'b0 ;
  assign n11345 = n10403 ^ n7003 ^ n6528 ;
  assign n11348 = n11347 ^ n11345 ^ n9045 ;
  assign n11351 = n269 & ~n2056 ;
  assign n11352 = x198 | n11351 ;
  assign n11353 = n11352 ^ n7632 ^ 1'b0 ;
  assign n11349 = n8309 ^ n5226 ^ n2715 ;
  assign n11350 = n11349 ^ n7368 ^ n3109 ;
  assign n11354 = n11353 ^ n11350 ^ 1'b0 ;
  assign n11355 = n3015 & ~n11354 ;
  assign n11356 = n9632 & n10842 ;
  assign n11357 = n11356 ^ n5836 ^ 1'b0 ;
  assign n11358 = ( x85 & n2173 ) | ( x85 & n3391 ) | ( n2173 & n3391 ) ;
  assign n11359 = ~n7320 & n11358 ;
  assign n11360 = n941 & n3736 ;
  assign n11361 = n11360 ^ n1844 ^ 1'b0 ;
  assign n11362 = n9062 ^ n2903 ^ 1'b0 ;
  assign n11363 = n1229 ^ n341 ^ 1'b0 ;
  assign n11364 = n7279 & n11363 ;
  assign n11365 = n675 & n11364 ;
  assign n11366 = n9174 ^ n6720 ^ 1'b0 ;
  assign n11367 = ( x241 & n11365 ) | ( x241 & n11366 ) | ( n11365 & n11366 ) ;
  assign n11368 = ~n2986 & n4611 ;
  assign n11369 = n2863 & n11368 ;
  assign n11370 = n11369 ^ n3314 ^ 1'b0 ;
  assign n11371 = n11370 ^ n8756 ^ n5344 ;
  assign n11372 = n2025 ^ x101 ^ 1'b0 ;
  assign n11373 = n11372 ^ n952 ^ 1'b0 ;
  assign n11374 = n8544 & n8623 ;
  assign n11375 = ~n6627 & n11374 ;
  assign n11376 = n2070 & ~n5257 ;
  assign n11377 = n2823 | n6031 ;
  assign n11378 = n3934 & ~n11377 ;
  assign n11379 = n11376 & n11378 ;
  assign n11380 = ~n922 & n9188 ;
  assign n11381 = ( x95 & x214 ) | ( x95 & ~x239 ) | ( x214 & ~x239 ) ;
  assign n11382 = ~n5032 & n5316 ;
  assign n11383 = ~n11381 & n11382 ;
  assign n11384 = ( n928 & n1736 ) | ( n928 & ~n11383 ) | ( n1736 & ~n11383 ) ;
  assign n11385 = n8104 ^ n1933 ^ 1'b0 ;
  assign n11386 = n11384 | n11385 ;
  assign n11387 = n11380 & ~n11386 ;
  assign n11388 = n6810 ^ n5513 ^ 1'b0 ;
  assign n11389 = ~n4314 & n11388 ;
  assign n11390 = ~n9934 & n11389 ;
  assign n11391 = ( n7764 & ~n9200 ) | ( n7764 & n9741 ) | ( ~n9200 & n9741 ) ;
  assign n11392 = n10179 ^ n7661 ^ 1'b0 ;
  assign n11393 = n1441 ^ n1351 ^ n807 ;
  assign n11394 = n4111 & n9694 ;
  assign n11395 = n11393 & n11394 ;
  assign n11396 = n569 | n11395 ;
  assign n11397 = n11396 ^ n2362 ^ 1'b0 ;
  assign n11399 = ( n362 & ~n2494 ) | ( n362 & n7289 ) | ( ~n2494 & n7289 ) ;
  assign n11398 = ( n3040 & ~n3398 ) | ( n3040 & n4987 ) | ( ~n3398 & n4987 ) ;
  assign n11400 = n11399 ^ n11398 ^ n8299 ;
  assign n11401 = n11400 ^ n3496 ^ 1'b0 ;
  assign n11403 = n5106 ^ n4747 ^ 1'b0 ;
  assign n11404 = ~n8181 & n11403 ;
  assign n11405 = n11404 ^ n7646 ^ 1'b0 ;
  assign n11402 = ~n5429 & n7883 ;
  assign n11406 = n11405 ^ n11402 ^ 1'b0 ;
  assign n11407 = n4070 ^ n1653 ^ 1'b0 ;
  assign n11408 = ( x160 & n3599 ) | ( x160 & ~n5710 ) | ( n3599 & ~n5710 ) ;
  assign n11409 = ( n7235 & n11407 ) | ( n7235 & n11408 ) | ( n11407 & n11408 ) ;
  assign n11415 = ( n945 & n2023 ) | ( n945 & ~n5992 ) | ( n2023 & ~n5992 ) ;
  assign n11416 = n5754 ^ n374 ^ 1'b0 ;
  assign n11417 = n11416 ^ n1593 ^ 1'b0 ;
  assign n11418 = n11415 & n11417 ;
  assign n11410 = n1434 | n2515 ;
  assign n11411 = n6305 & n11410 ;
  assign n11412 = n11411 ^ n7560 ^ 1'b0 ;
  assign n11413 = ~n9478 & n11412 ;
  assign n11414 = n4189 & n11413 ;
  assign n11419 = n11418 ^ n11414 ^ 1'b0 ;
  assign n11420 = n10571 | n11419 ;
  assign n11421 = n5947 ^ n3674 ^ 1'b0 ;
  assign n11422 = n6450 & ~n11421 ;
  assign n11423 = n845 & n2832 ;
  assign n11424 = ~n11422 & n11423 ;
  assign n11425 = ~n10595 & n11424 ;
  assign n11426 = n490 | n6411 ;
  assign n11427 = n1323 | n7774 ;
  assign n11428 = n11426 & ~n11427 ;
  assign n11429 = n6417 & ~n11428 ;
  assign n11430 = n5412 ^ n379 ^ 1'b0 ;
  assign n11431 = n11430 ^ n2607 ^ n1810 ;
  assign n11434 = ( n1617 & n2266 ) | ( n1617 & ~n2386 ) | ( n2266 & ~n2386 ) ;
  assign n11432 = ( n2836 & n3652 ) | ( n2836 & n6133 ) | ( n3652 & n6133 ) ;
  assign n11433 = n4334 & ~n11432 ;
  assign n11435 = n11434 ^ n11433 ^ 1'b0 ;
  assign n11436 = n4144 ^ n2355 ^ 1'b0 ;
  assign n11437 = n3547 & ~n11436 ;
  assign n11438 = n2397 & n11437 ;
  assign n11439 = n3231 & n11438 ;
  assign n11440 = ( n6774 & n11435 ) | ( n6774 & n11439 ) | ( n11435 & n11439 ) ;
  assign n11441 = n6999 ^ n1890 ^ 1'b0 ;
  assign n11442 = n11441 ^ n9173 ^ 1'b0 ;
  assign n11443 = ~n1900 & n7068 ;
  assign n11444 = n11443 ^ n7442 ^ 1'b0 ;
  assign n11445 = n1489 | n4258 ;
  assign n11446 = n11445 ^ n1409 ^ 1'b0 ;
  assign n11447 = n11446 ^ n9329 ^ n3777 ;
  assign n11448 = n11447 ^ n4522 ^ 1'b0 ;
  assign n11449 = n4134 | n7417 ;
  assign n11450 = n10390 ^ n8089 ^ 1'b0 ;
  assign n11451 = n4816 & n11450 ;
  assign n11452 = ( n320 & ~n11449 ) | ( n320 & n11451 ) | ( ~n11449 & n11451 ) ;
  assign n11453 = n1405 & ~n9861 ;
  assign n11454 = n3404 & n11453 ;
  assign n11455 = ( ~n3072 & n4889 ) | ( ~n3072 & n9869 ) | ( n4889 & n9869 ) ;
  assign n11456 = ( n1562 & n1780 ) | ( n1562 & n11455 ) | ( n1780 & n11455 ) ;
  assign n11457 = n5778 ^ n1685 ^ n1397 ;
  assign n11458 = ~n2363 & n9643 ;
  assign n11459 = n11458 ^ n6316 ^ 1'b0 ;
  assign n11460 = n4838 & n11459 ;
  assign n11461 = n11460 ^ n6708 ^ 1'b0 ;
  assign n11462 = n11461 ^ n3869 ^ 1'b0 ;
  assign n11463 = ~n1505 & n7051 ;
  assign n11464 = ~n6988 & n11463 ;
  assign n11465 = n11462 & n11464 ;
  assign n11466 = ( n7471 & ~n8386 ) | ( n7471 & n9755 ) | ( ~n8386 & n9755 ) ;
  assign n11467 = x21 & n5255 ;
  assign n11471 = n3191 & ~n4031 ;
  assign n11468 = n4598 & n5786 ;
  assign n11469 = n4176 & n11468 ;
  assign n11470 = n11469 ^ n1190 ^ 1'b0 ;
  assign n11472 = n11471 ^ n11470 ^ x136 ;
  assign n11473 = ~n5762 & n7271 ;
  assign n11474 = n11472 & n11473 ;
  assign n11475 = ( n8945 & ~n11467 ) | ( n8945 & n11474 ) | ( ~n11467 & n11474 ) ;
  assign n11476 = n4565 & ~n6165 ;
  assign n11477 = n11475 & n11476 ;
  assign n11478 = x67 & n5782 ;
  assign n11479 = n2541 & n11478 ;
  assign n11480 = n1890 & n5119 ;
  assign n11481 = ( n2102 & n3458 ) | ( n2102 & n3529 ) | ( n3458 & n3529 ) ;
  assign n11482 = n11481 ^ n8763 ^ 1'b0 ;
  assign n11483 = x144 | n11482 ;
  assign n11485 = n3376 | n10011 ;
  assign n11484 = n2443 ^ n2038 ^ 1'b0 ;
  assign n11486 = n11485 ^ n11484 ^ 1'b0 ;
  assign n11487 = x244 & ~n5582 ;
  assign n11488 = n8818 & n11487 ;
  assign n11489 = n11488 ^ n7042 ^ n4172 ;
  assign n11490 = ( ~n3685 & n4330 ) | ( ~n3685 & n11489 ) | ( n4330 & n11489 ) ;
  assign n11491 = n5857 ^ n5361 ^ 1'b0 ;
  assign n11492 = n952 & ~n4806 ;
  assign n11493 = n11492 ^ n3351 ^ 1'b0 ;
  assign n11494 = n3049 & ~n3796 ;
  assign n11495 = n3735 & n11494 ;
  assign n11496 = n11495 ^ x73 ^ 1'b0 ;
  assign n11497 = n10032 & ~n11496 ;
  assign n11498 = n11497 ^ n11229 ^ 1'b0 ;
  assign n11499 = ~n4346 & n11498 ;
  assign n11500 = n2697 ^ x119 ^ 1'b0 ;
  assign n11501 = n435 & ~n11500 ;
  assign n11502 = n9800 ^ n517 ^ 1'b0 ;
  assign n11503 = n11502 ^ x89 ^ 1'b0 ;
  assign n11504 = n10999 & n11503 ;
  assign n11505 = n6469 ^ x229 ^ 1'b0 ;
  assign n11506 = n9665 ^ n6437 ^ 1'b0 ;
  assign n11508 = n3418 & ~n4472 ;
  assign n11509 = ~n7582 & n11508 ;
  assign n11507 = n3596 & ~n7160 ;
  assign n11510 = n11509 ^ n11507 ^ 1'b0 ;
  assign n11511 = n505 & n8399 ;
  assign n11512 = ~n5878 & n11511 ;
  assign n11513 = n11512 ^ n7015 ^ 1'b0 ;
  assign n11514 = n1705 & ~n8398 ;
  assign n11515 = n11514 ^ n9185 ^ 1'b0 ;
  assign n11516 = n1152 & ~n11515 ;
  assign n11517 = n7391 & ~n11516 ;
  assign n11518 = n2780 & ~n11517 ;
  assign n11519 = ( ~n3970 & n11513 ) | ( ~n3970 & n11518 ) | ( n11513 & n11518 ) ;
  assign n11520 = n4080 | n10777 ;
  assign n11521 = n11520 ^ n7929 ^ n1666 ;
  assign n11522 = ( n1802 & n3532 ) | ( n1802 & n11521 ) | ( n3532 & n11521 ) ;
  assign n11523 = ( x192 & ~n5761 ) | ( x192 & n11522 ) | ( ~n5761 & n11522 ) ;
  assign n11524 = n5638 | n9620 ;
  assign n11525 = n11524 ^ n6847 ^ 1'b0 ;
  assign n11526 = n6486 ^ n6039 ^ 1'b0 ;
  assign n11527 = n4575 & ~n11526 ;
  assign n11528 = n11527 ^ n9997 ^ 1'b0 ;
  assign n11529 = n11525 & ~n11528 ;
  assign n11530 = n3514 ^ n1126 ^ 1'b0 ;
  assign n11531 = ( ~n1187 & n3207 ) | ( ~n1187 & n5372 ) | ( n3207 & n5372 ) ;
  assign n11532 = n11531 ^ n3608 ^ 1'b0 ;
  assign n11533 = n11532 ^ n1890 ^ 1'b0 ;
  assign n11534 = ~n11530 & n11533 ;
  assign n11535 = n10529 ^ n6530 ^ n5462 ;
  assign n11536 = ( n2005 & ~n8429 ) | ( n2005 & n11535 ) | ( ~n8429 & n11535 ) ;
  assign n11537 = ~n1888 & n2178 ;
  assign n11538 = n11537 ^ n2145 ^ 1'b0 ;
  assign n11539 = n8091 ^ n5650 ^ n1809 ;
  assign n11540 = ~n11538 & n11539 ;
  assign n11544 = n6439 ^ n5655 ^ 1'b0 ;
  assign n11545 = ~n6041 & n11544 ;
  assign n11543 = n3631 & n4863 ;
  assign n11546 = n11545 ^ n11543 ^ 1'b0 ;
  assign n11547 = ~n1890 & n11546 ;
  assign n11548 = n11547 ^ n6393 ^ 1'b0 ;
  assign n11541 = n2174 & ~n8538 ;
  assign n11542 = ~n3758 & n11541 ;
  assign n11549 = n11548 ^ n11542 ^ 1'b0 ;
  assign n11550 = n426 | n6375 ;
  assign n11551 = n1434 & n11550 ;
  assign n11552 = n3037 & ~n11551 ;
  assign n11553 = n1455 & ~n8971 ;
  assign n11554 = n4695 & n11553 ;
  assign n11555 = n1202 | n11554 ;
  assign n11556 = x112 & ~n6777 ;
  assign n11557 = n11556 ^ n4206 ^ 1'b0 ;
  assign n11558 = n5357 | n11557 ;
  assign n11559 = n580 | n11558 ;
  assign n11560 = n9601 ^ n4016 ^ 1'b0 ;
  assign n11561 = n11559 & n11560 ;
  assign n11562 = n11561 ^ n8280 ^ n7777 ;
  assign n11563 = ( ~n5389 & n7032 ) | ( ~n5389 & n7468 ) | ( n7032 & n7468 ) ;
  assign n11564 = n11563 ^ n1910 ^ 1'b0 ;
  assign n11565 = n5215 & n11564 ;
  assign n11566 = n11565 ^ n345 ^ 1'b0 ;
  assign n11567 = n9098 ^ n5815 ^ 1'b0 ;
  assign n11568 = n11567 ^ n9333 ^ n1865 ;
  assign n11569 = n11568 ^ n7317 ^ 1'b0 ;
  assign n11570 = n2939 & n11569 ;
  assign n11571 = n5253 ^ n3494 ^ 1'b0 ;
  assign n11572 = ~n4876 & n11571 ;
  assign n11574 = n9933 ^ n9251 ^ 1'b0 ;
  assign n11573 = n8807 & ~n9802 ;
  assign n11575 = n11574 ^ n11573 ^ 1'b0 ;
  assign n11576 = ~n1270 & n5610 ;
  assign n11577 = ( n612 & n1050 ) | ( n612 & n11576 ) | ( n1050 & n11576 ) ;
  assign n11578 = n2583 | n5702 ;
  assign n11580 = ( ~x240 & n1651 ) | ( ~x240 & n1913 ) | ( n1651 & n1913 ) ;
  assign n11581 = ( ~n1034 & n1934 ) | ( ~n1034 & n11580 ) | ( n1934 & n11580 ) ;
  assign n11582 = n11581 ^ n1993 ^ 1'b0 ;
  assign n11583 = n11582 ^ n7058 ^ n6471 ;
  assign n11579 = n1516 | n2677 ;
  assign n11584 = n11583 ^ n11579 ^ n8934 ;
  assign n11585 = n11584 ^ n9511 ^ 1'b0 ;
  assign n11586 = ( n363 & ~n1510 ) | ( n363 & n2678 ) | ( ~n1510 & n2678 ) ;
  assign n11587 = n402 & n3370 ;
  assign n11588 = n11587 ^ x178 ^ 1'b0 ;
  assign n11589 = n571 | n1900 ;
  assign n11590 = ~n389 & n11589 ;
  assign n11591 = n11590 ^ n6167 ^ 1'b0 ;
  assign n11592 = n11591 ^ n3516 ^ 1'b0 ;
  assign n11593 = n1076 | n1123 ;
  assign n11594 = n8404 | n11593 ;
  assign n11595 = n317 & ~n11594 ;
  assign n11596 = x78 & n11595 ;
  assign n11597 = n8521 ^ x235 ^ 1'b0 ;
  assign n11598 = n1472 | n3062 ;
  assign n11599 = ( n3944 & n5104 ) | ( n3944 & ~n11598 ) | ( n5104 & ~n11598 ) ;
  assign n11600 = ( x142 & n2565 ) | ( x142 & ~n11599 ) | ( n2565 & ~n11599 ) ;
  assign n11601 = ( n11596 & n11597 ) | ( n11596 & n11600 ) | ( n11597 & n11600 ) ;
  assign n11602 = ~n2888 & n7233 ;
  assign n11603 = n11602 ^ n6413 ^ 1'b0 ;
  assign n11604 = n8939 & n11215 ;
  assign n11605 = n7855 | n10194 ;
  assign n11606 = n11605 ^ n4014 ^ 1'b0 ;
  assign n11607 = n10310 & ~n11606 ;
  assign n11608 = n11607 ^ n1869 ^ 1'b0 ;
  assign n11609 = n462 & ~n9180 ;
  assign n11610 = n11609 ^ n6708 ^ 1'b0 ;
  assign n11611 = n4669 & ~n7916 ;
  assign n11612 = n7892 ^ n2243 ^ n402 ;
  assign n11613 = n5170 ^ n2019 ^ n1583 ;
  assign n11614 = n4518 & n10267 ;
  assign n11615 = ~n11613 & n11614 ;
  assign n11616 = n10776 ^ n6749 ^ 1'b0 ;
  assign n11617 = ~n11615 & n11616 ;
  assign n11618 = n599 & n4117 ;
  assign n11619 = ~n2453 & n8715 ;
  assign n11623 = ~n9622 & n10122 ;
  assign n11620 = n5190 ^ n2504 ^ n838 ;
  assign n11621 = n11620 ^ n5677 ^ 1'b0 ;
  assign n11622 = n8802 & ~n11621 ;
  assign n11624 = n11623 ^ n11622 ^ n7172 ;
  assign n11625 = ( n3719 & n7697 ) | ( n3719 & n8987 ) | ( n7697 & n8987 ) ;
  assign n11626 = ( n678 & n4085 ) | ( n678 & n11625 ) | ( n4085 & n11625 ) ;
  assign n11627 = n11626 ^ n6555 ^ n1561 ;
  assign n11628 = n5761 ^ n936 ^ 1'b0 ;
  assign n11629 = n11628 ^ n8827 ^ n5105 ;
  assign n11630 = n3418 & ~n11629 ;
  assign n11631 = n11630 ^ n2199 ^ 1'b0 ;
  assign n11632 = n9266 & n10428 ;
  assign n11633 = n11632 ^ n1593 ^ 1'b0 ;
  assign n11634 = n1936 & n3318 ;
  assign n11635 = ( x42 & ~n11633 ) | ( x42 & n11634 ) | ( ~n11633 & n11634 ) ;
  assign n11636 = n7812 & ~n11635 ;
  assign n11640 = n323 & n573 ;
  assign n11641 = ~n573 & n11640 ;
  assign n11642 = n547 & ~n684 ;
  assign n11643 = ~n547 & n11642 ;
  assign n11644 = n11641 | n11643 ;
  assign n11645 = n11641 & ~n11644 ;
  assign n11646 = n3708 & ~n11645 ;
  assign n11647 = ~n3708 & n11646 ;
  assign n11637 = n1778 & n1976 ;
  assign n11638 = ~n1976 & n11637 ;
  assign n11639 = n4625 & ~n11638 ;
  assign n11648 = n11647 ^ n11639 ^ 1'b0 ;
  assign n11649 = n3327 | n6157 ;
  assign n11650 = ~n4561 & n10185 ;
  assign n11651 = n11650 ^ n3071 ^ 1'b0 ;
  assign n11652 = n11651 ^ n10968 ^ 1'b0 ;
  assign n11653 = ( ~n464 & n1336 ) | ( ~n464 & n1609 ) | ( n1336 & n1609 ) ;
  assign n11654 = n8585 & n11653 ;
  assign n11655 = n11654 ^ x194 ^ 1'b0 ;
  assign n11656 = ~n3726 & n7248 ;
  assign n11657 = n7750 & n11656 ;
  assign n11658 = n4013 | n11657 ;
  assign n11661 = ~n402 & n1799 ;
  assign n11662 = ~n3119 & n4690 ;
  assign n11663 = ~n320 & n11662 ;
  assign n11664 = n11663 ^ n11511 ^ n853 ;
  assign n11665 = ( n3974 & ~n11661 ) | ( n3974 & n11664 ) | ( ~n11661 & n11664 ) ;
  assign n11659 = n7990 ^ n7288 ^ n2613 ;
  assign n11660 = n2106 & n11659 ;
  assign n11666 = n11665 ^ n11660 ^ 1'b0 ;
  assign n11667 = n2141 ^ n1206 ^ x6 ;
  assign n11668 = ( n2976 & n6135 ) | ( n2976 & n11667 ) | ( n6135 & n11667 ) ;
  assign n11669 = n3009 ^ x46 ^ 1'b0 ;
  assign n11678 = n3700 & n9941 ;
  assign n11670 = n2216 & ~n7072 ;
  assign n11672 = n1943 & n3843 ;
  assign n11673 = ~x243 & n11672 ;
  assign n11674 = ( ~n6444 & n8571 ) | ( ~n6444 & n11673 ) | ( n8571 & n11673 ) ;
  assign n11671 = n5155 & ~n9187 ;
  assign n11675 = n11674 ^ n11671 ^ 1'b0 ;
  assign n11676 = n9062 | n11675 ;
  assign n11677 = n11670 & ~n11676 ;
  assign n11679 = n11678 ^ n11677 ^ 1'b0 ;
  assign n11680 = n10181 ^ n6377 ^ n3578 ;
  assign n11681 = n3220 | n11680 ;
  assign n11682 = n11681 ^ n5645 ^ 1'b0 ;
  assign n11683 = n4930 & n9099 ;
  assign n11684 = n11683 ^ n6010 ^ 1'b0 ;
  assign n11685 = n3508 & ~n11684 ;
  assign n11686 = n4515 & n11685 ;
  assign n11687 = ( n3725 & n4612 ) | ( n3725 & ~n11686 ) | ( n4612 & ~n11686 ) ;
  assign n11688 = x159 & ~n11687 ;
  assign n11689 = n5386 & n11688 ;
  assign n11690 = n2041 & n9700 ;
  assign n11691 = n11690 ^ n10947 ^ 1'b0 ;
  assign n11692 = n11691 ^ n1030 ^ 1'b0 ;
  assign n11693 = ~n5426 & n7591 ;
  assign n11694 = n11693 ^ n3644 ^ n3152 ;
  assign n11695 = n2518 & n4945 ;
  assign n11696 = n11695 ^ n2459 ^ 1'b0 ;
  assign n11697 = n9847 | n11696 ;
  assign n11698 = n1359 & n3600 ;
  assign n11699 = n11698 ^ n4638 ^ 1'b0 ;
  assign n11700 = n11699 ^ n11416 ^ 1'b0 ;
  assign n11701 = n10041 & n11700 ;
  assign n11702 = n2955 & ~n4805 ;
  assign n11703 = n11702 ^ n6515 ^ 1'b0 ;
  assign n11704 = ( n3190 & n5025 ) | ( n3190 & ~n11593 ) | ( n5025 & ~n11593 ) ;
  assign n11705 = ~n11703 & n11704 ;
  assign n11706 = ~n11701 & n11705 ;
  assign n11707 = n5251 & ~n8856 ;
  assign n11708 = n2527 & ~n11707 ;
  assign n11709 = ( n2405 & ~n8276 ) | ( n2405 & n11708 ) | ( ~n8276 & n11708 ) ;
  assign n11710 = ( n7062 & ~n8279 ) | ( n7062 & n11709 ) | ( ~n8279 & n11709 ) ;
  assign n11711 = n9477 ^ n9246 ^ n5949 ;
  assign n11712 = ( n4050 & n7932 ) | ( n4050 & n11711 ) | ( n7932 & n11711 ) ;
  assign n11713 = n9364 ^ n2990 ^ 1'b0 ;
  assign n11714 = n1232 & ~n11713 ;
  assign n11715 = n11714 ^ n4720 ^ x155 ;
  assign n11716 = n11715 ^ n4974 ^ 1'b0 ;
  assign n11717 = n3590 ^ x179 ^ 1'b0 ;
  assign n11718 = n7407 & n11717 ;
  assign n11719 = ~n10024 & n11718 ;
  assign n11720 = ~n5638 & n11719 ;
  assign n11721 = n11720 ^ n7780 ^ 1'b0 ;
  assign n11722 = n2169 ^ n1359 ^ 1'b0 ;
  assign n11725 = ~n5058 & n5328 ;
  assign n11726 = n11725 ^ n5996 ^ 1'b0 ;
  assign n11727 = n11726 ^ n3591 ^ 1'b0 ;
  assign n11728 = ~n10443 & n11727 ;
  assign n11723 = ( n1365 & n2857 ) | ( n1365 & ~n7653 ) | ( n2857 & ~n7653 ) ;
  assign n11724 = n5107 | n11723 ;
  assign n11729 = n11728 ^ n11724 ^ 1'b0 ;
  assign n11730 = n11529 ^ n5611 ^ 1'b0 ;
  assign n11731 = n2724 | n11730 ;
  assign n11732 = n6999 ^ n1810 ^ 1'b0 ;
  assign n11733 = n4542 & n11732 ;
  assign n11734 = n8792 ^ n2718 ^ 1'b0 ;
  assign n11735 = n438 | n11734 ;
  assign n11736 = n11735 ^ n10323 ^ n7885 ;
  assign n11737 = n3255 & n9426 ;
  assign n11738 = n7543 ^ n7305 ^ 1'b0 ;
  assign n11739 = n11737 & ~n11738 ;
  assign n11740 = n6461 | n10960 ;
  assign n11741 = n11740 ^ x198 ^ 1'b0 ;
  assign n11742 = x87 & n11741 ;
  assign n11743 = ~n11739 & n11742 ;
  assign n11744 = n11301 ^ n10851 ^ 1'b0 ;
  assign n11747 = n647 & ~n6046 ;
  assign n11745 = n7641 ^ n5914 ^ 1'b0 ;
  assign n11746 = n3736 & n11745 ;
  assign n11748 = n11747 ^ n11746 ^ 1'b0 ;
  assign n11749 = n11748 ^ n610 ^ 1'b0 ;
  assign n11750 = n3062 | n5671 ;
  assign n11751 = ~n1641 & n11750 ;
  assign n11752 = n5014 ^ n4531 ^ 1'b0 ;
  assign n11753 = ~n5121 & n11752 ;
  assign n11754 = ( n6400 & n9536 ) | ( n6400 & n11753 ) | ( n9536 & n11753 ) ;
  assign n11755 = n11751 & n11754 ;
  assign n11756 = ~n5692 & n11755 ;
  assign n11757 = x141 & n515 ;
  assign n11758 = ( n442 & ~n7741 ) | ( n442 & n11757 ) | ( ~n7741 & n11757 ) ;
  assign n11759 = n4548 & n11758 ;
  assign n11760 = ( n4419 & n8201 ) | ( n4419 & n11759 ) | ( n8201 & n11759 ) ;
  assign n11764 = ~n3997 & n4696 ;
  assign n11765 = ( n1775 & n6430 ) | ( n1775 & n11764 ) | ( n6430 & n11764 ) ;
  assign n11761 = n1423 ^ n1006 ^ 1'b0 ;
  assign n11762 = n11761 ^ n8540 ^ 1'b0 ;
  assign n11763 = n2435 | n11762 ;
  assign n11766 = n11765 ^ n11763 ^ 1'b0 ;
  assign n11767 = n2032 & n3166 ;
  assign n11768 = n4214 | n11767 ;
  assign n11769 = n11768 ^ n5740 ^ n4338 ;
  assign n11773 = n4395 & n5934 ;
  assign n11774 = n11773 ^ n5991 ^ 1'b0 ;
  assign n11770 = x131 & ~n6435 ;
  assign n11771 = n11770 ^ n1685 ^ 1'b0 ;
  assign n11772 = ( ~x118 & n557 ) | ( ~x118 & n11771 ) | ( n557 & n11771 ) ;
  assign n11775 = n11774 ^ n11772 ^ 1'b0 ;
  assign n11780 = n3922 & n4049 ;
  assign n11781 = n5053 & n11780 ;
  assign n11782 = n11781 ^ n7412 ^ n4985 ;
  assign n11783 = n11782 ^ n3812 ^ n1696 ;
  assign n11776 = n2412 & ~n4155 ;
  assign n11777 = ~n1451 & n11776 ;
  assign n11778 = ( n6408 & n6649 ) | ( n6408 & ~n11777 ) | ( n6649 & ~n11777 ) ;
  assign n11779 = n11778 ^ n10727 ^ n2958 ;
  assign n11784 = n11783 ^ n11779 ^ n6581 ;
  assign n11785 = n11784 ^ n4007 ^ 1'b0 ;
  assign n11786 = n5033 | n11785 ;
  assign n11787 = n4065 & ~n11028 ;
  assign n11788 = n11787 ^ x212 ^ 1'b0 ;
  assign n11791 = ( ~n6551 & n7730 ) | ( ~n6551 & n7892 ) | ( n7730 & n7892 ) ;
  assign n11789 = x81 ^ x4 ^ 1'b0 ;
  assign n11790 = n11789 ^ n5494 ^ 1'b0 ;
  assign n11792 = n11791 ^ n11790 ^ n8207 ;
  assign n11793 = ( n848 & n2017 ) | ( n848 & ~n2639 ) | ( n2017 & ~n2639 ) ;
  assign n11794 = n3381 & ~n5572 ;
  assign n11795 = n11794 ^ n11659 ^ 1'b0 ;
  assign n11796 = ( n8794 & n9754 ) | ( n8794 & n11432 ) | ( n9754 & n11432 ) ;
  assign n11797 = n1199 & n6627 ;
  assign n11798 = n8801 & n11797 ;
  assign n11799 = n3208 | n11798 ;
  assign n11800 = n11796 & ~n11799 ;
  assign n11801 = n2164 & ~n11800 ;
  assign n11802 = n2663 ^ n887 ^ 1'b0 ;
  assign n11803 = n936 ^ n807 ^ 1'b0 ;
  assign n11804 = ( n3696 & ~n11802 ) | ( n3696 & n11803 ) | ( ~n11802 & n11803 ) ;
  assign n11805 = ( n1452 & n3188 ) | ( n1452 & ~n8929 ) | ( n3188 & ~n8929 ) ;
  assign n11806 = n9000 ^ n3620 ^ x67 ;
  assign n11807 = n11805 & ~n11806 ;
  assign n11808 = n11807 ^ n10149 ^ 1'b0 ;
  assign n11809 = ( n806 & ~n936 ) | ( n806 & n6353 ) | ( ~n936 & n6353 ) ;
  assign n11810 = n7070 & ~n11809 ;
  assign n11811 = n11810 ^ n3617 ^ 1'b0 ;
  assign n11812 = n9232 ^ n7813 ^ 1'b0 ;
  assign n11813 = n11811 & n11812 ;
  assign n11814 = n11813 ^ n10796 ^ 1'b0 ;
  assign n11815 = n1074 & n7732 ;
  assign n11816 = n5584 ^ n2162 ^ 1'b0 ;
  assign n11817 = n11815 & ~n11816 ;
  assign n11818 = n10356 ^ n5629 ^ 1'b0 ;
  assign n11819 = n11817 & n11818 ;
  assign n11821 = n1427 | n2622 ;
  assign n11822 = n11821 ^ n1486 ^ 1'b0 ;
  assign n11820 = x56 & ~n4273 ;
  assign n11823 = n11822 ^ n11820 ^ 1'b0 ;
  assign n11831 = ~n1138 & n3639 ;
  assign n11832 = ~n3639 & n11831 ;
  assign n11833 = n1709 & ~n11832 ;
  assign n11824 = n572 | n667 ;
  assign n11825 = n667 & ~n11824 ;
  assign n11826 = ~n1395 & n4979 ;
  assign n11827 = n11825 & n11826 ;
  assign n11828 = ~n1450 & n11827 ;
  assign n11829 = n8589 & n11828 ;
  assign n11830 = n1359 & n11829 ;
  assign n11834 = n11833 ^ n11830 ^ 1'b0 ;
  assign n11835 = ~n3027 & n11834 ;
  assign n11837 = ( n2009 & n4417 ) | ( n2009 & n9378 ) | ( n4417 & n9378 ) ;
  assign n11836 = ~n6848 & n9337 ;
  assign n11838 = n11837 ^ n11836 ^ 1'b0 ;
  assign n11839 = n11838 ^ n9919 ^ n435 ;
  assign n11840 = ( n4404 & n5637 ) | ( n4404 & n11839 ) | ( n5637 & n11839 ) ;
  assign n11841 = n7293 ^ n3592 ^ 1'b0 ;
  assign n11842 = ( n3403 & ~n10707 ) | ( n3403 & n11651 ) | ( ~n10707 & n11651 ) ;
  assign n11843 = n7899 ^ n2674 ^ 1'b0 ;
  assign n11844 = ~n447 & n4580 ;
  assign n11845 = ( n7051 & ~n11843 ) | ( n7051 & n11844 ) | ( ~n11843 & n11844 ) ;
  assign n11846 = n11845 ^ n10516 ^ 1'b0 ;
  assign n11847 = n10138 ^ n5229 ^ 1'b0 ;
  assign n11848 = n5624 & n11847 ;
  assign n11849 = ~n3360 & n11848 ;
  assign n11850 = n853 & n5763 ;
  assign n11851 = n11850 ^ x76 ^ 1'b0 ;
  assign n11852 = n11851 ^ n1899 ^ n284 ;
  assign n11853 = n11852 ^ n3750 ^ 1'b0 ;
  assign n11854 = n11853 ^ n5987 ^ 1'b0 ;
  assign n11855 = n3068 & n4086 ;
  assign n11856 = n7562 ^ n3605 ^ 1'b0 ;
  assign n11857 = ( n457 & n713 ) | ( n457 & ~n5078 ) | ( n713 & ~n5078 ) ;
  assign n11858 = n7622 ^ n7266 ^ 1'b0 ;
  assign n11859 = n951 & ~n1524 ;
  assign n11860 = n11859 ^ n631 ^ 1'b0 ;
  assign n11861 = n5185 ^ n3351 ^ 1'b0 ;
  assign n11862 = n1291 & n3314 ;
  assign n11863 = ~n11861 & n11862 ;
  assign n11864 = n11860 & ~n11863 ;
  assign n11865 = n11864 ^ n1439 ^ 1'b0 ;
  assign n11866 = n2171 & ~n7650 ;
  assign n11867 = n401 | n4454 ;
  assign n11872 = n3624 & n7528 ;
  assign n11873 = n11872 ^ n2860 ^ 1'b0 ;
  assign n11870 = n5919 & n9775 ;
  assign n11871 = n973 & ~n11870 ;
  assign n11874 = n11873 ^ n11871 ^ 1'b0 ;
  assign n11869 = ~n795 & n1010 ;
  assign n11875 = n11874 ^ n11869 ^ 1'b0 ;
  assign n11868 = n1672 & n6127 ;
  assign n11876 = n11875 ^ n11868 ^ x235 ;
  assign n11877 = ( n8631 & n9085 ) | ( n8631 & ~n11876 ) | ( n9085 & ~n11876 ) ;
  assign n11878 = ( n3312 & ~n9608 ) | ( n3312 & n9966 ) | ( ~n9608 & n9966 ) ;
  assign n11879 = n1388 & ~n2726 ;
  assign n11880 = n11879 ^ n3126 ^ 1'b0 ;
  assign n11881 = n9296 ^ n8526 ^ 1'b0 ;
  assign n11882 = n2375 & n11881 ;
  assign n11883 = ( n2976 & ~n10044 ) | ( n2976 & n11882 ) | ( ~n10044 & n11882 ) ;
  assign n11884 = n11880 & n11883 ;
  assign n11885 = n3109 & n8269 ;
  assign n11886 = n11885 ^ n1063 ^ 1'b0 ;
  assign n11887 = n1290 | n2453 ;
  assign n11888 = n6587 & ~n11887 ;
  assign n11889 = n3456 & n11888 ;
  assign n11890 = n11889 ^ n11540 ^ 1'b0 ;
  assign n11891 = n8167 ^ n797 ^ x92 ;
  assign n11892 = n10597 & n11891 ;
  assign n11893 = ( n5172 & ~n6517 ) | ( n5172 & n9198 ) | ( ~n6517 & n9198 ) ;
  assign n11894 = ~n3567 & n6878 ;
  assign n11895 = ~n1598 & n11894 ;
  assign n11896 = n8045 ^ n4176 ^ 1'b0 ;
  assign n11897 = ~n11895 & n11896 ;
  assign n11898 = ( n2678 & n11893 ) | ( n2678 & ~n11897 ) | ( n11893 & ~n11897 ) ;
  assign n11899 = n4886 ^ n3857 ^ 1'b0 ;
  assign n11900 = n10407 & ~n11899 ;
  assign n11901 = n8067 ^ n2760 ^ 1'b0 ;
  assign n11902 = n3479 & ~n11901 ;
  assign n11903 = n2722 ^ n2515 ^ n901 ;
  assign n11904 = n2611 | n11903 ;
  assign n11905 = n11902 | n11904 ;
  assign n11906 = ~n4696 & n11905 ;
  assign n11907 = ~n4870 & n11906 ;
  assign n11908 = n1794 & ~n3590 ;
  assign n11909 = ( n4862 & n7697 ) | ( n4862 & n11908 ) | ( n7697 & n11908 ) ;
  assign n11910 = ( n2154 & ~n5460 ) | ( n2154 & n11909 ) | ( ~n5460 & n11909 ) ;
  assign n11911 = n9509 & ~n11910 ;
  assign n11912 = ~n1995 & n11911 ;
  assign n11913 = n11912 ^ n9857 ^ n5627 ;
  assign n11914 = n1542 & n5602 ;
  assign n11915 = ~n10230 & n11914 ;
  assign n11916 = n4032 | n9222 ;
  assign n11917 = n11916 ^ n2770 ^ 1'b0 ;
  assign n11918 = x27 | n11917 ;
  assign n11919 = ~n7026 & n8705 ;
  assign n11920 = n11919 ^ n8913 ^ 1'b0 ;
  assign n11921 = ( n559 & ~n7173 ) | ( n559 & n11920 ) | ( ~n7173 & n11920 ) ;
  assign n11922 = n7686 & ~n11858 ;
  assign n11923 = n1037 & n11922 ;
  assign n11924 = x78 & n6260 ;
  assign n11925 = n4739 & n11924 ;
  assign n11926 = n11925 ^ n4013 ^ x94 ;
  assign n11931 = n5984 ^ n3798 ^ 1'b0 ;
  assign n11927 = n6105 ^ x131 ^ 1'b0 ;
  assign n11928 = ~n2937 & n11927 ;
  assign n11929 = n11928 ^ n8772 ^ 1'b0 ;
  assign n11930 = ~n2326 & n11929 ;
  assign n11932 = n11931 ^ n11930 ^ n2433 ;
  assign n11933 = ( n6200 & n8978 ) | ( n6200 & n11932 ) | ( n8978 & n11932 ) ;
  assign n11934 = n11933 ^ n1500 ^ x72 ;
  assign n11935 = ( ~n1622 & n2755 ) | ( ~n1622 & n4299 ) | ( n2755 & n4299 ) ;
  assign n11936 = n11935 ^ n5768 ^ n2828 ;
  assign n11937 = ~n257 & n11936 ;
  assign n11938 = n11937 ^ n7561 ^ 1'b0 ;
  assign n11939 = ( n1124 & ~n5764 ) | ( n1124 & n8465 ) | ( ~n5764 & n8465 ) ;
  assign n11940 = ~n6482 & n11939 ;
  assign n11941 = n11940 ^ n2092 ^ n1022 ;
  assign n11942 = n2294 ^ n1241 ^ 1'b0 ;
  assign n11943 = n3151 & ~n11942 ;
  assign n11944 = n11943 ^ n3217 ^ 1'b0 ;
  assign n11945 = n5535 ^ n2448 ^ 1'b0 ;
  assign n11946 = n11118 ^ n8454 ^ 1'b0 ;
  assign n11947 = ( n1341 & n11945 ) | ( n1341 & ~n11946 ) | ( n11945 & ~n11946 ) ;
  assign n11948 = n5374 & ~n11947 ;
  assign n11949 = n8231 & n11948 ;
  assign n11950 = n11303 ^ n1142 ^ 1'b0 ;
  assign n11951 = n1460 | n11950 ;
  assign n11952 = n4004 ^ n449 ^ 1'b0 ;
  assign n11953 = n2085 | n11952 ;
  assign n11954 = ( ~n520 & n8658 ) | ( ~n520 & n11953 ) | ( n8658 & n11953 ) ;
  assign n11955 = n7305 ^ n652 ^ 1'b0 ;
  assign n11956 = n1882 | n7345 ;
  assign n11957 = n11956 ^ n6209 ^ 1'b0 ;
  assign n11958 = n7759 ^ n4830 ^ 1'b0 ;
  assign n11959 = n3375 & n11958 ;
  assign n11960 = n5183 & ~n5466 ;
  assign n11961 = n11960 ^ n1709 ^ 1'b0 ;
  assign n11962 = n11961 ^ n11873 ^ 1'b0 ;
  assign n11963 = n1828 | n11962 ;
  assign n11967 = n4299 ^ n3984 ^ 1'b0 ;
  assign n11964 = n1832 | n7391 ;
  assign n11965 = n3950 & ~n11964 ;
  assign n11966 = n11965 ^ n5344 ^ 1'b0 ;
  assign n11968 = n11967 ^ n11966 ^ 1'b0 ;
  assign n11969 = n3219 ^ n1813 ^ 1'b0 ;
  assign n11970 = n11969 ^ n3592 ^ n2219 ;
  assign n11971 = n11970 ^ x157 ^ 1'b0 ;
  assign n11972 = n1882 | n11971 ;
  assign n11973 = n8600 & ~n11972 ;
  assign n11974 = n4104 | n8788 ;
  assign n11975 = ~n4007 & n5838 ;
  assign n11976 = n8052 & n11975 ;
  assign n11977 = ~n1244 & n4583 ;
  assign n11978 = n5742 | n7005 ;
  assign n11979 = n11978 ^ n7238 ^ 1'b0 ;
  assign n11980 = ~n11977 & n11979 ;
  assign n11981 = ~n7305 & n11980 ;
  assign n11982 = ( ~n1586 & n3071 ) | ( ~n1586 & n4552 ) | ( n3071 & n4552 ) ;
  assign n11983 = n11982 ^ n5907 ^ 1'b0 ;
  assign n11984 = ( n10023 & n11981 ) | ( n10023 & ~n11983 ) | ( n11981 & ~n11983 ) ;
  assign n11985 = n6406 & n7804 ;
  assign n11986 = n5528 | n11985 ;
  assign n11987 = n3159 | n11986 ;
  assign n11988 = x150 & n577 ;
  assign n11989 = n9860 ^ n4676 ^ 1'b0 ;
  assign n11990 = ( n9041 & n11988 ) | ( n9041 & ~n11989 ) | ( n11988 & ~n11989 ) ;
  assign n11996 = n6467 ^ n6129 ^ 1'b0 ;
  assign n11997 = ~n3406 & n11996 ;
  assign n11994 = ~n8365 & n9010 ;
  assign n11995 = ~n4121 & n11994 ;
  assign n11998 = n11997 ^ n11995 ^ 1'b0 ;
  assign n11999 = n7979 & ~n11998 ;
  assign n12000 = ~n807 & n11999 ;
  assign n12001 = n9916 ^ n8750 ^ 1'b0 ;
  assign n12002 = n12000 | n12001 ;
  assign n11991 = n6827 | n7282 ;
  assign n11992 = n11991 ^ x5 ^ 1'b0 ;
  assign n11993 = n3552 & n11992 ;
  assign n12003 = n12002 ^ n11993 ^ 1'b0 ;
  assign n12004 = ( n928 & n6393 ) | ( n928 & n7182 ) | ( n6393 & n7182 ) ;
  assign n12005 = n1865 | n4720 ;
  assign n12006 = ( x77 & n8449 ) | ( x77 & ~n12005 ) | ( n8449 & ~n12005 ) ;
  assign n12007 = ~n12004 & n12006 ;
  assign n12008 = n10974 & n12007 ;
  assign n12009 = ~n630 & n8709 ;
  assign n12010 = n12009 ^ n11903 ^ 1'b0 ;
  assign n12011 = ~n3923 & n9070 ;
  assign n12012 = n12011 ^ n7289 ^ n3449 ;
  assign n12013 = n1240 | n5996 ;
  assign n12014 = n12013 ^ n8801 ^ 1'b0 ;
  assign n12015 = n5938 ^ n3360 ^ n271 ;
  assign n12016 = n12015 ^ n8403 ^ 1'b0 ;
  assign n12017 = n2706 | n12016 ;
  assign n12018 = n3515 & n10639 ;
  assign n12019 = n12017 & n12018 ;
  assign n12020 = n12019 ^ n802 ^ 1'b0 ;
  assign n12021 = n12014 | n12020 ;
  assign n12022 = ~n11925 & n12021 ;
  assign n12023 = n10529 ^ n4557 ^ 1'b0 ;
  assign n12024 = n6571 ^ n6417 ^ 1'b0 ;
  assign n12025 = n2162 ^ x71 ^ 1'b0 ;
  assign n12026 = n748 & n12025 ;
  assign n12027 = n3163 | n12026 ;
  assign n12028 = n6493 | n12027 ;
  assign n12029 = n12028 ^ n9417 ^ 1'b0 ;
  assign n12030 = ~n2482 & n12029 ;
  assign n12031 = ~n5515 & n12030 ;
  assign n12032 = ~n9420 & n12031 ;
  assign n12034 = ~x194 & n4291 ;
  assign n12033 = n3396 | n9818 ;
  assign n12035 = n12034 ^ n12033 ^ 1'b0 ;
  assign n12036 = n12035 ^ n3327 ^ n1301 ;
  assign n12037 = n11598 ^ n6585 ^ n4589 ;
  assign n12038 = n12036 & ~n12037 ;
  assign n12039 = n1413 & ~n2369 ;
  assign n12040 = ~n12038 & n12039 ;
  assign n12041 = n3325 & ~n8128 ;
  assign n12042 = n9161 ^ n8732 ^ n4097 ;
  assign n12043 = n8837 ^ n1331 ^ n888 ;
  assign n12044 = ~n8202 & n12043 ;
  assign n12045 = ~n12043 & n12044 ;
  assign n12048 = n8024 ^ n4292 ^ 1'b0 ;
  assign n12046 = x176 & ~n4833 ;
  assign n12047 = n7827 | n12046 ;
  assign n12049 = n12048 ^ n12047 ^ 1'b0 ;
  assign n12050 = ~n7381 & n7506 ;
  assign n12051 = n1722 | n12050 ;
  assign n12052 = ( n1229 & n3211 ) | ( n1229 & n7715 ) | ( n3211 & n7715 ) ;
  assign n12053 = ~n11506 & n12052 ;
  assign n12054 = n661 & ~n7147 ;
  assign n12055 = n12054 ^ n2255 ^ 1'b0 ;
  assign n12056 = ~n1197 & n3029 ;
  assign n12057 = n1775 & n12056 ;
  assign n12058 = n12057 ^ n8657 ^ 1'b0 ;
  assign n12059 = n12055 & n12058 ;
  assign n12060 = x123 | n441 ;
  assign n12061 = n12060 ^ n9681 ^ n4008 ;
  assign n12062 = ~n2610 & n3475 ;
  assign n12063 = n12062 ^ n1711 ^ 1'b0 ;
  assign n12064 = n12061 | n12063 ;
  assign n12065 = n8682 ^ n6310 ^ n2289 ;
  assign n12066 = n3775 & n7215 ;
  assign n12067 = n1996 | n2658 ;
  assign n12068 = n12067 ^ n5801 ^ 1'b0 ;
  assign n12069 = n6236 | n12068 ;
  assign n12070 = n3581 & ~n12069 ;
  assign n12071 = n2736 ^ n1755 ^ 1'b0 ;
  assign n12072 = ( ~n12066 & n12070 ) | ( ~n12066 & n12071 ) | ( n12070 & n12071 ) ;
  assign n12073 = ~n9877 & n12072 ;
  assign n12074 = n12073 ^ n5855 ^ 1'b0 ;
  assign n12075 = n5458 & ~n12074 ;
  assign n12076 = n3406 & n12075 ;
  assign n12077 = n5844 ^ n1563 ^ n381 ;
  assign n12078 = n4379 ^ n978 ^ 1'b0 ;
  assign n12079 = ( n3217 & n10108 ) | ( n3217 & n12078 ) | ( n10108 & n12078 ) ;
  assign n12080 = ( n10667 & ~n11032 ) | ( n10667 & n12079 ) | ( ~n11032 & n12079 ) ;
  assign n12081 = ( ~n8675 & n12077 ) | ( ~n8675 & n12080 ) | ( n12077 & n12080 ) ;
  assign n12082 = x35 & n12081 ;
  assign n12083 = n1596 | n3068 ;
  assign n12084 = n12083 ^ n3338 ^ 1'b0 ;
  assign n12085 = n9086 & n12084 ;
  assign n12086 = ~n2120 & n12085 ;
  assign n12087 = n12086 ^ n5978 ^ x203 ;
  assign n12090 = n3145 & n5975 ;
  assign n12088 = x74 & ~n7242 ;
  assign n12089 = n2759 & n12088 ;
  assign n12091 = n12090 ^ n12089 ^ n3180 ;
  assign n12092 = ( n3184 & n4063 ) | ( n3184 & ~n10620 ) | ( n4063 & ~n10620 ) ;
  assign n12093 = n6796 ^ n5004 ^ 1'b0 ;
  assign n12094 = n7321 | n12093 ;
  assign n12095 = n12094 ^ n9803 ^ 1'b0 ;
  assign n12096 = n12092 & n12095 ;
  assign n12097 = n12096 ^ n10906 ^ 1'b0 ;
  assign n12098 = n9884 ^ n4600 ^ n2777 ;
  assign n12099 = n7321 | n12098 ;
  assign n12100 = ~n6565 & n12099 ;
  assign n12101 = n3743 & n5307 ;
  assign n12102 = n12101 ^ n9366 ^ 1'b0 ;
  assign n12103 = n5156 & n12102 ;
  assign n12104 = n2261 & n12103 ;
  assign n12105 = x2 & ~n4285 ;
  assign n12106 = ( n3100 & ~n3719 ) | ( n3100 & n5937 ) | ( ~n3719 & n5937 ) ;
  assign n12107 = n12105 & n12106 ;
  assign n12108 = n5805 ^ n2006 ^ 1'b0 ;
  assign n12109 = ~n4343 & n12108 ;
  assign n12110 = ( ~n2426 & n9773 ) | ( ~n2426 & n12109 ) | ( n9773 & n12109 ) ;
  assign n12111 = n1079 & ~n12110 ;
  assign n12112 = n4700 ^ n2957 ^ 1'b0 ;
  assign n12113 = n3453 | n7296 ;
  assign n12114 = ~n737 & n2356 ;
  assign n12119 = n3412 & ~n10739 ;
  assign n12120 = n12119 ^ n6045 ^ 1'b0 ;
  assign n12115 = n7322 ^ n3862 ^ 1'b0 ;
  assign n12116 = n556 & ~n12115 ;
  assign n12117 = n12116 ^ n3389 ^ 1'b0 ;
  assign n12118 = n1482 | n12117 ;
  assign n12121 = n12120 ^ n12118 ^ n11135 ;
  assign n12122 = ( n2526 & n3062 ) | ( n2526 & n8286 ) | ( n3062 & n8286 ) ;
  assign n12123 = ( n5146 & ~n7622 ) | ( n5146 & n12122 ) | ( ~n7622 & n12122 ) ;
  assign n12126 = x218 & ~n6127 ;
  assign n12124 = n8346 ^ n7016 ^ n3578 ;
  assign n12125 = n3237 & ~n12124 ;
  assign n12127 = n12126 ^ n12125 ^ 1'b0 ;
  assign n12130 = ( ~n7621 & n8217 ) | ( ~n7621 & n8908 ) | ( n8217 & n8908 ) ;
  assign n12128 = n10978 ^ n6138 ^ 1'b0 ;
  assign n12129 = n6888 & ~n12128 ;
  assign n12131 = n12130 ^ n12129 ^ 1'b0 ;
  assign n12132 = n6626 ^ n5657 ^ 1'b0 ;
  assign n12133 = ~n3726 & n12132 ;
  assign n12134 = n1600 | n5705 ;
  assign n12135 = n12134 ^ n8202 ^ 1'b0 ;
  assign n12136 = n12133 & n12135 ;
  assign n12137 = n12136 ^ n2680 ^ n1145 ;
  assign n12138 = ( x44 & ~x152 ) | ( x44 & n1213 ) | ( ~x152 & n1213 ) ;
  assign n12139 = n12138 ^ n6791 ^ 1'b0 ;
  assign n12140 = ~n682 & n6361 ;
  assign n12141 = n12140 ^ n8404 ^ 1'b0 ;
  assign n12142 = n625 & ~n12141 ;
  assign n12143 = ~n8616 & n12142 ;
  assign n12144 = n12139 & n12143 ;
  assign n12145 = n9385 ^ n5314 ^ 1'b0 ;
  assign n12146 = n8140 ^ n1820 ^ 1'b0 ;
  assign n12147 = ~n544 & n12146 ;
  assign n12148 = n9823 & n12147 ;
  assign n12149 = ~n12145 & n12148 ;
  assign n12150 = n1496 & ~n8878 ;
  assign n12151 = n12150 ^ n2192 ^ 1'b0 ;
  assign n12152 = n3619 ^ n1665 ^ n1423 ;
  assign n12153 = n2257 & ~n4016 ;
  assign n12154 = n1773 & ~n7831 ;
  assign n12155 = n12154 ^ n3095 ^ 1'b0 ;
  assign n12156 = n1698 & n5967 ;
  assign n12157 = n12156 ^ n11723 ^ n10055 ;
  assign n12158 = ( n12153 & n12155 ) | ( n12153 & ~n12157 ) | ( n12155 & ~n12157 ) ;
  assign n12159 = n12158 ^ n4007 ^ n2827 ;
  assign n12160 = n5057 ^ n2015 ^ n1320 ;
  assign n12161 = ~n9296 & n12160 ;
  assign n12162 = n12161 ^ n436 ^ 1'b0 ;
  assign n12163 = x68 & ~n12027 ;
  assign n12164 = n12163 ^ x240 ^ 1'b0 ;
  assign n12165 = ( n4725 & n12162 ) | ( n4725 & ~n12164 ) | ( n12162 & ~n12164 ) ;
  assign n12166 = n12165 ^ n4824 ^ 1'b0 ;
  assign n12167 = n12159 & n12166 ;
  assign n12168 = n8191 ^ n1327 ^ 1'b0 ;
  assign n12169 = n8965 & n11202 ;
  assign n12170 = n2574 | n7434 ;
  assign n12171 = n12170 ^ n11749 ^ 1'b0 ;
  assign n12172 = ( n2086 & n2790 ) | ( n2086 & ~n10355 ) | ( n2790 & ~n10355 ) ;
  assign n12177 = n9863 ^ n8171 ^ n3402 ;
  assign n12178 = n3044 & n9177 ;
  assign n12179 = ~n1451 & n12178 ;
  assign n12180 = ( n2105 & ~n12177 ) | ( n2105 & n12179 ) | ( ~n12177 & n12179 ) ;
  assign n12173 = n4039 | n7774 ;
  assign n12174 = n4648 & ~n12173 ;
  assign n12175 = n11242 ^ n5657 ^ 1'b0 ;
  assign n12176 = n12174 | n12175 ;
  assign n12181 = n12180 ^ n12176 ^ 1'b0 ;
  assign n12182 = n2546 ^ x199 ^ 1'b0 ;
  assign n12183 = n1214 | n12182 ;
  assign n12184 = ( ~n2713 & n4490 ) | ( ~n2713 & n12183 ) | ( n4490 & n12183 ) ;
  assign n12185 = n7004 | n12184 ;
  assign n12186 = n12185 ^ n8716 ^ 1'b0 ;
  assign n12189 = n7784 ^ n7655 ^ n3000 ;
  assign n12187 = x128 & ~n7805 ;
  assign n12188 = n12187 ^ n3853 ^ 1'b0 ;
  assign n12190 = n12189 ^ n12188 ^ n1856 ;
  assign n12191 = ( n3447 & n6602 ) | ( n3447 & ~n7502 ) | ( n6602 & ~n7502 ) ;
  assign n12192 = n5324 & ~n5326 ;
  assign n12193 = n4741 & n12192 ;
  assign n12196 = n5677 ^ n3656 ^ n1098 ;
  assign n12194 = ( ~n835 & n2245 ) | ( ~n835 & n3873 ) | ( n2245 & n3873 ) ;
  assign n12195 = n4898 & n12194 ;
  assign n12197 = n12196 ^ n12195 ^ 1'b0 ;
  assign n12198 = ~n12193 & n12197 ;
  assign n12199 = n8843 | n12198 ;
  assign n12200 = n12199 ^ n10998 ^ 1'b0 ;
  assign n12201 = ( ~n1365 & n5077 ) | ( ~n1365 & n5796 ) | ( n5077 & n5796 ) ;
  assign n12202 = ( ~n2186 & n4899 ) | ( ~n2186 & n12201 ) | ( n4899 & n12201 ) ;
  assign n12205 = x73 & ~n3110 ;
  assign n12206 = n1934 & n12205 ;
  assign n12203 = n9399 ^ n2796 ^ 1'b0 ;
  assign n12204 = n12203 ^ n4072 ^ 1'b0 ;
  assign n12207 = n12206 ^ n12204 ^ n7760 ;
  assign n12208 = n12193 ^ n914 ^ 1'b0 ;
  assign n12209 = n2722 | n12208 ;
  assign n12210 = n9367 | n11152 ;
  assign n12211 = n7983 & n10753 ;
  assign n12212 = n3212 & n12211 ;
  assign n12213 = n2491 | n4485 ;
  assign n12214 = n12213 ^ n802 ^ 1'b0 ;
  assign n12215 = n12212 | n12214 ;
  assign n12216 = n4282 ^ n2042 ^ 1'b0 ;
  assign n12217 = ~n8806 & n12216 ;
  assign n12218 = n12217 ^ n9323 ^ n8399 ;
  assign n12224 = n9608 ^ n3145 ^ 1'b0 ;
  assign n12225 = n10322 & n12224 ;
  assign n12219 = n725 | n10413 ;
  assign n12220 = n10076 ^ n1786 ^ x96 ;
  assign n12221 = n10464 | n12220 ;
  assign n12222 = n12219 & ~n12221 ;
  assign n12223 = n433 & ~n12222 ;
  assign n12226 = n12225 ^ n12223 ^ 1'b0 ;
  assign n12227 = n12226 ^ n6716 ^ 1'b0 ;
  assign n12228 = ( ~n906 & n2189 ) | ( ~n906 & n11570 ) | ( n2189 & n11570 ) ;
  assign n12229 = n389 | n7446 ;
  assign n12230 = n2822 | n12229 ;
  assign n12231 = n3328 | n6879 ;
  assign n12232 = n8993 ^ n6908 ^ 1'b0 ;
  assign n12233 = n12232 ^ n1527 ^ 1'b0 ;
  assign n12238 = n9061 ^ n5741 ^ 1'b0 ;
  assign n12239 = n9958 & ~n12238 ;
  assign n12234 = n3700 ^ n3100 ^ 1'b0 ;
  assign n12235 = ( ~n4983 & n7019 ) | ( ~n4983 & n7638 ) | ( n7019 & n7638 ) ;
  assign n12236 = ( n5937 & n7140 ) | ( n5937 & n12235 ) | ( n7140 & n12235 ) ;
  assign n12237 = n12234 | n12236 ;
  assign n12240 = n12239 ^ n12237 ^ 1'b0 ;
  assign n12241 = ( n1013 & ~n1993 ) | ( n1013 & n2818 ) | ( ~n1993 & n2818 ) ;
  assign n12242 = ~n3383 & n12241 ;
  assign n12243 = n259 | n1341 ;
  assign n12244 = n12243 ^ n6505 ^ n675 ;
  assign n12245 = n6776 & ~n10782 ;
  assign n12246 = n4712 & ~n12245 ;
  assign n12247 = n845 & n3255 ;
  assign n12248 = n11839 & n12247 ;
  assign n12249 = n12248 ^ n3087 ^ 1'b0 ;
  assign n12250 = n10348 ^ n6207 ^ 1'b0 ;
  assign n12251 = n11517 & n11944 ;
  assign n12252 = n6353 | n12067 ;
  assign n12253 = n5265 | n7425 ;
  assign n12254 = x188 & ~n12253 ;
  assign n12255 = ~n12252 & n12254 ;
  assign n12256 = n1452 & ~n2854 ;
  assign n12257 = n3753 | n12256 ;
  assign n12258 = n4747 & ~n12257 ;
  assign n12259 = n8608 ^ n7568 ^ 1'b0 ;
  assign n12260 = n4240 | n12259 ;
  assign n12261 = n10739 | n12260 ;
  assign n12262 = x162 | n9366 ;
  assign n12263 = n5325 & ~n12262 ;
  assign n12264 = n3261 ^ n2882 ^ x250 ;
  assign n12265 = ~n6056 & n8524 ;
  assign n12266 = n12264 & n12265 ;
  assign n12267 = ~n5872 & n12266 ;
  assign n12268 = ( n5530 & ~n12263 ) | ( n5530 & n12267 ) | ( ~n12263 & n12267 ) ;
  assign n12269 = n12147 ^ n7366 ^ 1'b0 ;
  assign n12271 = n6896 ^ n4150 ^ n3858 ;
  assign n12272 = n8411 | n12271 ;
  assign n12270 = n3302 ^ n2191 ^ 1'b0 ;
  assign n12273 = n12272 ^ n12270 ^ n7564 ;
  assign n12274 = n6610 & n9711 ;
  assign n12275 = n9700 ^ n7769 ^ 1'b0 ;
  assign n12276 = n12275 ^ n5942 ^ 1'b0 ;
  assign n12277 = n10877 | n12276 ;
  assign n12278 = n3063 | n12277 ;
  assign n12279 = n12278 ^ n2937 ^ 1'b0 ;
  assign n12280 = ~n7919 & n8556 ;
  assign n12281 = n12279 & n12280 ;
  assign n12282 = ~n9415 & n12281 ;
  assign n12283 = n4633 & ~n11005 ;
  assign n12284 = ( n288 & ~n1211 ) | ( n288 & n1350 ) | ( ~n1211 & n1350 ) ;
  assign n12288 = ( n678 & n4602 ) | ( n678 & ~n6611 ) | ( n4602 & ~n6611 ) ;
  assign n12286 = n7254 ^ n3455 ^ 1'b0 ;
  assign n12287 = ~n11035 & n12286 ;
  assign n12289 = n12288 ^ n12287 ^ n10632 ;
  assign n12285 = ~n2160 & n12068 ;
  assign n12290 = n12289 ^ n12285 ^ n8257 ;
  assign n12291 = ~n3632 & n6832 ;
  assign n12292 = n12291 ^ n11007 ^ 1'b0 ;
  assign n12293 = n1200 & ~n9802 ;
  assign n12294 = ~n9306 & n12293 ;
  assign n12295 = n2323 ^ n530 ^ 1'b0 ;
  assign n12296 = n2736 & n12295 ;
  assign n12297 = n12296 ^ n4512 ^ n3066 ;
  assign n12298 = n2510 & ~n2998 ;
  assign n12299 = x124 & n12298 ;
  assign n12300 = n9139 ^ n7873 ^ n4614 ;
  assign n12301 = ~n4174 & n10495 ;
  assign n12302 = ( n8093 & n9555 ) | ( n8093 & n12301 ) | ( n9555 & n12301 ) ;
  assign n12305 = x22 | n708 ;
  assign n12303 = n6711 | n7885 ;
  assign n12304 = n1249 & ~n12303 ;
  assign n12306 = n12305 ^ n12304 ^ 1'b0 ;
  assign n12307 = n3578 & n7075 ;
  assign n12308 = n8913 & n12307 ;
  assign n12309 = n5264 ^ n3289 ^ 1'b0 ;
  assign n12310 = n12309 ^ x103 ^ 1'b0 ;
  assign n12311 = n8695 & ~n12310 ;
  assign n12312 = n4678 | n4947 ;
  assign n12313 = n12312 ^ n11931 ^ n11245 ;
  assign n12314 = n6200 ^ n4322 ^ 1'b0 ;
  assign n12315 = n2462 & n4801 ;
  assign n12316 = n5098 | n12315 ;
  assign n12317 = n12314 & ~n12316 ;
  assign n12318 = ( n2333 & n3756 ) | ( n2333 & ~n12317 ) | ( n3756 & ~n12317 ) ;
  assign n12319 = n10407 & ~n11949 ;
  assign n12320 = n12319 ^ n6650 ^ 1'b0 ;
  assign n12321 = n6439 ^ n2560 ^ n332 ;
  assign n12322 = n5433 ^ n5049 ^ 1'b0 ;
  assign n12323 = ~n12321 & n12322 ;
  assign n12324 = ~n7308 & n12323 ;
  assign n12325 = n10608 ^ n4439 ^ 1'b0 ;
  assign n12326 = ~n2214 & n12325 ;
  assign n12327 = x224 & ~n7381 ;
  assign n12337 = ~n1410 & n1543 ;
  assign n12338 = n12337 ^ n2846 ^ 1'b0 ;
  assign n12339 = n1550 & ~n3866 ;
  assign n12340 = ~n12338 & n12339 ;
  assign n12336 = n2754 | n4695 ;
  assign n12341 = n12340 ^ n12336 ^ 1'b0 ;
  assign n12342 = n12341 ^ n6445 ^ n4598 ;
  assign n12343 = n12342 ^ n6319 ^ n2339 ;
  assign n12328 = ( n2247 & ~n4520 ) | ( n2247 & n5737 ) | ( ~n4520 & n5737 ) ;
  assign n12329 = n12328 ^ n4084 ^ 1'b0 ;
  assign n12330 = n718 & ~n12329 ;
  assign n12331 = n639 & n12330 ;
  assign n12332 = n426 | n1170 ;
  assign n12333 = n1729 | n12332 ;
  assign n12334 = n481 | n10937 ;
  assign n12335 = ( n12331 & ~n12333 ) | ( n12331 & n12334 ) | ( ~n12333 & n12334 ) ;
  assign n12344 = n12343 ^ n12335 ^ 1'b0 ;
  assign n12345 = n8810 ^ n1453 ^ 1'b0 ;
  assign n12346 = n1572 & n12345 ;
  assign n12348 = n6417 ^ n3472 ^ 1'b0 ;
  assign n12347 = n8100 & ~n9641 ;
  assign n12349 = n12348 ^ n12347 ^ 1'b0 ;
  assign n12350 = n3609 ^ n3336 ^ 1'b0 ;
  assign n12351 = ( ~n6649 & n8281 ) | ( ~n6649 & n12350 ) | ( n8281 & n12350 ) ;
  assign n12352 = n11667 ^ n1983 ^ 1'b0 ;
  assign n12353 = n1254 | n1769 ;
  assign n12354 = n9831 & ~n12353 ;
  assign n12355 = n9692 | n11687 ;
  assign n12356 = n6866 | n12355 ;
  assign n12357 = ( n11055 & n12354 ) | ( n11055 & n12356 ) | ( n12354 & n12356 ) ;
  assign n12358 = n2720 & ~n8932 ;
  assign n12359 = n7124 ^ n5974 ^ n5065 ;
  assign n12360 = ( n2822 & ~n5394 ) | ( n2822 & n12359 ) | ( ~n5394 & n12359 ) ;
  assign n12365 = n4304 & ~n7520 ;
  assign n12362 = n803 ^ n300 ^ 1'b0 ;
  assign n12361 = n8991 ^ n8182 ^ n5376 ;
  assign n12363 = n12362 ^ n12361 ^ 1'b0 ;
  assign n12364 = ~n750 & n12363 ;
  assign n12366 = n12365 ^ n12364 ^ 1'b0 ;
  assign n12367 = n4767 ^ n957 ^ 1'b0 ;
  assign n12368 = n9650 ^ n6447 ^ 1'b0 ;
  assign n12369 = n2551 ^ n1265 ^ 1'b0 ;
  assign n12370 = n3200 & n11334 ;
  assign n12371 = n1994 | n4672 ;
  assign n12372 = n12371 ^ n4881 ^ 1'b0 ;
  assign n12373 = n3064 | n7333 ;
  assign n12374 = n10205 ^ n4539 ^ 1'b0 ;
  assign n12375 = n12374 ^ n2966 ^ 1'b0 ;
  assign n12376 = n12373 | n12375 ;
  assign n12377 = n3891 | n12376 ;
  assign n12378 = ( n2133 & ~n7001 ) | ( n2133 & n8718 ) | ( ~n7001 & n8718 ) ;
  assign n12379 = n11431 | n12378 ;
  assign n12380 = n12379 ^ n8986 ^ 1'b0 ;
  assign n12381 = n6048 ^ n1064 ^ 1'b0 ;
  assign n12382 = n10034 | n12381 ;
  assign n12383 = n7415 ^ n5189 ^ 1'b0 ;
  assign n12384 = n6200 & ~n12383 ;
  assign n12385 = ( ~n1254 & n2584 ) | ( ~n1254 & n12384 ) | ( n2584 & n12384 ) ;
  assign n12386 = ~n4244 & n12385 ;
  assign n12387 = n12386 ^ n6216 ^ 1'b0 ;
  assign n12388 = n12382 | n12387 ;
  assign n12389 = n2871 & n7554 ;
  assign n12390 = n6355 | n6510 ;
  assign n12391 = n9419 ^ n3447 ^ n2754 ;
  assign n12392 = n660 | n9875 ;
  assign n12393 = n2171 | n12392 ;
  assign n12394 = n8502 | n12393 ;
  assign n12395 = n12394 ^ n5796 ^ n4756 ;
  assign n12396 = n4840 & ~n8128 ;
  assign n12397 = n4973 ^ n2123 ^ n1611 ;
  assign n12398 = n12397 ^ n9103 ^ 1'b0 ;
  assign n12399 = n12398 ^ n6149 ^ 1'b0 ;
  assign n12400 = ~n976 & n12399 ;
  assign n12401 = n305 | n8898 ;
  assign n12402 = ( n1914 & n3081 ) | ( n1914 & ~n12401 ) | ( n3081 & ~n12401 ) ;
  assign n12403 = n3512 & n4367 ;
  assign n12404 = n12403 ^ n3316 ^ 1'b0 ;
  assign n12405 = ( ~x143 & n5045 ) | ( ~x143 & n12404 ) | ( n5045 & n12404 ) ;
  assign n12406 = n1366 & ~n2721 ;
  assign n12407 = n6788 & n12406 ;
  assign n12408 = n834 | n6913 ;
  assign n12409 = n11087 & ~n11379 ;
  assign n12410 = n12409 ^ n5393 ^ 1'b0 ;
  assign n12411 = ( n12407 & n12408 ) | ( n12407 & n12410 ) | ( n12408 & n12410 ) ;
  assign n12412 = n9346 ^ n672 ^ 1'b0 ;
  assign n12413 = n12412 ^ n4672 ^ n4350 ;
  assign n12414 = n5751 & n6536 ;
  assign n12415 = n2042 & n12414 ;
  assign n12416 = n8083 | n12415 ;
  assign n12417 = ( ~n8755 & n12413 ) | ( ~n8755 & n12416 ) | ( n12413 & n12416 ) ;
  assign n12418 = n2924 ^ n729 ^ x226 ;
  assign n12419 = n5602 | n12418 ;
  assign n12420 = n6531 ^ n6509 ^ 1'b0 ;
  assign n12423 = ~n1549 & n3378 ;
  assign n12424 = n3425 ^ n1542 ^ 1'b0 ;
  assign n12425 = n5391 & ~n12424 ;
  assign n12426 = n2311 & n12425 ;
  assign n12427 = ~n6516 & n12426 ;
  assign n12428 = n12427 ^ n7676 ^ 1'b0 ;
  assign n12429 = ~n12423 & n12428 ;
  assign n12421 = n4518 ^ x131 ^ 1'b0 ;
  assign n12422 = n6015 | n12421 ;
  assign n12430 = n12429 ^ n12422 ^ n1053 ;
  assign n12431 = n1222 & n1741 ;
  assign n12432 = x187 ^ x41 ^ 1'b0 ;
  assign n12433 = ~n12431 & n12432 ;
  assign n12434 = n6589 ^ n358 ^ 1'b0 ;
  assign n12435 = ( n741 & n3691 ) | ( n741 & ~n5929 ) | ( n3691 & ~n5929 ) ;
  assign n12436 = n10443 ^ n5381 ^ 1'b0 ;
  assign n12437 = n1605 & n12436 ;
  assign n12438 = n12435 & n12437 ;
  assign n12439 = n6868 ^ n4570 ^ n2073 ;
  assign n12440 = n12439 ^ n2678 ^ 1'b0 ;
  assign n12441 = n12142 & ~n12440 ;
  assign n12442 = n12441 ^ n9552 ^ 1'b0 ;
  assign n12457 = n4343 ^ n2611 ^ 1'b0 ;
  assign n12458 = n10780 | n12457 ;
  assign n12459 = n12458 ^ n978 ^ 1'b0 ;
  assign n12443 = ( n329 & ~n1201 ) | ( n329 & n10503 ) | ( ~n1201 & n10503 ) ;
  assign n12446 = n1283 & ~n5588 ;
  assign n12447 = ~n1243 & n12446 ;
  assign n12444 = ~n2199 & n6487 ;
  assign n12445 = n12444 ^ n3047 ^ 1'b0 ;
  assign n12448 = n12447 ^ n12445 ^ 1'b0 ;
  assign n12449 = n12443 & ~n12448 ;
  assign n12450 = n12449 ^ n1666 ^ 1'b0 ;
  assign n12451 = n982 & n12450 ;
  assign n12452 = n1413 & n5359 ;
  assign n12453 = n12452 ^ n7549 ^ 1'b0 ;
  assign n12454 = ( n7625 & ~n8354 ) | ( n7625 & n12453 ) | ( ~n8354 & n12453 ) ;
  assign n12455 = n7883 & ~n12454 ;
  assign n12456 = n12451 & n12455 ;
  assign n12460 = n12459 ^ n12456 ^ 1'b0 ;
  assign n12461 = n1229 | n1409 ;
  assign n12462 = n10089 ^ n7353 ^ n3368 ;
  assign n12465 = n603 & n7586 ;
  assign n12466 = n12465 ^ x206 ^ 1'b0 ;
  assign n12463 = n4875 ^ n4154 ^ n2915 ;
  assign n12464 = n12463 ^ n5114 ^ n2966 ;
  assign n12467 = n12466 ^ n12464 ^ 1'b0 ;
  assign n12468 = n12467 ^ n8891 ^ 1'b0 ;
  assign n12469 = n332 | n12468 ;
  assign n12470 = ( n8222 & n12462 ) | ( n8222 & n12469 ) | ( n12462 & n12469 ) ;
  assign n12471 = n2268 & n7549 ;
  assign n12472 = n9653 ^ n5795 ^ 1'b0 ;
  assign n12473 = ( n3046 & n8307 ) | ( n3046 & n11741 ) | ( n8307 & n11741 ) ;
  assign n12476 = ( n1791 & n4472 ) | ( n1791 & ~n6381 ) | ( n4472 & ~n6381 ) ;
  assign n12474 = n10387 ^ n8483 ^ n4924 ;
  assign n12475 = ~n4176 & n12474 ;
  assign n12477 = n12476 ^ n12475 ^ 1'b0 ;
  assign n12478 = n12477 ^ n1164 ^ 1'b0 ;
  assign n12479 = n4875 & n5486 ;
  assign n12480 = n1156 & ~n3557 ;
  assign n12481 = x150 | n10757 ;
  assign n12482 = x87 & n12481 ;
  assign n12483 = n10170 ^ n1386 ^ 1'b0 ;
  assign n12484 = n4912 ^ n4164 ^ 1'b0 ;
  assign n12485 = ~n530 & n12484 ;
  assign n12486 = n9831 ^ n4689 ^ 1'b0 ;
  assign n12487 = ( ~n4350 & n4536 ) | ( ~n4350 & n12486 ) | ( n4536 & n12486 ) ;
  assign n12488 = ( ~n2662 & n12485 ) | ( ~n2662 & n12487 ) | ( n12485 & n12487 ) ;
  assign n12489 = x211 & ~n2354 ;
  assign n12490 = n12489 ^ n2159 ^ 1'b0 ;
  assign n12491 = n10230 | n12490 ;
  assign n12493 = n10201 ^ n2820 ^ n802 ;
  assign n12492 = ( n1010 & n2106 ) | ( n1010 & ~n6839 ) | ( n2106 & ~n6839 ) ;
  assign n12494 = n12493 ^ n12492 ^ 1'b0 ;
  assign n12495 = n11461 | n12494 ;
  assign n12496 = n12495 ^ n9902 ^ 1'b0 ;
  assign n12497 = n789 & ~n12496 ;
  assign n12502 = x219 & ~n1452 ;
  assign n12501 = x242 & n2619 ;
  assign n12503 = n12502 ^ n12501 ^ 1'b0 ;
  assign n12504 = n12503 ^ n1039 ^ 1'b0 ;
  assign n12498 = n1447 ^ n902 ^ x113 ;
  assign n12499 = ( n2838 & n10914 ) | ( n2838 & ~n12498 ) | ( n10914 & ~n12498 ) ;
  assign n12500 = n12499 ^ n2543 ^ 1'b0 ;
  assign n12505 = n12504 ^ n12500 ^ 1'b0 ;
  assign n12506 = n8372 ^ n5948 ^ n4767 ;
  assign n12507 = n12506 ^ n3170 ^ 1'b0 ;
  assign n12508 = n5865 | n12507 ;
  assign n12509 = n8122 ^ n3360 ^ 1'b0 ;
  assign n12510 = x242 & n12509 ;
  assign n12511 = ( n2007 & n2568 ) | ( n2007 & ~n7923 ) | ( n2568 & ~n7923 ) ;
  assign n12512 = n12510 & ~n12511 ;
  assign n12513 = n5646 ^ n1823 ^ 1'b0 ;
  assign n12514 = n9430 ^ n4263 ^ 1'b0 ;
  assign n12515 = n12514 ^ n256 ^ 1'b0 ;
  assign n12516 = n8883 ^ n2022 ^ 1'b0 ;
  assign n12523 = n10547 ^ n3208 ^ 1'b0 ;
  assign n12524 = n6032 | n12523 ;
  assign n12525 = n1040 | n12524 ;
  assign n12526 = n12525 ^ n3690 ^ n3083 ;
  assign n12521 = n8908 ^ n2645 ^ n1711 ;
  assign n12518 = ~n8030 & n9048 ;
  assign n12519 = n12518 ^ n5412 ^ 1'b0 ;
  assign n12517 = n2121 & n6251 ;
  assign n12520 = n12519 ^ n12517 ^ 1'b0 ;
  assign n12522 = n12521 ^ n12520 ^ n323 ;
  assign n12527 = n12526 ^ n12522 ^ 1'b0 ;
  assign n12528 = n1603 & ~n5045 ;
  assign n12529 = n4865 & ~n12528 ;
  assign n12530 = ( n332 & n7957 ) | ( n332 & n12529 ) | ( n7957 & n12529 ) ;
  assign n12531 = ~n7831 & n10888 ;
  assign n12532 = n12531 ^ n6592 ^ 1'b0 ;
  assign n12533 = n11893 ^ n9997 ^ n5379 ;
  assign n12534 = n399 & ~n1999 ;
  assign n12535 = n3016 ^ x208 ^ 1'b0 ;
  assign n12536 = ~n2701 & n12535 ;
  assign n12537 = ~n5525 & n12536 ;
  assign n12538 = n12537 ^ n5039 ^ 1'b0 ;
  assign n12539 = n2995 ^ n807 ^ 1'b0 ;
  assign n12540 = n2606 ^ x169 ^ 1'b0 ;
  assign n12541 = n12540 ^ n287 ^ 1'b0 ;
  assign n12542 = n621 & n1243 ;
  assign n12543 = n12542 ^ n5095 ^ n2566 ;
  assign n12544 = n12543 ^ n3208 ^ 1'b0 ;
  assign n12545 = n9749 & n12544 ;
  assign n12546 = n12545 ^ n5781 ^ 1'b0 ;
  assign n12547 = n7404 ^ n7132 ^ n3523 ;
  assign n12548 = n12547 ^ n5584 ^ n2770 ;
  assign n12549 = n5146 & ~n12548 ;
  assign n12550 = ( n3095 & n4448 ) | ( n3095 & n5797 ) | ( n4448 & n5797 ) ;
  assign n12551 = ~n401 & n1284 ;
  assign n12552 = n12550 & n12551 ;
  assign n12553 = ( n853 & n1795 ) | ( n853 & n6574 ) | ( n1795 & n6574 ) ;
  assign n12554 = ( n1807 & ~n4978 ) | ( n1807 & n12553 ) | ( ~n4978 & n12553 ) ;
  assign n12555 = n1327 & ~n5502 ;
  assign n12556 = n1420 & n12555 ;
  assign n12557 = n12556 ^ n2047 ^ 1'b0 ;
  assign n12558 = ~n12554 & n12557 ;
  assign n12559 = ~n7753 & n9201 ;
  assign n12560 = n1324 & ~n3891 ;
  assign n12561 = n12560 ^ n8900 ^ 1'b0 ;
  assign n12562 = ( n1455 & n9961 ) | ( n1455 & n10216 ) | ( n9961 & n10216 ) ;
  assign n12563 = n11455 ^ n9198 ^ 1'b0 ;
  assign n12564 = n2268 & ~n12563 ;
  assign n12565 = n11188 ^ n6807 ^ 1'b0 ;
  assign n12573 = n4874 ^ x175 ^ 1'b0 ;
  assign n12574 = n4615 & n12573 ;
  assign n12575 = n12574 ^ n2991 ^ 1'b0 ;
  assign n12566 = ( ~n777 & n3853 ) | ( ~n777 & n3878 ) | ( n3853 & n3878 ) ;
  assign n12567 = n7758 ^ n7741 ^ n6831 ;
  assign n12568 = n12566 & n12567 ;
  assign n12569 = n4330 & n12568 ;
  assign n12570 = n747 & n12569 ;
  assign n12571 = n6828 & n12570 ;
  assign n12572 = ~n3314 & n12571 ;
  assign n12576 = n12575 ^ n12572 ^ 1'b0 ;
  assign n12577 = n7616 ^ x139 ^ 1'b0 ;
  assign n12578 = n2150 & ~n12577 ;
  assign n12579 = n3966 & n12578 ;
  assign n12580 = x109 & ~n2742 ;
  assign n12581 = n9045 & n12580 ;
  assign n12582 = ( x2 & ~n12579 ) | ( x2 & n12581 ) | ( ~n12579 & n12581 ) ;
  assign n12583 = n6371 ^ n727 ^ 1'b0 ;
  assign n12584 = n6744 & n12583 ;
  assign n12586 = n507 | n11580 ;
  assign n12587 = n2070 & ~n12586 ;
  assign n12588 = n589 & ~n7262 ;
  assign n12589 = n12588 ^ n1328 ^ 1'b0 ;
  assign n12590 = n4282 ^ n2092 ^ 1'b0 ;
  assign n12591 = ~n2900 & n12590 ;
  assign n12592 = ( n2116 & ~n12589 ) | ( n2116 & n12591 ) | ( ~n12589 & n12591 ) ;
  assign n12593 = n12592 ^ x246 ^ 1'b0 ;
  assign n12594 = ( n5485 & n12587 ) | ( n5485 & ~n12593 ) | ( n12587 & ~n12593 ) ;
  assign n12585 = n12271 ^ n7677 ^ n6948 ;
  assign n12595 = n12594 ^ n12585 ^ n10973 ;
  assign n12596 = n334 | n2471 ;
  assign n12597 = n2484 & ~n12596 ;
  assign n12598 = n1512 & ~n4740 ;
  assign n12599 = n10771 & n12598 ;
  assign n12600 = n12597 & n12599 ;
  assign n12601 = ( n932 & ~n1741 ) | ( n932 & n7551 ) | ( ~n1741 & n7551 ) ;
  assign n12602 = n4274 ^ n3766 ^ 1'b0 ;
  assign n12603 = ~n12079 & n12602 ;
  assign n12604 = n2804 & n12603 ;
  assign n12605 = n6634 & ~n9899 ;
  assign n12606 = n12605 ^ n12190 ^ 1'b0 ;
  assign n12607 = ( n2786 & n3366 ) | ( n2786 & n12004 ) | ( n3366 & n12004 ) ;
  assign n12608 = ~n7290 & n11420 ;
  assign n12609 = n10306 & n12608 ;
  assign n12610 = n8128 ^ n7758 ^ 1'b0 ;
  assign n12614 = n2962 ^ n2099 ^ 1'b0 ;
  assign n12615 = n12614 ^ n11874 ^ n7439 ;
  assign n12611 = n5506 ^ n4448 ^ 1'b0 ;
  assign n12612 = n10202 & n12611 ;
  assign n12613 = n12612 ^ n1116 ^ 1'b0 ;
  assign n12616 = n12615 ^ n12613 ^ 1'b0 ;
  assign n12617 = n12616 ^ n9507 ^ 1'b0 ;
  assign n12618 = n1827 | n3617 ;
  assign n12619 = n6910 & ~n12618 ;
  assign n12620 = n1959 | n12619 ;
  assign n12621 = n12620 ^ n4340 ^ 1'b0 ;
  assign n12622 = n8416 ^ n1766 ^ 1'b0 ;
  assign n12623 = ~n10525 & n12622 ;
  assign n12624 = n12621 & n12623 ;
  assign n12625 = n5023 ^ n697 ^ 1'b0 ;
  assign n12626 = n2334 & n12625 ;
  assign n12627 = ( n804 & ~n4823 ) | ( n804 & n12626 ) | ( ~n4823 & n12626 ) ;
  assign n12628 = n12374 ^ n9792 ^ 1'b0 ;
  assign n12629 = ~n12627 & n12628 ;
  assign n12630 = n6425 | n9777 ;
  assign n12631 = n12630 ^ n10456 ^ n326 ;
  assign n12632 = n12078 ^ n667 ^ 1'b0 ;
  assign n12633 = n5412 & n12632 ;
  assign n12634 = n3721 & n7680 ;
  assign n12635 = ( n3823 & n5099 ) | ( n3823 & ~n12634 ) | ( n5099 & ~n12634 ) ;
  assign n12636 = ( n1220 & n1462 ) | ( n1220 & ~n12635 ) | ( n1462 & ~n12635 ) ;
  assign n12637 = n6828 ^ n3732 ^ 1'b0 ;
  assign n12638 = n12636 & ~n12637 ;
  assign n12639 = n1462 & ~n8116 ;
  assign n12640 = n1653 & n12639 ;
  assign n12641 = n5288 & n9738 ;
  assign n12642 = ~n7130 & n12641 ;
  assign n12643 = n1262 & n1444 ;
  assign n12644 = ~x33 & n12643 ;
  assign n12645 = n5317 & n12644 ;
  assign n12646 = ( n3630 & n7785 ) | ( n3630 & n12645 ) | ( n7785 & n12645 ) ;
  assign n12647 = ~n5627 & n11187 ;
  assign n12648 = ~n4970 & n12647 ;
  assign n12649 = ( n6394 & ~n6845 ) | ( n6394 & n12648 ) | ( ~n6845 & n12648 ) ;
  assign n12650 = ( n2980 & n6242 ) | ( n2980 & n12649 ) | ( n6242 & n12649 ) ;
  assign n12651 = n12650 ^ n9077 ^ 1'b0 ;
  assign n12653 = n9780 ^ n8332 ^ 1'b0 ;
  assign n12652 = n4791 | n5868 ;
  assign n12654 = n12653 ^ n12652 ^ 1'b0 ;
  assign n12655 = ( n2662 & n4276 ) | ( n2662 & ~n6795 ) | ( n4276 & ~n6795 ) ;
  assign n12656 = n12655 ^ n7366 ^ n5056 ;
  assign n12657 = ( x72 & ~n3242 ) | ( x72 & n5307 ) | ( ~n3242 & n5307 ) ;
  assign n12658 = ~n8979 & n12657 ;
  assign n12659 = ~n12656 & n12658 ;
  assign n12660 = n12090 ^ n7230 ^ 1'b0 ;
  assign n12661 = ~n1852 & n12660 ;
  assign n12662 = n12661 ^ n9761 ^ n7353 ;
  assign n12663 = n603 & ~n2733 ;
  assign n12664 = n2990 & ~n12663 ;
  assign n12671 = n10421 ^ x150 ^ 1'b0 ;
  assign n12665 = ~n777 & n5025 ;
  assign n12666 = n5521 & n12665 ;
  assign n12667 = n12666 ^ n1141 ^ 1'b0 ;
  assign n12668 = ( n1226 & ~n1718 ) | ( n1226 & n12667 ) | ( ~n1718 & n12667 ) ;
  assign n12669 = n12668 ^ n8951 ^ 1'b0 ;
  assign n12670 = ~n949 & n12669 ;
  assign n12672 = n12671 ^ n12670 ^ 1'b0 ;
  assign n12673 = n12672 ^ n11243 ^ 1'b0 ;
  assign n12674 = n2919 & ~n5198 ;
  assign n12675 = n1484 & n12674 ;
  assign n12676 = n11406 ^ n7361 ^ 1'b0 ;
  assign n12677 = ( n1164 & ~n10429 ) | ( n1164 & n11221 ) | ( ~n10429 & n11221 ) ;
  assign n12678 = n7621 ^ x166 ^ 1'b0 ;
  assign n12679 = n12677 & n12678 ;
  assign n12680 = n4283 & n8508 ;
  assign n12681 = n12680 ^ n6473 ^ 1'b0 ;
  assign n12682 = n6164 & ~n9568 ;
  assign n12683 = n774 & n4363 ;
  assign n12684 = ~n5834 & n12683 ;
  assign n12685 = ~n3454 & n5854 ;
  assign n12686 = ~n8893 & n12685 ;
  assign n12687 = n12686 ^ n512 ^ 1'b0 ;
  assign n12688 = n1766 & ~n12687 ;
  assign n12689 = x59 & n12688 ;
  assign n12690 = n859 | n4909 ;
  assign n12691 = n7746 ^ n3096 ^ 1'b0 ;
  assign n12692 = n12691 ^ n1497 ^ 1'b0 ;
  assign n12693 = n5153 & ~n12692 ;
  assign n12694 = ~n4292 & n7248 ;
  assign n12695 = n987 & n12694 ;
  assign n12696 = n12695 ^ n1727 ^ 1'b0 ;
  assign n12697 = n3336 & ~n3793 ;
  assign n12698 = ~n6765 & n12697 ;
  assign n12699 = n4579 ^ n365 ^ 1'b0 ;
  assign n12700 = n8821 | n12699 ;
  assign n12701 = n8836 | n12700 ;
  assign n12702 = n12701 ^ n8137 ^ n2980 ;
  assign n12703 = ( n6672 & n12698 ) | ( n6672 & n12702 ) | ( n12698 & n12702 ) ;
  assign n12704 = n11169 ^ n4851 ^ 1'b0 ;
  assign n12705 = ~n6587 & n10365 ;
  assign n12706 = n12705 ^ n11128 ^ 1'b0 ;
  assign n12707 = n12506 ^ n9525 ^ 1'b0 ;
  assign n12708 = ~n11152 & n12483 ;
  assign n12709 = n5548 & ~n5925 ;
  assign n12710 = n10568 & ~n12709 ;
  assign n12711 = n6228 & ~n9043 ;
  assign n12712 = n12711 ^ n5486 ^ 1'b0 ;
  assign n12713 = n12710 & n12712 ;
  assign n12715 = n702 & n848 ;
  assign n12716 = n12715 ^ n4827 ^ 1'b0 ;
  assign n12714 = ( n1403 & n6103 ) | ( n1403 & ~n7894 ) | ( n6103 & ~n7894 ) ;
  assign n12717 = n12716 ^ n12714 ^ n5797 ;
  assign n12718 = n9529 ^ n8179 ^ 1'b0 ;
  assign n12719 = n2557 | n12718 ;
  assign n12720 = n12719 ^ n7715 ^ 1'b0 ;
  assign n12721 = n12720 ^ n1068 ^ 1'b0 ;
  assign n12722 = n2915 & ~n8272 ;
  assign n12723 = ~n589 & n12722 ;
  assign n12724 = n5301 & ~n12723 ;
  assign n12725 = n11430 ^ n814 ^ 1'b0 ;
  assign n12726 = n2939 & ~n12725 ;
  assign n12727 = n12726 ^ n7980 ^ 1'b0 ;
  assign n12728 = n3237 & ~n12727 ;
  assign n12729 = n8540 ^ n6102 ^ 1'b0 ;
  assign n12730 = ~n3075 & n12729 ;
  assign n12731 = n12730 ^ n11863 ^ n4723 ;
  assign n12733 = n2107 | n3422 ;
  assign n12732 = n4157 & n4304 ;
  assign n12734 = n12733 ^ n12732 ^ 1'b0 ;
  assign n12735 = ( ~n817 & n4490 ) | ( ~n817 & n6240 ) | ( n4490 & n6240 ) ;
  assign n12736 = n12491 ^ n8993 ^ 1'b0 ;
  assign n12737 = n5023 ^ n1176 ^ 1'b0 ;
  assign n12738 = n2683 & n12737 ;
  assign n12739 = ~n1922 & n12738 ;
  assign n12740 = n12739 ^ n7591 ^ 1'b0 ;
  assign n12741 = n6228 ^ n1030 ^ 1'b0 ;
  assign n12742 = n5821 & ~n12741 ;
  assign n12743 = n5725 ^ n4807 ^ n3416 ;
  assign n12744 = n11723 ^ n1321 ^ n472 ;
  assign n12745 = ~n12743 & n12744 ;
  assign n12746 = n1806 & n12745 ;
  assign n12747 = n12746 ^ x200 ^ 1'b0 ;
  assign n12748 = n8281 & ~n12747 ;
  assign n12749 = n2125 | n8667 ;
  assign n12750 = n6795 & n12749 ;
  assign n12751 = ~n1197 & n7697 ;
  assign n12752 = n12751 ^ n1746 ^ 1'b0 ;
  assign n12753 = ( n5148 & n10140 ) | ( n5148 & ~n12752 ) | ( n10140 & ~n12752 ) ;
  assign n12754 = ( n3724 & ~n4840 ) | ( n3724 & n12753 ) | ( ~n4840 & n12753 ) ;
  assign n12755 = n7298 | n12754 ;
  assign n12756 = n12750 | n12755 ;
  assign n12757 = n3309 & n6430 ;
  assign n12758 = n2490 & ~n5702 ;
  assign n12761 = n6302 ^ n2516 ^ x158 ;
  assign n12759 = n1060 ^ n275 ^ 1'b0 ;
  assign n12760 = n12759 ^ n6897 ^ 1'b0 ;
  assign n12762 = n12761 ^ n12760 ^ n4130 ;
  assign n12763 = n6236 | n12762 ;
  assign n12764 = n5706 | n12763 ;
  assign n12765 = n12764 ^ n3768 ^ 1'b0 ;
  assign n12766 = n9566 & n12765 ;
  assign n12767 = n8500 ^ n1463 ^ 1'b0 ;
  assign n12768 = ~n1096 & n12767 ;
  assign n12769 = n12768 ^ n7071 ^ n6316 ;
  assign n12770 = n12521 ^ n3085 ^ 1'b0 ;
  assign n12771 = n7512 | n12770 ;
  assign n12772 = n7859 ^ n6742 ^ n5797 ;
  assign n12773 = n2938 & n12772 ;
  assign n12774 = n12773 ^ n1064 ^ 1'b0 ;
  assign n12775 = n6399 & ~n12774 ;
  assign n12779 = n2259 & n6320 ;
  assign n12776 = n616 | n1309 ;
  assign n12777 = n4245 & n12776 ;
  assign n12778 = n12777 ^ n3894 ^ 1'b0 ;
  assign n12780 = n12779 ^ n12778 ^ 1'b0 ;
  assign n12781 = n3068 | n12780 ;
  assign n12782 = n9712 & ~n11925 ;
  assign n12783 = x132 & ~n2201 ;
  assign n12784 = n1110 | n12783 ;
  assign n12785 = n7189 & ~n12784 ;
  assign n12786 = n7232 ^ n4544 ^ 1'b0 ;
  assign n12787 = n8083 & ~n12786 ;
  assign n12788 = n12615 | n12787 ;
  assign n12789 = n1402 | n11895 ;
  assign n12790 = n12789 ^ n6942 ^ 1'b0 ;
  assign n12791 = n8202 ^ n718 ^ 1'b0 ;
  assign n12792 = n1755 | n12791 ;
  assign n12793 = n2498 & ~n12792 ;
  assign n12794 = n12793 ^ n2441 ^ 1'b0 ;
  assign n12795 = n7099 & n12794 ;
  assign n12796 = n12795 ^ n10744 ^ 1'b0 ;
  assign n12797 = n11007 ^ n10348 ^ n8753 ;
  assign n12798 = n2992 | n7952 ;
  assign n12799 = n2822 & ~n12798 ;
  assign n12800 = n2056 & n3370 ;
  assign n12801 = n4313 & n9398 ;
  assign n12807 = n5263 ^ n711 ^ 1'b0 ;
  assign n12808 = ~n6904 & n12807 ;
  assign n12804 = n3439 ^ n898 ^ 1'b0 ;
  assign n12802 = ~n5326 & n6930 ;
  assign n12803 = n5302 & n12802 ;
  assign n12805 = n12804 ^ n12803 ^ n6278 ;
  assign n12806 = n738 & n12805 ;
  assign n12809 = n12808 ^ n12806 ^ 1'b0 ;
  assign n12810 = n257 & ~n11180 ;
  assign n12811 = ( n931 & n2468 ) | ( n931 & n9286 ) | ( n2468 & n9286 ) ;
  assign n12812 = ( n3494 & n6250 ) | ( n3494 & n8201 ) | ( n6250 & n8201 ) ;
  assign n12813 = n1347 & ~n12812 ;
  assign n12814 = ~n8929 & n12813 ;
  assign n12815 = n1166 ^ n403 ^ 1'b0 ;
  assign n12816 = n7652 & n12815 ;
  assign n12817 = ~n4713 & n12816 ;
  assign n12818 = ( ~n2409 & n12814 ) | ( ~n2409 & n12817 ) | ( n12814 & n12817 ) ;
  assign n12819 = n2645 & ~n5053 ;
  assign n12820 = n1415 & n12819 ;
  assign n12821 = n6914 & ~n12820 ;
  assign n12822 = n12821 ^ n806 ^ 1'b0 ;
  assign n12823 = ( ~n3833 & n7542 ) | ( ~n3833 & n12822 ) | ( n7542 & n12822 ) ;
  assign n12824 = n5017 | n6280 ;
  assign n12825 = n12824 ^ n6191 ^ 1'b0 ;
  assign n12826 = n5522 & ~n6012 ;
  assign n12827 = ( n9351 & n10968 ) | ( n9351 & ~n12826 ) | ( n10968 & ~n12826 ) ;
  assign n12828 = n5872 ^ x226 ^ 1'b0 ;
  assign n12829 = n12828 ^ n1881 ^ 1'b0 ;
  assign n12830 = n5814 | n12008 ;
  assign n12831 = n5173 | n12830 ;
  assign n12832 = ( n4818 & n5582 ) | ( n4818 & n6351 ) | ( n5582 & n6351 ) ;
  assign n12833 = n430 & n12832 ;
  assign n12834 = ~n5226 & n12833 ;
  assign n12835 = n10398 ^ n5925 ^ 1'b0 ;
  assign n12836 = ~n12834 & n12835 ;
  assign n12837 = n7904 ^ n5393 ^ 1'b0 ;
  assign n12841 = n3688 ^ n1199 ^ n992 ;
  assign n12842 = ( ~n3681 & n4857 ) | ( ~n3681 & n12841 ) | ( n4857 & n12841 ) ;
  assign n12838 = n2111 & n2208 ;
  assign n12839 = n12838 ^ n1983 ^ 1'b0 ;
  assign n12840 = ~n816 & n12839 ;
  assign n12843 = n12842 ^ n12840 ^ 1'b0 ;
  assign n12844 = n3905 & n4253 ;
  assign n12845 = n12844 ^ n6812 ^ 1'b0 ;
  assign n12846 = n12807 ^ n7232 ^ 1'b0 ;
  assign n12847 = ( ~n1323 & n5017 ) | ( ~n1323 & n9732 ) | ( n5017 & n9732 ) ;
  assign n12848 = ( x98 & ~n702 ) | ( x98 & n782 ) | ( ~n702 & n782 ) ;
  assign n12849 = ( n3814 & n12847 ) | ( n3814 & n12848 ) | ( n12847 & n12848 ) ;
  assign n12850 = n12849 ^ n5283 ^ 1'b0 ;
  assign n12851 = ~n12846 & n12850 ;
  assign n12852 = n12851 ^ n6023 ^ 1'b0 ;
  assign n12853 = n7915 ^ n5624 ^ 1'b0 ;
  assign n12854 = ( n2217 & n10767 ) | ( n2217 & ~n12853 ) | ( n10767 & ~n12853 ) ;
  assign n12855 = n5549 & n9532 ;
  assign n12856 = n12855 ^ n7046 ^ 1'b0 ;
  assign n12857 = n12856 ^ n6706 ^ 1'b0 ;
  assign n12858 = n1961 | n2386 ;
  assign n12859 = n12858 ^ n6307 ^ 1'b0 ;
  assign n12860 = n12859 ^ n7806 ^ n5619 ;
  assign n12861 = n1280 & n6015 ;
  assign n12862 = n10729 ^ n3208 ^ 1'b0 ;
  assign n12863 = n1727 & n12862 ;
  assign n12864 = n12861 & n12863 ;
  assign n12865 = n5296 & n12864 ;
  assign n12866 = ( n7988 & ~n11628 ) | ( n7988 & n12092 ) | ( ~n11628 & n12092 ) ;
  assign n12867 = n12866 ^ n5075 ^ 1'b0 ;
  assign n12868 = n3828 ^ n1403 ^ n1331 ;
  assign n12869 = n12089 | n12868 ;
  assign n12870 = n12869 ^ n1936 ^ 1'b0 ;
  assign n12872 = n11056 ^ n5014 ^ 1'b0 ;
  assign n12871 = n6474 | n10780 ;
  assign n12873 = n12872 ^ n12871 ^ 1'b0 ;
  assign n12874 = n627 & ~n2481 ;
  assign n12875 = ( x49 & n5364 ) | ( x49 & n6723 ) | ( n5364 & n6723 ) ;
  assign n12876 = n3755 & ~n12875 ;
  assign n12877 = n12876 ^ n7840 ^ 1'b0 ;
  assign n12878 = ( ~n2296 & n12874 ) | ( ~n2296 & n12877 ) | ( n12874 & n12877 ) ;
  assign n12879 = n12878 ^ n11966 ^ 1'b0 ;
  assign n12880 = n11173 ^ n9899 ^ 1'b0 ;
  assign n12881 = n10777 & n12880 ;
  assign n12882 = n12881 ^ n11437 ^ 1'b0 ;
  assign n12883 = n10380 ^ n4095 ^ 1'b0 ;
  assign n12885 = n4838 & ~n6003 ;
  assign n12884 = ~n1339 & n5156 ;
  assign n12886 = n12885 ^ n12884 ^ 1'b0 ;
  assign n12887 = n12886 ^ n4589 ^ 1'b0 ;
  assign n12889 = n3959 ^ n2764 ^ 1'b0 ;
  assign n12888 = n6373 ^ n1185 ^ 1'b0 ;
  assign n12890 = n12889 ^ n12888 ^ 1'b0 ;
  assign n12891 = n8578 & n12890 ;
  assign n12892 = n7675 ^ n2397 ^ 1'b0 ;
  assign n12893 = n3381 & ~n12892 ;
  assign n12894 = ~n10443 & n12893 ;
  assign n12895 = n12894 ^ n5812 ^ 1'b0 ;
  assign n12896 = ~n5773 & n12895 ;
  assign n12897 = n4920 & ~n5494 ;
  assign n12898 = ~n7753 & n12897 ;
  assign n12899 = ( n10636 & ~n11163 ) | ( n10636 & n12898 ) | ( ~n11163 & n12898 ) ;
  assign n12900 = n12899 ^ n6650 ^ 1'b0 ;
  assign n12901 = n12896 & n12900 ;
  assign n12902 = n3795 ^ n2799 ^ n644 ;
  assign n12903 = n12519 & ~n12902 ;
  assign n12905 = n2908 & ~n10745 ;
  assign n12906 = ~n1552 & n12905 ;
  assign n12904 = n10976 ^ n5660 ^ 1'b0 ;
  assign n12907 = n12906 ^ n12904 ^ n3252 ;
  assign n12908 = n6159 ^ n5480 ^ 1'b0 ;
  assign n12909 = n12908 ^ n6241 ^ 1'b0 ;
  assign n12910 = ( ~n1519 & n5801 ) | ( ~n1519 & n9665 ) | ( n5801 & n9665 ) ;
  assign n12911 = n12910 ^ n5483 ^ 1'b0 ;
  assign n12912 = n12911 ^ n3393 ^ n2471 ;
  assign n12913 = n12912 ^ n10036 ^ n7772 ;
  assign n12914 = n1120 | n2354 ;
  assign n12915 = n7426 ^ n2840 ^ 1'b0 ;
  assign n12916 = ~n8282 & n12915 ;
  assign n12917 = ( n4271 & ~n5391 ) | ( n4271 & n6540 ) | ( ~n5391 & n6540 ) ;
  assign n12918 = n12917 ^ n3110 ^ 1'b0 ;
  assign n12919 = ( n2548 & n3894 ) | ( n2548 & ~n8520 ) | ( n3894 & ~n8520 ) ;
  assign n12920 = n12919 ^ n7136 ^ n580 ;
  assign n12921 = n4593 & ~n6404 ;
  assign n12922 = n7037 ^ n3866 ^ 1'b0 ;
  assign n12923 = n9681 ^ n4288 ^ 1'b0 ;
  assign n12924 = n12922 & ~n12923 ;
  assign n12925 = n5363 & n12924 ;
  assign n12928 = ~n2509 & n4027 ;
  assign n12929 = n12928 ^ n1183 ^ 1'b0 ;
  assign n12926 = ~n9068 & n9885 ;
  assign n12927 = ~n8902 & n12926 ;
  assign n12930 = n12929 ^ n12927 ^ 1'b0 ;
  assign n12931 = n12253 & n12930 ;
  assign n12932 = n2843 & ~n3015 ;
  assign n12933 = ~n8163 & n12493 ;
  assign n12934 = n2927 & n12933 ;
  assign n12935 = n12934 ^ n6805 ^ 1'b0 ;
  assign n12936 = ~n12932 & n12935 ;
  assign n12937 = ~n6605 & n12936 ;
  assign n12938 = ~n1149 & n12937 ;
  assign n12939 = n12443 ^ n7113 ^ n310 ;
  assign n12940 = n12939 ^ n5437 ^ 1'b0 ;
  assign n12941 = n6571 & ~n12940 ;
  assign n12942 = ( n4332 & n6699 ) | ( n4332 & n12941 ) | ( n6699 & n12941 ) ;
  assign n12943 = ~n801 & n8569 ;
  assign n12944 = n12943 ^ n6313 ^ n398 ;
  assign n12945 = n12944 ^ n9103 ^ 1'b0 ;
  assign n12946 = n10789 & n12945 ;
  assign n12947 = ( n7369 & n12942 ) | ( n7369 & n12946 ) | ( n12942 & n12946 ) ;
  assign n12948 = ( n1226 & n8181 ) | ( n1226 & n12947 ) | ( n8181 & n12947 ) ;
  assign n12949 = n6776 & ~n11431 ;
  assign n12950 = ~n4487 & n12949 ;
  assign n12951 = ~n2856 & n8521 ;
  assign n12952 = n1034 & n12951 ;
  assign n12953 = n10848 ^ n10509 ^ n2047 ;
  assign n12954 = ~n9018 & n12953 ;
  assign n12955 = ( n4209 & n12952 ) | ( n4209 & n12954 ) | ( n12952 & n12954 ) ;
  assign n12956 = n6174 ^ n4078 ^ n3345 ;
  assign n12957 = n5679 & ~n12956 ;
  assign n12958 = n12957 ^ n3800 ^ x52 ;
  assign n12959 = n12005 ^ n743 ^ 1'b0 ;
  assign n12960 = n9447 ^ n5503 ^ x198 ;
  assign n12961 = n12362 ^ n4736 ^ 1'b0 ;
  assign n12962 = n6613 & n12961 ;
  assign n12963 = n2895 | n12962 ;
  assign n12964 = ( n2791 & n4616 ) | ( n2791 & n7446 ) | ( n4616 & n7446 ) ;
  assign n12965 = n12964 ^ n8331 ^ 1'b0 ;
  assign n12966 = n9149 | n12965 ;
  assign n12967 = n268 | n3204 ;
  assign n12968 = n12449 ^ n10732 ^ n4187 ;
  assign n12969 = ~n3207 & n12968 ;
  assign n12970 = n4314 ^ n2822 ^ 1'b0 ;
  assign n12971 = n6284 ^ n3187 ^ n381 ;
  assign n12972 = n12971 ^ n4359 ^ n1269 ;
  assign n12973 = n4625 | n7564 ;
  assign n12974 = n4261 ^ x12 ^ 1'b0 ;
  assign n12975 = n12973 & n12974 ;
  assign n12976 = x217 & ~n12975 ;
  assign n12977 = ~n3147 & n6271 ;
  assign n12978 = n12977 ^ n4200 ^ 1'b0 ;
  assign n12979 = n12976 | n12978 ;
  assign n12980 = n2068 & ~n12979 ;
  assign n12986 = n1557 | n2024 ;
  assign n12987 = ~n4928 & n8735 ;
  assign n12988 = n12986 | n12987 ;
  assign n12989 = n11076 | n12988 ;
  assign n12981 = n7338 ^ n1617 ^ 1'b0 ;
  assign n12982 = n12981 ^ n10900 ^ 1'b0 ;
  assign n12983 = n2244 & ~n12982 ;
  assign n12984 = n2884 & n12983 ;
  assign n12985 = n2133 & n12984 ;
  assign n12990 = n12989 ^ n12985 ^ 1'b0 ;
  assign n12991 = n12421 & ~n12990 ;
  assign n12992 = ~n2491 & n7260 ;
  assign n12993 = ~n1190 & n12992 ;
  assign n12994 = n12993 ^ x187 ^ 1'b0 ;
  assign n12995 = n5791 | n12994 ;
  assign n12996 = n1687 | n12995 ;
  assign n12997 = n12996 ^ n5546 ^ 1'b0 ;
  assign n12998 = n5052 & n12997 ;
  assign n12999 = n12244 ^ n11028 ^ n9545 ;
  assign n13000 = n8999 & ~n11203 ;
  assign n13001 = n4457 & n13000 ;
  assign n13002 = n7974 & n13001 ;
  assign n13003 = n6747 ^ n4417 ^ 1'b0 ;
  assign n13004 = ( ~n260 & n3798 ) | ( ~n260 & n13003 ) | ( n3798 & n13003 ) ;
  assign n13005 = n7852 | n12815 ;
  assign n13006 = n7026 & ~n8760 ;
  assign n13007 = n11018 & n13006 ;
  assign n13008 = n9676 ^ n2453 ^ n958 ;
  assign n13009 = n13008 ^ n9306 ^ 1'b0 ;
  assign n13010 = n8626 ^ n8381 ^ n327 ;
  assign n13011 = n10185 & ~n13010 ;
  assign n13012 = n13011 ^ n5655 ^ 1'b0 ;
  assign n13013 = n13012 ^ n5969 ^ 1'b0 ;
  assign n13014 = n13009 & ~n13013 ;
  assign n13015 = n7909 ^ n1493 ^ x81 ;
  assign n13016 = n13015 ^ n10623 ^ n9475 ;
  assign n13017 = ~n335 & n2220 ;
  assign n13018 = n13017 ^ n3097 ^ 1'b0 ;
  assign n13019 = n5057 & n13018 ;
  assign n13020 = ~n5888 & n9237 ;
  assign n13021 = ( n8052 & n13019 ) | ( n8052 & ~n13020 ) | ( n13019 & ~n13020 ) ;
  assign n13022 = n6846 ^ n5439 ^ 1'b0 ;
  assign n13023 = n11181 & n13022 ;
  assign n13024 = ~n599 & n3936 ;
  assign n13025 = n6898 & n10728 ;
  assign n13026 = n2282 | n3409 ;
  assign n13027 = n13026 ^ n8743 ^ 1'b0 ;
  assign n13028 = n1407 & ~n13027 ;
  assign n13032 = n6324 ^ n2251 ^ 1'b0 ;
  assign n13029 = ~n6028 & n8682 ;
  assign n13030 = n8515 & ~n13029 ;
  assign n13031 = ~n1890 & n13030 ;
  assign n13033 = n13032 ^ n13031 ^ 1'b0 ;
  assign n13034 = n384 | n5115 ;
  assign n13035 = n834 | n13034 ;
  assign n13036 = n9338 & n13035 ;
  assign n13038 = ~x117 & n2136 ;
  assign n13039 = ( ~n2075 & n5060 ) | ( ~n2075 & n13038 ) | ( n5060 & n13038 ) ;
  assign n13037 = x82 & ~n5253 ;
  assign n13040 = n13039 ^ n13037 ^ 1'b0 ;
  assign n13041 = ( n2085 & n2217 ) | ( n2085 & ~n13040 ) | ( n2217 & ~n13040 ) ;
  assign n13042 = n13041 ^ n11017 ^ n929 ;
  assign n13043 = ( n890 & n2052 ) | ( n890 & ~n3773 ) | ( n2052 & ~n3773 ) ;
  assign n13044 = n5289 | n13043 ;
  assign n13045 = n13044 ^ n1249 ^ 1'b0 ;
  assign n13046 = n8582 & ~n13045 ;
  assign n13047 = n13046 ^ n8243 ^ x90 ;
  assign n13050 = n2262 | n4122 ;
  assign n13048 = n3753 ^ n1256 ^ 1'b0 ;
  assign n13049 = x247 & ~n13048 ;
  assign n13051 = n13050 ^ n13049 ^ 1'b0 ;
  assign n13052 = ( ~n2962 & n6580 ) | ( ~n2962 & n13051 ) | ( n6580 & n13051 ) ;
  assign n13053 = n9976 ^ n1409 ^ 1'b0 ;
  assign n13054 = n3387 & n13053 ;
  assign n13055 = n4347 & ~n10859 ;
  assign n13056 = n13055 ^ n8781 ^ 1'b0 ;
  assign n13057 = ( n3037 & ~n3680 ) | ( n3037 & n6229 ) | ( ~n3680 & n6229 ) ;
  assign n13058 = ~n7912 & n13057 ;
  assign n13059 = n13058 ^ n10509 ^ 1'b0 ;
  assign n13060 = ~n13056 & n13059 ;
  assign n13061 = n11684 ^ n5446 ^ n588 ;
  assign n13062 = ~n5556 & n13061 ;
  assign n13063 = n12004 & ~n13062 ;
  assign n13065 = ( ~n1948 & n2047 ) | ( ~n1948 & n2702 ) | ( n2047 & n2702 ) ;
  assign n13064 = ~n987 & n1213 ;
  assign n13066 = n13065 ^ n13064 ^ n11691 ;
  assign n13067 = n6386 ^ x67 ^ 1'b0 ;
  assign n13068 = n3021 & n13067 ;
  assign n13069 = ~n13066 & n13068 ;
  assign n13070 = n9393 ^ n6620 ^ n5827 ;
  assign n13071 = n5065 & ~n12019 ;
  assign n13072 = n13070 & n13071 ;
  assign n13073 = ( n777 & n2562 ) | ( n777 & n13072 ) | ( n2562 & n13072 ) ;
  assign n13074 = n519 | n4302 ;
  assign n13075 = n7827 | n13074 ;
  assign n13076 = n13075 ^ n11584 ^ 1'b0 ;
  assign n13077 = n5153 ^ n1005 ^ 1'b0 ;
  assign n13079 = n7613 ^ n5833 ^ n2798 ;
  assign n13082 = n11467 ^ n5382 ^ n1543 ;
  assign n13080 = ~n4861 & n12413 ;
  assign n13081 = ~n7347 & n13080 ;
  assign n13083 = n13082 ^ n13081 ^ 1'b0 ;
  assign n13084 = n13079 | n13083 ;
  assign n13078 = ( n1134 & ~n2731 ) | ( n1134 & n8936 ) | ( ~n2731 & n8936 ) ;
  assign n13085 = n13084 ^ n13078 ^ 1'b0 ;
  assign n13086 = ( n2722 & n8505 ) | ( n2722 & n12941 ) | ( n8505 & n12941 ) ;
  assign n13087 = ~n8775 & n10247 ;
  assign n13094 = n9917 ^ n8183 ^ 1'b0 ;
  assign n13089 = n3314 ^ n2032 ^ n627 ;
  assign n13088 = n1374 | n12502 ;
  assign n13090 = n13089 ^ n13088 ^ 1'b0 ;
  assign n13091 = n887 & ~n13090 ;
  assign n13092 = n13091 ^ n2835 ^ 1'b0 ;
  assign n13093 = ~n604 & n13092 ;
  assign n13095 = n13094 ^ n13093 ^ 1'b0 ;
  assign n13096 = n3851 & n5045 ;
  assign n13097 = ( ~n407 & n4121 ) | ( ~n407 & n13096 ) | ( n4121 & n13096 ) ;
  assign n13105 = n2182 & ~n6728 ;
  assign n13101 = n520 | n1737 ;
  assign n13102 = n13101 ^ n1759 ^ 1'b0 ;
  assign n13103 = n4052 & ~n13102 ;
  assign n13104 = n13103 ^ n6791 ^ 1'b0 ;
  assign n13106 = n13105 ^ n13104 ^ 1'b0 ;
  assign n13098 = n2614 ^ n1306 ^ 1'b0 ;
  assign n13099 = n13098 ^ n6507 ^ 1'b0 ;
  assign n13100 = ( n2560 & ~n5020 ) | ( n2560 & n13099 ) | ( ~n5020 & n13099 ) ;
  assign n13107 = n13106 ^ n13100 ^ n3941 ;
  assign n13108 = ( n11969 & n13097 ) | ( n11969 & n13107 ) | ( n13097 & n13107 ) ;
  assign n13109 = n9934 ^ n1103 ^ 1'b0 ;
  assign n13112 = ~x151 & n3191 ;
  assign n13113 = n13112 ^ n4968 ^ n2421 ;
  assign n13114 = ( n8873 & n11048 ) | ( n8873 & n13113 ) | ( n11048 & n13113 ) ;
  assign n13110 = n3389 | n3421 ;
  assign n13111 = n852 | n13110 ;
  assign n13115 = n13114 ^ n13111 ^ 1'b0 ;
  assign n13116 = n675 | n1969 ;
  assign n13117 = x226 & n12886 ;
  assign n13118 = ( n4983 & n13116 ) | ( n4983 & ~n13117 ) | ( n13116 & ~n13117 ) ;
  assign n13119 = ( n389 & n4659 ) | ( n389 & ~n13118 ) | ( n4659 & ~n13118 ) ;
  assign n13120 = ( n1189 & ~n2791 ) | ( n1189 & n7430 ) | ( ~n2791 & n7430 ) ;
  assign n13122 = n451 & ~n5436 ;
  assign n13123 = ~n5801 & n13122 ;
  assign n13121 = ~n2449 & n3494 ;
  assign n13124 = n13123 ^ n13121 ^ n10582 ;
  assign n13125 = n13120 | n13124 ;
  assign n13126 = n12813 | n13125 ;
  assign n13127 = ~n3285 & n4431 ;
  assign n13128 = n12524 | n13127 ;
  assign n13129 = n1294 | n13128 ;
  assign n13130 = n13129 ^ n12338 ^ n8488 ;
  assign n13131 = n3238 | n9375 ;
  assign n13132 = n6891 | n13131 ;
  assign n13133 = n13132 ^ n8525 ^ n345 ;
  assign n13134 = n2024 & ~n5686 ;
  assign n13135 = n13134 ^ n7606 ^ 1'b0 ;
  assign n13136 = n1487 | n13135 ;
  assign n13137 = n13136 ^ n2496 ^ 1'b0 ;
  assign n13138 = n9134 ^ n8266 ^ n4451 ;
  assign n13139 = n9103 ^ n5209 ^ 1'b0 ;
  assign n13140 = n5778 & n9010 ;
  assign n13141 = n13140 ^ n2066 ^ 1'b0 ;
  assign n13142 = n13139 | n13141 ;
  assign n13143 = n2030 & ~n6927 ;
  assign n13144 = n13143 ^ n10275 ^ 1'b0 ;
  assign n13145 = ~n2437 & n6093 ;
  assign n13146 = n13145 ^ n12079 ^ 1'b0 ;
  assign n13147 = n13146 ^ n7354 ^ 1'b0 ;
  assign n13148 = n958 & n2257 ;
  assign n13149 = n13148 ^ n1472 ^ 1'b0 ;
  assign n13150 = n5087 & ~n13149 ;
  assign n13151 = ( n2740 & n7200 ) | ( n2740 & ~n13150 ) | ( n7200 & ~n13150 ) ;
  assign n13152 = ~n10122 & n13151 ;
  assign n13153 = ~n4670 & n4984 ;
  assign n13154 = ~n1865 & n2439 ;
  assign n13155 = n13154 ^ n3712 ^ 1'b0 ;
  assign n13156 = ( n537 & ~n5463 ) | ( n537 & n13155 ) | ( ~n5463 & n13155 ) ;
  assign n13157 = n13156 ^ n1405 ^ 1'b0 ;
  assign n13158 = n9393 & ~n13157 ;
  assign n13159 = ( n3810 & ~n13153 ) | ( n3810 & n13158 ) | ( ~n13153 & n13158 ) ;
  assign n13160 = ( n3322 & n12541 ) | ( n3322 & n13159 ) | ( n12541 & n13159 ) ;
  assign n13161 = n5405 ^ n4390 ^ 1'b0 ;
  assign n13162 = n6056 & n13161 ;
  assign n13163 = n5565 | n13162 ;
  assign n13164 = n2331 ^ n727 ^ x122 ;
  assign n13165 = n844 & ~n13164 ;
  assign n13166 = ~n13163 & n13165 ;
  assign n13167 = n10558 & ~n12969 ;
  assign n13168 = n1566 & ~n4244 ;
  assign n13169 = n8821 ^ n2505 ^ 1'b0 ;
  assign n13170 = x160 & ~n13169 ;
  assign n13171 = n13170 ^ n2575 ^ 1'b0 ;
  assign n13172 = ( n3747 & n10650 ) | ( n3747 & n13171 ) | ( n10650 & n13171 ) ;
  assign n13173 = ( n4104 & n13168 ) | ( n4104 & n13172 ) | ( n13168 & n13172 ) ;
  assign n13174 = n716 & n2538 ;
  assign n13175 = ( n953 & ~n5826 ) | ( n953 & n9630 ) | ( ~n5826 & n9630 ) ;
  assign n13176 = n3356 & ~n3599 ;
  assign n13177 = n7176 ^ n2421 ^ 1'b0 ;
  assign n13178 = n773 & ~n13177 ;
  assign n13179 = n9020 & n13178 ;
  assign n13180 = n4542 & n10861 ;
  assign n13181 = n4371 ^ n4223 ^ 1'b0 ;
  assign n13182 = n11125 & ~n13181 ;
  assign n13183 = n13182 ^ n6686 ^ 1'b0 ;
  assign n13184 = n3527 | n13183 ;
  assign n13185 = n13184 ^ n10183 ^ 1'b0 ;
  assign n13186 = n4690 & ~n13185 ;
  assign n13187 = n3282 | n9576 ;
  assign n13188 = n12474 ^ n12296 ^ 1'b0 ;
  assign n13189 = n2230 ^ n1576 ^ 1'b0 ;
  assign n13190 = n3324 | n9578 ;
  assign n13191 = n13189 | n13190 ;
  assign n13196 = n5255 ^ n5241 ^ 1'b0 ;
  assign n13195 = n2283 | n8296 ;
  assign n13197 = n13196 ^ n13195 ^ n3984 ;
  assign n13192 = ~n895 & n1936 ;
  assign n13193 = n455 & n13192 ;
  assign n13194 = n4197 & ~n13193 ;
  assign n13198 = n13197 ^ n13194 ^ 1'b0 ;
  assign n13199 = n6147 & n13198 ;
  assign n13200 = ~n12511 & n13199 ;
  assign n13201 = n3181 ^ n2878 ^ n1051 ;
  assign n13202 = n9316 ^ n8376 ^ n3381 ;
  assign n13203 = n10914 | n13202 ;
  assign n13204 = n13203 ^ n6264 ^ 1'b0 ;
  assign n13206 = n9561 ^ n7779 ^ 1'b0 ;
  assign n13205 = n1755 ^ x139 ^ 1'b0 ;
  assign n13207 = n13206 ^ n13205 ^ 1'b0 ;
  assign n13208 = n10542 ^ n7415 ^ x71 ;
  assign n13209 = n4522 ^ n2275 ^ 1'b0 ;
  assign n13210 = n11043 ^ n898 ^ 1'b0 ;
  assign n13211 = n3264 & ~n5922 ;
  assign n13212 = n10536 & ~n13211 ;
  assign n13213 = ( n7279 & ~n9632 ) | ( n7279 & n11047 ) | ( ~n9632 & n11047 ) ;
  assign n13214 = n13213 ^ n11152 ^ n9721 ;
  assign n13215 = n2387 ^ x188 ^ 1'b0 ;
  assign n13216 = n13215 ^ n12602 ^ n640 ;
  assign n13217 = n9144 & ~n13216 ;
  assign n13218 = n13217 ^ n1898 ^ 1'b0 ;
  assign n13219 = n3542 ^ n3256 ^ n1842 ;
  assign n13220 = ( n6371 & ~n8049 ) | ( n6371 & n13219 ) | ( ~n8049 & n13219 ) ;
  assign n13221 = n13220 ^ n5990 ^ n5381 ;
  assign n13222 = n4071 & n13221 ;
  assign n13223 = n3439 & n13222 ;
  assign n13224 = n9472 ^ n544 ^ 1'b0 ;
  assign n13225 = ~n7195 & n13224 ;
  assign n13226 = ( n1096 & n3679 ) | ( n1096 & n6706 ) | ( n3679 & n6706 ) ;
  assign n13227 = n2769 ^ n1051 ^ 1'b0 ;
  assign n13228 = ~n5386 & n13227 ;
  assign n13229 = ~n2873 & n13228 ;
  assign n13230 = n13226 | n13229 ;
  assign n13231 = n7235 & ~n13230 ;
  assign n13232 = n800 & ~n13231 ;
  assign n13233 = ~n13225 & n13232 ;
  assign n13234 = n11171 ^ n7064 ^ 1'b0 ;
  assign n13235 = ( n2454 & n3289 ) | ( n2454 & ~n3338 ) | ( n3289 & ~n3338 ) ;
  assign n13236 = n13235 ^ n2804 ^ 1'b0 ;
  assign n13237 = n13234 | n13236 ;
  assign n13238 = ~n5376 & n11046 ;
  assign n13239 = ~n5754 & n13238 ;
  assign n13240 = n10519 ^ n4948 ^ 1'b0 ;
  assign n13241 = n3238 | n13240 ;
  assign n13242 = ~n604 & n4154 ;
  assign n13243 = n4039 & n13242 ;
  assign n13246 = ~n2116 & n6031 ;
  assign n13247 = n13246 ^ n1653 ^ 1'b0 ;
  assign n13248 = n9141 & n13247 ;
  assign n13244 = n6291 ^ n4970 ^ 1'b0 ;
  assign n13245 = n4746 & ~n13244 ;
  assign n13249 = n13248 ^ n13245 ^ 1'b0 ;
  assign n13250 = n10269 ^ n9626 ^ 1'b0 ;
  assign n13251 = n884 | n1797 ;
  assign n13252 = ( n259 & ~n709 ) | ( n259 & n990 ) | ( ~n709 & n990 ) ;
  assign n13253 = n349 | n13074 ;
  assign n13254 = n13252 | n13253 ;
  assign n13256 = n7157 ^ n2605 ^ 1'b0 ;
  assign n13255 = n13216 ^ n3387 ^ n3100 ;
  assign n13257 = n13256 ^ n13255 ^ n1429 ;
  assign n13258 = n1651 & n7400 ;
  assign n13259 = n13258 ^ n3262 ^ 1'b0 ;
  assign n13260 = n12086 ^ n1776 ^ 1'b0 ;
  assign n13261 = n298 & ~n4943 ;
  assign n13262 = ~x40 & n1343 ;
  assign n13263 = ( ~n4950 & n13261 ) | ( ~n4950 & n13262 ) | ( n13261 & n13262 ) ;
  assign n13264 = n13263 ^ n5641 ^ 1'b0 ;
  assign n13265 = n13118 | n13264 ;
  assign n13266 = n5974 ^ n303 ^ 1'b0 ;
  assign n13267 = ~n5230 & n13266 ;
  assign n13268 = ~n1082 & n13267 ;
  assign n13270 = n1306 & n7448 ;
  assign n13271 = n13270 ^ n3369 ^ n2880 ;
  assign n13272 = n5495 ^ n4858 ^ 1'b0 ;
  assign n13273 = x158 & n13272 ;
  assign n13274 = ~n13271 & n13273 ;
  assign n13269 = ~n3640 & n12627 ;
  assign n13275 = n13274 ^ n13269 ^ n2808 ;
  assign n13276 = n5204 ^ n1448 ^ 1'b0 ;
  assign n13277 = n13276 ^ n10885 ^ 1'b0 ;
  assign n13278 = ~n3305 & n7215 ;
  assign n13279 = n4140 & n13278 ;
  assign n13280 = ( n8867 & n12487 ) | ( n8867 & n13279 ) | ( n12487 & n13279 ) ;
  assign n13281 = n7755 & n9176 ;
  assign n13282 = n1389 & n6688 ;
  assign n13283 = n13282 ^ n8428 ^ 1'b0 ;
  assign n13284 = ( ~x244 & n783 ) | ( ~x244 & n7044 ) | ( n783 & n7044 ) ;
  assign n13285 = n557 & n2742 ;
  assign n13286 = ( n4397 & n5320 ) | ( n4397 & n6853 ) | ( n5320 & n6853 ) ;
  assign n13287 = n3444 & n9581 ;
  assign n13288 = n13287 ^ n409 ^ 1'b0 ;
  assign n13289 = n13288 ^ n7863 ^ 1'b0 ;
  assign n13290 = n1047 & n13289 ;
  assign n13291 = ( ~n2517 & n13286 ) | ( ~n2517 & n13290 ) | ( n13286 & n13290 ) ;
  assign n13292 = x2 & ~n5569 ;
  assign n13293 = n13292 ^ n13263 ^ 1'b0 ;
  assign n13294 = n2942 & n7339 ;
  assign n13295 = n13294 ^ n7641 ^ 1'b0 ;
  assign n13296 = n3146 & n3727 ;
  assign n13297 = n13296 ^ n4122 ^ 1'b0 ;
  assign n13298 = n13297 ^ n11012 ^ 1'b0 ;
  assign n13299 = ~n5631 & n13298 ;
  assign n13300 = n6310 & n7066 ;
  assign n13301 = ~n4714 & n10349 ;
  assign n13302 = ~n4561 & n10644 ;
  assign n13303 = n13301 & n13302 ;
  assign n13304 = ( n1635 & ~n6431 ) | ( n1635 & n7257 ) | ( ~n6431 & n7257 ) ;
  assign n13305 = ~n629 & n3099 ;
  assign n13306 = n4273 & n13305 ;
  assign n13307 = x146 & n1055 ;
  assign n13308 = n13307 ^ n4476 ^ 1'b0 ;
  assign n13309 = n13308 ^ n475 ^ 1'b0 ;
  assign n13310 = n13306 | n13309 ;
  assign n13311 = n1707 | n13310 ;
  assign n13312 = n4433 | n13311 ;
  assign n13313 = n6997 ^ n6077 ^ n3299 ;
  assign n13314 = n292 | n2135 ;
  assign n13315 = n13314 ^ x225 ^ 1'b0 ;
  assign n13316 = n13313 & ~n13315 ;
  assign n13317 = n10448 ^ n1532 ^ 1'b0 ;
  assign n13318 = ~n4353 & n4544 ;
  assign n13319 = n7973 & ~n13318 ;
  assign n13320 = n500 & n5672 ;
  assign n13321 = n13320 ^ n9351 ^ 1'b0 ;
  assign n13322 = n3464 ^ x240 ^ 1'b0 ;
  assign n13323 = n6093 & n13322 ;
  assign n13324 = ~n1709 & n13323 ;
  assign n13325 = n3009 ^ n807 ^ 1'b0 ;
  assign n13326 = n1149 & n13325 ;
  assign n13327 = n7988 ^ n2830 ^ 1'b0 ;
  assign n13328 = n13326 & ~n13327 ;
  assign n13329 = n2051 & n13328 ;
  assign n13330 = n2645 & n9714 ;
  assign n13331 = x172 & n13330 ;
  assign n13332 = n12361 ^ n5361 ^ 1'b0 ;
  assign n13333 = ~n10949 & n13332 ;
  assign n13334 = ~n2267 & n4868 ;
  assign n13335 = n13334 ^ n2783 ^ 1'b0 ;
  assign n13336 = x110 & ~n2726 ;
  assign n13337 = n13336 ^ n3233 ^ 1'b0 ;
  assign n13338 = ~n2764 & n13337 ;
  assign n13339 = n4013 & n13338 ;
  assign n13340 = n13335 & n13339 ;
  assign n13341 = n4052 & ~n13227 ;
  assign n13342 = n13341 ^ n4932 ^ n2688 ;
  assign n13343 = n11771 ^ n10191 ^ n5368 ;
  assign n13344 = n13343 ^ n12902 ^ n1352 ;
  assign n13345 = ( n10961 & n11196 ) | ( n10961 & n13040 ) | ( n11196 & n13040 ) ;
  assign n13346 = ( n3891 & n4878 ) | ( n3891 & ~n5591 ) | ( n4878 & ~n5591 ) ;
  assign n13347 = n720 | n7562 ;
  assign n13348 = n3375 | n13347 ;
  assign n13349 = ~n4139 & n13348 ;
  assign n13350 = ~n13346 & n13349 ;
  assign n13351 = n12328 ^ n1921 ^ 1'b0 ;
  assign n13352 = x172 & ~n13351 ;
  assign n13353 = n11283 & n13352 ;
  assign n13354 = n8911 ^ n7813 ^ n6653 ;
  assign n13355 = n4925 ^ n826 ^ 1'b0 ;
  assign n13356 = n9174 & n13355 ;
  assign n13357 = n13356 ^ n9100 ^ n6661 ;
  assign n13358 = n13357 ^ n9096 ^ 1'b0 ;
  assign n13359 = n5246 & n10708 ;
  assign n13360 = x209 & n2736 ;
  assign n13361 = ~n13176 & n13360 ;
  assign n13362 = n12967 ^ n7927 ^ n1000 ;
  assign n13363 = ( n3567 & n5287 ) | ( n3567 & ~n10365 ) | ( n5287 & ~n10365 ) ;
  assign n13364 = n2354 | n5848 ;
  assign n13365 = n4243 & ~n13364 ;
  assign n13366 = n13363 | n13365 ;
  assign n13367 = n13366 ^ n5507 ^ 1'b0 ;
  assign n13372 = n2041 | n3487 ;
  assign n13373 = n13372 ^ n5608 ^ 1'b0 ;
  assign n13374 = ( ~n9148 & n10332 ) | ( ~n9148 & n13373 ) | ( n10332 & n13373 ) ;
  assign n13368 = ( n329 & ~n1655 ) | ( n329 & n5947 ) | ( ~n1655 & n5947 ) ;
  assign n13369 = n8067 ^ n5491 ^ n1746 ;
  assign n13370 = ( ~n1562 & n13368 ) | ( ~n1562 & n13369 ) | ( n13368 & n13369 ) ;
  assign n13371 = n6471 & ~n13370 ;
  assign n13375 = n13374 ^ n13371 ^ 1'b0 ;
  assign n13376 = ( n3379 & n5855 ) | ( n3379 & n13375 ) | ( n5855 & n13375 ) ;
  assign n13378 = n9240 ^ n5429 ^ 1'b0 ;
  assign n13379 = ~n4067 & n13378 ;
  assign n13380 = n13379 ^ n12768 ^ 1'b0 ;
  assign n13381 = n7932 ^ n1308 ^ 1'b0 ;
  assign n13382 = n13380 | n13381 ;
  assign n13377 = n2990 ^ n1572 ^ n440 ;
  assign n13383 = n13382 ^ n13377 ^ 1'b0 ;
  assign n13384 = n5279 & n13383 ;
  assign n13385 = ( n4048 & n12288 ) | ( n4048 & n13384 ) | ( n12288 & n13384 ) ;
  assign n13386 = n12566 ^ n4754 ^ 1'b0 ;
  assign n13387 = ~n316 & n6874 ;
  assign n13388 = ~n13386 & n13387 ;
  assign n13389 = n2023 | n7131 ;
  assign n13390 = n384 & ~n3689 ;
  assign n13391 = n6045 & ~n13390 ;
  assign n13392 = n7259 & n7956 ;
  assign n13393 = ~n6080 & n13392 ;
  assign n13394 = n7369 ^ n3690 ^ 1'b0 ;
  assign n13395 = n6313 | n13394 ;
  assign n13396 = n2169 & ~n13395 ;
  assign n13397 = ( n10559 & ~n12123 ) | ( n10559 & n13396 ) | ( ~n12123 & n13396 ) ;
  assign n13398 = ~n3283 & n3797 ;
  assign n13399 = ( n6817 & ~n8292 ) | ( n6817 & n13398 ) | ( ~n8292 & n13398 ) ;
  assign n13400 = ~n8251 & n13399 ;
  assign n13401 = n2778 | n5927 ;
  assign n13402 = n13401 ^ n1682 ^ 1'b0 ;
  assign n13403 = n13402 ^ n6302 ^ n1639 ;
  assign n13404 = n13403 ^ n4999 ^ 1'b0 ;
  assign n13405 = n8483 | n10120 ;
  assign n13406 = n7402 ^ n1858 ^ 1'b0 ;
  assign n13407 = n4298 & n13406 ;
  assign n13408 = n2974 & n13407 ;
  assign n13409 = n13408 ^ n11201 ^ 1'b0 ;
  assign n13410 = n6678 | n13409 ;
  assign n13411 = n13410 ^ n859 ^ 1'b0 ;
  assign n13413 = ~n7081 & n8256 ;
  assign n13414 = ~n3831 & n13413 ;
  assign n13412 = ~n2005 & n11510 ;
  assign n13415 = n13414 ^ n13412 ^ 1'b0 ;
  assign n13416 = ( n4143 & ~n7983 ) | ( n4143 & n11465 ) | ( ~n7983 & n11465 ) ;
  assign n13417 = ( n722 & ~n7476 ) | ( n722 & n10631 ) | ( ~n7476 & n10631 ) ;
  assign n13418 = n10298 ^ n4128 ^ n350 ;
  assign n13419 = n5133 & ~n8419 ;
  assign n13420 = n13419 ^ n5437 ^ 1'b0 ;
  assign n13421 = n3439 & ~n9051 ;
  assign n13422 = ~n8582 & n13421 ;
  assign n13424 = ( n540 & n4179 ) | ( n540 & n4891 ) | ( n4179 & n4891 ) ;
  assign n13423 = n471 & n9967 ;
  assign n13425 = n13424 ^ n13423 ^ n8718 ;
  assign n13426 = n1244 | n8050 ;
  assign n13427 = n4984 | n13426 ;
  assign n13428 = n8069 & n13427 ;
  assign n13429 = ~n13425 & n13428 ;
  assign n13430 = n5830 | n10121 ;
  assign n13431 = n2297 | n13430 ;
  assign n13432 = n13431 ^ n9168 ^ n6310 ;
  assign n13433 = n1925 & ~n8244 ;
  assign n13434 = n2058 | n9929 ;
  assign n13435 = n13433 & ~n13434 ;
  assign n13436 = ~n2819 & n6973 ;
  assign n13437 = n4189 & ~n5126 ;
  assign n13438 = n13437 ^ n3145 ^ x147 ;
  assign n13439 = n10281 ^ n4895 ^ n4461 ;
  assign n13440 = ~n13438 & n13439 ;
  assign n13441 = n5713 & n6082 ;
  assign n13442 = ~n8047 & n13441 ;
  assign n13443 = n3842 | n13442 ;
  assign n13444 = ( n1133 & n3192 ) | ( n1133 & ~n12634 ) | ( n3192 & ~n12634 ) ;
  assign n13445 = ~n3305 & n13444 ;
  assign n13446 = ~n1454 & n13445 ;
  assign n13447 = n8955 & ~n13446 ;
  assign n13448 = n13447 ^ n5402 ^ 1'b0 ;
  assign n13449 = ( x46 & n10501 ) | ( x46 & ~n13448 ) | ( n10501 & ~n13448 ) ;
  assign n13450 = n8327 ^ n6858 ^ 1'b0 ;
  assign n13451 = n8808 ^ n1061 ^ 1'b0 ;
  assign n13452 = n7342 ^ n4016 ^ n2708 ;
  assign n13453 = ~n2919 & n13452 ;
  assign n13454 = ( n1197 & ~n2165 ) | ( n1197 & n6248 ) | ( ~n2165 & n6248 ) ;
  assign n13455 = n9251 & ~n13454 ;
  assign n13456 = n13455 ^ n8672 ^ 1'b0 ;
  assign n13457 = n13456 ^ n5834 ^ 1'b0 ;
  assign n13458 = n13453 & ~n13457 ;
  assign n13459 = n13458 ^ n6552 ^ n2971 ;
  assign n13460 = n599 & ~n7427 ;
  assign n13461 = n3252 & n13460 ;
  assign n13462 = n5717 | n13461 ;
  assign n13463 = n11521 | n13462 ;
  assign n13464 = n7802 & ~n13463 ;
  assign n13465 = n9336 ^ n500 ^ 1'b0 ;
  assign n13466 = n5953 ^ n5330 ^ 1'b0 ;
  assign n13467 = n4050 ^ n3065 ^ 1'b0 ;
  assign n13468 = n12285 | n13467 ;
  assign n13469 = n1956 & ~n2914 ;
  assign n13470 = ~n1956 & n13469 ;
  assign n13471 = n974 & n13470 ;
  assign n13472 = n5118 & n13471 ;
  assign n13473 = n2107 & n13472 ;
  assign n13474 = ~n4925 & n13473 ;
  assign n13475 = n4514 ^ n1511 ^ n606 ;
  assign n13476 = n13475 ^ n8634 ^ 1'b0 ;
  assign n13477 = n13474 | n13476 ;
  assign n13478 = n2851 ^ n1727 ^ 1'b0 ;
  assign n13479 = n13478 ^ n12709 ^ 1'b0 ;
  assign n13480 = n13479 ^ n4979 ^ 1'b0 ;
  assign n13481 = n4006 ^ n966 ^ 1'b0 ;
  assign n13482 = ~n2050 & n6981 ;
  assign n13483 = n13482 ^ n9574 ^ 1'b0 ;
  assign n13484 = x55 & ~n13483 ;
  assign n13485 = n13481 & n13484 ;
  assign n13487 = ~n6994 & n9447 ;
  assign n13488 = ~n3140 & n13487 ;
  assign n13486 = n9933 | n10505 ;
  assign n13489 = n13488 ^ n13486 ^ 1'b0 ;
  assign n13490 = ( n2412 & n5879 ) | ( n2412 & ~n7874 ) | ( n5879 & ~n7874 ) ;
  assign n13491 = n6313 ^ n5171 ^ 1'b0 ;
  assign n13492 = n13490 & n13491 ;
  assign n13493 = n13492 ^ n9653 ^ 1'b0 ;
  assign n13501 = n1505 ^ n1247 ^ 1'b0 ;
  assign n13498 = n9378 ^ n7726 ^ 1'b0 ;
  assign n13494 = n2095 | n4991 ;
  assign n13495 = ( n5072 & ~n5665 ) | ( n5072 & n13494 ) | ( ~n5665 & n13494 ) ;
  assign n13496 = n1904 & ~n7942 ;
  assign n13497 = n13495 & n13496 ;
  assign n13499 = n13498 ^ n13497 ^ n8553 ;
  assign n13500 = ~n8867 & n13499 ;
  assign n13502 = n13501 ^ n13500 ^ 1'b0 ;
  assign n13503 = ( ~n3814 & n7238 ) | ( ~n3814 & n12382 ) | ( n7238 & n12382 ) ;
  assign n13504 = n4299 ^ n3015 ^ 1'b0 ;
  assign n13505 = ~n13503 & n13504 ;
  assign n13506 = ( x57 & n678 ) | ( x57 & n3371 ) | ( n678 & n3371 ) ;
  assign n13507 = n6272 | n13506 ;
  assign n13510 = n4416 & n5687 ;
  assign n13511 = ~n7569 & n13510 ;
  assign n13512 = n13511 ^ n8286 ^ n3012 ;
  assign n13513 = n13512 ^ n6892 ^ 1'b0 ;
  assign n13514 = ~n9668 & n10925 ;
  assign n13515 = n13513 & n13514 ;
  assign n13508 = n8454 ^ n3816 ^ n3770 ;
  assign n13509 = n888 & ~n13508 ;
  assign n13516 = n13515 ^ n13509 ^ 1'b0 ;
  assign n13517 = n6628 ^ n3383 ^ 1'b0 ;
  assign n13518 = n7801 | n13517 ;
  assign n13519 = n1206 & n3517 ;
  assign n13520 = n1116 & ~n6249 ;
  assign n13521 = n10191 & n13520 ;
  assign n13522 = n8579 & n11813 ;
  assign n13523 = n13521 & n13522 ;
  assign n13524 = ( ~n992 & n13519 ) | ( ~n992 & n13523 ) | ( n13519 & n13523 ) ;
  assign n13525 = n3409 ^ n1684 ^ n1063 ;
  assign n13526 = n13525 ^ n10169 ^ 1'b0 ;
  assign n13527 = n5034 & ~n6376 ;
  assign n13528 = n1284 & n1963 ;
  assign n13529 = n13528 ^ n13283 ^ 1'b0 ;
  assign n13530 = n11988 ^ n9345 ^ n4101 ;
  assign n13531 = n5263 & n13530 ;
  assign n13532 = n4139 | n6001 ;
  assign n13533 = n13532 ^ n757 ^ 1'b0 ;
  assign n13534 = ( ~n6905 & n12313 ) | ( ~n6905 & n13533 ) | ( n12313 & n13533 ) ;
  assign n13535 = ( n1727 & n2859 ) | ( n1727 & n7280 ) | ( n2859 & n7280 ) ;
  assign n13536 = n12769 ^ x147 ^ 1'b0 ;
  assign n13537 = n13535 | n13536 ;
  assign n13538 = ~n3351 & n9496 ;
  assign n13542 = ~x156 & n3855 ;
  assign n13539 = ~n8491 & n8702 ;
  assign n13540 = n12402 & n13539 ;
  assign n13541 = x153 & ~n13540 ;
  assign n13543 = n13542 ^ n13541 ^ 1'b0 ;
  assign n13544 = n5479 & n6944 ;
  assign n13545 = n1724 & n13544 ;
  assign n13546 = n3304 | n13545 ;
  assign n13547 = n12897 & ~n13033 ;
  assign n13548 = n13546 & n13547 ;
  assign n13549 = n1187 ^ n453 ^ 1'b0 ;
  assign n13550 = n2955 & ~n13549 ;
  assign n13551 = n1916 & ~n4681 ;
  assign n13552 = n12070 | n13551 ;
  assign n13553 = x166 | n13552 ;
  assign n13554 = n1413 & ~n13553 ;
  assign n13555 = n13554 ^ n3473 ^ 1'b0 ;
  assign n13556 = n4963 & n5920 ;
  assign n13557 = n557 & n3328 ;
  assign n13558 = ~n2618 & n13175 ;
  assign n13559 = ~n5975 & n13558 ;
  assign n13560 = n10773 | n11285 ;
  assign n13561 = ( ~n7627 & n8958 ) | ( ~n7627 & n9433 ) | ( n8958 & n9433 ) ;
  assign n13562 = n13561 ^ n10039 ^ n5627 ;
  assign n13563 = n6062 & ~n10180 ;
  assign n13568 = ~n7128 & n9102 ;
  assign n13569 = n5274 & n13568 ;
  assign n13564 = ( n375 & n801 ) | ( n375 & n4159 ) | ( n801 & n4159 ) ;
  assign n13565 = n13564 ^ n557 ^ 1'b0 ;
  assign n13566 = x1 & ~n13565 ;
  assign n13567 = ~n12846 & n13566 ;
  assign n13570 = n13569 ^ n13567 ^ 1'b0 ;
  assign n13571 = ( n4773 & n4997 ) | ( n4773 & ~n13570 ) | ( n4997 & ~n13570 ) ;
  assign n13572 = n5913 & n9653 ;
  assign n13573 = n13572 ^ n2692 ^ 1'b0 ;
  assign n13574 = n3325 & ~n13573 ;
  assign n13575 = n10937 ^ n3402 ^ 1'b0 ;
  assign n13576 = n11256 | n13575 ;
  assign n13577 = n7721 | n13373 ;
  assign n13578 = n4498 | n13577 ;
  assign n13579 = ( n7753 & n13576 ) | ( n7753 & n13578 ) | ( n13576 & n13578 ) ;
  assign n13584 = ( n6125 & n6408 ) | ( n6125 & n7067 ) | ( n6408 & n7067 ) ;
  assign n13581 = n7913 ^ n2007 ^ x85 ;
  assign n13580 = n2106 & ~n2152 ;
  assign n13582 = n13581 ^ n13580 ^ 1'b0 ;
  assign n13583 = ( n2688 & n9580 ) | ( n2688 & ~n13582 ) | ( n9580 & ~n13582 ) ;
  assign n13585 = n13584 ^ n13583 ^ 1'b0 ;
  assign n13586 = ~n4512 & n7629 ;
  assign n13587 = n7169 & n13586 ;
  assign n13589 = ~n2538 & n6982 ;
  assign n13588 = ~n7784 & n10414 ;
  assign n13590 = n13589 ^ n13588 ^ 1'b0 ;
  assign n13591 = n13587 & ~n13590 ;
  assign n13592 = n13591 ^ n4257 ^ 1'b0 ;
  assign n13593 = n12225 ^ n9360 ^ n3781 ;
  assign n13594 = n13593 ^ n2819 ^ 1'b0 ;
  assign n13595 = n11221 & ~n13594 ;
  assign n13596 = n7854 ^ n4857 ^ 1'b0 ;
  assign n13597 = n617 & n13596 ;
  assign n13598 = n2531 & ~n3354 ;
  assign n13599 = n6738 & ~n13598 ;
  assign n13600 = ~n13597 & n13599 ;
  assign n13601 = n2859 | n11631 ;
  assign n13602 = n13601 ^ n7212 ^ 1'b0 ;
  assign n13603 = n13513 ^ n8787 ^ 1'b0 ;
  assign n13604 = ~n821 & n1636 ;
  assign n13605 = n13604 ^ n7787 ^ n5135 ;
  assign n13606 = n7489 ^ n2639 ^ x51 ;
  assign n13607 = ~n1000 & n13606 ;
  assign n13608 = ~n2152 & n9089 ;
  assign n13609 = ~n2026 & n13608 ;
  assign n13610 = n6364 ^ n3910 ^ 1'b0 ;
  assign n13611 = n4330 | n12530 ;
  assign n13612 = n6058 & ~n13611 ;
  assign n13613 = n1283 & ~n3633 ;
  assign n13614 = n3666 & n13613 ;
  assign n13615 = n3773 ^ n2453 ^ 1'b0 ;
  assign n13616 = ~n13614 & n13615 ;
  assign n13617 = n9690 ^ n8951 ^ n7902 ;
  assign n13619 = n4370 ^ n1542 ^ n1107 ;
  assign n13620 = n11119 & ~n13619 ;
  assign n13618 = n1108 & ~n3342 ;
  assign n13621 = n13620 ^ n13618 ^ 1'b0 ;
  assign n13622 = n6724 ^ n4788 ^ 1'b0 ;
  assign n13623 = n1094 ^ x155 ^ 1'b0 ;
  assign n13624 = n11589 ^ n6368 ^ 1'b0 ;
  assign n13625 = ~n1636 & n13624 ;
  assign n13626 = n13625 ^ n12407 ^ 1'b0 ;
  assign n13627 = n7002 & n13354 ;
  assign n13631 = n3506 & ~n4884 ;
  assign n13632 = n13631 ^ n10820 ^ 1'b0 ;
  assign n13629 = x0 & x81 ;
  assign n13630 = n13629 ^ n9652 ^ n3896 ;
  assign n13628 = n3898 ^ n3645 ^ 1'b0 ;
  assign n13633 = n13632 ^ n13630 ^ n13628 ;
  assign n13634 = n11329 ^ n4493 ^ 1'b0 ;
  assign n13635 = n9163 & n13634 ;
  assign n13639 = n6901 ^ n4994 ^ 1'b0 ;
  assign n13640 = n3898 & n13639 ;
  assign n13641 = ~n9452 & n13640 ;
  assign n13642 = n13499 & n13641 ;
  assign n13636 = ~n8191 & n12239 ;
  assign n13637 = n1076 & n13636 ;
  assign n13638 = n1227 | n13637 ;
  assign n13643 = n13642 ^ n13638 ^ 1'b0 ;
  assign n13644 = n5858 ^ n2685 ^ 1'b0 ;
  assign n13645 = ( n1487 & ~n1896 ) | ( n1487 & n2724 ) | ( ~n1896 & n2724 ) ;
  assign n13646 = n6463 | n13645 ;
  assign n13647 = n13646 ^ n6321 ^ 1'b0 ;
  assign n13648 = n1316 & n13647 ;
  assign n13649 = ( n490 & ~n8338 ) | ( n490 & n13648 ) | ( ~n8338 & n13648 ) ;
  assign n13650 = n10757 ^ n3581 ^ 1'b0 ;
  assign n13651 = n11543 ^ n8538 ^ 1'b0 ;
  assign n13652 = ~n5685 & n13651 ;
  assign n13653 = n13652 ^ n3508 ^ 1'b0 ;
  assign n13654 = ~n12627 & n13653 ;
  assign n13655 = n4495 ^ n4162 ^ 1'b0 ;
  assign n13656 = ~n5554 & n13655 ;
  assign n13657 = n8922 ^ n7712 ^ 1'b0 ;
  assign n13658 = n13657 ^ n9238 ^ 1'b0 ;
  assign n13659 = n5653 ^ x92 ^ 1'b0 ;
  assign n13660 = n8644 & n13659 ;
  assign n13661 = n13660 ^ n9600 ^ 1'b0 ;
  assign n13662 = n4097 & n13661 ;
  assign n13663 = n1636 ^ n1564 ^ 1'b0 ;
  assign n13664 = n13662 & ~n13663 ;
  assign n13665 = n827 & ~n3750 ;
  assign n13666 = n12469 | n13665 ;
  assign n13667 = n5575 | n13666 ;
  assign n13668 = n861 & n12206 ;
  assign n13669 = n13668 ^ n11196 ^ n861 ;
  assign n13670 = ~x210 & n4577 ;
  assign n13671 = n5809 & ~n13670 ;
  assign n13672 = n4081 & n13671 ;
  assign n13673 = ( n6519 & ~n7932 ) | ( n6519 & n11385 ) | ( ~n7932 & n11385 ) ;
  assign n13674 = n3088 & n8935 ;
  assign n13675 = n13674 ^ n8688 ^ 1'b0 ;
  assign n13676 = n9953 & ~n13675 ;
  assign n13677 = ~n9311 & n13676 ;
  assign n13678 = n11053 ^ n5303 ^ 1'b0 ;
  assign n13679 = n13678 ^ n6319 ^ 1'b0 ;
  assign n13680 = n9824 | n13017 ;
  assign n13681 = ( n1769 & ~n13679 ) | ( n1769 & n13680 ) | ( ~n13679 & n13680 ) ;
  assign n13682 = ( n329 & n4086 ) | ( n329 & n12849 ) | ( n4086 & n12849 ) ;
  assign n13683 = n9902 ^ n3336 ^ 1'b0 ;
  assign n13684 = n13682 & n13683 ;
  assign n13685 = n11653 ^ n2867 ^ x95 ;
  assign n13686 = ( ~n6948 & n7740 ) | ( ~n6948 & n13685 ) | ( n7740 & n13685 ) ;
  assign n13687 = n13686 ^ n1197 ^ 1'b0 ;
  assign n13688 = ~n4767 & n13687 ;
  assign n13689 = n7871 & ~n13688 ;
  assign n13690 = n3403 & ~n4031 ;
  assign n13691 = n13690 ^ n9787 ^ 1'b0 ;
  assign n13692 = n6720 | n7987 ;
  assign n13693 = n13692 ^ n3714 ^ 1'b0 ;
  assign n13694 = n9906 ^ n4989 ^ 1'b0 ;
  assign n13695 = n1260 & ~n1506 ;
  assign n13696 = ~n6096 & n13695 ;
  assign n13697 = n1522 & ~n13696 ;
  assign n13698 = ~x77 & n13697 ;
  assign n13699 = n13698 ^ n2189 ^ 1'b0 ;
  assign n13700 = n13694 & ~n13699 ;
  assign n13701 = n9542 ^ n5787 ^ 1'b0 ;
  assign n13702 = n7509 & n13701 ;
  assign n13703 = n13702 ^ n2672 ^ 1'b0 ;
  assign n13704 = n11753 | n13703 ;
  assign n13705 = n13700 & ~n13704 ;
  assign n13706 = ~n12433 & n13705 ;
  assign n13711 = n2458 ^ n1145 ^ 1'b0 ;
  assign n13712 = n13711 ^ n3875 ^ n1524 ;
  assign n13713 = n13712 ^ n10075 ^ 1'b0 ;
  assign n13714 = ~n11116 & n13713 ;
  assign n13707 = x97 | n421 ;
  assign n13708 = n13707 ^ n6960 ^ 1'b0 ;
  assign n13709 = x80 & n13708 ;
  assign n13710 = ~n839 & n13709 ;
  assign n13715 = n13714 ^ n13710 ^ 1'b0 ;
  assign n13716 = n8264 ^ n5744 ^ 1'b0 ;
  assign n13717 = ( n2494 & n3545 ) | ( n2494 & n9910 ) | ( n3545 & n9910 ) ;
  assign n13718 = ( n2977 & n13716 ) | ( n2977 & n13717 ) | ( n13716 & n13717 ) ;
  assign n13732 = n7366 ^ n2229 ^ 1'b0 ;
  assign n13733 = n997 & n13732 ;
  assign n13724 = n1979 & n2279 ;
  assign n13725 = n13724 ^ n451 ^ 1'b0 ;
  assign n13726 = x158 | n13725 ;
  assign n13727 = n1768 & n8638 ;
  assign n13728 = n2680 & n13727 ;
  assign n13729 = ( n3952 & ~n13726 ) | ( n3952 & n13728 ) | ( ~n13726 & n13728 ) ;
  assign n13723 = x77 & ~n8911 ;
  assign n13730 = n13729 ^ n13723 ^ 1'b0 ;
  assign n13731 = n7661 | n13730 ;
  assign n13720 = ~n2349 & n8340 ;
  assign n13721 = n13720 ^ n9314 ^ 1'b0 ;
  assign n13719 = ~n5041 & n7915 ;
  assign n13722 = n13721 ^ n13719 ^ 1'b0 ;
  assign n13734 = n13733 ^ n13731 ^ n13722 ;
  assign n13735 = ( n4405 & n6613 ) | ( n4405 & ~n6640 ) | ( n6613 & ~n6640 ) ;
  assign n13736 = n11104 & ~n13735 ;
  assign n13737 = n10665 & ~n13736 ;
  assign n13738 = ~n6130 & n13737 ;
  assign n13742 = n4875 ^ n509 ^ 1'b0 ;
  assign n13743 = n4496 & n13742 ;
  assign n13744 = n13743 ^ n3800 ^ 1'b0 ;
  assign n13739 = ~n4492 & n4598 ;
  assign n13740 = n13739 ^ n9869 ^ 1'b0 ;
  assign n13741 = n13740 ^ n1231 ^ 1'b0 ;
  assign n13745 = n13744 ^ n13741 ^ 1'b0 ;
  assign n13746 = n3185 & ~n5837 ;
  assign n13747 = ~n1489 & n13746 ;
  assign n13748 = n8952 ^ n4277 ^ n4203 ;
  assign n13749 = n6080 & ~n13748 ;
  assign n13750 = n13749 ^ n7084 ^ 1'b0 ;
  assign n13751 = n13747 | n13750 ;
  assign n13752 = n3986 | n8468 ;
  assign n13753 = n13752 ^ n5728 ^ 1'b0 ;
  assign n13754 = n3275 | n7663 ;
  assign n13755 = n8235 & n10854 ;
  assign n13756 = n13755 ^ n3322 ^ 1'b0 ;
  assign n13757 = n13756 ^ n5746 ^ n3308 ;
  assign n13758 = n13757 ^ n656 ^ 1'b0 ;
  assign n13759 = n10356 ^ n2133 ^ 1'b0 ;
  assign n13760 = n3932 & ~n8784 ;
  assign n13761 = ~n1605 & n13760 ;
  assign n13762 = ~n410 & n13761 ;
  assign n13763 = ( n1083 & n6068 ) | ( n1083 & n8660 ) | ( n6068 & n8660 ) ;
  assign n13764 = n4979 | n5565 ;
  assign n13765 = x37 | n9143 ;
  assign n13766 = n2396 | n13765 ;
  assign n13767 = n13766 ^ n5975 ^ 1'b0 ;
  assign n13768 = ~n13764 & n13767 ;
  assign n13769 = n7014 ^ n2878 ^ 1'b0 ;
  assign n13770 = n13768 & ~n13769 ;
  assign n13771 = n10804 ^ n8422 ^ 1'b0 ;
  assign n13772 = n292 & ~n4836 ;
  assign n13773 = n13771 & n13772 ;
  assign n13774 = x155 & ~x198 ;
  assign n13775 = ( n3032 & n4477 ) | ( n3032 & ~n13774 ) | ( n4477 & ~n13774 ) ;
  assign n13776 = n13775 ^ n8094 ^ 1'b0 ;
  assign n13777 = n12158 ^ n4498 ^ 1'b0 ;
  assign n13778 = ~n2075 & n13777 ;
  assign n13779 = n13778 ^ n3210 ^ 1'b0 ;
  assign n13780 = n13779 ^ n11758 ^ 1'b0 ;
  assign n13781 = n9634 | n13780 ;
  assign n13782 = x164 & n1453 ;
  assign n13783 = ~n3273 & n13782 ;
  assign n13784 = ~n5148 & n12617 ;
  assign n13785 = n13783 & n13784 ;
  assign n13786 = n7145 | n8469 ;
  assign n13787 = n13786 ^ n11535 ^ 1'b0 ;
  assign n13788 = ~n13785 & n13787 ;
  assign n13789 = n2955 | n10949 ;
  assign n13790 = n13789 ^ n6899 ^ 1'b0 ;
  assign n13791 = n5646 & n13790 ;
  assign n13792 = n13791 ^ n2577 ^ n1521 ;
  assign n13793 = ~n1682 & n3609 ;
  assign n13794 = n4130 & n5982 ;
  assign n13795 = n13794 ^ n6403 ^ 1'b0 ;
  assign n13796 = n7214 & ~n13795 ;
  assign n13798 = n5339 ^ n3354 ^ n2886 ;
  assign n13797 = n3856 ^ n2955 ^ 1'b0 ;
  assign n13799 = n13798 ^ n13797 ^ 1'b0 ;
  assign n13800 = n12078 | n13799 ;
  assign n13801 = n4580 ^ n2555 ^ 1'b0 ;
  assign n13802 = n6989 ^ n3138 ^ 1'b0 ;
  assign n13803 = n8553 & n13802 ;
  assign n13807 = n6015 ^ n3810 ^ n1508 ;
  assign n13804 = n6260 | n12627 ;
  assign n13805 = n1253 & ~n9396 ;
  assign n13806 = ~n13804 & n13805 ;
  assign n13808 = n13807 ^ n13806 ^ n8043 ;
  assign n13809 = n1862 & n6524 ;
  assign n13810 = n13809 ^ n7741 ^ n2174 ;
  assign n13811 = n6314 & n10127 ;
  assign n13812 = n13811 ^ n6071 ^ 1'b0 ;
  assign n13813 = n3816 | n10205 ;
  assign n13814 = n1173 & ~n3004 ;
  assign n13815 = x46 & ~n2997 ;
  assign n13816 = ~n13814 & n13815 ;
  assign n13817 = n3445 ^ n823 ^ 1'b0 ;
  assign n13818 = ~n1727 & n13817 ;
  assign n13819 = n593 & n13818 ;
  assign n13820 = ~n7839 & n13819 ;
  assign n13821 = n2243 ^ n462 ^ 1'b0 ;
  assign n13822 = n13821 ^ x38 ^ 1'b0 ;
  assign n13823 = ~n1433 & n3546 ;
  assign n13824 = ~x85 & n6776 ;
  assign n13825 = n1462 & ~n13824 ;
  assign n13826 = n13825 ^ n2783 ^ 1'b0 ;
  assign n13832 = x201 & ~n5151 ;
  assign n13833 = n13832 ^ n6334 ^ 1'b0 ;
  assign n13834 = n11105 & n13833 ;
  assign n13835 = n8909 & n13834 ;
  assign n13836 = n6046 ^ n4220 ^ 1'b0 ;
  assign n13837 = n8941 & n13836 ;
  assign n13838 = ~n3755 & n13837 ;
  assign n13839 = n13835 & n13838 ;
  assign n13829 = x127 & n7825 ;
  assign n13830 = n13829 ^ n2859 ^ 1'b0 ;
  assign n13827 = n5436 & n6660 ;
  assign n13828 = n13827 ^ n11902 ^ 1'b0 ;
  assign n13831 = n13830 ^ n13828 ^ 1'b0 ;
  assign n13840 = n13839 ^ n13831 ^ 1'b0 ;
  assign n13841 = n7293 & n13840 ;
  assign n13842 = n13572 ^ n1106 ^ 1'b0 ;
  assign n13843 = n5758 & n7370 ;
  assign n13844 = x120 & n13843 ;
  assign n13845 = n386 & n8626 ;
  assign n13846 = ~n10075 & n13845 ;
  assign n13847 = ( n476 & n1729 ) | ( n476 & n1805 ) | ( n1729 & n1805 ) ;
  assign n13848 = ( n3512 & ~n7382 ) | ( n3512 & n9624 ) | ( ~n7382 & n9624 ) ;
  assign n13849 = ~n9209 & n13848 ;
  assign n13850 = n5017 & n13849 ;
  assign n13851 = n1910 & ~n13850 ;
  assign n13852 = n6992 & n13851 ;
  assign n13853 = n13847 & n13852 ;
  assign n13854 = ( x113 & n13846 ) | ( x113 & n13853 ) | ( n13846 & n13853 ) ;
  assign n13859 = n4070 ^ n673 ^ 1'b0 ;
  assign n13860 = n2247 & n13859 ;
  assign n13861 = ( n1155 & n1592 ) | ( n1155 & ~n13860 ) | ( n1592 & ~n13860 ) ;
  assign n13855 = n3363 ^ n3338 ^ x177 ;
  assign n13856 = n4924 & ~n6415 ;
  assign n13857 = ( n5918 & ~n13855 ) | ( n5918 & n13856 ) | ( ~n13855 & n13856 ) ;
  assign n13858 = ~n2919 & n13857 ;
  assign n13862 = n13861 ^ n13858 ^ n12361 ;
  assign n13866 = n11777 ^ n1380 ^ 1'b0 ;
  assign n13863 = n9360 ^ n6472 ^ n394 ;
  assign n13864 = n13863 ^ n4932 ^ 1'b0 ;
  assign n13865 = n5699 & ~n13864 ;
  assign n13867 = n13866 ^ n13865 ^ 1'b0 ;
  assign n13868 = n5844 & n10565 ;
  assign n13869 = n13868 ^ n9841 ^ 1'b0 ;
  assign n13871 = n3105 & ~n4454 ;
  assign n13872 = ~x200 & n13871 ;
  assign n13873 = ~n13678 & n13872 ;
  assign n13874 = x170 & n13873 ;
  assign n13870 = n1969 & ~n7364 ;
  assign n13875 = n13874 ^ n13870 ^ 1'b0 ;
  assign n13876 = n10416 ^ n6945 ^ n5042 ;
  assign n13877 = n13876 ^ n1296 ^ 1'b0 ;
  assign n13878 = n7140 ^ n4755 ^ 1'b0 ;
  assign n13879 = n13877 & ~n13878 ;
  assign n13880 = ~n1103 & n3899 ;
  assign n13881 = ( ~n4011 & n13322 ) | ( ~n4011 & n13880 ) | ( n13322 & n13880 ) ;
  assign n13882 = n13881 ^ n3175 ^ 1'b0 ;
  assign n13883 = n1185 & ~n13882 ;
  assign n13884 = n11045 ^ n3615 ^ 1'b0 ;
  assign n13885 = n12885 & ~n13884 ;
  assign n13886 = n13885 ^ n13824 ^ n11789 ;
  assign n13887 = n9347 & n10584 ;
  assign n13888 = n4589 ^ n3878 ^ 1'b0 ;
  assign n13889 = n673 & ~n13888 ;
  assign n13890 = ~n567 & n13889 ;
  assign n13891 = n10504 ^ n797 ^ 1'b0 ;
  assign n13892 = n12004 ^ n9652 ^ 1'b0 ;
  assign n13893 = n522 | n4651 ;
  assign n13894 = n13893 ^ n6607 ^ 1'b0 ;
  assign n13895 = n1593 & n12743 ;
  assign n13896 = n5842 ^ n4257 ^ 1'b0 ;
  assign n13897 = ~n5526 & n13896 ;
  assign n13898 = n10063 ^ n2312 ^ 1'b0 ;
  assign n13899 = n10644 & n13898 ;
  assign n13900 = n610 & n5425 ;
  assign n13901 = n3636 & n13900 ;
  assign n13902 = ( n8051 & n10322 ) | ( n8051 & n13901 ) | ( n10322 & n13901 ) ;
  assign n13903 = n10881 & ~n11851 ;
  assign n13904 = n7100 & n8340 ;
  assign n13905 = n12396 & n13904 ;
  assign n13906 = n5909 ^ n573 ^ 1'b0 ;
  assign n13907 = ~n651 & n13906 ;
  assign n13908 = n4086 & ~n8984 ;
  assign n13909 = n5828 & n13908 ;
  assign n13910 = ( ~n967 & n9331 ) | ( ~n967 & n13909 ) | ( n9331 & n13909 ) ;
  assign n13911 = ( n2568 & n8890 ) | ( n2568 & ~n11941 ) | ( n8890 & ~n11941 ) ;
  assign n13912 = n6988 | n13911 ;
  assign n13913 = n13912 ^ n1074 ^ 1'b0 ;
  assign n13914 = ~n4441 & n11572 ;
  assign n13915 = ~n7509 & n13914 ;
  assign n13916 = n4138 | n4282 ;
  assign n13917 = n13916 ^ n4408 ^ 1'b0 ;
  assign n13918 = ~n10889 & n13917 ;
  assign n13920 = n11880 ^ n10262 ^ x104 ;
  assign n13919 = x129 & n1812 ;
  assign n13921 = n13920 ^ n13919 ^ 1'b0 ;
  assign n13922 = n13736 ^ n3756 ^ 1'b0 ;
  assign n13923 = ( ~x18 & n3510 ) | ( ~x18 & n9682 ) | ( n3510 & n9682 ) ;
  assign n13924 = n6528 | n8548 ;
  assign n13925 = n13924 ^ n5357 ^ 1'b0 ;
  assign n13926 = n13925 ^ n857 ^ 1'b0 ;
  assign n13927 = n6319 & n6808 ;
  assign n13928 = ~n6188 & n13927 ;
  assign n13931 = ~n2914 & n11851 ;
  assign n13929 = x150 & ~n4280 ;
  assign n13930 = ~n7840 & n13929 ;
  assign n13932 = n13931 ^ n13930 ^ 1'b0 ;
  assign n13933 = n13928 | n13932 ;
  assign n13934 = n6693 ^ n5075 ^ 1'b0 ;
  assign n13935 = n13933 | n13934 ;
  assign n13936 = n13521 ^ x123 ^ 1'b0 ;
  assign n13937 = n13935 | n13936 ;
  assign n13938 = n8896 ^ n6640 ^ 1'b0 ;
  assign n13939 = n13449 & n13938 ;
  assign n13940 = ~n5225 & n13939 ;
  assign n13941 = ~n3056 & n4797 ;
  assign n13942 = n10076 & n13941 ;
  assign n13943 = ( n3371 & ~n12081 ) | ( n3371 & n13942 ) | ( ~n12081 & n13942 ) ;
  assign n13944 = n10660 & n13665 ;
  assign n13945 = n13944 ^ n4879 ^ 1'b0 ;
  assign n13946 = n13716 & ~n13945 ;
  assign n13947 = n5083 ^ n2943 ^ n1671 ;
  assign n13948 = n12239 & ~n13116 ;
  assign n13949 = n13947 & n13948 ;
  assign n13950 = n1521 ^ n1200 ^ 1'b0 ;
  assign n13951 = n6916 & n13950 ;
  assign n13952 = n557 & ~n979 ;
  assign n13953 = n5690 ^ n4519 ^ 1'b0 ;
  assign n13954 = n881 | n13953 ;
  assign n13955 = n13952 | n13954 ;
  assign n13956 = n13955 ^ n10017 ^ 1'b0 ;
  assign n13958 = n2634 & ~n3413 ;
  assign n13959 = n13958 ^ n935 ^ 1'b0 ;
  assign n13960 = ~n2017 & n13959 ;
  assign n13957 = n5789 & n9444 ;
  assign n13961 = n13960 ^ n13957 ^ n9181 ;
  assign n13962 = n2362 & n6972 ;
  assign n13963 = n12812 | n13824 ;
  assign n13964 = n13962 | n13963 ;
  assign n13969 = n460 & ~n1602 ;
  assign n13970 = n13969 ^ n3316 ^ 1'b0 ;
  assign n13971 = n13970 ^ n11187 ^ 1'b0 ;
  assign n13972 = n1064 & ~n13971 ;
  assign n13966 = n2205 | n3473 ;
  assign n13967 = n691 | n13966 ;
  assign n13968 = n13967 ^ n9861 ^ n1696 ;
  assign n13973 = n13972 ^ n13968 ^ n616 ;
  assign n13974 = ( n1429 & n2989 ) | ( n1429 & ~n13973 ) | ( n2989 & ~n13973 ) ;
  assign n13975 = ( n12275 & n12738 ) | ( n12275 & n13974 ) | ( n12738 & n13974 ) ;
  assign n13965 = n1413 & ~n10167 ;
  assign n13976 = n13975 ^ n13965 ^ 1'b0 ;
  assign n13981 = ( x205 & ~n731 ) | ( x205 & n3100 ) | ( ~n731 & n3100 ) ;
  assign n13982 = n4574 ^ n3764 ^ 1'b0 ;
  assign n13983 = n13981 & ~n13982 ;
  assign n13984 = n13983 ^ n7839 ^ 1'b0 ;
  assign n13985 = n5762 | n13984 ;
  assign n13986 = n13985 ^ n5923 ^ 1'b0 ;
  assign n13977 = ( n3990 & n4052 ) | ( n3990 & ~n9050 ) | ( n4052 & ~n9050 ) ;
  assign n13978 = ~n6253 & n13977 ;
  assign n13979 = n2901 & n13978 ;
  assign n13980 = n6452 & ~n13979 ;
  assign n13987 = n13986 ^ n13980 ^ 1'b0 ;
  assign n13988 = ~n6588 & n7616 ;
  assign n13989 = n1360 | n4019 ;
  assign n13990 = n13988 | n13989 ;
  assign n13991 = ~n11118 & n13990 ;
  assign n13992 = n1880 & n13991 ;
  assign n13993 = n13017 | n13984 ;
  assign n13994 = n1799 ^ n1751 ^ 1'b0 ;
  assign n13995 = n13994 ^ n428 ^ 1'b0 ;
  assign n13996 = n295 & ~n13995 ;
  assign n13997 = ~n9664 & n13996 ;
  assign n13998 = n13997 ^ n9246 ^ n4833 ;
  assign n13999 = n13512 ^ n9188 ^ n6211 ;
  assign n14000 = n12749 ^ n2879 ^ n1115 ;
  assign n14004 = x147 & n4219 ;
  assign n14002 = ~n3808 & n8213 ;
  assign n14001 = n4327 & n4733 ;
  assign n14003 = n14002 ^ n14001 ^ 1'b0 ;
  assign n14005 = n14004 ^ n14003 ^ 1'b0 ;
  assign n14006 = n4766 | n14005 ;
  assign n14007 = n14000 & ~n14006 ;
  assign n14008 = n6679 & ~n10543 ;
  assign n14009 = ~n11513 & n14008 ;
  assign n14010 = n12758 & n14009 ;
  assign n14011 = n8578 ^ n1624 ^ n777 ;
  assign n14012 = n7629 | n14011 ;
  assign n14016 = n6270 & ~n7246 ;
  assign n14013 = ( n1150 & ~n2516 ) | ( n1150 & n6420 ) | ( ~n2516 & n6420 ) ;
  assign n14014 = n14013 ^ n848 ^ 1'b0 ;
  assign n14015 = ~n4067 & n14014 ;
  assign n14017 = n14016 ^ n14015 ^ 1'b0 ;
  assign n14018 = n6027 ^ n2294 ^ 1'b0 ;
  assign n14019 = n442 & ~n14018 ;
  assign n14020 = ( n305 & n10045 ) | ( n305 & n13360 ) | ( n10045 & n13360 ) ;
  assign n14021 = n3410 ^ n2786 ^ 1'b0 ;
  assign n14022 = ( ~n1000 & n3117 ) | ( ~n1000 & n14021 ) | ( n3117 & n14021 ) ;
  assign n14023 = n14022 ^ n6783 ^ n6320 ;
  assign n14024 = n11225 & ~n14023 ;
  assign n14025 = n14020 & n14024 ;
  assign n14026 = ~n3640 & n9787 ;
  assign n14027 = ( n2989 & n5223 ) | ( n2989 & n14026 ) | ( n5223 & n14026 ) ;
  assign n14028 = ~n3498 & n13674 ;
  assign n14029 = ~n7404 & n14028 ;
  assign n14030 = n14029 ^ n4861 ^ 1'b0 ;
  assign n14032 = n5985 ^ n1813 ^ x250 ;
  assign n14033 = ~n1155 & n14032 ;
  assign n14031 = ( ~n3231 & n3659 ) | ( ~n3231 & n4567 ) | ( n3659 & n4567 ) ;
  assign n14034 = n14033 ^ n14031 ^ n8299 ;
  assign n14035 = ( n1202 & n3024 ) | ( n1202 & n13640 ) | ( n3024 & n13640 ) ;
  assign n14036 = n14035 ^ n12550 ^ 1'b0 ;
  assign n14037 = n4498 & ~n14036 ;
  assign n14038 = n2823 & ~n10462 ;
  assign n14039 = n14038 ^ n536 ^ 1'b0 ;
  assign n14040 = n5681 & n14039 ;
  assign n14041 = n3806 | n14040 ;
  assign n14042 = n8114 | n12479 ;
  assign n14043 = n14042 ^ n5472 ^ 1'b0 ;
  assign n14044 = ( ~x206 & n433 ) | ( ~x206 & n4236 ) | ( n433 & n4236 ) ;
  assign n14045 = ~n587 & n3543 ;
  assign n14046 = n13135 ^ n4614 ^ n2494 ;
  assign n14047 = n2425 & ~n3358 ;
  assign n14048 = n1597 & n14047 ;
  assign n14049 = n14048 ^ n1832 ^ n992 ;
  assign n14050 = n14049 ^ n1701 ^ 1'b0 ;
  assign n14051 = n8149 | n14050 ;
  assign n14052 = n14051 ^ n2997 ^ 1'b0 ;
  assign n14055 = n851 | n1744 ;
  assign n14053 = n4251 & n5014 ;
  assign n14054 = n14053 ^ x21 ^ 1'b0 ;
  assign n14056 = n14055 ^ n14054 ^ 1'b0 ;
  assign n14057 = n3771 & n12026 ;
  assign n14058 = n814 | n14057 ;
  assign n14059 = n4766 & n8444 ;
  assign n14060 = n14059 ^ n3578 ^ 1'b0 ;
  assign n14061 = n540 | n14060 ;
  assign n14062 = x66 & ~n5254 ;
  assign n14063 = n2538 & n14062 ;
  assign n14064 = n2702 | n14063 ;
  assign n14065 = n7580 ^ n7549 ^ n1401 ;
  assign n14066 = n13887 ^ n9577 ^ 1'b0 ;
  assign n14067 = n14065 & n14066 ;
  assign n14068 = n10392 ^ n5441 ^ n5058 ;
  assign n14069 = ~n7309 & n10963 ;
  assign n14070 = ~n440 & n6392 ;
  assign n14071 = n14070 ^ n9944 ^ n4128 ;
  assign n14072 = ~n7508 & n14071 ;
  assign n14073 = n14069 & n14072 ;
  assign n14074 = n14068 & ~n14073 ;
  assign n14075 = n5680 & n14074 ;
  assign n14076 = ( n3447 & n7006 ) | ( n3447 & ~n8263 ) | ( n7006 & ~n8263 ) ;
  assign n14077 = n14076 ^ n6088 ^ 1'b0 ;
  assign n14078 = n11451 ^ n1331 ^ 1'b0 ;
  assign n14079 = n6358 & n8051 ;
  assign n14080 = n3442 | n14079 ;
  assign n14081 = n14080 ^ n6322 ^ 1'b0 ;
  assign n14082 = n6965 & n8277 ;
  assign n14083 = n14082 ^ n7723 ^ 1'b0 ;
  assign n14084 = n11449 ^ n659 ^ 1'b0 ;
  assign n14085 = n8026 | n14084 ;
  assign n14086 = n4118 & ~n8653 ;
  assign n14087 = n4816 ^ n1158 ^ 1'b0 ;
  assign n14088 = n3781 & n14087 ;
  assign n14089 = n13483 ^ n3490 ^ n1671 ;
  assign n14090 = x48 & ~n8193 ;
  assign n14091 = ~n1224 & n14090 ;
  assign n14092 = n9497 ^ n7044 ^ 1'b0 ;
  assign n14093 = ~n2453 & n14092 ;
  assign n14094 = ( n1877 & ~n10595 ) | ( n1877 & n14093 ) | ( ~n10595 & n14093 ) ;
  assign n14095 = ( ~n4451 & n14091 ) | ( ~n4451 & n14094 ) | ( n14091 & n14094 ) ;
  assign n14096 = ( n10814 & n12967 ) | ( n10814 & ~n14095 ) | ( n12967 & ~n14095 ) ;
  assign n14097 = ( n3830 & ~n7238 ) | ( n3830 & n8507 ) | ( ~n7238 & n8507 ) ;
  assign n14098 = ~n6473 & n14097 ;
  assign n14099 = n8492 & n14098 ;
  assign n14100 = ~n7883 & n14099 ;
  assign n14101 = n8675 ^ x49 ^ 1'b0 ;
  assign n14102 = n14100 & n14101 ;
  assign n14103 = n9391 | n11388 ;
  assign n14104 = ( n2677 & n6433 ) | ( n2677 & n14103 ) | ( n6433 & n14103 ) ;
  assign n14105 = n4890 | n14104 ;
  assign n14106 = n10101 ^ n9761 ^ 1'b0 ;
  assign n14107 = ~n14105 & n14106 ;
  assign n14108 = n531 & ~n12458 ;
  assign n14109 = n14108 ^ n2174 ^ 1'b0 ;
  assign n14110 = n3046 | n14109 ;
  assign n14111 = n6857 & n12264 ;
  assign n14112 = n14110 & n14111 ;
  assign n14113 = n10042 & ~n14112 ;
  assign n14115 = n2266 & ~n6875 ;
  assign n14116 = n14115 ^ n8924 ^ 1'b0 ;
  assign n14114 = n2978 & n7176 ;
  assign n14117 = n14116 ^ n14114 ^ 1'b0 ;
  assign n14118 = n13000 ^ n11753 ^ n4317 ;
  assign n14119 = ( n1166 & n12060 ) | ( n1166 & ~n14118 ) | ( n12060 & ~n14118 ) ;
  assign n14121 = n3328 & ~n9088 ;
  assign n14120 = n5528 & n12003 ;
  assign n14122 = n14121 ^ n14120 ^ n424 ;
  assign n14125 = ( n425 & ~n2354 ) | ( n425 & n6933 ) | ( ~n2354 & n6933 ) ;
  assign n14123 = n9092 ^ n584 ^ 1'b0 ;
  assign n14124 = ~n5842 & n14123 ;
  assign n14126 = n14125 ^ n14124 ^ n8620 ;
  assign n14127 = n11257 | n14126 ;
  assign n14128 = n2841 | n12655 ;
  assign n14129 = n14128 ^ n6234 ^ 1'b0 ;
  assign n14130 = ~n7067 & n14129 ;
  assign n14131 = n1702 ^ n493 ^ 1'b0 ;
  assign n14132 = n14130 & n14131 ;
  assign n14133 = ~n13688 & n14132 ;
  assign n14135 = n5742 ^ n1439 ^ 1'b0 ;
  assign n14134 = ( n3759 & ~n3932 ) | ( n3759 & n5291 ) | ( ~n3932 & n5291 ) ;
  assign n14136 = n14135 ^ n14134 ^ n10454 ;
  assign n14137 = n14136 ^ n3774 ^ 1'b0 ;
  assign n14138 = ( ~n1301 & n5685 ) | ( ~n1301 & n13977 ) | ( n5685 & n13977 ) ;
  assign n14139 = ( ~n460 & n1007 ) | ( ~n460 & n3188 ) | ( n1007 & n3188 ) ;
  assign n14140 = ( n4924 & n14138 ) | ( n4924 & n14139 ) | ( n14138 & n14139 ) ;
  assign n14142 = n3439 ^ n2603 ^ 1'b0 ;
  assign n14143 = n1827 | n1987 ;
  assign n14144 = n14142 | n14143 ;
  assign n14145 = n1980 | n14144 ;
  assign n14141 = ~n7777 & n8807 ;
  assign n14146 = n14145 ^ n14141 ^ 1'b0 ;
  assign n14147 = n5643 & n9483 ;
  assign n14148 = ~n4191 & n7963 ;
  assign n14149 = n917 | n2323 ;
  assign n14150 = n9010 | n14149 ;
  assign n14151 = ( ~n3260 & n14148 ) | ( ~n3260 & n14150 ) | ( n14148 & n14150 ) ;
  assign n14152 = n13968 ^ n11898 ^ 1'b0 ;
  assign n14153 = n14151 & n14152 ;
  assign n14154 = n14153 ^ n10852 ^ 1'b0 ;
  assign n14155 = n14147 & ~n14154 ;
  assign n14156 = n1061 & n5807 ;
  assign n14157 = n3196 & ~n12431 ;
  assign n14158 = n13226 ^ n3691 ^ x54 ;
  assign n14159 = ( n11108 & n14157 ) | ( n11108 & ~n14158 ) | ( n14157 & ~n14158 ) ;
  assign n14160 = n9264 ^ n7998 ^ 1'b0 ;
  assign n14161 = ~n14159 & n14160 ;
  assign n14162 = n3140 & ~n12021 ;
  assign n14163 = n14162 ^ n10106 ^ 1'b0 ;
  assign n14164 = n12546 ^ n5909 ^ n3961 ;
  assign n14165 = n5433 ^ n1006 ^ 1'b0 ;
  assign n14166 = n14164 & ~n14165 ;
  assign n14167 = n10114 ^ n9258 ^ 1'b0 ;
  assign n14168 = n12488 | n14167 ;
  assign n14169 = n5441 ^ n2341 ^ 1'b0 ;
  assign n14170 = n6086 ^ n1962 ^ 1'b0 ;
  assign n14171 = ( x38 & n2720 ) | ( x38 & n4357 ) | ( n2720 & n4357 ) ;
  assign n14172 = ( n11320 & n14170 ) | ( n11320 & n14171 ) | ( n14170 & n14171 ) ;
  assign n14173 = ~n13818 & n14131 ;
  assign n14174 = n11401 ^ n5622 ^ 1'b0 ;
  assign n14175 = n3786 ^ n3532 ^ 1'b0 ;
  assign n14176 = n7754 & ~n14175 ;
  assign n14177 = n561 & ~n5619 ;
  assign n14178 = n1182 & ~n8063 ;
  assign n14179 = n12757 & n14178 ;
  assign n14180 = n13467 ^ n6062 ^ 1'b0 ;
  assign n14181 = n7821 & n13170 ;
  assign n14182 = ~n11342 & n14181 ;
  assign n14183 = ~n8412 & n13803 ;
  assign n14184 = n495 & n8862 ;
  assign n14185 = n5905 & n14184 ;
  assign n14186 = ( ~n3464 & n9077 ) | ( ~n3464 & n14185 ) | ( n9077 & n14185 ) ;
  assign n14187 = n14186 ^ n1576 ^ 1'b0 ;
  assign n14188 = n5134 & ~n14187 ;
  assign n14189 = n12657 ^ n3729 ^ n2589 ;
  assign n14190 = n14189 ^ n597 ^ 1'b0 ;
  assign n14191 = n8772 & ~n14190 ;
  assign n14192 = n8621 & ~n10134 ;
  assign n14193 = ~n3242 & n14192 ;
  assign n14194 = n14193 ^ n5615 ^ 1'b0 ;
  assign n14195 = n14191 & ~n14194 ;
  assign n14196 = n11765 & n14195 ;
  assign n14197 = n1013 | n14196 ;
  assign n14198 = n14197 ^ n10793 ^ 1'b0 ;
  assign n14199 = n2645 & ~n9501 ;
  assign n14200 = n13255 ^ x155 ^ 1'b0 ;
  assign n14201 = n10517 & n14200 ;
  assign n14202 = ~n3312 & n7619 ;
  assign n14203 = n733 & n14202 ;
  assign n14204 = n2912 | n14203 ;
  assign n14205 = ~n4751 & n11184 ;
  assign n14206 = n3052 ^ n2212 ^ 1'b0 ;
  assign n14207 = n5827 ^ x109 ^ 1'b0 ;
  assign n14208 = n12466 | n14207 ;
  assign n14209 = ~n1327 & n14208 ;
  assign n14210 = ~n1298 & n14209 ;
  assign n14211 = n14206 & n14210 ;
  assign n14212 = n8102 & n14211 ;
  assign n14213 = n7860 ^ n6627 ^ n3952 ;
  assign n14214 = n4417 ^ n4115 ^ 1'b0 ;
  assign n14215 = ~n5480 & n14214 ;
  assign n14216 = ( ~n1965 & n2831 ) | ( ~n1965 & n6065 ) | ( n2831 & n6065 ) ;
  assign n14217 = n14216 ^ n8637 ^ 1'b0 ;
  assign n14218 = ( n260 & n14215 ) | ( n260 & n14217 ) | ( n14215 & n14217 ) ;
  assign n14219 = ~n1018 & n14218 ;
  assign n14220 = n2219 ^ n1160 ^ 1'b0 ;
  assign n14221 = n5787 & n14220 ;
  assign n14222 = n8496 & n10646 ;
  assign n14223 = ~n14221 & n14222 ;
  assign n14224 = n5710 ^ n2440 ^ n333 ;
  assign n14225 = ( n485 & n6523 ) | ( n485 & ~n14224 ) | ( n6523 & ~n14224 ) ;
  assign n14226 = n9111 ^ n2541 ^ 1'b0 ;
  assign n14227 = n14226 ^ n12360 ^ n6868 ;
  assign n14228 = ( ~n2005 & n4577 ) | ( ~n2005 & n10367 ) | ( n4577 & n10367 ) ;
  assign n14229 = n1023 & n14228 ;
  assign n14230 = n14229 ^ n1527 ^ 1'b0 ;
  assign n14231 = n269 | n6389 ;
  assign n14232 = n14230 & ~n14231 ;
  assign n14235 = n6919 ^ n271 ^ 1'b0 ;
  assign n14233 = n2356 ^ n2253 ^ 1'b0 ;
  assign n14234 = n2121 & n14233 ;
  assign n14236 = n14235 ^ n14234 ^ n13452 ;
  assign n14237 = ( n6141 & n7855 ) | ( n6141 & ~n14236 ) | ( n7855 & ~n14236 ) ;
  assign n14238 = ~n500 & n6585 ;
  assign n14239 = n14238 ^ n6842 ^ 1'b0 ;
  assign n14240 = ~n14237 & n14239 ;
  assign n14241 = n14240 ^ n3999 ^ 1'b0 ;
  assign n14242 = ( ~n485 & n4416 ) | ( ~n485 & n11992 ) | ( n4416 & n11992 ) ;
  assign n14243 = n6389 & ~n8794 ;
  assign n14244 = ~n832 & n14243 ;
  assign n14245 = n12521 ^ n1450 ^ 1'b0 ;
  assign n14246 = ~n5277 & n14245 ;
  assign n14247 = ~n9342 & n14246 ;
  assign n14248 = ~n14244 & n14247 ;
  assign n14249 = n3237 & ~n4293 ;
  assign n14250 = ~x194 & n14249 ;
  assign n14251 = n14250 ^ n13598 ^ n3288 ;
  assign n14252 = n13342 ^ n8039 ^ 1'b0 ;
  assign n14253 = n10147 ^ n9287 ^ n3176 ;
  assign n14254 = n8676 & ~n13545 ;
  assign n14255 = n14254 ^ n3261 ^ 1'b0 ;
  assign n14256 = n12260 | n13467 ;
  assign n14257 = n2339 | n14256 ;
  assign n14258 = n14257 ^ n989 ^ 1'b0 ;
  assign n14259 = n9158 | n14258 ;
  assign n14260 = n1434 ^ n483 ^ 1'b0 ;
  assign n14262 = n4150 ^ x189 ^ 1'b0 ;
  assign n14261 = ~n2071 & n2146 ;
  assign n14263 = n14262 ^ n14261 ^ 1'b0 ;
  assign n14264 = n5391 & ~n14263 ;
  assign n14265 = ( n3173 & n3947 ) | ( n3173 & ~n11583 ) | ( n3947 & ~n11583 ) ;
  assign n14266 = n2802 ^ n1705 ^ 1'b0 ;
  assign n14267 = n2639 & n8967 ;
  assign n14268 = n14267 ^ n1467 ^ 1'b0 ;
  assign n14269 = n2301 & ~n7545 ;
  assign n14270 = n10531 & n14269 ;
  assign n14271 = n4514 & n14270 ;
  assign n14272 = n2133 | n2998 ;
  assign n14273 = n5556 & ~n14272 ;
  assign n14274 = ( n798 & ~n1329 ) | ( n798 & n3099 ) | ( ~n1329 & n3099 ) ;
  assign n14275 = ( n1199 & n4317 ) | ( n1199 & n14274 ) | ( n4317 & n14274 ) ;
  assign n14276 = n14275 ^ n5102 ^ x82 ;
  assign n14277 = ( n1018 & n14273 ) | ( n1018 & ~n14276 ) | ( n14273 & ~n14276 ) ;
  assign n14278 = n14271 | n14277 ;
  assign n14279 = n14278 ^ n2748 ^ 1'b0 ;
  assign n14280 = ~n756 & n1671 ;
  assign n14281 = ~n12694 & n14280 ;
  assign n14282 = n8578 ^ n7160 ^ n2038 ;
  assign n14283 = n3535 ^ n1636 ^ x177 ;
  assign n14284 = ~n1585 & n7956 ;
  assign n14285 = n14283 & n14284 ;
  assign n14286 = ~n5053 & n8794 ;
  assign n14287 = n14286 ^ n11412 ^ 1'b0 ;
  assign n14288 = n14285 | n14287 ;
  assign n14289 = n10449 ^ n3542 ^ 1'b0 ;
  assign n14290 = n14289 ^ x203 ^ 1'b0 ;
  assign n14291 = n807 & ~n14290 ;
  assign n14292 = n2759 ^ n1368 ^ 1'b0 ;
  assign n14293 = n6307 | n14292 ;
  assign n14294 = n861 | n14293 ;
  assign n14295 = n4253 ^ n3341 ^ x38 ;
  assign n14296 = n14295 ^ n4529 ^ 1'b0 ;
  assign n14297 = n14294 & n14296 ;
  assign n14298 = n1680 & n2106 ;
  assign n14299 = n14298 ^ n7131 ^ 1'b0 ;
  assign n14300 = n8836 ^ n6433 ^ n5618 ;
  assign n14301 = n11557 | n14300 ;
  assign n14302 = n14299 & ~n14301 ;
  assign n14303 = n1470 ^ n991 ^ 1'b0 ;
  assign n14304 = n11358 & ~n14303 ;
  assign n14305 = n4473 & ~n14304 ;
  assign n14306 = n2385 & n14305 ;
  assign n14307 = ( x33 & n1401 ) | ( x33 & n8595 ) | ( n1401 & n8595 ) ;
  assign n14308 = n12672 ^ n11315 ^ 1'b0 ;
  assign n14309 = ~n13069 & n14308 ;
  assign n14314 = n544 & n3245 ;
  assign n14310 = n11440 ^ n496 ^ 1'b0 ;
  assign n14311 = n7880 | n14310 ;
  assign n14312 = n2637 & ~n14311 ;
  assign n14313 = n7929 & n14312 ;
  assign n14315 = n14314 ^ n14313 ^ n10729 ;
  assign n14316 = n12849 ^ n10011 ^ 1'b0 ;
  assign n14317 = n964 | n3414 ;
  assign n14318 = ( n6477 & ~n14316 ) | ( n6477 & n14317 ) | ( ~n14316 & n14317 ) ;
  assign n14319 = n9561 ^ n377 ^ n307 ;
  assign n14320 = x193 & ~n14319 ;
  assign n14321 = n14320 ^ n1046 ^ 1'b0 ;
  assign n14322 = n14321 ^ n432 ^ 1'b0 ;
  assign n14323 = n12060 ^ n464 ^ 1'b0 ;
  assign n14324 = n14322 & ~n14323 ;
  assign n14325 = n14324 ^ n6384 ^ 1'b0 ;
  assign n14326 = ( ~n8367 & n10042 ) | ( ~n8367 & n11422 ) | ( n10042 & n11422 ) ;
  assign n14327 = ( n419 & n13319 ) | ( n419 & n14326 ) | ( n13319 & n14326 ) ;
  assign n14328 = n13380 ^ n3304 ^ n2706 ;
  assign n14329 = n8201 ^ n2791 ^ 1'b0 ;
  assign n14330 = n10182 | n13233 ;
  assign n14331 = n9149 & ~n14330 ;
  assign n14332 = n4391 | n6511 ;
  assign n14333 = n14332 ^ n6652 ^ 1'b0 ;
  assign n14335 = n5118 ^ n3814 ^ n1196 ;
  assign n14334 = n4422 & n8622 ;
  assign n14336 = n14335 ^ n14334 ^ n7079 ;
  assign n14337 = n13120 & n14336 ;
  assign n14338 = n1702 & ~n12762 ;
  assign n14339 = n14338 ^ n3439 ^ 1'b0 ;
  assign n14340 = n12160 & ~n12663 ;
  assign n14341 = n14340 ^ n6555 ^ 1'b0 ;
  assign n14342 = n14341 ^ n12294 ^ n409 ;
  assign n14343 = n4664 & ~n5124 ;
  assign n14344 = n14343 ^ n2715 ^ 1'b0 ;
  assign n14345 = n14344 ^ n3017 ^ 1'b0 ;
  assign n14346 = n9181 & n14345 ;
  assign n14347 = n5153 & n9426 ;
  assign n14348 = n14347 ^ n3744 ^ 1'b0 ;
  assign n14349 = n8927 & n11302 ;
  assign n14350 = n14348 & n14349 ;
  assign n14351 = ~n14346 & n14350 ;
  assign n14352 = n1196 & n7189 ;
  assign n14353 = n9366 & n9406 ;
  assign n14354 = n787 | n4719 ;
  assign n14355 = n9741 & ~n14354 ;
  assign n14357 = n371 | n4927 ;
  assign n14358 = n2756 | n3136 ;
  assign n14359 = n14358 ^ n7699 ^ 1'b0 ;
  assign n14360 = n14357 & n14359 ;
  assign n14356 = n5732 ^ n2155 ^ 1'b0 ;
  assign n14361 = n14360 ^ n14356 ^ 1'b0 ;
  assign n14362 = ~n4394 & n8760 ;
  assign n14363 = ( n2001 & n9369 ) | ( n2001 & n14362 ) | ( n9369 & n14362 ) ;
  assign n14364 = n14363 ^ n6459 ^ n1555 ;
  assign n14365 = n12906 ^ n4952 ^ 1'b0 ;
  assign n14371 = n459 | n1803 ;
  assign n14372 = n1064 | n14371 ;
  assign n14373 = n4154 & n14372 ;
  assign n14374 = n14373 ^ n7686 ^ 1'b0 ;
  assign n14366 = ( n5171 & ~n7396 ) | ( n5171 & n10011 ) | ( ~n7396 & n10011 ) ;
  assign n14367 = n3281 | n14366 ;
  assign n14368 = n14367 ^ n5888 ^ 1'b0 ;
  assign n14369 = n14368 ^ n9366 ^ 1'b0 ;
  assign n14370 = n1827 | n14369 ;
  assign n14375 = n14374 ^ n14370 ^ 1'b0 ;
  assign n14376 = ~n1322 & n14375 ;
  assign n14377 = ( n2311 & ~n10308 ) | ( n2311 & n14100 ) | ( ~n10308 & n14100 ) ;
  assign n14378 = ( x172 & n6310 ) | ( x172 & n12019 ) | ( n6310 & n12019 ) ;
  assign n14379 = n8106 | n14378 ;
  assign n14380 = ( n6127 & ~n10271 ) | ( n6127 & n14379 ) | ( ~n10271 & n14379 ) ;
  assign n14381 = ~n3428 & n14372 ;
  assign n14382 = ( n3203 & ~n11822 ) | ( n3203 & n14381 ) | ( ~n11822 & n14381 ) ;
  assign n14383 = n14382 ^ n6603 ^ 1'b0 ;
  assign n14384 = n8571 & ~n14383 ;
  assign n14385 = n2917 & ~n5428 ;
  assign n14386 = n14385 ^ n4223 ^ 1'b0 ;
  assign n14390 = n287 ^ x217 ^ 1'b0 ;
  assign n14391 = n1650 & n14390 ;
  assign n14387 = n362 & n5209 ;
  assign n14388 = n5070 | n14387 ;
  assign n14389 = n14388 ^ n5433 ^ 1'b0 ;
  assign n14392 = n14391 ^ n14389 ^ 1'b0 ;
  assign n14393 = n2787 & ~n14392 ;
  assign n14394 = ~n354 & n14393 ;
  assign n14395 = ~n14386 & n14394 ;
  assign n14396 = ( n8942 & n11803 ) | ( n8942 & ~n14395 ) | ( n11803 & ~n14395 ) ;
  assign n14397 = n14396 ^ n5882 ^ n4806 ;
  assign n14398 = n1013 ^ n887 ^ 1'b0 ;
  assign n14399 = n10633 ^ n2895 ^ 1'b0 ;
  assign n14400 = n10323 & ~n14399 ;
  assign n14401 = ~x231 & n1838 ;
  assign n14402 = n14401 ^ n12326 ^ 1'b0 ;
  assign n14403 = n13887 ^ n3112 ^ 1'b0 ;
  assign n14404 = n1958 & ~n14163 ;
  assign n14405 = n13844 ^ n6430 ^ n4637 ;
  assign n14406 = n12360 ^ n2240 ^ 1'b0 ;
  assign n14407 = n1875 ^ n878 ^ n411 ;
  assign n14408 = x205 & n14407 ;
  assign n14409 = n14327 ^ n11355 ^ n2750 ;
  assign n14410 = n13659 ^ n4851 ^ n1768 ;
  assign n14412 = n11192 ^ n2850 ^ 1'b0 ;
  assign n14411 = n8069 & ~n8597 ;
  assign n14413 = n14412 ^ n14411 ^ 1'b0 ;
  assign n14414 = n14410 & ~n14413 ;
  assign n14415 = n14414 ^ n9759 ^ 1'b0 ;
  assign n14416 = n5677 | n13098 ;
  assign n14417 = n14416 ^ n2590 ^ 1'b0 ;
  assign n14418 = n14417 ^ n7252 ^ 1'b0 ;
  assign n14419 = n8006 ^ n3080 ^ 1'b0 ;
  assign n14420 = n3986 | n14419 ;
  assign n14421 = n14420 ^ n10969 ^ 1'b0 ;
  assign n14422 = n9721 ^ n3507 ^ 1'b0 ;
  assign n14423 = ( ~n5717 & n13343 ) | ( ~n5717 & n14422 ) | ( n13343 & n14422 ) ;
  assign n14426 = n6520 ^ n2608 ^ 1'b0 ;
  assign n14427 = ~n440 & n14426 ;
  assign n14424 = n8036 ^ n2225 ^ n1501 ;
  assign n14425 = n13970 | n14424 ;
  assign n14428 = n14427 ^ n14425 ^ 1'b0 ;
  assign n14429 = n14428 ^ n7665 ^ 1'b0 ;
  assign n14430 = n8102 ^ n1030 ^ x247 ;
  assign n14431 = n6581 ^ n5536 ^ 1'b0 ;
  assign n14432 = n14430 | n14431 ;
  assign n14433 = n14163 | n14432 ;
  assign n14434 = n2662 & n4518 ;
  assign n14435 = ~n9793 & n14434 ;
  assign n14436 = n286 | n905 ;
  assign n14437 = ( n5316 & n9879 ) | ( n5316 & n14436 ) | ( n9879 & n14436 ) ;
  assign n14438 = n8839 ^ n987 ^ 1'b0 ;
  assign n14439 = ( x63 & ~n5532 ) | ( x63 & n14208 ) | ( ~n5532 & n14208 ) ;
  assign n14440 = ( ~n5801 & n11415 ) | ( ~n5801 & n14439 ) | ( n11415 & n14439 ) ;
  assign n14441 = n14440 ^ n4070 ^ 1'b0 ;
  assign n14442 = ( n6339 & n14349 ) | ( n6339 & n14441 ) | ( n14349 & n14441 ) ;
  assign n14443 = ~n326 & n14442 ;
  assign n14444 = ( n1759 & n4544 ) | ( n1759 & n5408 ) | ( n4544 & n5408 ) ;
  assign n14445 = x229 & ~n14444 ;
  assign n14446 = n14445 ^ n6863 ^ 1'b0 ;
  assign n14448 = n6827 & n8531 ;
  assign n14449 = n1578 & n7266 ;
  assign n14450 = n4837 & ~n14449 ;
  assign n14451 = ~n4983 & n14450 ;
  assign n14452 = n14448 | n14451 ;
  assign n14447 = n1555 | n3285 ;
  assign n14453 = n14452 ^ n14447 ^ 1'b0 ;
  assign n14454 = n2538 & n10470 ;
  assign n14455 = n5107 | n12572 ;
  assign n14456 = n14455 ^ n8446 ^ 1'b0 ;
  assign n14457 = n9731 ^ n4243 ^ 1'b0 ;
  assign n14458 = n2705 & n14457 ;
  assign n14459 = n2507 ^ n385 ^ 1'b0 ;
  assign n14460 = n288 | n14459 ;
  assign n14461 = n4922 & n8331 ;
  assign n14462 = n2748 & n14461 ;
  assign n14463 = ~n8301 & n10981 ;
  assign n14464 = ~n1326 & n14463 ;
  assign n14469 = ( n1523 & ~n9051 ) | ( n1523 & n12754 ) | ( ~n9051 & n12754 ) ;
  assign n14465 = n11800 ^ n11445 ^ 1'b0 ;
  assign n14466 = n8061 ^ n4837 ^ 1'b0 ;
  assign n14467 = n14466 ^ n6631 ^ n2019 ;
  assign n14468 = ~n14465 & n14467 ;
  assign n14470 = n14469 ^ n14468 ^ 1'b0 ;
  assign n14471 = n1402 & ~n12506 ;
  assign n14472 = n14471 ^ n3568 ^ 1'b0 ;
  assign n14473 = n8883 | n14472 ;
  assign n14474 = n13221 ^ n8201 ^ 1'b0 ;
  assign n14475 = ~n14389 & n14474 ;
  assign n14478 = n6795 | n11863 ;
  assign n14479 = ( x66 & ~n11581 ) | ( x66 & n14478 ) | ( ~n11581 & n14478 ) ;
  assign n14480 = n9653 & n14479 ;
  assign n14476 = ~n2958 & n3690 ;
  assign n14477 = n6477 | n14476 ;
  assign n14481 = n14480 ^ n14477 ^ 1'b0 ;
  assign n14482 = n12470 ^ n4602 ^ 1'b0 ;
  assign n14483 = n7296 & n7484 ;
  assign n14484 = n1257 ^ n1148 ^ 1'b0 ;
  assign n14485 = n10075 ^ n5215 ^ 1'b0 ;
  assign n14486 = n3767 & n8341 ;
  assign n14487 = ( n435 & ~n3256 ) | ( n435 & n4033 ) | ( ~n3256 & n4033 ) ;
  assign n14488 = n890 & n3507 ;
  assign n14489 = n14488 ^ n13382 ^ 1'b0 ;
  assign n14490 = n4540 & ~n14489 ;
  assign n14491 = n14490 ^ n7436 ^ 1'b0 ;
  assign n14492 = n14487 | n14491 ;
  assign n14495 = ~n3808 & n6137 ;
  assign n14493 = n7393 & n8858 ;
  assign n14494 = n14493 ^ n11665 ^ 1'b0 ;
  assign n14496 = n14495 ^ n14494 ^ x180 ;
  assign n14497 = n5903 & ~n14105 ;
  assign n14498 = n14497 ^ n2370 ^ n2215 ;
  assign n14499 = ~n4159 & n12807 ;
  assign n14500 = n14499 ^ n9421 ^ 1'b0 ;
  assign n14506 = n4435 & n5840 ;
  assign n14501 = n1451 & n2299 ;
  assign n14502 = n14501 ^ n3264 ^ 1'b0 ;
  assign n14503 = n3740 & ~n5686 ;
  assign n14504 = n8015 | n14503 ;
  assign n14505 = n14502 & ~n14504 ;
  assign n14507 = n14506 ^ n14505 ^ 1'b0 ;
  assign n14508 = n4318 | n14507 ;
  assign n14509 = n12314 | n13659 ;
  assign n14512 = ~n2964 & n4811 ;
  assign n14513 = n5434 | n12079 ;
  assign n14514 = n14512 | n14513 ;
  assign n14515 = n14514 ^ n3146 ^ 1'b0 ;
  assign n14511 = n6267 & ~n11178 ;
  assign n14516 = n14515 ^ n14511 ^ 1'b0 ;
  assign n14510 = n7039 ^ n1022 ^ 1'b0 ;
  assign n14517 = n14516 ^ n14510 ^ 1'b0 ;
  assign n14518 = n5687 & n8616 ;
  assign n14519 = n3059 & n14518 ;
  assign n14520 = n11976 ^ n9482 ^ 1'b0 ;
  assign n14521 = n9181 & ~n14520 ;
  assign n14522 = ~n1226 & n12787 ;
  assign n14523 = n11178 & n14522 ;
  assign n14524 = ( ~n11867 & n14509 ) | ( ~n11867 & n14523 ) | ( n14509 & n14523 ) ;
  assign n14526 = ~n440 & n1383 ;
  assign n14527 = n7672 & n14526 ;
  assign n14525 = n1994 & n4901 ;
  assign n14528 = n14527 ^ n14525 ^ 1'b0 ;
  assign n14529 = ~n1269 & n14528 ;
  assign n14530 = n4308 ^ n3414 ^ 1'b0 ;
  assign n14531 = ~n14529 & n14530 ;
  assign n14532 = n5310 & n12591 ;
  assign n14533 = ~n11936 & n14532 ;
  assign n14534 = ~n5190 & n8787 ;
  assign n14535 = ~n12111 & n14534 ;
  assign n14536 = n1492 & n14535 ;
  assign n14537 = n2174 & ~n10860 ;
  assign n14538 = n12168 ^ n9581 ^ 1'b0 ;
  assign n14539 = n14538 ^ n6337 ^ n4763 ;
  assign n14540 = ( ~n888 & n12589 ) | ( ~n888 & n13947 ) | ( n12589 & n13947 ) ;
  assign n14541 = ~n5070 & n9345 ;
  assign n14542 = n14541 ^ n9237 ^ 1'b0 ;
  assign n14543 = n4101 ^ n2513 ^ n1754 ;
  assign n14544 = ~n4302 & n14543 ;
  assign n14545 = n3874 ^ x146 ^ 1'b0 ;
  assign n14546 = n14544 & n14545 ;
  assign n14547 = n2860 | n10429 ;
  assign n14548 = n14547 ^ n2062 ^ 1'b0 ;
  assign n14549 = ( n3036 & ~n4928 ) | ( n3036 & n14548 ) | ( ~n4928 & n14548 ) ;
  assign n14550 = ( n8903 & n14546 ) | ( n8903 & ~n14549 ) | ( n14546 & ~n14549 ) ;
  assign n14551 = n14550 ^ n5292 ^ n3102 ;
  assign n14552 = ~n2523 & n5456 ;
  assign n14553 = n14552 ^ n5706 ^ 1'b0 ;
  assign n14554 = ~n4244 & n6973 ;
  assign n14555 = n14553 & n14554 ;
  assign n14556 = ( n14542 & ~n14551 ) | ( n14542 & n14555 ) | ( ~n14551 & n14555 ) ;
  assign n14557 = n9539 & ~n14556 ;
  assign n14558 = n14557 ^ n4019 ^ 1'b0 ;
  assign n14559 = n11589 ^ n2426 ^ 1'b0 ;
  assign n14560 = n6137 ^ x45 ^ 1'b0 ;
  assign n14561 = ~n14559 & n14560 ;
  assign n14562 = n14561 ^ n8106 ^ 1'b0 ;
  assign n14563 = n8129 ^ n6558 ^ n5999 ;
  assign n14564 = n8669 & ~n14563 ;
  assign n14565 = n14564 ^ n3581 ^ 1'b0 ;
  assign n14566 = n12866 ^ n11759 ^ 1'b0 ;
  assign n14567 = ( ~n1409 & n11764 ) | ( ~n1409 & n13277 ) | ( n11764 & n13277 ) ;
  assign n14568 = n13494 ^ n12963 ^ x31 ;
  assign n14569 = n2210 & n4700 ;
  assign n14570 = n4085 & n14569 ;
  assign n14571 = n1185 & n12655 ;
  assign n14572 = n14571 ^ n2682 ^ 1'b0 ;
  assign n14573 = n14570 | n14572 ;
  assign n14575 = n2050 & ~n4754 ;
  assign n14574 = n3227 | n7887 ;
  assign n14576 = n14575 ^ n14574 ^ 1'b0 ;
  assign n14577 = ( n7843 & n12983 ) | ( n7843 & n14576 ) | ( n12983 & n14576 ) ;
  assign n14578 = n4395 ^ n3514 ^ 1'b0 ;
  assign n14579 = n9332 & ~n14578 ;
  assign n14580 = n14277 & n14579 ;
  assign n14581 = n887 & n8317 ;
  assign n14582 = n6818 ^ n5499 ^ n4305 ;
  assign n14583 = ( n7008 & n9882 ) | ( n7008 & n12160 ) | ( n9882 & n12160 ) ;
  assign n14587 = n300 & n8528 ;
  assign n14585 = ~n3557 & n3798 ;
  assign n14584 = n4108 | n6438 ;
  assign n14586 = n14585 ^ n14584 ^ 1'b0 ;
  assign n14588 = n14587 ^ n14586 ^ 1'b0 ;
  assign n14589 = ( n2875 & ~n14583 ) | ( n2875 & n14588 ) | ( ~n14583 & n14588 ) ;
  assign n14590 = x165 & ~n6133 ;
  assign n14591 = n333 & n14590 ;
  assign n14592 = n1881 | n8997 ;
  assign n14593 = n12644 & ~n14592 ;
  assign n14594 = n14593 ^ n5174 ^ 1'b0 ;
  assign n14595 = ~n14591 & n14594 ;
  assign n14596 = n14595 ^ n6458 ^ n407 ;
  assign n14597 = n10990 ^ n10852 ^ 1'b0 ;
  assign n14598 = ~n9593 & n14597 ;
  assign n14599 = n13968 ^ n6679 ^ 1'b0 ;
  assign n14600 = ( n840 & n11634 ) | ( n840 & ~n14401 ) | ( n11634 & ~n14401 ) ;
  assign n14601 = n11998 | n14600 ;
  assign n14602 = n14601 ^ n5073 ^ 1'b0 ;
  assign n14603 = ~n2522 & n4952 ;
  assign n14604 = ~n9497 & n14603 ;
  assign n14605 = n14559 ^ n12271 ^ n9365 ;
  assign n14606 = ( ~n6138 & n7046 ) | ( ~n6138 & n14605 ) | ( n7046 & n14605 ) ;
  assign n14607 = n10456 | n14606 ;
  assign n14608 = n14607 ^ n4212 ^ 1'b0 ;
  assign n14609 = n7451 ^ n4515 ^ 1'b0 ;
  assign n14611 = n1580 ^ n922 ^ n826 ;
  assign n14612 = ( ~n3056 & n6064 ) | ( ~n3056 & n14611 ) | ( n6064 & n14611 ) ;
  assign n14610 = n2995 & n6669 ;
  assign n14613 = n14612 ^ n14610 ^ 1'b0 ;
  assign n14614 = n2117 & n14613 ;
  assign n14615 = n14614 ^ n3538 ^ 1'b0 ;
  assign n14616 = n4653 & ~n6032 ;
  assign n14617 = n14616 ^ n3239 ^ 1'b0 ;
  assign n14618 = ( n10953 & ~n11686 ) | ( n10953 & n14617 ) | ( ~n11686 & n14617 ) ;
  assign n14619 = n14618 ^ n9803 ^ n7136 ;
  assign n14620 = n4616 & ~n14619 ;
  assign n14621 = ~n9224 & n14620 ;
  assign n14622 = n3339 & ~n4725 ;
  assign n14623 = n14622 ^ n1750 ^ 1'b0 ;
  assign n14624 = n14623 ^ n5070 ^ 1'b0 ;
  assign n14625 = n10306 & ~n14624 ;
  assign n14626 = ( n1005 & n1148 ) | ( n1005 & ~n10724 ) | ( n1148 & ~n10724 ) ;
  assign n14627 = x70 & n6477 ;
  assign n14628 = n4514 ^ n4448 ^ 1'b0 ;
  assign n14629 = n14628 ^ n5236 ^ n1770 ;
  assign n14630 = n14629 ^ n4653 ^ 1'b0 ;
  assign n14631 = n4351 | n14020 ;
  assign n14632 = n1949 & ~n14631 ;
  assign n14633 = ~n8020 & n8858 ;
  assign n14634 = n12540 & n14633 ;
  assign n14635 = n14632 & ~n14634 ;
  assign n14636 = n716 & n3557 ;
  assign n14637 = ~n9498 & n14636 ;
  assign n14638 = ( n9376 & n9890 ) | ( n9376 & ~n14637 ) | ( n9890 & ~n14637 ) ;
  assign n14639 = ( n1063 & n1067 ) | ( n1063 & ~n9605 ) | ( n1067 & ~n9605 ) ;
  assign n14640 = x226 & ~n14639 ;
  assign n14641 = n14640 ^ n2648 ^ 1'b0 ;
  assign n14642 = ( n6077 & ~n6767 ) | ( n6077 & n10857 ) | ( ~n6767 & n10857 ) ;
  assign n14643 = n14642 ^ n4579 ^ 1'b0 ;
  assign n14644 = ~n11504 & n14643 ;
  assign n14645 = n5591 | n10180 ;
  assign n14646 = n10826 & ~n14645 ;
  assign n14648 = n8217 ^ n6588 ^ n1499 ;
  assign n14647 = ~n9012 & n14307 ;
  assign n14649 = n14648 ^ n14647 ^ n2600 ;
  assign n14651 = n1258 ^ n847 ^ 1'b0 ;
  assign n14650 = ~n2624 & n7113 ;
  assign n14652 = n14651 ^ n14650 ^ 1'b0 ;
  assign n14653 = n3150 ^ x159 ^ 1'b0 ;
  assign n14654 = ~n1081 & n14653 ;
  assign n14655 = n14654 ^ n12889 ^ n1274 ;
  assign n14656 = n14655 ^ n10794 ^ 1'b0 ;
  assign n14657 = n14652 & ~n14656 ;
  assign n14658 = ( n1258 & n7968 ) | ( n1258 & ~n8593 ) | ( n7968 & ~n8593 ) ;
  assign n14659 = n5024 & ~n9602 ;
  assign n14660 = n14659 ^ n9525 ^ n8722 ;
  assign n14661 = ( n3957 & n14658 ) | ( n3957 & n14660 ) | ( n14658 & n14660 ) ;
  assign n14662 = n7294 ^ n5672 ^ 1'b0 ;
  assign n14663 = ~n5655 & n14662 ;
  assign n14664 = x104 & ~n9295 ;
  assign n14665 = n10252 & n14664 ;
  assign n14666 = n14665 ^ n4773 ^ 1'b0 ;
  assign n14667 = n14663 | n14666 ;
  assign n14668 = n12550 ^ n6846 ^ 1'b0 ;
  assign n14669 = n11330 & n14668 ;
  assign n14670 = n771 & ~n1076 ;
  assign n14671 = n3492 & n14670 ;
  assign n14672 = ~n14669 & n14671 ;
  assign n14673 = n6986 & ~n14672 ;
  assign n14682 = ~n12034 & n12084 ;
  assign n14683 = ~n10267 & n14682 ;
  assign n14684 = n14683 ^ n4847 ^ 1'b0 ;
  assign n14680 = n9278 ^ n2680 ^ 1'b0 ;
  assign n14681 = n994 | n14680 ;
  assign n14674 = n5257 | n14274 ;
  assign n14675 = n7682 & ~n14674 ;
  assign n14676 = n1932 ^ n1335 ^ 1'b0 ;
  assign n14677 = n14675 | n14676 ;
  assign n14678 = n3203 | n14677 ;
  assign n14679 = n14678 ^ n1481 ^ 1'b0 ;
  assign n14685 = n14684 ^ n14681 ^ n14679 ;
  assign n14687 = n8151 ^ n6642 ^ 1'b0 ;
  assign n14686 = n1018 & ~n4971 ;
  assign n14688 = n14687 ^ n14686 ^ n4595 ;
  assign n14689 = n12847 ^ n11620 ^ n5156 ;
  assign n14690 = n14689 ^ n3255 ^ 1'b0 ;
  assign n14704 = n660 ^ n442 ^ 1'b0 ;
  assign n14703 = n1860 & ~n8703 ;
  assign n14691 = n8368 ^ n3212 ^ 1'b0 ;
  assign n14692 = n1657 & n6249 ;
  assign n14693 = x202 | n14692 ;
  assign n14694 = n14691 & ~n14693 ;
  assign n14695 = n10489 | n14694 ;
  assign n14696 = n14695 ^ n1672 ^ 1'b0 ;
  assign n14697 = n6938 ^ n2335 ^ 1'b0 ;
  assign n14698 = ~n5018 & n14697 ;
  assign n14699 = ~n8208 & n14698 ;
  assign n14700 = n14699 ^ n13189 ^ 1'b0 ;
  assign n14701 = n14700 ^ n5699 ^ 1'b0 ;
  assign n14702 = ~n14696 & n14701 ;
  assign n14705 = n14704 ^ n14703 ^ n14702 ;
  assign n14706 = n8753 & ~n10034 ;
  assign n14707 = n493 & n14706 ;
  assign n14708 = n14401 ^ n13737 ^ 1'b0 ;
  assign n14714 = n4286 ^ n2626 ^ 1'b0 ;
  assign n14715 = n14714 ^ n11489 ^ n2378 ;
  assign n14711 = n1350 | n8588 ;
  assign n14712 = n14711 ^ n11502 ^ n2128 ;
  assign n14709 = n5810 | n8013 ;
  assign n14710 = n1107 & ~n14709 ;
  assign n14713 = n14712 ^ n14710 ^ 1'b0 ;
  assign n14716 = n14715 ^ n14713 ^ 1'b0 ;
  assign n14717 = n8926 & n14716 ;
  assign n14718 = n6037 | n12721 ;
  assign n14719 = n14718 ^ x244 ^ 1'b0 ;
  assign n14720 = n9511 ^ n2983 ^ 1'b0 ;
  assign n14721 = n8273 | n14720 ;
  assign n14722 = n14721 ^ n12231 ^ n7386 ;
  assign n14723 = x32 & ~n9567 ;
  assign n14724 = n13096 & n14723 ;
  assign n14725 = n4247 ^ n637 ^ 1'b0 ;
  assign n14726 = n12374 ^ n3132 ^ 1'b0 ;
  assign n14727 = n14726 ^ n2317 ^ 1'b0 ;
  assign n14728 = n8753 & ~n14727 ;
  assign n14729 = n5805 ^ n487 ^ 1'b0 ;
  assign n14730 = n13288 | n14729 ;
  assign n14731 = n12726 | n14730 ;
  assign n14732 = n1026 | n1214 ;
  assign n14733 = n2972 | n3791 ;
  assign n14734 = n14733 ^ n5077 ^ 1'b0 ;
  assign n14735 = n14734 ^ n8481 ^ 1'b0 ;
  assign n14736 = n4931 ^ n1713 ^ 1'b0 ;
  assign n14737 = ~n5446 & n14736 ;
  assign n14738 = n4999 & n14737 ;
  assign n14739 = n14738 ^ n1769 ^ 1'b0 ;
  assign n14740 = x200 & n9694 ;
  assign n14741 = ~n14739 & n14740 ;
  assign n14742 = n14741 ^ n6833 ^ n921 ;
  assign n14743 = n3335 | n14742 ;
  assign n14744 = n1970 & ~n8272 ;
  assign n14745 = ~n7244 & n13618 ;
  assign n14746 = ~n11372 & n14745 ;
  assign n14747 = ( n2731 & n5327 ) | ( n2731 & ~n9255 ) | ( n5327 & ~n9255 ) ;
  assign n14748 = n14747 ^ n1140 ^ 1'b0 ;
  assign n14749 = n1503 & ~n11530 ;
  assign n14750 = n7222 | n8775 ;
  assign n14751 = n14749 | n14750 ;
  assign n14752 = n12140 ^ n7240 ^ 1'b0 ;
  assign n14753 = n6546 ^ n1888 ^ 1'b0 ;
  assign n14754 = n14753 ^ n14262 ^ n7746 ;
  assign n14755 = ( n1846 & n14752 ) | ( n1846 & n14754 ) | ( n14752 & n14754 ) ;
  assign n14756 = n1016 | n8993 ;
  assign n14757 = n8902 ^ n7174 ^ n2693 ;
  assign n14758 = n4324 & n8580 ;
  assign n14759 = n4079 ^ n1711 ^ 1'b0 ;
  assign n14760 = ( n1304 & n14758 ) | ( n1304 & ~n14759 ) | ( n14758 & ~n14759 ) ;
  assign n14761 = n1734 | n5965 ;
  assign n14762 = n14761 ^ n8476 ^ 1'b0 ;
  assign n14763 = n1527 ^ n512 ^ 1'b0 ;
  assign n14764 = n1427 | n14763 ;
  assign n14765 = ~x209 & n14764 ;
  assign n14766 = n10327 & ~n13806 ;
  assign n14767 = n14498 ^ n6618 ^ 1'b0 ;
  assign n14768 = n14766 | n14767 ;
  assign n14769 = ~n5684 & n12265 ;
  assign n14770 = n3051 & n14769 ;
  assign n14771 = n2835 & ~n2906 ;
  assign n14772 = ~n9436 & n14771 ;
  assign n14773 = n5137 & n11997 ;
  assign n14774 = ~n9438 & n14773 ;
  assign n14775 = n10356 & ~n11242 ;
  assign n14776 = n14774 & ~n14775 ;
  assign n14777 = ~n8613 & n14714 ;
  assign n14778 = n14777 ^ n3700 ^ 1'b0 ;
  assign n14779 = ( n4013 & ~n5166 ) | ( n4013 & n5355 ) | ( ~n5166 & n5355 ) ;
  assign n14780 = ~n4355 & n4827 ;
  assign n14781 = n6967 ^ n3924 ^ n3072 ;
  assign n14782 = ~n10364 & n14781 ;
  assign n14783 = ~n2860 & n10768 ;
  assign n14784 = ~n11817 & n14783 ;
  assign n14785 = n922 & n2204 ;
  assign n14786 = n12678 | n14785 ;
  assign n14788 = n3557 & ~n4357 ;
  assign n14789 = n14788 ^ n6965 ^ 1'b0 ;
  assign n14787 = n3255 & ~n3475 ;
  assign n14790 = n14789 ^ n14787 ^ n5928 ;
  assign n14791 = ( n1442 & ~n4523 ) | ( n1442 & n6032 ) | ( ~n4523 & n6032 ) ;
  assign n14792 = n3959 & ~n14791 ;
  assign n14793 = n14792 ^ n10493 ^ 1'b0 ;
  assign n14794 = n10145 | n14793 ;
  assign n14795 = n3955 | n14794 ;
  assign n14796 = n3068 ^ n2217 ^ 1'b0 ;
  assign n14797 = n4493 ^ n4278 ^ 1'b0 ;
  assign n14798 = ~n14796 & n14797 ;
  assign n14799 = ~n2280 & n14798 ;
  assign n14800 = ~n11815 & n14799 ;
  assign n14801 = ( n1784 & ~n3790 ) | ( n1784 & n14800 ) | ( ~n3790 & n14800 ) ;
  assign n14802 = n3994 & n12333 ;
  assign n14803 = ~n2362 & n14802 ;
  assign n14804 = n14803 ^ n6820 ^ 1'b0 ;
  assign n14805 = n5411 ^ n2678 ^ 1'b0 ;
  assign n14806 = n3523 | n14805 ;
  assign n14807 = n14806 ^ n8948 ^ 1'b0 ;
  assign n14808 = n4696 | n14807 ;
  assign n14809 = n10796 & ~n14808 ;
  assign n14810 = n14809 ^ n9601 ^ n9158 ;
  assign n14811 = ( ~n303 & n3953 ) | ( ~n303 & n4286 ) | ( n3953 & n4286 ) ;
  assign n14812 = n14811 ^ n4591 ^ 1'b0 ;
  assign n14813 = n12817 | n14812 ;
  assign n14814 = n14766 ^ n9704 ^ 1'b0 ;
  assign n14815 = n12720 & ~n14814 ;
  assign n14816 = ( ~n4922 & n10862 ) | ( ~n4922 & n14815 ) | ( n10862 & n14815 ) ;
  assign n14823 = n3259 & ~n12674 ;
  assign n14824 = n14823 ^ n3060 ^ 1'b0 ;
  assign n14818 = x207 & n1022 ;
  assign n14819 = n4676 ^ n4522 ^ n4298 ;
  assign n14820 = ~n14818 & n14819 ;
  assign n14821 = n6936 & n14820 ;
  assign n14817 = n6557 & n8315 ;
  assign n14822 = n14821 ^ n14817 ^ 1'b0 ;
  assign n14825 = n14824 ^ n14822 ^ n10941 ;
  assign n14830 = x205 & n4326 ;
  assign n14831 = n396 & n14830 ;
  assign n14832 = n14831 ^ n5985 ^ n5135 ;
  assign n14826 = ~n1748 & n3677 ;
  assign n14827 = n14826 ^ n5405 ^ 1'b0 ;
  assign n14828 = n3267 & ~n4553 ;
  assign n14829 = ~n14827 & n14828 ;
  assign n14833 = n14832 ^ n14829 ^ 1'b0 ;
  assign n14834 = n6390 & n9332 ;
  assign n14835 = ~n4299 & n14834 ;
  assign n14836 = n7954 | n14835 ;
  assign n14837 = n14836 ^ n651 ^ 1'b0 ;
  assign n14838 = n2808 & ~n14837 ;
  assign n14839 = ~n3113 & n5239 ;
  assign n14840 = ( ~n3373 & n9073 ) | ( ~n3373 & n14839 ) | ( n9073 & n14839 ) ;
  assign n14841 = n3759 ^ n3742 ^ n269 ;
  assign n14842 = n14841 ^ n7677 ^ 1'b0 ;
  assign n14843 = n6632 ^ x35 ^ 1'b0 ;
  assign n14844 = n14549 | n14843 ;
  assign n14845 = n14844 ^ n10398 ^ n619 ;
  assign n14846 = n9090 ^ n8282 ^ n1755 ;
  assign n14847 = n8387 ^ n2235 ^ n337 ;
  assign n14848 = n14847 ^ n4009 ^ 1'b0 ;
  assign n14849 = n10614 ^ n7716 ^ n1264 ;
  assign n14850 = ( n5639 & n11217 ) | ( n5639 & n14849 ) | ( n11217 & n14849 ) ;
  assign n14851 = ( n4123 & n14848 ) | ( n4123 & ~n14850 ) | ( n14848 & ~n14850 ) ;
  assign n14852 = ( n9653 & n14846 ) | ( n9653 & ~n14851 ) | ( n14846 & ~n14851 ) ;
  assign n14853 = n754 & ~n9388 ;
  assign n14854 = n14853 ^ n2766 ^ 1'b0 ;
  assign n14855 = n14854 ^ n10258 ^ n2229 ;
  assign n14856 = n14855 ^ n523 ^ 1'b0 ;
  assign n14857 = n14856 ^ n9483 ^ 1'b0 ;
  assign n14858 = n9161 | n14857 ;
  assign n14863 = n12140 ^ n545 ^ 1'b0 ;
  assign n14862 = ~n433 & n10311 ;
  assign n14859 = n1836 | n8818 ;
  assign n14860 = n2859 | n14859 ;
  assign n14861 = n14860 ^ n3640 ^ 1'b0 ;
  assign n14864 = n14863 ^ n14862 ^ n14861 ;
  assign n14866 = n4928 ^ n4164 ^ n711 ;
  assign n14870 = n4550 ^ n3892 ^ n3883 ;
  assign n14867 = ( n1220 & n2920 ) | ( n1220 & ~n9536 ) | ( n2920 & ~n9536 ) ;
  assign n14868 = n14867 ^ n3256 ^ 1'b0 ;
  assign n14869 = n5193 & n14868 ;
  assign n14871 = n14870 ^ n14869 ^ n3328 ;
  assign n14872 = n14866 & ~n14871 ;
  assign n14873 = n14872 ^ n6613 ^ 1'b0 ;
  assign n14865 = n13326 & n14150 ;
  assign n14874 = n14873 ^ n14865 ^ 1'b0 ;
  assign n14875 = n1247 & n8003 ;
  assign n14876 = n14306 & n14875 ;
  assign n14877 = n9670 ^ n1895 ^ 1'b0 ;
  assign n14878 = n12595 ^ n4844 ^ n2418 ;
  assign n14879 = n2482 & ~n5105 ;
  assign n14880 = n14879 ^ n13068 ^ 1'b0 ;
  assign n14881 = n4053 & n11412 ;
  assign n14882 = ~n3409 & n14881 ;
  assign n14883 = n7540 & n14882 ;
  assign n14884 = n3519 & ~n10172 ;
  assign n14885 = n9537 & ~n14884 ;
  assign n14886 = n14885 ^ n9086 ^ 1'b0 ;
  assign n14888 = n4979 & ~n5672 ;
  assign n14889 = ( n3342 & n6075 ) | ( n3342 & ~n14888 ) | ( n6075 & ~n14888 ) ;
  assign n14887 = n4455 & ~n5359 ;
  assign n14890 = n14889 ^ n14887 ^ 1'b0 ;
  assign n14891 = ~n14886 & n14890 ;
  assign n14892 = ~n6921 & n9050 ;
  assign n14894 = ( n1629 & n1770 ) | ( n1629 & n1975 ) | ( n1770 & n1975 ) ;
  assign n14893 = n6954 & n9631 ;
  assign n14895 = n14894 ^ n14893 ^ 1'b0 ;
  assign n14896 = n11251 ^ n7176 ^ n813 ;
  assign n14897 = n14896 ^ n8374 ^ 1'b0 ;
  assign n14898 = ( n1140 & ~n8431 ) | ( n1140 & n14897 ) | ( ~n8431 & n14897 ) ;
  assign n14899 = n3100 & n14898 ;
  assign n14900 = ( ~n7878 & n7994 ) | ( ~n7878 & n9485 ) | ( n7994 & n9485 ) ;
  assign n14912 = n8254 ^ n5438 ^ n4159 ;
  assign n14913 = n14912 ^ x123 ^ 1'b0 ;
  assign n14914 = n4512 | n14913 ;
  assign n14904 = n1564 & ~n5326 ;
  assign n14905 = n14904 ^ n4155 ^ 1'b0 ;
  assign n14906 = n14905 ^ n13089 ^ n5662 ;
  assign n14907 = ~x102 & n5206 ;
  assign n14908 = n14907 ^ n10084 ^ n4059 ;
  assign n14909 = ( ~n1407 & n5089 ) | ( ~n1407 & n14908 ) | ( n5089 & n14908 ) ;
  assign n14910 = ~n12929 & n14909 ;
  assign n14911 = ~n14906 & n14910 ;
  assign n14915 = n14914 ^ n14911 ^ 1'b0 ;
  assign n14916 = ~n12772 & n14915 ;
  assign n14917 = ~n6482 & n14916 ;
  assign n14918 = ~n14049 & n14917 ;
  assign n14901 = x124 & n263 ;
  assign n14902 = n9408 & n14901 ;
  assign n14903 = n2522 & n14902 ;
  assign n14919 = n14918 ^ n14903 ^ 1'b0 ;
  assign n14924 = ( ~n966 & n1189 ) | ( ~n966 & n3813 ) | ( n1189 & n3813 ) ;
  assign n14925 = n4761 | n14924 ;
  assign n14926 = n13511 & ~n14925 ;
  assign n14921 = ( n4600 & ~n6211 ) | ( n4600 & n8266 ) | ( ~n6211 & n8266 ) ;
  assign n14920 = ~n691 & n11201 ;
  assign n14922 = n14921 ^ n14920 ^ 1'b0 ;
  assign n14923 = n3153 & n14922 ;
  assign n14927 = n14926 ^ n14923 ^ n12565 ;
  assign n14928 = n6585 & ~n7789 ;
  assign n14929 = n3359 & n14928 ;
  assign n14930 = n14929 ^ n12413 ^ n3796 ;
  assign n14931 = ~n6717 & n14930 ;
  assign n14932 = ~n12735 & n14931 ;
  assign n14933 = n4359 | n12193 ;
  assign n14934 = n14932 & ~n14933 ;
  assign n14935 = n4097 ^ n1958 ^ 1'b0 ;
  assign n14936 = n365 & n14935 ;
  assign n14937 = ~n713 & n1580 ;
  assign n14938 = n14937 ^ n5483 ^ 1'b0 ;
  assign n14939 = n2780 | n14938 ;
  assign n14940 = n14936 | n14939 ;
  assign n14941 = n2152 | n14940 ;
  assign n14942 = ~n4879 & n6685 ;
  assign n14943 = ( n5653 & ~n10829 ) | ( n5653 & n12425 ) | ( ~n10829 & n12425 ) ;
  assign n14944 = n14943 ^ n7908 ^ n5238 ;
  assign n14945 = n3728 ^ x250 ^ 1'b0 ;
  assign n14946 = n329 & n14945 ;
  assign n14947 = n14946 ^ n8388 ^ 1'b0 ;
  assign n14948 = ~n4427 & n14947 ;
  assign n14949 = n14948 ^ n7416 ^ n5318 ;
  assign n14950 = n14870 ^ n5976 ^ 1'b0 ;
  assign n14951 = n11080 & ~n14950 ;
  assign n14952 = n14951 ^ n11576 ^ 1'b0 ;
  assign n14953 = n9191 & ~n14952 ;
  assign n14954 = ( n1737 & n11772 ) | ( n1737 & n14953 ) | ( n11772 & n14953 ) ;
  assign n14955 = ~n13137 & n14954 ;
  assign n14956 = n6310 ^ n1540 ^ 1'b0 ;
  assign n14957 = n13252 | n14956 ;
  assign n14958 = ( x176 & n2182 ) | ( x176 & n14957 ) | ( n2182 & n14957 ) ;
  assign n14959 = n2953 ^ n358 ^ 1'b0 ;
  assign n14960 = ~n3307 & n14959 ;
  assign n14961 = n8552 | n14960 ;
  assign n14962 = n7578 ^ n5522 ^ 1'b0 ;
  assign n14963 = ~n1603 & n14962 ;
  assign n14968 = n5935 ^ n4234 ^ 1'b0 ;
  assign n14969 = ( n5766 & n8215 ) | ( n5766 & n14968 ) | ( n8215 & n14968 ) ;
  assign n14967 = n9085 ^ n6215 ^ n658 ;
  assign n14964 = ~n1019 & n2824 ;
  assign n14965 = ~n3909 & n14964 ;
  assign n14966 = ( n6189 & n6732 ) | ( n6189 & n14965 ) | ( n6732 & n14965 ) ;
  assign n14970 = n14969 ^ n14967 ^ n14966 ;
  assign n14971 = ~n904 & n14970 ;
  assign n14972 = n12274 & ~n14255 ;
  assign n14973 = n14972 ^ n4902 ^ 1'b0 ;
  assign n14976 = n3426 ^ n3173 ^ n773 ;
  assign n14974 = n6574 ^ n1199 ^ 1'b0 ;
  assign n14975 = n14974 ^ n6531 ^ 1'b0 ;
  assign n14977 = n14976 ^ n14975 ^ n5631 ;
  assign n14978 = n8646 ^ n6453 ^ 1'b0 ;
  assign n14979 = n12820 | n14978 ;
  assign n14980 = n1006 | n14979 ;
  assign n14981 = ( x123 & n335 ) | ( x123 & ~n2117 ) | ( n335 & ~n2117 ) ;
  assign n14982 = n14981 ^ n6398 ^ 1'b0 ;
  assign n14983 = ~n6990 & n14261 ;
  assign n14984 = ~n2843 & n6188 ;
  assign n14985 = ( ~n2204 & n2892 ) | ( ~n2204 & n14984 ) | ( n2892 & n14984 ) ;
  assign n14986 = n14985 ^ n7869 ^ 1'b0 ;
  assign n14987 = n6691 & ~n10691 ;
  assign n14988 = n8138 & n14987 ;
  assign n14989 = ( x113 & n2138 ) | ( x113 & ~n8180 ) | ( n2138 & ~n8180 ) ;
  assign n14990 = n14909 ^ n13907 ^ n11543 ;
  assign n14991 = n4428 & ~n5155 ;
  assign n14992 = n14991 ^ n691 ^ 1'b0 ;
  assign n14993 = ( n4163 & n4215 ) | ( n4163 & ~n14992 ) | ( n4215 & ~n14992 ) ;
  assign n14994 = n4143 & ~n14993 ;
  assign n14995 = n14994 ^ n1781 ^ 1'b0 ;
  assign n14996 = ~n4207 & n7228 ;
  assign n14997 = ~n932 & n14996 ;
  assign n14998 = n5524 & ~n14997 ;
  assign n14999 = n7641 ^ x149 ^ 1'b0 ;
  assign n15000 = n14999 ^ n7469 ^ n1944 ;
  assign n15001 = n6836 ^ n2090 ^ 1'b0 ;
  assign n15002 = n9869 | n15001 ;
  assign n15003 = n15002 ^ n6669 ^ 1'b0 ;
  assign n15004 = n9276 | n10957 ;
  assign n15005 = n15003 & ~n15004 ;
  assign n15006 = n6379 & n15005 ;
  assign n15007 = n7396 ^ n5894 ^ 1'b0 ;
  assign n15010 = n5427 ^ n968 ^ 1'b0 ;
  assign n15011 = n15010 ^ n4242 ^ 1'b0 ;
  assign n15012 = n4274 & n15011 ;
  assign n15013 = ( n6962 & ~n10657 ) | ( n6962 & n15012 ) | ( ~n10657 & n15012 ) ;
  assign n15009 = n1252 & ~n12885 ;
  assign n15008 = n4659 | n9711 ;
  assign n15014 = n15013 ^ n15009 ^ n15008 ;
  assign n15015 = n15014 ^ n11062 ^ n4854 ;
  assign n15016 = n4925 | n8030 ;
  assign n15017 = n13630 | n15016 ;
  assign n15018 = n6370 ^ n3910 ^ 1'b0 ;
  assign n15019 = n12102 & ~n14168 ;
  assign n15020 = n13362 & n15019 ;
  assign n15021 = n6382 & n8494 ;
  assign n15022 = n8268 & n15021 ;
  assign n15023 = n8626 ^ n7115 ^ 1'b0 ;
  assign n15024 = ~n3279 & n15023 ;
  assign n15025 = n3967 ^ n1452 ^ 1'b0 ;
  assign n15026 = ~n6023 & n15025 ;
  assign n15027 = ( ~n943 & n2294 ) | ( ~n943 & n15026 ) | ( n2294 & n15026 ) ;
  assign n15028 = n1675 & ~n8467 ;
  assign n15029 = ~n15027 & n15028 ;
  assign n15030 = x114 | n5653 ;
  assign n15031 = n8381 & ~n15030 ;
  assign n15032 = n7942 ^ n1476 ^ x48 ;
  assign n15033 = ~n10955 & n15032 ;
  assign n15034 = n15033 ^ n13346 ^ 1'b0 ;
  assign n15035 = ~n7736 & n15034 ;
  assign n15036 = n15031 & n15035 ;
  assign n15037 = n15029 & n15036 ;
  assign n15038 = n5326 & ~n5548 ;
  assign n15039 = ~n3550 & n15038 ;
  assign n15040 = n12378 ^ n5898 ^ n2945 ;
  assign n15041 = n15039 & ~n15040 ;
  assign n15042 = n4747 & n15041 ;
  assign n15043 = n6981 ^ n2763 ^ 1'b0 ;
  assign n15044 = n4740 & n15043 ;
  assign n15045 = n15044 ^ n5258 ^ n3693 ;
  assign n15049 = n4457 ^ n264 ^ 1'b0 ;
  assign n15046 = ( n1508 & n2124 ) | ( n1508 & n3546 ) | ( n2124 & n3546 ) ;
  assign n15047 = n1076 | n15046 ;
  assign n15048 = n4752 | n15047 ;
  assign n15050 = n15049 ^ n15048 ^ 1'b0 ;
  assign n15051 = n11842 ^ n9675 ^ 1'b0 ;
  assign n15052 = ~n5664 & n11174 ;
  assign n15053 = n7199 & n13988 ;
  assign n15054 = ~n15052 & n15053 ;
  assign n15055 = n1047 | n6860 ;
  assign n15056 = n15054 & ~n15055 ;
  assign n15057 = ~n472 & n495 ;
  assign n15058 = n7376 ^ n1540 ^ n574 ;
  assign n15059 = n15058 ^ n9948 ^ 1'b0 ;
  assign n15060 = n12814 | n15059 ;
  assign n15061 = ~n330 & n15060 ;
  assign n15062 = n15061 ^ n11663 ^ 1'b0 ;
  assign n15063 = n6195 ^ n2638 ^ n2459 ;
  assign n15064 = n15062 & ~n15063 ;
  assign n15065 = ~n15057 & n15064 ;
  assign n15068 = n2200 ^ n1537 ^ 1'b0 ;
  assign n15066 = n633 | n3615 ;
  assign n15067 = n15066 ^ n487 ^ 1'b0 ;
  assign n15069 = n15068 ^ n15067 ^ n12474 ;
  assign n15070 = ~n802 & n15069 ;
  assign n15071 = n11435 ^ n8015 ^ 1'b0 ;
  assign n15072 = n15071 ^ n1835 ^ 1'b0 ;
  assign n15073 = n4398 & ~n15072 ;
  assign n15074 = n10346 | n15073 ;
  assign n15081 = ( n6511 & n6516 ) | ( n6511 & n6664 ) | ( n6516 & n6664 ) ;
  assign n15075 = n3470 & ~n5206 ;
  assign n15076 = n2663 & ~n15075 ;
  assign n15077 = n2220 | n11488 ;
  assign n15078 = n15077 ^ n6938 ^ 1'b0 ;
  assign n15079 = n15078 ^ n1995 ^ 1'b0 ;
  assign n15080 = n15076 & n15079 ;
  assign n15082 = n15081 ^ n15080 ^ 1'b0 ;
  assign n15083 = n12220 ^ n4920 ^ 1'b0 ;
  assign n15084 = n6776 ^ n2290 ^ x24 ;
  assign n15085 = n9650 & ~n14588 ;
  assign n15086 = n14018 ^ n6065 ^ 1'b0 ;
  assign n15087 = n3312 & n15086 ;
  assign n15088 = n15085 & n15087 ;
  assign n15089 = n12608 ^ n9859 ^ n1519 ;
  assign n15090 = n4404 & ~n14051 ;
  assign n15091 = n4454 & n7131 ;
  assign n15092 = n15091 ^ n2230 ^ n1185 ;
  assign n15093 = n9795 ^ n8999 ^ 1'b0 ;
  assign n15094 = n453 & n1486 ;
  assign n15095 = ( n7006 & n13117 ) | ( n7006 & ~n13155 ) | ( n13117 & ~n13155 ) ;
  assign n15096 = ( n2546 & n6752 ) | ( n2546 & ~n8418 ) | ( n6752 & ~n8418 ) ;
  assign n15097 = ( ~n2529 & n12903 ) | ( ~n2529 & n15096 ) | ( n12903 & n15096 ) ;
  assign n15098 = ( n1641 & n5144 ) | ( n1641 & n12008 ) | ( n5144 & n12008 ) ;
  assign n15099 = ( n861 & ~n12531 ) | ( n861 & n15098 ) | ( ~n12531 & n15098 ) ;
  assign n15100 = ~n1320 & n7454 ;
  assign n15101 = ~n7746 & n15100 ;
  assign n15102 = ~n6931 & n15101 ;
  assign n15103 = n11062 & n14268 ;
  assign n15104 = ~n12050 & n15103 ;
  assign n15105 = n12309 | n15104 ;
  assign n15106 = n15105 ^ n725 ^ 1'b0 ;
  assign n15107 = n7939 ^ n4405 ^ n1493 ;
  assign n15108 = n4351 | n15107 ;
  assign n15109 = n269 | n3719 ;
  assign n15110 = ( n2098 & n10613 ) | ( n2098 & n15109 ) | ( n10613 & n15109 ) ;
  assign n15111 = n9739 ^ n3609 ^ 1'b0 ;
  assign n15112 = n15110 | n15111 ;
  assign n15113 = n15108 & ~n15112 ;
  assign n15114 = n10375 ^ n9611 ^ 1'b0 ;
  assign n15115 = ~n2570 & n15114 ;
  assign n15116 = ( ~n2003 & n9099 ) | ( ~n2003 & n15115 ) | ( n9099 & n15115 ) ;
  assign n15117 = n11188 ^ n11044 ^ 1'b0 ;
  assign n15118 = n10332 & ~n15117 ;
  assign n15119 = n5628 | n9160 ;
  assign n15120 = n15118 | n15119 ;
  assign n15121 = n4071 ^ n352 ^ 1'b0 ;
  assign n15122 = n3705 | n6913 ;
  assign n15123 = n15121 | n15122 ;
  assign n15124 = n4689 ^ n1956 ^ 1'b0 ;
  assign n15125 = n1071 | n15124 ;
  assign n15126 = ( n1382 & n5050 ) | ( n1382 & n15125 ) | ( n5050 & n15125 ) ;
  assign n15129 = ~n7425 & n11100 ;
  assign n15130 = n1586 & n15129 ;
  assign n15131 = n6091 & n15130 ;
  assign n15132 = n15131 ^ n8250 ^ 1'b0 ;
  assign n15128 = n10683 ^ n8331 ^ 1'b0 ;
  assign n15127 = n9566 ^ n2363 ^ 1'b0 ;
  assign n15133 = n15132 ^ n15128 ^ n15127 ;
  assign n15134 = n15133 ^ n9745 ^ n3433 ;
  assign n15135 = x84 | n7196 ;
  assign n15136 = n15135 ^ n8228 ^ 1'b0 ;
  assign n15137 = n2799 & n5316 ;
  assign n15139 = n3191 ^ n1314 ^ 1'b0 ;
  assign n15140 = n15139 ^ n2155 ^ 1'b0 ;
  assign n15141 = n5133 & ~n15140 ;
  assign n15138 = n11972 ^ n10072 ^ n3640 ;
  assign n15142 = n15141 ^ n15138 ^ n2362 ;
  assign n15143 = n12425 & n12842 ;
  assign n15144 = n3517 ^ n2909 ^ 1'b0 ;
  assign n15145 = x42 & n15144 ;
  assign n15146 = n9859 & n15145 ;
  assign n15147 = n15146 ^ n14986 ^ 1'b0 ;
  assign n15152 = n14243 ^ n1536 ^ 1'b0 ;
  assign n15153 = n3020 & n15152 ;
  assign n15154 = n15153 ^ n7707 ^ 1'b0 ;
  assign n15148 = ( n2769 & n9257 ) | ( n2769 & n11099 ) | ( n9257 & n11099 ) ;
  assign n15149 = n15148 ^ n966 ^ 1'b0 ;
  assign n15150 = n2418 ^ n915 ^ 1'b0 ;
  assign n15151 = n15149 & ~n15150 ;
  assign n15155 = n15154 ^ n15151 ^ 1'b0 ;
  assign n15156 = n14553 ^ n8626 ^ x209 ;
  assign n15157 = n3899 | n15156 ;
  assign n15158 = n8073 & n12632 ;
  assign n15159 = n15158 ^ n12315 ^ 1'b0 ;
  assign n15160 = ~n10616 & n15159 ;
  assign n15161 = ( n4677 & n9378 ) | ( n4677 & ~n15160 ) | ( n9378 & ~n15160 ) ;
  assign n15162 = n3500 ^ n3054 ^ n1895 ;
  assign n15163 = n763 & n15162 ;
  assign n15164 = ( ~n7028 & n8780 ) | ( ~n7028 & n15163 ) | ( n8780 & n15163 ) ;
  assign n15165 = n9682 ^ n374 ^ 1'b0 ;
  assign n15166 = ~n8500 & n15165 ;
  assign n15167 = ~n5666 & n10836 ;
  assign n15168 = n4061 ^ n1149 ^ 1'b0 ;
  assign n15169 = n3096 & ~n13246 ;
  assign n15170 = ( n2169 & ~n6191 ) | ( n2169 & n13634 ) | ( ~n6191 & n13634 ) ;
  assign n15171 = ( n308 & n5181 ) | ( n308 & n11152 ) | ( n5181 & n11152 ) ;
  assign n15172 = n9879 & ~n15171 ;
  assign n15173 = n2921 & n15172 ;
  assign n15174 = n10058 ^ n5686 ^ 1'b0 ;
  assign n15175 = n15174 ^ n13890 ^ 1'b0 ;
  assign n15183 = n549 | n5949 ;
  assign n15176 = n3738 & ~n3865 ;
  assign n15177 = n4709 & n15176 ;
  assign n15178 = n10888 | n15177 ;
  assign n15179 = n15178 ^ n3398 ^ 1'b0 ;
  assign n15180 = n15179 ^ n10757 ^ n1142 ;
  assign n15181 = ~n6223 & n15180 ;
  assign n15182 = n15181 ^ n3474 ^ 1'b0 ;
  assign n15184 = n15183 ^ n15182 ^ 1'b0 ;
  assign n15185 = n3021 & ~n5156 ;
  assign n15186 = n15185 ^ n6386 ^ n3235 ;
  assign n15187 = n5157 | n15186 ;
  assign n15188 = n14030 ^ n11203 ^ n9795 ;
  assign n15189 = ( n3444 & n4592 ) | ( n3444 & n15188 ) | ( n4592 & n15188 ) ;
  assign n15190 = ~n1115 & n5110 ;
  assign n15191 = n15190 ^ n2336 ^ 1'b0 ;
  assign n15192 = n15191 ^ n14869 ^ 1'b0 ;
  assign n15194 = n5199 & n14936 ;
  assign n15195 = ~n4184 & n15194 ;
  assign n15193 = n4501 | n12312 ;
  assign n15196 = n15195 ^ n15193 ^ 1'b0 ;
  assign n15197 = n7796 & n15132 ;
  assign n15198 = n15196 & n15197 ;
  assign n15201 = n6854 ^ n3692 ^ 1'b0 ;
  assign n15199 = n2670 & n6832 ;
  assign n15200 = n15199 ^ n5935 ^ 1'b0 ;
  assign n15202 = n15201 ^ n15200 ^ n1370 ;
  assign n15203 = n10046 ^ n4971 ^ n4285 ;
  assign n15204 = n15203 ^ n13987 ^ n4162 ;
  assign n15205 = n737 | n8323 ;
  assign n15206 = ( n906 & n9149 ) | ( n906 & ~n13104 ) | ( n9149 & ~n13104 ) ;
  assign n15207 = ~n269 & n14381 ;
  assign n15208 = n15207 ^ n5021 ^ 1'b0 ;
  assign n15209 = n3108 ^ n2878 ^ 1'b0 ;
  assign n15210 = n15208 | n15209 ;
  assign n15211 = n2367 ^ n1446 ^ 1'b0 ;
  assign n15212 = n6292 ^ n2319 ^ 1'b0 ;
  assign n15213 = ~n1209 & n15212 ;
  assign n15214 = ~n6710 & n15213 ;
  assign n15215 = n15211 & n15214 ;
  assign n15216 = ~n10304 & n15215 ;
  assign n15217 = n15216 ^ n9381 ^ 1'b0 ;
  assign n15220 = n794 & n5138 ;
  assign n15221 = ~n6145 & n15220 ;
  assign n15222 = n15221 ^ n6430 ^ x86 ;
  assign n15218 = n11347 ^ n7734 ^ 1'b0 ;
  assign n15219 = n15218 ^ n2733 ^ 1'b0 ;
  assign n15223 = n15222 ^ n15219 ^ 1'b0 ;
  assign n15224 = n3674 ^ n2697 ^ 1'b0 ;
  assign n15229 = x57 & x224 ;
  assign n15225 = ( n3316 & n7848 ) | ( n3316 & ~n11979 ) | ( n7848 & ~n11979 ) ;
  assign n15226 = n15225 ^ n15027 ^ n2807 ;
  assign n15227 = n11105 & n15226 ;
  assign n15228 = n9158 & n15227 ;
  assign n15230 = n15229 ^ n15228 ^ 1'b0 ;
  assign n15231 = n3422 & n5723 ;
  assign n15232 = ~n5723 & n15231 ;
  assign n15233 = x37 & x226 ;
  assign n15234 = ~x226 & n15233 ;
  assign n15235 = n15234 ^ n6728 ^ 1'b0 ;
  assign n15237 = ~n5226 & n5945 ;
  assign n15238 = n2702 & n15237 ;
  assign n15239 = ~x24 & n15238 ;
  assign n15236 = n5025 & n5612 ;
  assign n15240 = n15239 ^ n15236 ^ 1'b0 ;
  assign n15241 = ~n15235 & n15240 ;
  assign n15242 = n15232 & n15241 ;
  assign n15243 = n11203 | n15242 ;
  assign n15244 = n11203 & ~n15243 ;
  assign n15245 = n2418 & ~n8407 ;
  assign n15246 = n15245 ^ n4011 ^ 1'b0 ;
  assign n15247 = n7697 & ~n15246 ;
  assign n15248 = ~n1007 & n15247 ;
  assign n15249 = n3148 & ~n6103 ;
  assign n15250 = n1757 & n15249 ;
  assign n15251 = n13888 ^ n10854 ^ 1'b0 ;
  assign n15252 = n12569 | n15251 ;
  assign n15253 = n15250 | n15252 ;
  assign n15254 = n15253 ^ n4518 ^ 1'b0 ;
  assign n15255 = n15014 ^ n7694 ^ 1'b0 ;
  assign n15256 = n2509 ^ x77 ^ 1'b0 ;
  assign n15257 = ( n6050 & n13606 ) | ( n6050 & n15256 ) | ( n13606 & n15256 ) ;
  assign n15258 = ( ~n5345 & n14449 ) | ( ~n5345 & n15257 ) | ( n14449 & n15257 ) ;
  assign n15259 = n663 & n2974 ;
  assign n15260 = n11462 & n15259 ;
  assign n15261 = n15260 ^ n13592 ^ n6571 ;
  assign n15262 = n3083 ^ x187 ^ 1'b0 ;
  assign n15263 = x102 & ~n15262 ;
  assign n15264 = n6776 ^ n989 ^ 1'b0 ;
  assign n15265 = ~n3409 & n12194 ;
  assign n15266 = n2723 & n15265 ;
  assign n15267 = ( n5928 & n15264 ) | ( n5928 & n15266 ) | ( n15264 & n15266 ) ;
  assign n15268 = n15267 ^ n284 ^ 1'b0 ;
  assign n15269 = n15263 & ~n15268 ;
  assign n15270 = n15269 ^ n14960 ^ 1'b0 ;
  assign n15271 = n12630 ^ n1084 ^ 1'b0 ;
  assign n15272 = n4516 & n4621 ;
  assign n15273 = ~n663 & n9245 ;
  assign n15274 = n15273 ^ n14654 ^ n5172 ;
  assign n15275 = n6493 & n12385 ;
  assign n15276 = n280 | n2826 ;
  assign n15277 = x236 & ~n14382 ;
  assign n15278 = ~n7978 & n15277 ;
  assign n15279 = n15278 ^ n3984 ^ 1'b0 ;
  assign n15280 = n3059 & n5342 ;
  assign n15281 = n9115 | n12911 ;
  assign n15282 = n15281 ^ n7711 ^ 1'b0 ;
  assign n15283 = ( n3342 & n15280 ) | ( n3342 & n15282 ) | ( n15280 & n15282 ) ;
  assign n15284 = n15283 ^ n5412 ^ 1'b0 ;
  assign n15285 = n4701 & n15284 ;
  assign n15286 = n4729 | n8465 ;
  assign n15287 = n1463 & ~n15286 ;
  assign n15288 = n11426 | n15287 ;
  assign n15289 = ( n800 & n8467 ) | ( n800 & ~n9643 ) | ( n8467 & ~n9643 ) ;
  assign n15291 = ~n978 & n6618 ;
  assign n15290 = n14112 ^ n6556 ^ 1'b0 ;
  assign n15292 = n15291 ^ n15290 ^ 1'b0 ;
  assign n15293 = ( n4233 & n14116 ) | ( n4233 & ~n15292 ) | ( n14116 & ~n15292 ) ;
  assign n15294 = n7839 ^ n3331 ^ n1327 ;
  assign n15295 = n861 | n12886 ;
  assign n15296 = ~n2372 & n12121 ;
  assign n15297 = ~n1079 & n1921 ;
  assign n15298 = ~n3796 & n15297 ;
  assign n15299 = n12801 & n15298 ;
  assign n15300 = ( ~n848 & n4419 ) | ( ~n848 & n7047 ) | ( n4419 & n7047 ) ;
  assign n15301 = ~n7225 & n15300 ;
  assign n15302 = ~n7550 & n15301 ;
  assign n15303 = ( ~n1934 & n8213 ) | ( ~n1934 & n15302 ) | ( n8213 & n15302 ) ;
  assign n15304 = n2219 & n8837 ;
  assign n15305 = n15304 ^ n561 ^ 1'b0 ;
  assign n15306 = n15305 ^ n14815 ^ 1'b0 ;
  assign n15307 = ( n1736 & n11486 ) | ( n1736 & n14164 ) | ( n11486 & n14164 ) ;
  assign n15308 = n5199 & n11173 ;
  assign n15309 = n15308 ^ n14911 ^ 1'b0 ;
  assign n15311 = n7317 ^ n391 ^ 1'b0 ;
  assign n15310 = n3317 | n7604 ;
  assign n15312 = n15311 ^ n15310 ^ 1'b0 ;
  assign n15313 = n3051 & ~n10659 ;
  assign n15314 = n15313 ^ n3677 ^ 1'b0 ;
  assign n15315 = n15312 & ~n15314 ;
  assign n15320 = n2448 ^ n402 ^ x171 ;
  assign n15316 = n9967 ^ n6926 ^ 1'b0 ;
  assign n15317 = n1134 & n4189 ;
  assign n15318 = n15316 | n15317 ;
  assign n15319 = ~n14634 & n15318 ;
  assign n15321 = n15320 ^ n15319 ^ 1'b0 ;
  assign n15322 = ~n9261 & n12872 ;
  assign n15323 = n15322 ^ n12402 ^ 1'b0 ;
  assign n15324 = n1940 & ~n7307 ;
  assign n15325 = ~n6188 & n15324 ;
  assign n15326 = n15325 ^ n14946 ^ n8524 ;
  assign n15327 = n10894 & ~n14351 ;
  assign n15329 = n2914 & ~n6863 ;
  assign n15328 = n1951 | n8486 ;
  assign n15330 = n15329 ^ n15328 ^ 1'b0 ;
  assign n15331 = n7484 ^ n5993 ^ 1'b0 ;
  assign n15332 = n12693 & n15331 ;
  assign n15333 = n15332 ^ n8696 ^ 1'b0 ;
  assign n15334 = ~n3738 & n4572 ;
  assign n15335 = n8212 & n11972 ;
  assign n15336 = ( n1725 & ~n2754 ) | ( n1725 & n15335 ) | ( ~n2754 & n15335 ) ;
  assign n15337 = n1766 & n15336 ;
  assign n15338 = n15334 & n15337 ;
  assign n15339 = ~x157 & n12474 ;
  assign n15340 = n15339 ^ n2572 ^ 1'b0 ;
  assign n15341 = n15340 ^ n1661 ^ 1'b0 ;
  assign n15342 = n3705 | n8947 ;
  assign n15343 = ~x153 & n6294 ;
  assign n15344 = n15343 ^ n4616 ^ n3358 ;
  assign n15345 = ~n11680 & n15344 ;
  assign n15346 = n11422 ^ n9642 ^ 1'b0 ;
  assign n15348 = n5500 | n13665 ;
  assign n15347 = ( ~n1898 & n3188 ) | ( ~n1898 & n3700 ) | ( n3188 & n3700 ) ;
  assign n15349 = n15348 ^ n15347 ^ 1'b0 ;
  assign n15350 = ~n15346 & n15349 ;
  assign n15352 = n660 & n11758 ;
  assign n15353 = n15352 ^ n1363 ^ 1'b0 ;
  assign n15351 = n8609 ^ n1709 ^ x82 ;
  assign n15354 = n15353 ^ n15351 ^ 1'b0 ;
  assign n15355 = n5860 & ~n15354 ;
  assign n15356 = n11381 & ~n15355 ;
  assign n15357 = n11985 | n15356 ;
  assign n15358 = n5947 ^ n1035 ^ 1'b0 ;
  assign n15359 = n9924 & n15358 ;
  assign n15360 = n15359 ^ n7971 ^ 1'b0 ;
  assign n15361 = n15360 ^ n15356 ^ n1090 ;
  assign n15362 = n4193 | n15361 ;
  assign n15363 = n4901 | n15362 ;
  assign n15364 = ~n13548 & n15363 ;
  assign n15365 = n8278 ^ n6358 ^ 1'b0 ;
  assign n15366 = n13414 | n15365 ;
  assign n15367 = n15366 ^ n4561 ^ 1'b0 ;
  assign n15368 = n3148 & n15367 ;
  assign n15369 = n1088 & ~n11798 ;
  assign n15370 = n11100 ^ n4705 ^ n3941 ;
  assign n15371 = n15370 ^ n10659 ^ n944 ;
  assign n15372 = n15371 ^ n339 ^ 1'b0 ;
  assign n15373 = n12544 & n15372 ;
  assign n15374 = n5536 | n6941 ;
  assign n15375 = n2192 | n15374 ;
  assign n15376 = n13756 ^ n7235 ^ 1'b0 ;
  assign n15377 = n14563 ^ n8812 ^ 1'b0 ;
  assign n15378 = ~n15376 & n15377 ;
  assign n15379 = n15378 ^ n7522 ^ n3669 ;
  assign n15380 = ( n1321 & n2787 ) | ( n1321 & ~n15379 ) | ( n2787 & ~n15379 ) ;
  assign n15381 = x123 & n9430 ;
  assign n15382 = n3615 & n15381 ;
  assign n15383 = n7956 ^ n6588 ^ 1'b0 ;
  assign n15384 = n4217 & n11332 ;
  assign n15385 = n1058 & n6950 ;
  assign n15386 = n447 & ~n3401 ;
  assign n15387 = ~n13398 & n15386 ;
  assign n15388 = n12853 ^ n9444 ^ 1'b0 ;
  assign n15389 = ~n5749 & n8763 ;
  assign n15390 = ~n391 & n15389 ;
  assign n15392 = n2032 | n6275 ;
  assign n15391 = n9163 ^ n8026 ^ 1'b0 ;
  assign n15393 = n15392 ^ n15391 ^ n7975 ;
  assign n15394 = n9569 ^ n843 ^ 1'b0 ;
  assign n15395 = n15394 ^ n4512 ^ n1987 ;
  assign n15400 = n8409 | n8932 ;
  assign n15401 = x194 | n15400 ;
  assign n15402 = n15401 ^ n6047 ^ 1'b0 ;
  assign n15396 = n4945 ^ n3123 ^ 1'b0 ;
  assign n15397 = n3358 | n15396 ;
  assign n15398 = ( n4260 & n4939 ) | ( n4260 & ~n15397 ) | ( n4939 & ~n15397 ) ;
  assign n15399 = n14967 & ~n15398 ;
  assign n15403 = n15402 ^ n15399 ^ 1'b0 ;
  assign n15404 = n7641 ^ n2055 ^ 1'b0 ;
  assign n15405 = n7238 & n15404 ;
  assign n15406 = ( n2502 & n5364 ) | ( n2502 & ~n14314 ) | ( n5364 & ~n14314 ) ;
  assign n15407 = ( n1285 & n3883 ) | ( n1285 & ~n6043 ) | ( n3883 & ~n6043 ) ;
  assign n15408 = n15407 ^ n9885 ^ 1'b0 ;
  assign n15409 = ~n14829 & n15408 ;
  assign n15410 = n1250 & ~n8149 ;
  assign n15411 = ( n3683 & n10298 ) | ( n3683 & n15410 ) | ( n10298 & n15410 ) ;
  assign n15412 = n15411 ^ n12597 ^ 1'b0 ;
  assign n15413 = n1981 | n15412 ;
  assign n15416 = n6121 & ~n14091 ;
  assign n15414 = ( n4754 & n9806 ) | ( n4754 & ~n14502 ) | ( n9806 & ~n14502 ) ;
  assign n15415 = ( n1505 & ~n8311 ) | ( n1505 & n15414 ) | ( ~n8311 & n15414 ) ;
  assign n15417 = n15416 ^ n15415 ^ n11008 ;
  assign n15418 = ~n5528 & n9799 ;
  assign n15419 = n8700 | n15418 ;
  assign n15420 = n3784 | n15419 ;
  assign n15421 = n8360 & ~n10330 ;
  assign n15422 = n4730 & n8341 ;
  assign n15423 = n15421 & n15422 ;
  assign n15424 = n2058 ^ n1487 ^ 1'b0 ;
  assign n15425 = n8828 ^ n3274 ^ 1'b0 ;
  assign n15426 = n5632 & ~n15425 ;
  assign n15427 = n5445 ^ n1999 ^ 1'b0 ;
  assign n15428 = n15426 & n15427 ;
  assign n15429 = n12175 ^ n3250 ^ 1'b0 ;
  assign n15430 = ~n4469 & n11822 ;
  assign n15431 = n15430 ^ n10839 ^ n967 ;
  assign n15432 = ( ~n15428 & n15429 ) | ( ~n15428 & n15431 ) | ( n15429 & n15431 ) ;
  assign n15433 = n7490 | n14089 ;
  assign n15434 = n10299 & ~n15433 ;
  assign n15435 = n15434 ^ n873 ^ 1'b0 ;
  assign n15436 = ( n3458 & n3731 ) | ( n3458 & n7760 ) | ( n3731 & n7760 ) ;
  assign n15437 = n15436 ^ n12343 ^ 1'b0 ;
  assign n15438 = n10542 & ~n15437 ;
  assign n15439 = n15438 ^ n7785 ^ 1'b0 ;
  assign n15440 = n6695 & ~n15439 ;
  assign n15441 = n12642 | n13769 ;
  assign n15442 = n4481 | n15441 ;
  assign n15444 = n3016 & n11128 ;
  assign n15445 = n15444 ^ n3880 ^ 1'b0 ;
  assign n15443 = n13833 ^ n5679 ^ 1'b0 ;
  assign n15446 = n15445 ^ n15443 ^ 1'b0 ;
  assign n15447 = n1909 & n15446 ;
  assign n15448 = ( n535 & n970 ) | ( n535 & ~n4515 ) | ( n970 & ~n4515 ) ;
  assign n15449 = n4067 | n14116 ;
  assign n15450 = ( x251 & n15448 ) | ( x251 & n15449 ) | ( n15448 & n15449 ) ;
  assign n15451 = n12111 ^ n472 ^ 1'b0 ;
  assign n15453 = n12919 & n13841 ;
  assign n15454 = ~n12919 & n15453 ;
  assign n15452 = n10767 & ~n14480 ;
  assign n15455 = n15454 ^ n15452 ^ 1'b0 ;
  assign n15456 = n1024 ^ n718 ^ 1'b0 ;
  assign n15457 = ( n2185 & ~n7484 ) | ( n2185 & n11651 ) | ( ~n7484 & n11651 ) ;
  assign n15458 = n4975 & ~n14807 ;
  assign n15459 = ~n15211 & n15458 ;
  assign n15460 = n14589 ^ n711 ^ 1'b0 ;
  assign n15461 = ~n6524 & n15460 ;
  assign n15462 = ( n3444 & n3938 ) | ( n3444 & n12877 ) | ( n3938 & n12877 ) ;
  assign n15463 = n13605 ^ n9014 ^ 1'b0 ;
  assign n15464 = n15462 | n15463 ;
  assign n15465 = ( n3157 & n8525 ) | ( n3157 & n12032 ) | ( n8525 & n12032 ) ;
  assign n15466 = ~n5875 & n15465 ;
  assign n15469 = n870 & ~n10629 ;
  assign n15467 = n7998 ^ n3804 ^ 1'b0 ;
  assign n15468 = ~n7378 & n15467 ;
  assign n15470 = n15469 ^ n15468 ^ 1'b0 ;
  assign n15471 = n7399 & n15470 ;
  assign n15472 = n12333 & n15471 ;
  assign n15473 = ( n1698 & ~n2004 ) | ( n1698 & n8937 ) | ( ~n2004 & n8937 ) ;
  assign n15474 = ( x183 & ~n4715 ) | ( x183 & n15473 ) | ( ~n4715 & n15473 ) ;
  assign n15475 = n3724 ^ n3121 ^ 1'b0 ;
  assign n15476 = n8041 ^ n5761 ^ 1'b0 ;
  assign n15477 = n13291 | n15476 ;
  assign n15478 = ~n2892 & n5725 ;
  assign n15479 = n15478 ^ n12792 ^ 1'b0 ;
  assign n15480 = n13270 & n15479 ;
  assign n15481 = ~n3324 & n7743 ;
  assign n15482 = n15481 ^ n8700 ^ 1'b0 ;
  assign n15483 = n4788 & n6511 ;
  assign n15484 = n15482 & ~n15483 ;
  assign n15485 = ( n6851 & ~n9086 ) | ( n6851 & n9582 ) | ( ~n9086 & n9582 ) ;
  assign n15486 = n12046 & ~n12575 ;
  assign n15487 = n15485 | n15486 ;
  assign n15488 = n9311 ^ n913 ^ 1'b0 ;
  assign n15489 = n12566 & ~n15488 ;
  assign n15490 = n10854 & ~n15489 ;
  assign n15491 = n4835 | n5118 ;
  assign n15492 = n10690 ^ n7851 ^ 1'b0 ;
  assign n15493 = n13357 & ~n15492 ;
  assign n15494 = n5381 ^ n2951 ^ 1'b0 ;
  assign n15495 = n9707 ^ n7732 ^ 1'b0 ;
  assign n15496 = n12674 | n15495 ;
  assign n15497 = ~n621 & n7457 ;
  assign n15498 = n5905 | n8085 ;
  assign n15499 = n15498 ^ n7736 ^ 1'b0 ;
  assign n15500 = n11500 ^ n7364 ^ 1'b0 ;
  assign n15501 = ~n15499 & n15500 ;
  assign n15502 = n4417 ^ n2939 ^ 1'b0 ;
  assign n15503 = n2083 & n15502 ;
  assign n15504 = n6295 ^ n838 ^ 1'b0 ;
  assign n15505 = n10662 ^ n8622 ^ n3256 ;
  assign n15506 = n14293 & ~n15505 ;
  assign n15507 = ( x141 & ~n3360 ) | ( x141 & n3589 ) | ( ~n3360 & n3589 ) ;
  assign n15508 = n6875 & n15507 ;
  assign n15509 = n11625 ^ n6375 ^ n3440 ;
  assign n15510 = n3731 & n15509 ;
  assign n15511 = n12648 & n15510 ;
  assign n15512 = n4519 & ~n10739 ;
  assign n15513 = n7480 ^ n2421 ^ 1'b0 ;
  assign n15514 = n2253 | n15513 ;
  assign n15515 = ~n3856 & n3994 ;
  assign n15516 = n15515 ^ n15373 ^ n2995 ;
  assign n15519 = ( n665 & n1809 ) | ( n665 & n13454 ) | ( n1809 & n13454 ) ;
  assign n15517 = ( n530 & n4614 ) | ( n530 & n8213 ) | ( n4614 & n8213 ) ;
  assign n15518 = n5569 | n15517 ;
  assign n15520 = n15519 ^ n15518 ^ 1'b0 ;
  assign n15521 = n9685 ^ n2463 ^ 1'b0 ;
  assign n15522 = ~n1893 & n15521 ;
  assign n15523 = n8103 ^ x37 ^ 1'b0 ;
  assign n15524 = n15522 & ~n15523 ;
  assign n15525 = ( ~n9108 & n15520 ) | ( ~n9108 & n15524 ) | ( n15520 & n15524 ) ;
  assign n15526 = n8991 ^ n4472 ^ 1'b0 ;
  assign n15527 = n15526 ^ n4767 ^ n2441 ;
  assign n15528 = n6028 & ~n15527 ;
  assign n15529 = n12312 ^ n9743 ^ n9008 ;
  assign n15530 = n15529 ^ n7839 ^ 1'b0 ;
  assign n15531 = n1893 | n4437 ;
  assign n15532 = n15531 ^ n12423 ^ 1'b0 ;
  assign n15534 = ~n6221 & n11774 ;
  assign n15533 = n8808 ^ n1529 ^ 1'b0 ;
  assign n15535 = n15534 ^ n15533 ^ 1'b0 ;
  assign n15536 = n2740 ^ n2092 ^ 1'b0 ;
  assign n15537 = n15536 ^ n11023 ^ n305 ;
  assign n15538 = n1257 | n3792 ;
  assign n15539 = n15538 ^ n8845 ^ 1'b0 ;
  assign n15540 = n15539 ^ n9379 ^ 1'b0 ;
  assign n15541 = n1061 & n9869 ;
  assign n15542 = n6364 & n15541 ;
  assign n15543 = ( n5376 & ~n15540 ) | ( n5376 & n15542 ) | ( ~n15540 & n15542 ) ;
  assign n15544 = n5451 & n7111 ;
  assign n15545 = n3083 & ~n15544 ;
  assign n15546 = n1265 & ~n11673 ;
  assign n15547 = n11368 ^ n2845 ^ n2375 ;
  assign n15548 = n15311 & n15547 ;
  assign n15549 = n1533 & n15548 ;
  assign n15550 = ( ~n1908 & n6114 ) | ( ~n1908 & n6983 ) | ( n6114 & n6983 ) ;
  assign n15551 = ~n642 & n7808 ;
  assign n15552 = ~n15550 & n15551 ;
  assign n15553 = ~n6610 & n15552 ;
  assign n15554 = n9325 | n10427 ;
  assign n15555 = n3254 & ~n15554 ;
  assign n15556 = n702 & n2722 ;
  assign n15557 = n8991 & ~n10178 ;
  assign n15558 = n6442 | n12848 ;
  assign n15559 = n14168 | n15558 ;
  assign n15560 = n15559 ^ n1197 ^ 1'b0 ;
  assign n15561 = n2439 & n5397 ;
  assign n15562 = n15561 ^ n2012 ^ 1'b0 ;
  assign n15563 = n15562 ^ n10313 ^ n8254 ;
  assign n15564 = n2114 ^ n1958 ^ n1514 ;
  assign n15565 = ( n2287 & n6786 ) | ( n2287 & n7335 ) | ( n6786 & n7335 ) ;
  assign n15566 = n1018 & ~n2682 ;
  assign n15567 = n489 & n15566 ;
  assign n15568 = n15567 ^ n10506 ^ n2499 ;
  assign n15569 = ( n2529 & n15565 ) | ( n2529 & ~n15568 ) | ( n15565 & ~n15568 ) ;
  assign n15577 = ( ~n1433 & n7077 ) | ( ~n1433 & n7674 ) | ( n7077 & n7674 ) ;
  assign n15575 = ~x133 & x171 ;
  assign n15576 = n15575 ^ n4544 ^ n2098 ;
  assign n15573 = n5151 ^ n4034 ^ 1'b0 ;
  assign n15574 = n15573 ^ n7317 ^ n3669 ;
  assign n15578 = n15577 ^ n15576 ^ n15574 ;
  assign n15571 = n4525 ^ n1634 ^ 1'b0 ;
  assign n15570 = n885 | n10424 ;
  assign n15572 = n15571 ^ n15570 ^ 1'b0 ;
  assign n15579 = n15578 ^ n15572 ^ n11093 ;
  assign n15580 = n15579 ^ n6524 ^ n2573 ;
  assign n15581 = n12134 | n12312 ;
  assign n15582 = n15581 ^ n3274 ^ 1'b0 ;
  assign n15588 = n981 & ~n6913 ;
  assign n15583 = ~n4946 & n5819 ;
  assign n15584 = n15583 ^ n6824 ^ 1'b0 ;
  assign n15585 = n2030 & ~n15584 ;
  assign n15586 = n15585 ^ n647 ^ 1'b0 ;
  assign n15587 = n8896 & ~n15586 ;
  assign n15589 = n15588 ^ n15587 ^ 1'b0 ;
  assign n15590 = n13947 ^ n1615 ^ 1'b0 ;
  assign n15591 = n6889 & ~n15590 ;
  assign n15592 = ( n11103 & n11469 ) | ( n11103 & n14804 ) | ( n11469 & n14804 ) ;
  assign n15593 = n6371 ^ n4148 ^ 1'b0 ;
  assign n15594 = n10080 & n15593 ;
  assign n15595 = ~n7502 & n9765 ;
  assign n15596 = ~n15594 & n15595 ;
  assign n15597 = ( n5949 & n13643 ) | ( n5949 & ~n15596 ) | ( n13643 & ~n15596 ) ;
  assign n15598 = n2854 & n13201 ;
  assign n15599 = n15598 ^ n13114 ^ 1'b0 ;
  assign n15600 = n6971 ^ n2292 ^ 1'b0 ;
  assign n15601 = n13626 & n15600 ;
  assign n15602 = ~n6256 & n15601 ;
  assign n15603 = n15602 ^ n2586 ^ 1'b0 ;
  assign n15607 = n3007 & ~n5609 ;
  assign n15604 = ~n2329 & n5685 ;
  assign n15605 = n10837 ^ n293 ^ 1'b0 ;
  assign n15606 = ~n15604 & n15605 ;
  assign n15608 = n15607 ^ n15606 ^ n1939 ;
  assign n15609 = n13789 & n15608 ;
  assign n15610 = n9929 & n13733 ;
  assign n15611 = n15610 ^ n4408 ^ 1'b0 ;
  assign n15612 = n3091 & n11229 ;
  assign n15613 = n10135 & n15612 ;
  assign n15614 = n4912 | n15613 ;
  assign n15615 = n513 | n4847 ;
  assign n15617 = n6989 ^ n1019 ^ n503 ;
  assign n15616 = ~n8798 & n14155 ;
  assign n15618 = n15617 ^ n15616 ^ 1'b0 ;
  assign n15619 = n12715 ^ n4303 ^ 1'b0 ;
  assign n15620 = n10052 ^ n2042 ^ 1'b0 ;
  assign n15621 = ( n288 & n425 ) | ( n288 & ~n8471 ) | ( n425 & ~n8471 ) ;
  assign n15622 = n15621 ^ n14206 ^ 1'b0 ;
  assign n15623 = n8909 | n15622 ;
  assign n15624 = n9620 | n15623 ;
  assign n15625 = n15624 ^ n11264 ^ 1'b0 ;
  assign n15626 = n14960 & ~n15625 ;
  assign n15627 = n6159 ^ n1626 ^ 1'b0 ;
  assign n15628 = n7985 & n15627 ;
  assign n15629 = n10510 ^ n3640 ^ 1'b0 ;
  assign n15630 = ~n1724 & n4502 ;
  assign n15631 = n1248 | n15630 ;
  assign n15632 = n10357 | n15631 ;
  assign n15633 = n15629 & n15632 ;
  assign n15634 = ~n9958 & n15633 ;
  assign n15635 = n13757 ^ n7502 ^ 1'b0 ;
  assign n15636 = ( n4937 & n9483 ) | ( n4937 & ~n15635 ) | ( n9483 & ~n15635 ) ;
  assign n15648 = n3404 | n8670 ;
  assign n15637 = n1392 | n8263 ;
  assign n15638 = n15637 ^ n5741 ^ 1'b0 ;
  assign n15639 = x18 & ~n15638 ;
  assign n15640 = n15639 ^ n9561 ^ 1'b0 ;
  assign n15644 = n4047 | n10346 ;
  assign n15645 = n15644 ^ n3328 ^ n1023 ;
  assign n15641 = n1156 | n7553 ;
  assign n15642 = n15641 ^ n545 ^ 1'b0 ;
  assign n15643 = n10514 & ~n15642 ;
  assign n15646 = n15645 ^ n15643 ^ 1'b0 ;
  assign n15647 = n15640 | n15646 ;
  assign n15649 = n15648 ^ n15647 ^ 1'b0 ;
  assign n15650 = n2578 & n9587 ;
  assign n15651 = n8582 ^ n2886 ^ 1'b0 ;
  assign n15652 = n5404 ^ n2945 ^ 1'b0 ;
  assign n15653 = n2687 & n13959 ;
  assign n15654 = ~n2001 & n15653 ;
  assign n15655 = n8553 & n8891 ;
  assign n15656 = n15655 ^ n14886 ^ 1'b0 ;
  assign n15657 = n15656 ^ n12818 ^ 1'b0 ;
  assign n15658 = n12820 | n15657 ;
  assign n15660 = n3683 & n4601 ;
  assign n15659 = n1067 & ~n1273 ;
  assign n15661 = n15660 ^ n15659 ^ 1'b0 ;
  assign n15662 = ( n10505 & ~n14128 ) | ( n10505 & n15661 ) | ( ~n14128 & n15661 ) ;
  assign n15663 = n6638 ^ n2414 ^ 1'b0 ;
  assign n15664 = n4947 | n15663 ;
  assign n15665 = n15664 ^ n3496 ^ 1'b0 ;
  assign n15666 = n6999 & n15568 ;
  assign n15667 = n5781 & n15666 ;
  assign n15668 = n15667 ^ n5056 ^ 1'b0 ;
  assign n15669 = n15668 ^ x131 ^ 1'b0 ;
  assign n15670 = ~n2133 & n5042 ;
  assign n15671 = n15670 ^ n2527 ^ 1'b0 ;
  assign n15672 = ( n2610 & n11527 ) | ( n2610 & ~n13326 ) | ( n11527 & ~n13326 ) ;
  assign n15673 = n15671 | n15672 ;
  assign n15674 = n15673 ^ n6627 ^ 1'b0 ;
  assign n15683 = n1472 & n7472 ;
  assign n15677 = n8028 ^ n5429 ^ 1'b0 ;
  assign n15678 = ( n2433 & n4255 ) | ( n2433 & n15677 ) | ( n4255 & n15677 ) ;
  assign n15679 = n15678 ^ n15130 ^ 1'b0 ;
  assign n15680 = ~n5642 & n15679 ;
  assign n15675 = ~n5642 & n9158 ;
  assign n15676 = n13163 & ~n15675 ;
  assign n15681 = n15680 ^ n15676 ^ 1'b0 ;
  assign n15682 = n4943 | n15681 ;
  assign n15684 = n15683 ^ n15682 ^ 1'b0 ;
  assign n15686 = n7426 ^ n2695 ^ n887 ;
  assign n15685 = ~n7627 & n12408 ;
  assign n15687 = n15686 ^ n15685 ^ 1'b0 ;
  assign n15688 = n8940 ^ n2068 ^ 1'b0 ;
  assign n15689 = ~n2282 & n15688 ;
  assign n15690 = ( ~n7028 & n15687 ) | ( ~n7028 & n15689 ) | ( n15687 & n15689 ) ;
  assign n15693 = n356 & n1685 ;
  assign n15694 = n6907 & n15693 ;
  assign n15695 = n15694 ^ n11488 ^ 1'b0 ;
  assign n15696 = n5420 & n15695 ;
  assign n15691 = ~n2847 & n6097 ;
  assign n15692 = n15691 ^ n10487 ^ 1'b0 ;
  assign n15697 = n15696 ^ n15692 ^ 1'b0 ;
  assign n15698 = n4326 | n15697 ;
  assign n15699 = n10734 ^ n1678 ^ 1'b0 ;
  assign n15700 = n3707 & ~n15699 ;
  assign n15701 = ~n4577 & n15700 ;
  assign n15702 = n6165 | n7280 ;
  assign n15703 = n1382 & ~n15702 ;
  assign n15704 = n15703 ^ n12670 ^ 1'b0 ;
  assign n15705 = n10101 | n11083 ;
  assign n15706 = n15704 & ~n15705 ;
  assign n15707 = n2468 & ~n6941 ;
  assign n15708 = ~n1501 & n15707 ;
  assign n15709 = n15708 ^ n8758 ^ 1'b0 ;
  assign n15710 = n469 | n10773 ;
  assign n15711 = n966 & ~n5115 ;
  assign n15712 = ~n10952 & n15711 ;
  assign n15713 = n14003 ^ n8025 ^ 1'b0 ;
  assign n15714 = n15712 | n15713 ;
  assign n15715 = ( n7958 & n15710 ) | ( n7958 & ~n15714 ) | ( n15710 & ~n15714 ) ;
  assign n15716 = n5438 ^ n1002 ^ 1'b0 ;
  assign n15717 = n3607 | n15716 ;
  assign n15718 = n3086 & n15717 ;
  assign n15723 = ~n4041 & n5374 ;
  assign n15724 = ~n8165 & n15723 ;
  assign n15722 = n11502 ^ n931 ^ 1'b0 ;
  assign n15719 = n8800 ^ n1598 ^ 1'b0 ;
  assign n15720 = n15719 ^ n7149 ^ 1'b0 ;
  assign n15721 = n15720 ^ n2661 ^ 1'b0 ;
  assign n15725 = n15724 ^ n15722 ^ n15721 ;
  assign n15730 = n1374 | n2319 ;
  assign n15731 = n13861 | n15730 ;
  assign n15726 = x133 & ~n322 ;
  assign n15727 = n15726 ^ n10990 ^ 1'b0 ;
  assign n15728 = ~n402 & n15727 ;
  assign n15729 = n2489 & n15728 ;
  assign n15732 = n15731 ^ n15729 ^ n8883 ;
  assign n15733 = n6106 ^ n1709 ^ 1'b0 ;
  assign n15734 = ~n2052 & n15733 ;
  assign n15735 = n15734 ^ n11940 ^ 1'b0 ;
  assign n15736 = n2052 & ~n3578 ;
  assign n15737 = n8654 & ~n10947 ;
  assign n15738 = n15737 ^ n13734 ^ 1'b0 ;
  assign n15739 = n2111 | n3404 ;
  assign n15740 = n2491 | n7695 ;
  assign n15741 = n15740 ^ n14512 ^ 1'b0 ;
  assign n15742 = ~n15739 & n15741 ;
  assign n15743 = n14490 & n15742 ;
  assign n15744 = ( n1161 & ~n4561 ) | ( n1161 & n6073 ) | ( ~n4561 & n6073 ) ;
  assign n15745 = n8248 & ~n15744 ;
  assign n15746 = ~n4210 & n7741 ;
  assign n15747 = ( n3727 & ~n7628 ) | ( n3727 & n15746 ) | ( ~n7628 & n15746 ) ;
  assign n15748 = ~n4112 & n15747 ;
  assign n15749 = n15745 & n15748 ;
  assign n15750 = ( x132 & n3071 ) | ( x132 & n15575 ) | ( n3071 & n15575 ) ;
  assign n15751 = ( ~n14386 & n14487 ) | ( ~n14386 & n15750 ) | ( n14487 & n15750 ) ;
  assign n15752 = n7720 ^ n2959 ^ 1'b0 ;
  assign n15753 = n13615 ^ n5791 ^ 1'b0 ;
  assign n15754 = n2468 & ~n15753 ;
  assign n15755 = n9232 ^ n6744 ^ n2466 ;
  assign n15756 = n2504 & n15755 ;
  assign n15757 = n15665 ^ n4919 ^ 1'b0 ;
  assign n15758 = n2709 & n6414 ;
  assign n15759 = n3821 & n15758 ;
  assign n15760 = n15759 ^ n13342 ^ 1'b0 ;
  assign n15761 = n2095 ^ n1213 ^ 1'b0 ;
  assign n15762 = n15761 ^ n10180 ^ 1'b0 ;
  assign n15763 = n15760 | n15762 ;
  assign n15764 = n15102 ^ n11115 ^ 1'b0 ;
  assign n15765 = n14108 & n15764 ;
  assign n15767 = n10970 ^ n9943 ^ 1'b0 ;
  assign n15766 = n3440 ^ n3331 ^ 1'b0 ;
  assign n15768 = n15767 ^ n15766 ^ 1'b0 ;
  assign n15771 = ~n3239 & n9866 ;
  assign n15772 = n15771 ^ n10940 ^ n879 ;
  assign n15769 = n6737 | n7840 ;
  assign n15770 = ( n1659 & ~n8760 ) | ( n1659 & n15769 ) | ( ~n8760 & n15769 ) ;
  assign n15773 = n15772 ^ n15770 ^ 1'b0 ;
  assign n15774 = ~n8505 & n15773 ;
  assign n15775 = n7830 & ~n12118 ;
  assign n15776 = n15775 ^ n7245 ^ 1'b0 ;
  assign n15777 = n745 & ~n2274 ;
  assign n15778 = n15777 ^ n13764 ^ 1'b0 ;
  assign n15779 = ( ~n7806 & n9500 ) | ( ~n7806 & n15778 ) | ( n9500 & n15778 ) ;
  assign n15780 = n3746 & n13111 ;
  assign n15781 = n2452 ^ x102 ^ 1'b0 ;
  assign n15782 = n3857 & ~n15781 ;
  assign n15783 = n3299 & n15782 ;
  assign n15784 = n15783 ^ n7464 ^ 1'b0 ;
  assign n15785 = n4056 ^ n554 ^ 1'b0 ;
  assign n15786 = n8431 & n15785 ;
  assign n15787 = n427 & n15786 ;
  assign n15788 = ( n5625 & ~n6467 ) | ( n5625 & n15787 ) | ( ~n6467 & n15787 ) ;
  assign n15789 = x68 & n15788 ;
  assign n15790 = n917 & n15789 ;
  assign n15791 = n831 | n3151 ;
  assign n15792 = n3466 | n15791 ;
  assign n15793 = n11891 ^ n1002 ^ 1'b0 ;
  assign n15794 = ( n3235 & n10902 ) | ( n3235 & n15793 ) | ( n10902 & n15793 ) ;
  assign n15795 = n11880 ^ n10323 ^ n4271 ;
  assign n15796 = n4308 & n6744 ;
  assign n15797 = ~n7976 & n12808 ;
  assign n15798 = n15797 ^ n326 ^ 1'b0 ;
  assign n15799 = n4430 ^ n3088 ^ n1639 ;
  assign n15802 = ( ~x122 & n3107 ) | ( ~x122 & n4022 ) | ( n3107 & n4022 ) ;
  assign n15800 = ( n2033 & ~n4390 ) | ( n2033 & n11953 ) | ( ~n4390 & n11953 ) ;
  assign n15801 = n5789 & ~n15800 ;
  assign n15803 = n15802 ^ n15801 ^ 1'b0 ;
  assign n15804 = ~n15799 & n15803 ;
  assign n15805 = n15804 ^ n10853 ^ 1'b0 ;
  assign n15806 = n2426 & ~n15805 ;
  assign n15807 = n4071 & n8181 ;
  assign n15808 = n7345 ^ n6283 ^ n2292 ;
  assign n15809 = n5318 & ~n15808 ;
  assign n15810 = n8247 & n15809 ;
  assign n15811 = ( ~n11753 & n15807 ) | ( ~n11753 & n15810 ) | ( n15807 & n15810 ) ;
  assign n15812 = n752 | n2226 ;
  assign n15813 = n5464 | n11533 ;
  assign n15814 = n15813 ^ n7535 ^ 1'b0 ;
  assign n15815 = n15812 & ~n15814 ;
  assign n15816 = n13089 ^ n6497 ^ n4425 ;
  assign n15817 = n292 & ~n922 ;
  assign n15818 = n15817 ^ n11663 ^ n1407 ;
  assign n15819 = ( ~n290 & n15816 ) | ( ~n290 & n15818 ) | ( n15816 & n15818 ) ;
  assign n15820 = ( n2571 & ~n4014 ) | ( n2571 & n15819 ) | ( ~n4014 & n15819 ) ;
  assign n15821 = n15820 ^ n11488 ^ 1'b0 ;
  assign n15822 = n1002 | n14133 ;
  assign n15823 = n15822 ^ n12733 ^ n4844 ;
  assign n15824 = n12225 ^ n5922 ^ 1'b0 ;
  assign n15825 = n766 & n15824 ;
  assign n15826 = n5985 ^ n2702 ^ 1'b0 ;
  assign n15827 = n2280 & n15826 ;
  assign n15828 = n9836 | n15171 ;
  assign n15829 = n402 | n15828 ;
  assign n15830 = n5306 ^ n4943 ^ 1'b0 ;
  assign n15831 = ~n2024 & n15830 ;
  assign n15832 = n2565 ^ n2558 ^ 1'b0 ;
  assign n15833 = ( n10524 & n12559 ) | ( n10524 & n15832 ) | ( n12559 & n15832 ) ;
  assign n15834 = n15831 & ~n15833 ;
  assign n15835 = ~n2162 & n15834 ;
  assign n15836 = n6917 & n11200 ;
  assign n15837 = n4863 ^ n4052 ^ 1'b0 ;
  assign n15838 = n396 & ~n15837 ;
  assign n15839 = n15838 ^ n10333 ^ 1'b0 ;
  assign n15840 = ( x114 & n6172 ) | ( x114 & n6673 ) | ( n6172 & n6673 ) ;
  assign n15841 = n15840 ^ n12155 ^ n1379 ;
  assign n15842 = n3139 | n15841 ;
  assign n15843 = n15839 & ~n15842 ;
  assign n15844 = ~n1053 & n2340 ;
  assign n15845 = n2112 | n9134 ;
  assign n15846 = n15845 ^ n6028 ^ 1'b0 ;
  assign n15847 = n14663 | n15448 ;
  assign n15848 = n13299 | n15847 ;
  assign n15851 = n1985 ^ n578 ^ 1'b0 ;
  assign n15852 = x116 & ~n15851 ;
  assign n15853 = n667 & n15852 ;
  assign n15854 = n2679 & ~n15853 ;
  assign n15849 = n10824 | n12875 ;
  assign n15850 = n1107 & ~n15849 ;
  assign n15855 = n15854 ^ n15850 ^ 1'b0 ;
  assign n15856 = n6102 ^ n1345 ^ 1'b0 ;
  assign n15857 = n13737 | n15856 ;
  assign n15858 = n8034 | n15857 ;
  assign n15859 = n597 | n1155 ;
  assign n15860 = n11983 | n15859 ;
  assign n15861 = n10412 & n13846 ;
  assign n15862 = n15861 ^ n11165 ^ 1'b0 ;
  assign n15863 = n13179 | n15862 ;
  assign n15864 = n11066 ^ n715 ^ 1'b0 ;
  assign n15865 = n853 & n15864 ;
  assign n15866 = n5972 ^ x115 ^ 1'b0 ;
  assign n15867 = ~n15865 & n15866 ;
  assign n15868 = n2854 & ~n6168 ;
  assign n15869 = x157 & n15868 ;
  assign n15870 = n12655 ^ n10764 ^ n7519 ;
  assign n15871 = ( n15867 & n15869 ) | ( n15867 & ~n15870 ) | ( n15869 & ~n15870 ) ;
  assign n15872 = ( n4822 & n7950 ) | ( n4822 & ~n14095 ) | ( n7950 & ~n14095 ) ;
  assign n15873 = n658 & n3329 ;
  assign n15874 = n11604 & n15873 ;
  assign n15875 = n15874 ^ n7551 ^ 1'b0 ;
  assign n15878 = n5984 & n9552 ;
  assign n15879 = n15878 ^ n11031 ^ 1'b0 ;
  assign n15876 = n6486 ^ n5283 ^ 1'b0 ;
  assign n15877 = n15876 ^ n9887 ^ n8357 ;
  assign n15880 = n15879 ^ n15877 ^ 1'b0 ;
  assign n15881 = n6667 ^ n4714 ^ n3156 ;
  assign n15882 = n15881 ^ n13243 ^ 1'b0 ;
  assign n15883 = n15264 & ~n15882 ;
  assign n15884 = ( ~x231 & n6515 ) | ( ~x231 & n14721 ) | ( n6515 & n14721 ) ;
  assign n15885 = n2775 & n2948 ;
  assign n15886 = ( n2908 & ~n7934 ) | ( n2908 & n15885 ) | ( ~n7934 & n15885 ) ;
  assign n15887 = ( n1849 & n5059 ) | ( n1849 & ~n15886 ) | ( n5059 & ~n15886 ) ;
  assign n15888 = n15887 ^ n2012 ^ 1'b0 ;
  assign n15889 = n4487 & ~n11439 ;
  assign n15890 = ~n1253 & n15889 ;
  assign n15891 = n15890 ^ n4159 ^ 1'b0 ;
  assign n15892 = n7161 & ~n9030 ;
  assign n15893 = n15892 ^ n4585 ^ 1'b0 ;
  assign n15894 = n15893 ^ n3825 ^ 1'b0 ;
  assign n15898 = n8784 ^ x159 ^ 1'b0 ;
  assign n15899 = x188 | n15898 ;
  assign n15900 = n5919 & n9138 ;
  assign n15901 = ~n15899 & n15900 ;
  assign n15895 = n1388 & n5143 ;
  assign n15896 = n6886 & n15895 ;
  assign n15897 = n15896 ^ n12649 ^ 1'b0 ;
  assign n15902 = n15901 ^ n15897 ^ n8399 ;
  assign n15903 = ~n10013 & n11304 ;
  assign n15904 = n13881 ^ n11099 ^ 1'b0 ;
  assign n15905 = n8556 & ~n15904 ;
  assign n15906 = n5985 & n15905 ;
  assign n15907 = n7787 | n13691 ;
  assign n15908 = n3146 ^ n717 ^ 1'b0 ;
  assign n15909 = n2909 & n15908 ;
  assign n15910 = n1766 & n5432 ;
  assign n15911 = n15910 ^ n11572 ^ 1'b0 ;
  assign n15912 = n15909 & n15911 ;
  assign n15913 = n935 & n7099 ;
  assign n15914 = n6321 ^ n5382 ^ 1'b0 ;
  assign n15915 = ( x148 & n15913 ) | ( x148 & n15914 ) | ( n15913 & n15914 ) ;
  assign n15916 = n3235 & n15915 ;
  assign n15918 = n15418 ^ x196 ^ 1'b0 ;
  assign n15919 = n5093 & ~n15918 ;
  assign n15917 = ( n1831 & ~n4628 ) | ( n1831 & n8807 ) | ( ~n4628 & n8807 ) ;
  assign n15920 = n15919 ^ n15917 ^ 1'b0 ;
  assign n15921 = n1376 | n9206 ;
  assign n15922 = n3198 | n15921 ;
  assign n15923 = n15922 ^ n5766 ^ 1'b0 ;
  assign n15924 = ~n1998 & n15923 ;
  assign n15925 = ~n6256 & n14151 ;
  assign n15926 = ~n15924 & n15925 ;
  assign n15930 = n9620 ^ n4024 ^ 1'b0 ;
  assign n15931 = n12528 | n15930 ;
  assign n15927 = n8907 ^ n902 ^ 1'b0 ;
  assign n15928 = x183 & ~n3342 ;
  assign n15929 = n15927 & n15928 ;
  assign n15932 = n15931 ^ n15929 ^ n3027 ;
  assign n15933 = n4163 ^ n1275 ^ x50 ;
  assign n15934 = n15933 ^ n9868 ^ n4059 ;
  assign n15935 = n11318 | n15934 ;
  assign n15936 = n15935 ^ n1156 ^ 1'b0 ;
  assign n15937 = ~n3533 & n8435 ;
  assign n15938 = n15936 & n15937 ;
  assign n15939 = n15938 ^ n6810 ^ 1'b0 ;
  assign n15940 = n13791 ^ n7772 ^ 1'b0 ;
  assign n15942 = n8054 ^ n4515 ^ n544 ;
  assign n15941 = n9378 ^ n4854 ^ 1'b0 ;
  assign n15943 = n15942 ^ n15941 ^ 1'b0 ;
  assign n15944 = n10206 | n14271 ;
  assign n15945 = n9250 | n15944 ;
  assign n15946 = n10411 & ~n15945 ;
  assign n15947 = ( ~n3102 & n7329 ) | ( ~n3102 & n7396 ) | ( n7329 & n7396 ) ;
  assign n15948 = ~n369 & n3800 ;
  assign n15949 = n15948 ^ n1658 ^ 1'b0 ;
  assign n15950 = n15949 ^ n10409 ^ 1'b0 ;
  assign n15951 = n1327 | n15468 ;
  assign n15952 = n3063 | n3878 ;
  assign n15953 = n5101 | n15952 ;
  assign n15954 = n9182 & n15953 ;
  assign n15955 = ( n5236 & n7416 ) | ( n5236 & ~n11180 ) | ( n7416 & ~n11180 ) ;
  assign n15956 = n15955 ^ n13017 ^ n4097 ;
  assign n15957 = ( x3 & ~n15954 ) | ( x3 & n15956 ) | ( ~n15954 & n15956 ) ;
  assign n15958 = n1813 & n8984 ;
  assign n15959 = n9054 ^ n1609 ^ 1'b0 ;
  assign n15960 = ~n15958 & n15959 ;
  assign n15961 = n13928 & n15960 ;
  assign n15962 = n15961 ^ n14478 ^ n1096 ;
  assign n15963 = n2994 & ~n15962 ;
  assign n15965 = n7252 | n7637 ;
  assign n15964 = n2532 & ~n3855 ;
  assign n15966 = n15965 ^ n15964 ^ 1'b0 ;
  assign n15969 = x146 & n2619 ;
  assign n15970 = n15969 ^ n7641 ^ 1'b0 ;
  assign n15971 = ~n8432 & n15970 ;
  assign n15972 = n9439 | n15971 ;
  assign n15967 = n9201 ^ n6489 ^ 1'b0 ;
  assign n15968 = ~n2346 & n15967 ;
  assign n15973 = n15972 ^ n15968 ^ 1'b0 ;
  assign n15974 = ( n15963 & n15966 ) | ( n15963 & n15973 ) | ( n15966 & n15973 ) ;
  assign n15986 = n9043 | n9839 ;
  assign n15987 = n6320 | n15986 ;
  assign n15980 = x165 & ~n1044 ;
  assign n15981 = n6227 & n15980 ;
  assign n15975 = x239 & ~n12619 ;
  assign n15976 = n15975 ^ n5313 ^ 1'b0 ;
  assign n15977 = n15976 ^ n1265 ^ 1'b0 ;
  assign n15978 = n8418 ^ n692 ^ 1'b0 ;
  assign n15979 = ~n15977 & n15978 ;
  assign n15982 = n15981 ^ n15979 ^ n4928 ;
  assign n15983 = ~n575 & n14116 ;
  assign n15984 = n15983 ^ n5576 ^ 1'b0 ;
  assign n15985 = n15982 | n15984 ;
  assign n15988 = n15987 ^ n15985 ^ 1'b0 ;
  assign n15989 = n10934 ^ n763 ^ 1'b0 ;
  assign n15990 = n7392 ^ n1884 ^ 1'b0 ;
  assign n15991 = n15989 | n15990 ;
  assign n15992 = n3604 & ~n15991 ;
  assign n15993 = n15992 ^ n7200 ^ 1'b0 ;
  assign n15994 = n2489 & ~n15993 ;
  assign n15995 = n7106 & ~n8015 ;
  assign n15996 = n15995 ^ n2441 ^ 1'b0 ;
  assign n15997 = n6009 ^ n2636 ^ n369 ;
  assign n15998 = ( n1455 & ~n15996 ) | ( n1455 & n15997 ) | ( ~n15996 & n15997 ) ;
  assign n15999 = ( n1653 & n14506 ) | ( n1653 & n15998 ) | ( n14506 & n15998 ) ;
  assign n16000 = n3786 & ~n7062 ;
  assign n16001 = n16000 ^ n3527 ^ 1'b0 ;
  assign n16002 = n16001 ^ n10165 ^ n702 ;
  assign n16003 = n3097 | n16002 ;
  assign n16005 = n1667 & ~n11634 ;
  assign n16004 = ~n1856 & n7161 ;
  assign n16006 = n16005 ^ n16004 ^ n2811 ;
  assign n16013 = n958 | n5451 ;
  assign n16014 = n1372 & ~n16013 ;
  assign n16007 = n4266 | n8418 ;
  assign n16008 = n16007 ^ n4832 ^ 1'b0 ;
  assign n16009 = n5844 & ~n16008 ;
  assign n16010 = n1299 & n9566 ;
  assign n16011 = ~n16009 & n16010 ;
  assign n16012 = ( n10515 & ~n12694 ) | ( n10515 & n16011 ) | ( ~n12694 & n16011 ) ;
  assign n16015 = n16014 ^ n16012 ^ 1'b0 ;
  assign n16016 = n2529 & n16015 ;
  assign n16017 = n15919 & n16016 ;
  assign n16018 = n16017 ^ n3322 ^ 1'b0 ;
  assign n16019 = ~n10662 & n16018 ;
  assign n16020 = ~n10483 & n14655 ;
  assign n16021 = n16020 ^ n12019 ^ n9318 ;
  assign n16022 = n13112 ^ n2447 ^ n577 ;
  assign n16023 = n12155 & n16022 ;
  assign n16024 = n12289 & n16023 ;
  assign n16025 = n8138 ^ n4343 ^ 1'b0 ;
  assign n16026 = x58 & n6946 ;
  assign n16027 = ~n16025 & n16026 ;
  assign n16028 = n9461 ^ n3768 ^ 1'b0 ;
  assign n16029 = ~n16027 & n16028 ;
  assign n16030 = n7835 & n11216 ;
  assign n16031 = n12378 & n16030 ;
  assign n16032 = n16031 ^ n14361 ^ 1'b0 ;
  assign n16033 = ( n5314 & ~n7015 ) | ( n5314 & n11800 ) | ( ~n7015 & n11800 ) ;
  assign n16034 = n13680 ^ n10432 ^ 1'b0 ;
  assign n16035 = n1031 ^ n856 ^ 1'b0 ;
  assign n16036 = n15279 | n16035 ;
  assign n16037 = ~n11048 & n12159 ;
  assign n16038 = n16037 ^ n1142 ^ 1'b0 ;
  assign n16039 = n13685 ^ n7991 ^ 1'b0 ;
  assign n16040 = n12896 & n16039 ;
  assign n16041 = n777 | n11474 ;
  assign n16042 = ~n14013 & n16041 ;
  assign n16045 = n1817 ^ n432 ^ 1'b0 ;
  assign n16046 = ~n5762 & n16045 ;
  assign n16043 = x19 & n8960 ;
  assign n16044 = n16043 ^ n8221 ^ 1'b0 ;
  assign n16047 = n16046 ^ n16044 ^ 1'b0 ;
  assign n16048 = ~n2295 & n16047 ;
  assign n16049 = n9596 ^ n9583 ^ 1'b0 ;
  assign n16055 = n10750 ^ n5655 ^ n4074 ;
  assign n16050 = n2317 | n2977 ;
  assign n16051 = n5217 & ~n16050 ;
  assign n16052 = n16051 ^ x77 ^ 1'b0 ;
  assign n16053 = n5988 | n16052 ;
  assign n16054 = n3198 | n16053 ;
  assign n16056 = n16055 ^ n16054 ^ 1'b0 ;
  assign n16057 = n5175 & n16056 ;
  assign n16058 = n16057 ^ n6998 ^ 1'b0 ;
  assign n16063 = n660 & n2767 ;
  assign n16059 = n5632 & ~n5931 ;
  assign n16060 = n3721 | n16059 ;
  assign n16061 = n8120 ^ n5118 ^ 1'b0 ;
  assign n16062 = n16060 | n16061 ;
  assign n16064 = n16063 ^ n16062 ^ 1'b0 ;
  assign n16065 = n338 & ~n5732 ;
  assign n16066 = ~n7542 & n16065 ;
  assign n16067 = n15849 | n16066 ;
  assign n16068 = n16067 ^ n8776 ^ n7329 ;
  assign n16069 = n12910 ^ n9300 ^ 1'b0 ;
  assign n16070 = n4090 & n5492 ;
  assign n16071 = n16070 ^ n7411 ^ 1'b0 ;
  assign n16072 = x219 & n8569 ;
  assign n16073 = n604 & n16072 ;
  assign n16074 = n5318 & ~n16073 ;
  assign n16075 = n16074 ^ n7481 ^ 1'b0 ;
  assign n16076 = n16071 & ~n16075 ;
  assign n16077 = n16076 ^ n2146 ^ 1'b0 ;
  assign n16078 = ( n7601 & n7814 ) | ( n7601 & ~n16077 ) | ( n7814 & ~n16077 ) ;
  assign n16082 = n835 | n8433 ;
  assign n16083 = n5991 & ~n16082 ;
  assign n16084 = ~n6983 & n15410 ;
  assign n16085 = n16083 & n16084 ;
  assign n16086 = ( n3830 & ~n5408 ) | ( n3830 & n16085 ) | ( ~n5408 & n16085 ) ;
  assign n16087 = n11365 | n16086 ;
  assign n16079 = n4595 ^ n1882 ^ 1'b0 ;
  assign n16080 = n403 | n16079 ;
  assign n16081 = n9358 & n16080 ;
  assign n16088 = n16087 ^ n16081 ^ 1'b0 ;
  assign n16089 = n7422 | n16088 ;
  assign n16090 = ( ~n7385 & n8101 ) | ( ~n7385 & n11784 ) | ( n8101 & n11784 ) ;
  assign n16091 = ~x33 & x232 ;
  assign n16092 = n901 | n16091 ;
  assign n16093 = n8827 ^ n4389 ^ 1'b0 ;
  assign n16094 = n1549 & ~n6865 ;
  assign n16095 = n16094 ^ n12139 ^ 1'b0 ;
  assign n16096 = n5427 ^ n3945 ^ n2071 ;
  assign n16097 = n4301 ^ n1448 ^ 1'b0 ;
  assign n16098 = n16096 & ~n16097 ;
  assign n16099 = n16095 & n16098 ;
  assign n16100 = ~n3779 & n6523 ;
  assign n16103 = n5004 ^ x41 ^ 1'b0 ;
  assign n16101 = n10002 ^ n3457 ^ n1406 ;
  assign n16102 = n9696 & n16101 ;
  assign n16104 = n16103 ^ n16102 ^ 1'b0 ;
  assign n16105 = n16104 ^ x20 ^ 1'b0 ;
  assign n16106 = n3731 | n12078 ;
  assign n16107 = ( n4745 & ~n5149 ) | ( n4745 & n6099 ) | ( ~n5149 & n6099 ) ;
  assign n16108 = n16107 ^ n7641 ^ n1530 ;
  assign n16109 = ( n2774 & ~n15772 ) | ( n2774 & n16108 ) | ( ~n15772 & n16108 ) ;
  assign n16110 = n302 | n11054 ;
  assign n16111 = n16110 ^ n14612 ^ 1'b0 ;
  assign n16112 = n5446 | n16111 ;
  assign n16113 = n8697 & ~n16112 ;
  assign n16114 = n3666 | n16113 ;
  assign n16115 = n16114 ^ x250 ^ 1'b0 ;
  assign n16116 = ~n8721 & n16115 ;
  assign n16117 = n8758 & n16116 ;
  assign n16118 = n10791 ^ n9271 ^ 1'b0 ;
  assign n16119 = n2372 & n6497 ;
  assign n16120 = n16118 & n16119 ;
  assign n16121 = n2529 ^ n1251 ^ 1'b0 ;
  assign n16122 = n8327 & ~n16121 ;
  assign n16123 = n8839 & ~n16122 ;
  assign n16124 = ( n402 & n8473 ) | ( n402 & n16123 ) | ( n8473 & n16123 ) ;
  assign n16125 = n9592 ^ n1593 ^ 1'b0 ;
  assign n16126 = n15599 ^ n6276 ^ n433 ;
  assign n16127 = n9857 ^ n3615 ^ 1'b0 ;
  assign n16128 = x90 | n16127 ;
  assign n16129 = n2688 & ~n3957 ;
  assign n16130 = n16129 ^ n2916 ^ 1'b0 ;
  assign n16131 = n10846 ^ n8895 ^ 1'b0 ;
  assign n16132 = ( n4685 & n16130 ) | ( n4685 & n16131 ) | ( n16130 & n16131 ) ;
  assign n16133 = ( n13708 & n16128 ) | ( n13708 & ~n16132 ) | ( n16128 & ~n16132 ) ;
  assign n16134 = ~n3317 & n9995 ;
  assign n16135 = n16134 ^ n12172 ^ 1'b0 ;
  assign n16136 = n1495 | n2005 ;
  assign n16137 = n6827 ^ n5097 ^ 1'b0 ;
  assign n16138 = ~n9986 & n16137 ;
  assign n16139 = n10368 & ~n16138 ;
  assign n16140 = n5276 & n16139 ;
  assign n16141 = n2962 & ~n12271 ;
  assign n16142 = ~n5709 & n16141 ;
  assign n16143 = n778 & ~n16142 ;
  assign n16144 = n2386 & n16143 ;
  assign n16145 = n8929 & ~n16144 ;
  assign n16146 = n16145 ^ n15771 ^ 1'b0 ;
  assign n16147 = n14210 ^ n13280 ^ 1'b0 ;
  assign n16148 = n6034 ^ n2493 ^ n519 ;
  assign n16149 = ( ~n3500 & n14410 ) | ( ~n3500 & n16148 ) | ( n14410 & n16148 ) ;
  assign n16150 = ( ~n2830 & n4314 ) | ( ~n2830 & n16149 ) | ( n4314 & n16149 ) ;
  assign n16151 = n808 & ~n7090 ;
  assign n16152 = ~n7754 & n16151 ;
  assign n16153 = n5923 ^ n4355 ^ 1'b0 ;
  assign n16154 = n1932 & ~n16153 ;
  assign n16155 = n16154 ^ n4043 ^ 1'b0 ;
  assign n16156 = n4129 & ~n7055 ;
  assign n16157 = n16156 ^ n4515 ^ 1'b0 ;
  assign n16158 = n3580 | n16152 ;
  assign n16159 = x244 | n16158 ;
  assign n16160 = n3770 ^ n2005 ^ 1'b0 ;
  assign n16161 = n2259 & n6632 ;
  assign n16162 = ~n16160 & n16161 ;
  assign n16163 = n16162 ^ n12004 ^ 1'b0 ;
  assign n16164 = n12029 ^ x243 ^ 1'b0 ;
  assign n16165 = n14618 & n16164 ;
  assign n16166 = n3025 & ~n7270 ;
  assign n16167 = n1350 | n16166 ;
  assign n16168 = ( n9344 & ~n13981 ) | ( n9344 & n16167 ) | ( ~n13981 & n16167 ) ;
  assign n16170 = n7484 ^ n5313 ^ 1'b0 ;
  assign n16171 = n8327 & ~n16170 ;
  assign n16169 = n1054 & n15509 ;
  assign n16172 = n16171 ^ n16169 ^ 1'b0 ;
  assign n16173 = ( n10934 & n15632 ) | ( n10934 & n16172 ) | ( n15632 & n16172 ) ;
  assign n16174 = n10122 ^ n5376 ^ 1'b0 ;
  assign n16175 = n6713 & n8004 ;
  assign n16176 = n16174 | n16175 ;
  assign n16177 = n16176 ^ n307 ^ 1'b0 ;
  assign n16182 = n6186 ^ n603 ^ x39 ;
  assign n16178 = n5751 & ~n11056 ;
  assign n16179 = n396 & n16178 ;
  assign n16180 = n14559 | n16179 ;
  assign n16181 = n4484 | n16180 ;
  assign n16183 = n16182 ^ n16181 ^ 1'b0 ;
  assign n16186 = n3865 ^ n2847 ^ 1'b0 ;
  assign n16184 = ~n1504 & n2461 ;
  assign n16185 = n16184 ^ n4396 ^ 1'b0 ;
  assign n16187 = n16186 ^ n16185 ^ n9781 ;
  assign n16188 = n6754 & ~n16187 ;
  assign n16189 = ~n16183 & n16188 ;
  assign n16190 = n9281 ^ n7197 ^ 1'b0 ;
  assign n16191 = ( n2769 & n13954 ) | ( n2769 & n14905 ) | ( n13954 & n14905 ) ;
  assign n16192 = n16190 & ~n16191 ;
  assign n16193 = n16192 ^ x140 ^ 1'b0 ;
  assign n16194 = n16193 ^ n10620 ^ 1'b0 ;
  assign n16195 = n7519 ^ n4300 ^ n3576 ;
  assign n16196 = x95 & n5909 ;
  assign n16197 = ~n12159 & n16196 ;
  assign n16198 = n6018 & ~n16197 ;
  assign n16199 = ~n16195 & n16198 ;
  assign n16200 = n2899 & n4764 ;
  assign n16201 = ~n4934 & n16200 ;
  assign n16202 = ~n13017 & n16201 ;
  assign n16203 = n5377 | n16202 ;
  assign n16204 = n11676 & ~n16203 ;
  assign n16205 = ( n1678 & ~n5865 ) | ( n1678 & n6192 ) | ( ~n5865 & n6192 ) ;
  assign n16206 = ( n3429 & n11936 ) | ( n3429 & n16205 ) | ( n11936 & n16205 ) ;
  assign n16207 = n10521 ^ n926 ^ 1'b0 ;
  assign n16208 = n2073 & ~n7080 ;
  assign n16209 = n16208 ^ x189 ^ 1'b0 ;
  assign n16210 = n10496 | n16209 ;
  assign n16211 = n16210 ^ n12567 ^ 1'b0 ;
  assign n16212 = ~n7417 & n8198 ;
  assign n16213 = n16212 ^ n3585 ^ 1'b0 ;
  assign n16214 = n16213 ^ n2847 ^ 1'b0 ;
  assign n16215 = ~n314 & n16214 ;
  assign n16216 = n16215 ^ n8257 ^ 1'b0 ;
  assign n16217 = n2994 & n10688 ;
  assign n16218 = n14444 & n16217 ;
  assign n16219 = n932 & n8567 ;
  assign n16220 = n16218 & n16219 ;
  assign n16221 = n2790 ^ n2090 ^ 1'b0 ;
  assign n16222 = n11318 ^ n5386 ^ 1'b0 ;
  assign n16223 = n587 | n10546 ;
  assign n16224 = n7145 & ~n7880 ;
  assign n16225 = ~n16223 & n16224 ;
  assign n16226 = n2223 | n13196 ;
  assign n16227 = n16225 & ~n16226 ;
  assign n16228 = ( n16221 & n16222 ) | ( n16221 & n16227 ) | ( n16222 & n16227 ) ;
  assign n16229 = ( n4804 & n7456 ) | ( n4804 & ~n16228 ) | ( n7456 & ~n16228 ) ;
  assign n16230 = n11108 ^ n7787 ^ n5279 ;
  assign n16231 = n16230 ^ x121 ^ 1'b0 ;
  assign n16232 = n5502 ^ n1962 ^ 1'b0 ;
  assign n16233 = ( x21 & n4869 ) | ( x21 & n9005 ) | ( n4869 & n9005 ) ;
  assign n16234 = n8801 ^ n4405 ^ 1'b0 ;
  assign n16235 = ~n2660 & n7399 ;
  assign n16236 = n16235 ^ x185 ^ 1'b0 ;
  assign n16237 = n4883 & n7285 ;
  assign n16238 = n16236 & n16237 ;
  assign n16239 = n5916 & n7029 ;
  assign n16242 = n12196 ^ n5881 ^ n4525 ;
  assign n16240 = ~n1476 & n14386 ;
  assign n16241 = n16240 ^ n5133 ^ 1'b0 ;
  assign n16243 = n16242 ^ n16241 ^ n6254 ;
  assign n16244 = n16243 ^ n14559 ^ n9534 ;
  assign n16245 = n11997 | n16244 ;
  assign n16246 = n16245 ^ n5539 ^ 1'b0 ;
  assign n16247 = ( n4833 & n13726 ) | ( n4833 & n16246 ) | ( n13726 & n16246 ) ;
  assign n16248 = ~n2831 & n15987 ;
  assign n16249 = n9484 & n16248 ;
  assign n16250 = n16249 ^ n14363 ^ 1'b0 ;
  assign n16251 = n2461 ^ n1571 ^ 1'b0 ;
  assign n16252 = n1760 & n16251 ;
  assign n16253 = n16252 ^ n13453 ^ n11110 ;
  assign n16254 = n16253 ^ n2172 ^ 1'b0 ;
  assign n16255 = n5576 ^ n5377 ^ n3555 ;
  assign n16256 = ~n13214 & n16255 ;
  assign n16257 = n6626 | n8962 ;
  assign n16258 = n12413 | n16257 ;
  assign n16259 = n4027 & n9187 ;
  assign n16260 = n888 & n16259 ;
  assign n16261 = n16260 ^ n15219 ^ 1'b0 ;
  assign n16262 = ~n12746 & n16261 ;
  assign n16263 = ~n9155 & n16262 ;
  assign n16264 = n8515 | n9955 ;
  assign n16265 = ( n3439 & n5949 ) | ( n3439 & ~n16264 ) | ( n5949 & ~n16264 ) ;
  assign n16266 = ( n7586 & ~n8275 ) | ( n7586 & n15940 ) | ( ~n8275 & n15940 ) ;
  assign n16269 = n8897 ^ n3115 ^ 1'b0 ;
  assign n16268 = ~n8420 & n9872 ;
  assign n16270 = n16269 ^ n16268 ^ 1'b0 ;
  assign n16267 = n10259 ^ n5520 ^ 1'b0 ;
  assign n16271 = n16270 ^ n16267 ^ n12299 ;
  assign n16275 = n8221 ^ n1145 ^ 1'b0 ;
  assign n16276 = n10442 & n16275 ;
  assign n16272 = n11802 | n12061 ;
  assign n16273 = n16272 ^ n3417 ^ 1'b0 ;
  assign n16274 = ~n16221 & n16273 ;
  assign n16277 = n16276 ^ n16274 ^ 1'b0 ;
  assign n16278 = ( n464 & n13206 ) | ( n464 & ~n15652 ) | ( n13206 & ~n15652 ) ;
  assign n16279 = n9125 & ~n11765 ;
  assign n16280 = ~n12888 & n16279 ;
  assign n16281 = n4695 & n16280 ;
  assign n16282 = n9180 & ~n10129 ;
  assign n16283 = n11331 & n14443 ;
  assign n16284 = n6649 & n16283 ;
  assign n16285 = x104 & ~n3636 ;
  assign n16286 = n1106 & n16285 ;
  assign n16287 = n16286 ^ n2891 ^ 1'b0 ;
  assign n16288 = n16287 ^ n11187 ^ 1'b0 ;
  assign n16289 = n540 | n16288 ;
  assign n16290 = n7426 & ~n12698 ;
  assign n16291 = n2868 & n4790 ;
  assign n16292 = ~n4197 & n16291 ;
  assign n16293 = ( n2823 & n3418 ) | ( n2823 & ~n16292 ) | ( n3418 & ~n16292 ) ;
  assign n16294 = n1778 | n15047 ;
  assign n16295 = n6489 & n10163 ;
  assign n16296 = ~n10463 & n16295 ;
  assign n16297 = n15494 ^ n6596 ^ 1'b0 ;
  assign n16298 = ~n2738 & n16297 ;
  assign n16299 = n4756 ^ n2708 ^ 1'b0 ;
  assign n16300 = n15091 ^ n13186 ^ 1'b0 ;
  assign n16301 = ~x215 & n10021 ;
  assign n16302 = n13420 & ~n16301 ;
  assign n16303 = n16302 ^ n2209 ^ 1'b0 ;
  assign n16305 = ( ~n6642 & n8597 ) | ( ~n6642 & n11242 ) | ( n8597 & n11242 ) ;
  assign n16304 = n1076 | n10536 ;
  assign n16306 = n16305 ^ n16304 ^ 1'b0 ;
  assign n16307 = n3333 & n9853 ;
  assign n16308 = n16307 ^ n7280 ^ 1'b0 ;
  assign n16309 = ( n9475 & n14985 ) | ( n9475 & n16308 ) | ( n14985 & n16308 ) ;
  assign n16310 = n2052 | n2993 ;
  assign n16311 = n3039 | n16310 ;
  assign n16312 = n16311 ^ n10063 ^ n4385 ;
  assign n16313 = n3521 ^ n2940 ^ 1'b0 ;
  assign n16314 = n9751 & ~n14464 ;
  assign n16315 = n16314 ^ n11676 ^ 1'b0 ;
  assign n16316 = n10781 ^ n6800 ^ 1'b0 ;
  assign n16317 = n6254 | n16316 ;
  assign n16318 = n8858 & ~n9884 ;
  assign n16319 = x198 | n14466 ;
  assign n16320 = n16318 | n16319 ;
  assign n16321 = ( ~n2339 & n4433 ) | ( ~n2339 & n11501 ) | ( n4433 & n11501 ) ;
  assign n16322 = n4324 & ~n9054 ;
  assign n16323 = n16322 ^ n14079 ^ 1'b0 ;
  assign n16324 = n4694 ^ n1470 ^ 1'b0 ;
  assign n16325 = n971 & n16324 ;
  assign n16326 = ~n2050 & n16325 ;
  assign n16327 = n16275 & n16326 ;
  assign n16328 = n15297 ^ n10524 ^ n10073 ;
  assign n16329 = n16328 ^ n2942 ^ 1'b0 ;
  assign n16330 = n7893 & ~n16329 ;
  assign n16332 = n4256 & ~n6583 ;
  assign n16333 = n16332 ^ n4756 ^ 1'b0 ;
  assign n16334 = ( n4118 & ~n9913 ) | ( n4118 & n16333 ) | ( ~n9913 & n16333 ) ;
  assign n16335 = n16334 ^ n12553 ^ n10753 ;
  assign n16331 = ~n3653 & n15512 ;
  assign n16336 = n16335 ^ n16331 ^ 1'b0 ;
  assign n16337 = n1394 | n7789 ;
  assign n16338 = ~n8603 & n13568 ;
  assign n16339 = n8356 ^ n3768 ^ n3393 ;
  assign n16340 = n16338 & n16339 ;
  assign n16341 = n11140 ^ n4697 ^ n1028 ;
  assign n16342 = n4911 & n16341 ;
  assign n16343 = n16342 ^ n8924 ^ 1'b0 ;
  assign n16344 = n5816 | n16343 ;
  assign n16345 = n7209 & ~n9492 ;
  assign n16346 = ~n16344 & n16345 ;
  assign n16351 = ( ~n4244 & n4280 ) | ( ~n4244 & n4858 ) | ( n4280 & n4858 ) ;
  assign n16347 = n8616 ^ x226 ^ x26 ;
  assign n16348 = n9806 & n16347 ;
  assign n16349 = ~n5818 & n16348 ;
  assign n16350 = n11431 & ~n16349 ;
  assign n16352 = n16351 ^ n16350 ^ x108 ;
  assign n16353 = ~n9235 & n15626 ;
  assign n16354 = ~n3510 & n16353 ;
  assign n16357 = n4558 ^ n4538 ^ n804 ;
  assign n16355 = n5782 & ~n10303 ;
  assign n16356 = n5027 & n16355 ;
  assign n16358 = n16357 ^ n16356 ^ n363 ;
  assign n16359 = n10165 & ~n12329 ;
  assign n16360 = ~x28 & n16359 ;
  assign n16361 = n12698 ^ n1124 ^ 1'b0 ;
  assign n16362 = ~n16360 & n16361 ;
  assign n16363 = n844 | n6152 ;
  assign n16364 = x11 & ~n2048 ;
  assign n16365 = n16364 ^ n1861 ^ 1'b0 ;
  assign n16366 = n16365 ^ n4826 ^ n2661 ;
  assign n16367 = x29 & ~n16366 ;
  assign n16368 = n7989 & n16367 ;
  assign n16369 = n7345 & ~n10860 ;
  assign n16370 = n16369 ^ n631 ^ 1'b0 ;
  assign n16371 = n16370 ^ n8164 ^ 1'b0 ;
  assign n16372 = n2727 | n6527 ;
  assign n16373 = n417 | n16372 ;
  assign n16374 = n1434 | n12624 ;
  assign n16375 = n16373 | n16374 ;
  assign n16376 = n16375 ^ n3475 ^ 1'b0 ;
  assign n16377 = n12828 & ~n16376 ;
  assign n16378 = ~n16371 & n16377 ;
  assign n16379 = n6796 ^ n4392 ^ 1'b0 ;
  assign n16380 = n5251 & ~n16379 ;
  assign n16381 = n2676 & n4883 ;
  assign n16382 = ~n3348 & n16381 ;
  assign n16383 = ( n1930 & n16380 ) | ( n1930 & n16382 ) | ( n16380 & n16382 ) ;
  assign n16384 = n4061 ^ n277 ^ 1'b0 ;
  assign n16385 = ~n11435 & n16384 ;
  assign n16386 = n2728 & n6968 ;
  assign n16387 = n6294 & n16386 ;
  assign n16388 = n12877 ^ n3892 ^ 1'b0 ;
  assign n16389 = n9475 & n14317 ;
  assign n16390 = n16389 ^ n10419 ^ 1'b0 ;
  assign n16391 = n16390 ^ n5417 ^ 1'b0 ;
  assign n16392 = x57 & n3680 ;
  assign n16393 = n13597 ^ n12450 ^ 1'b0 ;
  assign n16394 = ~n9971 & n16393 ;
  assign n16395 = n273 | n3122 ;
  assign n16396 = n16395 ^ n15348 ^ 1'b0 ;
  assign n16397 = n16396 ^ n5483 ^ 1'b0 ;
  assign n16403 = n9282 ^ n4685 ^ n3727 ;
  assign n16399 = x240 & ~n6374 ;
  assign n16400 = n16399 ^ n3057 ^ 1'b0 ;
  assign n16401 = n16400 ^ n5528 ^ 1'b0 ;
  assign n16402 = n16401 ^ n10160 ^ n9650 ;
  assign n16398 = n1362 & n1843 ;
  assign n16404 = n16403 ^ n16402 ^ n16398 ;
  assign n16405 = ~n8991 & n12903 ;
  assign n16406 = n3533 ^ x235 ^ 1'b0 ;
  assign n16407 = ( n8846 & n12576 ) | ( n8846 & ~n16406 ) | ( n12576 & ~n16406 ) ;
  assign n16408 = n14518 ^ n10675 ^ n547 ;
  assign n16409 = n2223 ^ n708 ^ n347 ;
  assign n16410 = n9005 & ~n16409 ;
  assign n16411 = ( n630 & n5244 ) | ( n630 & ~n8299 ) | ( n5244 & ~n8299 ) ;
  assign n16412 = n16411 ^ x44 ^ 1'b0 ;
  assign n16413 = n13112 ^ n1586 ^ x83 ;
  assign n16414 = n14544 & ~n16413 ;
  assign n16415 = n15334 & n16414 ;
  assign n16416 = ( n1719 & n3431 ) | ( n1719 & ~n8690 ) | ( n3431 & ~n8690 ) ;
  assign n16417 = n16415 & n16416 ;
  assign n16418 = ~n16328 & n16417 ;
  assign n16419 = n3742 ^ x4 ^ 1'b0 ;
  assign n16420 = n16419 ^ n7775 ^ 1'b0 ;
  assign n16421 = n11302 ^ n1261 ^ 1'b0 ;
  assign n16422 = n1554 | n16421 ;
  assign n16423 = n327 & n16422 ;
  assign n16424 = n552 & ~n16166 ;
  assign n16425 = n12197 & ~n16424 ;
  assign n16426 = n13625 & ~n16425 ;
  assign n16427 = n7549 & n16426 ;
  assign n16428 = n9590 | n16427 ;
  assign n16429 = n16428 ^ n308 ^ 1'b0 ;
  assign n16430 = n16429 ^ n13378 ^ 1'b0 ;
  assign n16431 = n1270 | n6989 ;
  assign n16432 = ~n15514 & n16431 ;
  assign n16433 = n16432 ^ n5582 ^ 1'b0 ;
  assign n16434 = n2292 | n8668 ;
  assign n16435 = n13901 ^ x94 ^ 1'b0 ;
  assign n16436 = n12415 & ~n16435 ;
  assign n16437 = n4556 ^ n3404 ^ 1'b0 ;
  assign n16438 = n6647 & ~n14407 ;
  assign n16439 = n16438 ^ n2728 ^ 1'b0 ;
  assign n16440 = n16439 ^ x61 ^ 1'b0 ;
  assign n16441 = n12493 ^ n6585 ^ 1'b0 ;
  assign n16442 = n4628 ^ n1347 ^ 1'b0 ;
  assign n16443 = n3854 & n16442 ;
  assign n16444 = n16443 ^ n15009 ^ 1'b0 ;
  assign n16445 = n9076 ^ n1128 ^ 1'b0 ;
  assign n16446 = n9201 & ~n16445 ;
  assign n16447 = n16444 & n16446 ;
  assign n16448 = ~n905 & n15414 ;
  assign n16449 = ~n4496 & n16448 ;
  assign n16450 = n8465 ^ n1161 ^ 1'b0 ;
  assign n16451 = n1290 | n2534 ;
  assign n16452 = n396 | n16451 ;
  assign n16453 = n16452 ^ n913 ^ 1'b0 ;
  assign n16454 = n8905 & ~n16453 ;
  assign n16455 = n7755 ^ n6678 ^ n3936 ;
  assign n16456 = n8225 ^ n7295 ^ n3353 ;
  assign n16468 = ( ~n941 & n1452 ) | ( ~n941 & n1956 ) | ( n1452 & n1956 ) ;
  assign n16467 = n5499 ^ n1140 ^ 1'b0 ;
  assign n16469 = n16468 ^ n16467 ^ 1'b0 ;
  assign n16460 = n6389 ^ n6018 ^ 1'b0 ;
  assign n16461 = n7192 & n16460 ;
  assign n16457 = n7660 ^ n6428 ^ 1'b0 ;
  assign n16458 = n9180 | n16457 ;
  assign n16459 = n2823 | n16458 ;
  assign n16462 = n16461 ^ n16459 ^ 1'b0 ;
  assign n16463 = ~n12279 & n16462 ;
  assign n16464 = ~n15509 & n16463 ;
  assign n16465 = n16464 ^ n1231 ^ 1'b0 ;
  assign n16466 = ~n3016 & n16465 ;
  assign n16470 = n16469 ^ n16466 ^ n1961 ;
  assign n16472 = ~n2349 & n4033 ;
  assign n16473 = n8818 & ~n16472 ;
  assign n16471 = n12808 ^ n1632 ^ n639 ;
  assign n16474 = n16473 ^ n16471 ^ 1'b0 ;
  assign n16475 = ~n5565 & n16474 ;
  assign n16476 = ~n3802 & n16475 ;
  assign n16477 = n1962 | n10798 ;
  assign n16478 = ~n4061 & n4868 ;
  assign n16479 = n16478 ^ n7708 ^ 1'b0 ;
  assign n16480 = n9393 & n16479 ;
  assign n16481 = n6705 & n9486 ;
  assign n16482 = ~n12589 & n16481 ;
  assign n16483 = n2268 ^ n1969 ^ n1354 ;
  assign n16484 = n6276 & ~n10670 ;
  assign n16485 = ~n7393 & n16484 ;
  assign n16486 = n8027 ^ n6392 ^ 1'b0 ;
  assign n16487 = n9269 & ~n16486 ;
  assign n16488 = ( n5807 & n7147 ) | ( n5807 & ~n16487 ) | ( n7147 & ~n16487 ) ;
  assign n16489 = n16488 ^ n13493 ^ 1'b0 ;
  assign n16490 = ( x137 & n1217 ) | ( x137 & ~n4422 ) | ( n1217 & ~n4422 ) ;
  assign n16491 = n5928 | n6791 ;
  assign n16492 = n8466 | n9196 ;
  assign n16493 = n16491 & ~n16492 ;
  assign n16494 = n4324 | n15573 ;
  assign n16495 = n16494 ^ n4916 ^ 1'b0 ;
  assign n16496 = n16493 & ~n16495 ;
  assign n16497 = n7291 ^ n1113 ^ 1'b0 ;
  assign n16498 = n16497 ^ n1600 ^ 1'b0 ;
  assign n16499 = ~n2598 & n16498 ;
  assign n16500 = n6488 ^ n5195 ^ 1'b0 ;
  assign n16501 = n8907 ^ n7222 ^ 1'b0 ;
  assign n16502 = ~n9319 & n16501 ;
  assign n16503 = ~n13335 & n16502 ;
  assign n16504 = n16503 ^ n5919 ^ 1'b0 ;
  assign n16505 = n16504 ^ n13390 ^ n1633 ;
  assign n16506 = n9896 | n14016 ;
  assign n16507 = n15720 ^ n1022 ^ 1'b0 ;
  assign n16508 = ~n16506 & n16507 ;
  assign n16509 = n3199 & n15364 ;
  assign n16510 = ~n1110 & n16509 ;
  assign n16511 = n5880 ^ n3636 ^ 1'b0 ;
  assign n16512 = ~n8984 & n16511 ;
  assign n16513 = n1923 & n11659 ;
  assign n16514 = ~n16512 & n16513 ;
  assign n16515 = n5443 ^ n5406 ^ 1'b0 ;
  assign n16516 = ~n8622 & n16515 ;
  assign n16517 = ~n10832 & n16516 ;
  assign n16518 = n16517 ^ n10021 ^ 1'b0 ;
  assign n16519 = n5768 ^ n5189 ^ x61 ;
  assign n16520 = n16519 ^ n706 ^ 1'b0 ;
  assign n16522 = n6994 ^ n1946 ^ 1'b0 ;
  assign n16521 = n3213 | n10044 ;
  assign n16523 = n16522 ^ n16521 ^ n13640 ;
  assign n16524 = x148 & n16523 ;
  assign n16525 = x130 & n11106 ;
  assign n16526 = n4314 | n16525 ;
  assign n16527 = n5665 & ~n16526 ;
  assign n16528 = ~n11419 & n15972 ;
  assign n16529 = n8909 ^ n1604 ^ 1'b0 ;
  assign n16530 = n15127 ^ n8986 ^ 1'b0 ;
  assign n16531 = n15397 ^ n7995 ^ 1'b0 ;
  assign n16532 = x109 & n16531 ;
  assign n16533 = n1234 & ~n16532 ;
  assign n16534 = ~n11054 & n11709 ;
  assign n16535 = n16534 ^ n16462 ^ 1'b0 ;
  assign n16536 = n7851 & ~n12184 ;
  assign n16537 = ~n4163 & n16536 ;
  assign n16538 = n16537 ^ n2024 ^ 1'b0 ;
  assign n16539 = ( n2295 & n15461 ) | ( n2295 & ~n16538 ) | ( n15461 & ~n16538 ) ;
  assign n16540 = n9969 ^ n4431 ^ n2827 ;
  assign n16541 = n11716 & ~n16540 ;
  assign n16542 = n16541 ^ n5778 ^ 1'b0 ;
  assign n16543 = ~n7883 & n10685 ;
  assign n16544 = n16543 ^ n11624 ^ n1261 ;
  assign n16545 = ~x117 & n10685 ;
  assign n16546 = n3169 | n13810 ;
  assign n16547 = n4014 ^ n3283 ^ 1'b0 ;
  assign n16548 = n16547 ^ n7549 ^ 1'b0 ;
  assign n16549 = n8642 ^ n6003 ^ 1'b0 ;
  assign n16550 = n16548 | n16549 ;
  assign n16551 = n8114 | n16550 ;
  assign n16552 = ~n2009 & n11447 ;
  assign n16553 = n6580 & n16552 ;
  assign n16554 = n6771 & ~n10581 ;
  assign n16555 = n16554 ^ n1326 ^ 1'b0 ;
  assign n16563 = n9967 ^ n5368 ^ 1'b0 ;
  assign n16564 = ~n2706 & n16563 ;
  assign n16565 = n16564 ^ n7774 ^ 1'b0 ;
  assign n16556 = n6745 ^ n1580 ^ n485 ;
  assign n16557 = n3983 ^ n3974 ^ 1'b0 ;
  assign n16558 = ~n16556 & n16557 ;
  assign n16559 = n16558 ^ x93 ^ 1'b0 ;
  assign n16560 = ~n980 & n11584 ;
  assign n16561 = n15958 & n16560 ;
  assign n16562 = n16559 | n16561 ;
  assign n16566 = n16565 ^ n16562 ^ 1'b0 ;
  assign n16567 = n16555 | n16566 ;
  assign n16568 = n13956 | n16567 ;
  assign n16569 = n957 & ~n13479 ;
  assign n16570 = n16569 ^ n8947 ^ 1'b0 ;
  assign n16571 = n1300 & n16570 ;
  assign n16572 = n12084 ^ n8471 ^ 1'b0 ;
  assign n16573 = ~n2405 & n16572 ;
  assign n16574 = n16573 ^ n4536 ^ 1'b0 ;
  assign n16575 = ~n12640 & n16574 ;
  assign n16576 = n13107 ^ n2782 ^ 1'b0 ;
  assign n16577 = n16354 ^ n11407 ^ n2157 ;
  assign n16578 = n1154 & n1350 ;
  assign n16579 = n13696 | n13761 ;
  assign n16580 = n16579 ^ n8800 ^ 1'b0 ;
  assign n16585 = n4690 & n12519 ;
  assign n16586 = n4543 & n16585 ;
  assign n16581 = ~n1470 & n5033 ;
  assign n16582 = n10157 ^ n1410 ^ 1'b0 ;
  assign n16583 = ~n7132 & n16582 ;
  assign n16584 = n16581 & n16583 ;
  assign n16587 = n16586 ^ n16584 ^ 1'b0 ;
  assign n16588 = ~n9507 & n16587 ;
  assign n16589 = ~n16580 & n16588 ;
  assign n16592 = n11809 ^ n3774 ^ n2247 ;
  assign n16590 = ~n3547 & n4703 ;
  assign n16591 = n2873 & n16590 ;
  assign n16593 = n16592 ^ n16591 ^ 1'b0 ;
  assign n16594 = ( ~x80 & n2954 ) | ( ~x80 & n3798 ) | ( n2954 & n3798 ) ;
  assign n16595 = n2690 & ~n4692 ;
  assign n16596 = n16595 ^ n9086 ^ 1'b0 ;
  assign n16597 = n16596 ^ n15592 ^ 1'b0 ;
  assign n16598 = n6014 & n16597 ;
  assign n16599 = n2571 ^ n1709 ^ n1388 ;
  assign n16600 = n5745 & n16599 ;
  assign n16601 = n5846 | n16600 ;
  assign n16602 = n8377 ^ n1709 ^ 1'b0 ;
  assign n16603 = n3239 & ~n16602 ;
  assign n16604 = n16603 ^ n1061 ^ 1'b0 ;
  assign n16605 = n4045 & ~n16604 ;
  assign n16606 = n6971 & n14528 ;
  assign n16607 = n16606 ^ n16046 ^ n8356 ;
  assign n16608 = ~n10616 & n16607 ;
  assign n16609 = n8110 & n16608 ;
  assign n16610 = ( ~n2251 & n16605 ) | ( ~n2251 & n16609 ) | ( n16605 & n16609 ) ;
  assign n16611 = ~n7222 & n10789 ;
  assign n16612 = n16480 ^ n5473 ^ 1'b0 ;
  assign n16613 = n6390 ^ n6248 ^ x98 ;
  assign n16614 = n789 & ~n3923 ;
  assign n16615 = ~n5809 & n16614 ;
  assign n16616 = n2516 & ~n14005 ;
  assign n16617 = n16616 ^ n884 ^ 1'b0 ;
  assign n16618 = n8204 ^ n2259 ^ 1'b0 ;
  assign n16619 = n8682 | n16618 ;
  assign n16620 = n2019 | n16619 ;
  assign n16621 = n16617 | n16620 ;
  assign n16622 = ( n16613 & n16615 ) | ( n16613 & ~n16621 ) | ( n16615 & ~n16621 ) ;
  assign n16623 = ( n8121 & n8622 ) | ( n8121 & ~n13860 ) | ( n8622 & ~n13860 ) ;
  assign n16624 = n8051 ^ n834 ^ 1'b0 ;
  assign n16625 = n3986 & ~n6944 ;
  assign n16626 = n16624 | n16625 ;
  assign n16627 = n16626 ^ n7394 ^ 1'b0 ;
  assign n16628 = n2005 & n16627 ;
  assign n16629 = n11221 & n13261 ;
  assign n16630 = n16629 ^ n1991 ^ 1'b0 ;
  assign n16631 = ( ~n396 & n5608 ) | ( ~n396 & n6843 ) | ( n5608 & n6843 ) ;
  assign n16632 = n16631 ^ n14079 ^ 1'b0 ;
  assign n16633 = n16630 & ~n16632 ;
  assign n16634 = n1123 | n4759 ;
  assign n16635 = n5687 | n16634 ;
  assign n16636 = n16635 ^ n1019 ^ 1'b0 ;
  assign n16637 = n8523 | n16636 ;
  assign n16638 = n16637 ^ n12086 ^ 1'b0 ;
  assign n16639 = n5261 ^ n2306 ^ 1'b0 ;
  assign n16640 = n5759 & ~n16639 ;
  assign n16641 = n365 & n16640 ;
  assign n16642 = n16641 ^ n9934 ^ 1'b0 ;
  assign n16643 = ( n1980 & n2532 ) | ( n1980 & n3122 ) | ( n2532 & n3122 ) ;
  assign n16644 = n16643 ^ n6448 ^ n1506 ;
  assign n16645 = n16644 ^ n8633 ^ n8294 ;
  assign n16646 = n6991 | n16645 ;
  assign n16647 = n15039 | n16646 ;
  assign n16648 = n4334 & n6486 ;
  assign n16649 = n16648 ^ n9882 ^ 1'b0 ;
  assign n16650 = n16649 ^ n13831 ^ 1'b0 ;
  assign n16652 = ( x97 & n6615 ) | ( x97 & n16643 ) | ( n6615 & n16643 ) ;
  assign n16651 = n1264 & n15509 ;
  assign n16653 = n16652 ^ n16651 ^ 1'b0 ;
  assign n16654 = n6465 & ~n7304 ;
  assign n16655 = n5143 & n14655 ;
  assign n16656 = n16655 ^ n3051 ^ 1'b0 ;
  assign n16657 = n2527 ^ x186 ^ 1'b0 ;
  assign n16658 = n16656 & n16657 ;
  assign n16659 = ~n2901 & n16658 ;
  assign n16660 = n16659 ^ n8670 ^ n1487 ;
  assign n16661 = n3080 | n9860 ;
  assign n16674 = n9972 ^ n4097 ^ 1'b0 ;
  assign n16662 = n1797 | n7733 ;
  assign n16663 = n16662 ^ n7816 ^ n976 ;
  assign n16664 = n1200 & ~n16663 ;
  assign n16665 = n16664 ^ n2315 ^ 1'b0 ;
  assign n16666 = n11232 & ~n16665 ;
  assign n16667 = ~n7987 & n10492 ;
  assign n16668 = n16667 ^ n3568 ^ 1'b0 ;
  assign n16669 = n10308 ^ n3485 ^ 1'b0 ;
  assign n16670 = n16668 | n16669 ;
  assign n16671 = n16666 & ~n16670 ;
  assign n16672 = n16671 ^ n4938 ^ 1'b0 ;
  assign n16673 = n13866 & ~n16672 ;
  assign n16675 = n16674 ^ n16673 ^ 1'b0 ;
  assign n16677 = ~n1832 & n11852 ;
  assign n16676 = n6041 | n8904 ;
  assign n16678 = n16677 ^ n16676 ^ 1'b0 ;
  assign n16679 = x117 & ~n6653 ;
  assign n16680 = n16679 ^ n13997 ^ 1'b0 ;
  assign n16681 = n6177 & n16680 ;
  assign n16682 = n5221 & n5901 ;
  assign n16683 = n16682 ^ n10695 ^ 1'b0 ;
  assign n16684 = n922 & ~n16683 ;
  assign n16685 = n1537 & ~n11759 ;
  assign n16686 = n6693 & ~n10603 ;
  assign n16687 = n16686 ^ n13094 ^ n8467 ;
  assign n16688 = n2603 & n16687 ;
  assign n16689 = n13691 ^ n9916 ^ n4893 ;
  assign n16690 = n4845 ^ n3812 ^ 1'b0 ;
  assign n16691 = n16690 ^ n7016 ^ 1'b0 ;
  assign n16692 = ~n5371 & n14638 ;
  assign n16693 = n13108 & n16692 ;
  assign n16697 = x44 & ~n4369 ;
  assign n16698 = ( n5475 & n13151 ) | ( n5475 & n16697 ) | ( n13151 & n16697 ) ;
  assign n16699 = n8209 & n16698 ;
  assign n16700 = n14623 & n16699 ;
  assign n16701 = n16700 ^ n8447 ^ n3622 ;
  assign n16702 = n10257 & ~n16701 ;
  assign n16694 = ( n1407 & ~n4078 ) | ( n1407 & n6723 ) | ( ~n4078 & n6723 ) ;
  assign n16695 = n11972 ^ n6202 ^ n2186 ;
  assign n16696 = n16694 & ~n16695 ;
  assign n16703 = n16702 ^ n16696 ^ n13331 ;
  assign n16704 = n16703 ^ n10092 ^ n8168 ;
  assign n16705 = ~n1122 & n1725 ;
  assign n16706 = n16705 ^ n14401 ^ 1'b0 ;
  assign n16707 = n509 & ~n5530 ;
  assign n16708 = n6060 & ~n16707 ;
  assign n16709 = ~n16706 & n16708 ;
  assign n16710 = ( n1367 & n3549 ) | ( n1367 & ~n16709 ) | ( n3549 & ~n16709 ) ;
  assign n16711 = ( n2334 & n5353 ) | ( n2334 & n16710 ) | ( n5353 & n16710 ) ;
  assign n16712 = n4585 | n5038 ;
  assign n16713 = n6292 | n16712 ;
  assign n16714 = n5358 & n7590 ;
  assign n16715 = ( ~n11426 & n15526 ) | ( ~n11426 & n16714 ) | ( n15526 & n16714 ) ;
  assign n16716 = n6071 & ~n16715 ;
  assign n16717 = ~n3297 & n16716 ;
  assign n16718 = ( n6431 & n16713 ) | ( n6431 & n16717 ) | ( n16713 & n16717 ) ;
  assign n16719 = ~n10157 & n14372 ;
  assign n16720 = n16718 & n16719 ;
  assign n16721 = ( n4117 & ~n11682 ) | ( n4117 & n12841 ) | ( ~n11682 & n12841 ) ;
  assign n16722 = n16721 ^ n6681 ^ n6147 ;
  assign n16723 = ~n3452 & n12362 ;
  assign n16724 = n617 & ~n7193 ;
  assign n16725 = n16723 & n16724 ;
  assign n16726 = n1452 & n16725 ;
  assign n16727 = n8315 & ~n13433 ;
  assign n16728 = ~n14372 & n16727 ;
  assign n16729 = n16728 ^ n8015 ^ 1'b0 ;
  assign n16730 = n9063 & n16729 ;
  assign n16731 = n6400 ^ n851 ^ 1'b0 ;
  assign n16732 = n16731 ^ n3262 ^ 1'b0 ;
  assign n16733 = n16732 ^ n14841 ^ 1'b0 ;
  assign n16734 = ~n7833 & n16733 ;
  assign n16735 = n5509 & ~n6215 ;
  assign n16736 = n11753 | n16735 ;
  assign n16739 = n7680 ^ n1620 ^ n927 ;
  assign n16737 = ( n495 & n4519 ) | ( n495 & n5740 ) | ( n4519 & n5740 ) ;
  assign n16738 = ( n3173 & n6381 ) | ( n3173 & n16737 ) | ( n6381 & n16737 ) ;
  assign n16740 = n16739 ^ n16738 ^ 1'b0 ;
  assign n16741 = n16740 ^ n3767 ^ 1'b0 ;
  assign n16742 = ~n16736 & n16741 ;
  assign n16743 = n731 & n7727 ;
  assign n16744 = ~n12165 & n16743 ;
  assign n16745 = n8642 ^ n5470 ^ 1'b0 ;
  assign n16746 = n16744 | n16745 ;
  assign n16747 = n12471 ^ n2651 ^ 1'b0 ;
  assign n16748 = n4416 & n16747 ;
  assign n16749 = ~n12271 & n15410 ;
  assign n16750 = ( n4993 & ~n8058 ) | ( n4993 & n10321 ) | ( ~n8058 & n10321 ) ;
  assign n16751 = ( n3719 & ~n7426 ) | ( n3719 & n16750 ) | ( ~n7426 & n16750 ) ;
  assign n16755 = ( n1415 & ~n12575 ) | ( n1415 & n14754 ) | ( ~n12575 & n14754 ) ;
  assign n16752 = n8374 ^ n675 ^ 1'b0 ;
  assign n16753 = n1999 & ~n16752 ;
  assign n16754 = n5989 & n16753 ;
  assign n16756 = n16755 ^ n16754 ^ 1'b0 ;
  assign n16757 = n10753 ^ n5815 ^ 1'b0 ;
  assign n16758 = n6862 & n16757 ;
  assign n16759 = n6972 ^ n3730 ^ n823 ;
  assign n16760 = n16759 ^ n7172 ^ 1'b0 ;
  assign n16761 = ~n4531 & n16760 ;
  assign n16762 = n2312 & n7200 ;
  assign n16763 = n16762 ^ n15424 ^ n1606 ;
  assign n16769 = n13346 ^ n10328 ^ 1'b0 ;
  assign n16764 = n16413 ^ n8057 ^ 1'b0 ;
  assign n16765 = ~n14265 & n16764 ;
  assign n16766 = ~n10948 & n13403 ;
  assign n16767 = n9240 & n16766 ;
  assign n16768 = n16765 & ~n16767 ;
  assign n16770 = n16769 ^ n16768 ^ 1'b0 ;
  assign n16771 = n13498 ^ n6555 ^ 1'b0 ;
  assign n16772 = n7218 & ~n14711 ;
  assign n16773 = n11895 & n16772 ;
  assign n16774 = n16773 ^ n1387 ^ 1'b0 ;
  assign n16776 = n8081 ^ n3753 ^ n3613 ;
  assign n16775 = n9370 & ~n16130 ;
  assign n16777 = n16776 ^ n16775 ^ 1'b0 ;
  assign n16778 = n16774 & ~n16777 ;
  assign n16779 = n5330 & n16778 ;
  assign n16780 = n2814 | n2943 ;
  assign n16781 = n16780 ^ n3457 ^ 1'b0 ;
  assign n16782 = n16781 ^ n8083 ^ 1'b0 ;
  assign n16783 = ~n16488 & n16782 ;
  assign n16784 = ~n16779 & n16783 ;
  assign n16785 = ~n2798 & n16784 ;
  assign n16786 = ~n7425 & n9312 ;
  assign n16787 = n16786 ^ n5839 ^ 1'b0 ;
  assign n16788 = n13806 | n16787 ;
  assign n16789 = n16788 ^ n8067 ^ n2471 ;
  assign n16790 = ~n2563 & n16767 ;
  assign n16791 = n7361 & ~n14382 ;
  assign n16792 = n16791 ^ n6968 ^ 1'b0 ;
  assign n16793 = n11046 & n16792 ;
  assign n16794 = n16793 ^ n9549 ^ 1'b0 ;
  assign n16795 = ( n8012 & n13809 ) | ( n8012 & ~n16424 ) | ( n13809 & ~n16424 ) ;
  assign n16796 = n1622 & n13050 ;
  assign n16797 = n3190 ^ n3156 ^ 1'b0 ;
  assign n16798 = ( n4095 & ~n4256 ) | ( n4095 & n16797 ) | ( ~n4256 & n16797 ) ;
  assign n16799 = n16798 ^ n4060 ^ 1'b0 ;
  assign n16800 = x69 & n16799 ;
  assign n16801 = ~n13584 & n16800 ;
  assign n16802 = n16801 ^ n16059 ^ 1'b0 ;
  assign n16803 = n5219 | n6428 ;
  assign n16804 = n1131 & ~n16803 ;
  assign n16805 = n8081 | n12814 ;
  assign n16806 = n9840 & ~n16805 ;
  assign n16807 = n16806 ^ n3821 ^ 1'b0 ;
  assign n16812 = ~n1504 & n2188 ;
  assign n16813 = n2357 ^ n1073 ^ 1'b0 ;
  assign n16814 = n16812 & ~n16813 ;
  assign n16808 = n1276 & ~n4454 ;
  assign n16809 = n16808 ^ n5018 ^ 1'b0 ;
  assign n16810 = n16809 ^ n4615 ^ 1'b0 ;
  assign n16811 = n1715 & ~n16810 ;
  assign n16815 = n16814 ^ n16811 ^ n16022 ;
  assign n16816 = n16815 ^ n2585 ^ n347 ;
  assign n16817 = x161 & ~n9360 ;
  assign n16818 = x172 & n3527 ;
  assign n16819 = ~n706 & n16818 ;
  assign n16820 = n9642 ^ n5736 ^ 1'b0 ;
  assign n16821 = ~n9454 & n16820 ;
  assign n16822 = n3494 ^ n1569 ^ 1'b0 ;
  assign n16823 = n6162 & ~n16822 ;
  assign n16824 = ( n6329 & n16821 ) | ( n6329 & n16823 ) | ( n16821 & n16823 ) ;
  assign n16825 = n16824 ^ n2412 ^ 1'b0 ;
  assign n16827 = ~n1392 & n9536 ;
  assign n16828 = n14886 | n16827 ;
  assign n16826 = n11747 ^ n8716 ^ n5907 ;
  assign n16829 = n16828 ^ n16826 ^ 1'b0 ;
  assign n16830 = n1220 & n5263 ;
  assign n16831 = n12145 & n16830 ;
  assign n16832 = n12878 & n16831 ;
  assign n16833 = n16832 ^ n15402 ^ n6231 ;
  assign n16834 = n3474 & n13350 ;
  assign n16835 = n11232 & n12273 ;
  assign n16836 = n16834 & n16835 ;
  assign n16837 = ( n576 & n1525 ) | ( n576 & ~n6503 ) | ( n1525 & ~n6503 ) ;
  assign n16838 = n9102 ^ n3965 ^ 1'b0 ;
  assign n16839 = ~n16837 & n16838 ;
  assign n16847 = n8257 | n12373 ;
  assign n16845 = n11488 ^ n2026 ^ 1'b0 ;
  assign n16846 = n16845 ^ n4784 ^ 1'b0 ;
  assign n16840 = ( ~n3619 & n10696 ) | ( ~n3619 & n13213 ) | ( n10696 & n13213 ) ;
  assign n16841 = n5506 ^ n1557 ^ 1'b0 ;
  assign n16842 = ~n4034 & n16841 ;
  assign n16843 = n16842 ^ n6961 ^ 1'b0 ;
  assign n16844 = n16840 | n16843 ;
  assign n16848 = n16847 ^ n16846 ^ n16844 ;
  assign n16849 = n4614 & ~n16848 ;
  assign n16850 = n544 | n6839 ;
  assign n16851 = n10007 & ~n16850 ;
  assign n16852 = ~n6352 & n9815 ;
  assign n16853 = n14786 | n16852 ;
  assign n16854 = n16853 ^ n1181 ^ 1'b0 ;
  assign n16855 = ~n405 & n8774 ;
  assign n16856 = n16855 ^ n10828 ^ 1'b0 ;
  assign n16857 = n4669 & n16856 ;
  assign n16858 = x18 | n16707 ;
  assign n16859 = ( n5572 & n12174 ) | ( n5572 & n16858 ) | ( n12174 & n16858 ) ;
  assign n16860 = ( n1383 & ~n2106 ) | ( n1383 & n4937 ) | ( ~n2106 & n4937 ) ;
  assign n16861 = ( n10429 & ~n13243 ) | ( n10429 & n16860 ) | ( ~n13243 & n16860 ) ;
  assign n16863 = n5715 ^ n5042 ^ n1412 ;
  assign n16864 = n6039 & ~n16863 ;
  assign n16862 = n1821 & ~n1860 ;
  assign n16865 = n16864 ^ n16862 ^ n2489 ;
  assign n16866 = n3527 & ~n9643 ;
  assign n16867 = ( n464 & ~n6467 ) | ( n464 & n7141 ) | ( ~n6467 & n7141 ) ;
  assign n16868 = n10432 ^ n3476 ^ 1'b0 ;
  assign n16869 = n6960 & n16868 ;
  assign n16870 = n16867 | n16869 ;
  assign n16871 = n16866 & ~n16870 ;
  assign n16872 = n11099 & n16871 ;
  assign n16873 = ~n2513 & n4987 ;
  assign n16874 = n2893 & n16873 ;
  assign n16875 = n16635 & ~n16874 ;
  assign n16876 = n16875 ^ n12828 ^ 1'b0 ;
  assign n16877 = ( n11308 & ~n12532 ) | ( n11308 & n16876 ) | ( ~n12532 & n16876 ) ;
  assign n16878 = ~n10495 & n16877 ;
  assign n16879 = n7766 | n16878 ;
  assign n16880 = n16879 ^ n5891 ^ 1'b0 ;
  assign n16881 = n11219 ^ n3740 ^ 1'b0 ;
  assign n16882 = n16881 ^ n9759 ^ n6835 ;
  assign n16883 = n16121 ^ n11571 ^ 1'b0 ;
  assign n16884 = n16883 ^ n3304 ^ 1'b0 ;
  assign n16885 = ~n13243 & n16884 ;
  assign n16886 = n4156 ^ n3497 ^ n2469 ;
  assign n16887 = n16425 ^ n377 ^ 1'b0 ;
  assign n16888 = n9976 & ~n16887 ;
  assign n16889 = ~n16886 & n16888 ;
  assign n16890 = n2677 ^ n1895 ^ x60 ;
  assign n16891 = ~n15863 & n16890 ;
  assign n16892 = n2825 ^ n2426 ^ 1'b0 ;
  assign n16893 = n2621 ^ n1257 ^ 1'b0 ;
  assign n16894 = ~n2154 & n3962 ;
  assign n16895 = n8987 & n16894 ;
  assign n16896 = n3475 | n16895 ;
  assign n16897 = n16412 & ~n16896 ;
  assign n16898 = n3599 | n6558 ;
  assign n16899 = n16898 ^ n8273 ^ 1'b0 ;
  assign n16900 = n13622 & ~n16899 ;
  assign n16901 = n16900 ^ n6989 ^ 1'b0 ;
  assign n16902 = n2394 | n5665 ;
  assign n16903 = n16902 ^ n1918 ^ 1'b0 ;
  assign n16904 = n6458 | n10168 ;
  assign n16905 = n4787 & ~n16904 ;
  assign n16906 = n5246 ^ n3556 ^ 1'b0 ;
  assign n16907 = n16380 ^ x202 ^ 1'b0 ;
  assign n16908 = ( n1532 & ~n3402 ) | ( n1532 & n9086 ) | ( ~n3402 & n9086 ) ;
  assign n16909 = n10577 & ~n16908 ;
  assign n16910 = n7267 & ~n7355 ;
  assign n16911 = n16910 ^ n6027 ^ 1'b0 ;
  assign n16912 = n16911 ^ n12314 ^ 1'b0 ;
  assign n16913 = n1999 & n12738 ;
  assign n16914 = n16912 & n16913 ;
  assign n16915 = n11070 ^ n4255 ^ n4151 ;
  assign n16927 = n9061 ^ n3069 ^ n1439 ;
  assign n16928 = n16927 ^ n13977 ^ n10777 ;
  assign n16925 = n10060 | n11179 ;
  assign n16916 = x237 & ~n5842 ;
  assign n16917 = ~n6718 & n16916 ;
  assign n16918 = n8046 ^ n1624 ^ 1'b0 ;
  assign n16919 = ~n6897 & n16918 ;
  assign n16920 = n1308 & n16919 ;
  assign n16921 = n16917 & n16920 ;
  assign n16922 = n8587 & n13635 ;
  assign n16923 = ( n5038 & n9125 ) | ( n5038 & n16922 ) | ( n9125 & n16922 ) ;
  assign n16924 = ~n16921 & n16923 ;
  assign n16926 = n16925 ^ n16924 ^ 1'b0 ;
  assign n16929 = n16928 ^ n16926 ^ 1'b0 ;
  assign n16930 = n4061 ^ n876 ^ 1'b0 ;
  assign n16931 = ( ~x75 & n7943 ) | ( ~x75 & n16930 ) | ( n7943 & n16930 ) ;
  assign n16932 = n11053 ^ n7788 ^ 1'b0 ;
  assign n16936 = ~n1322 & n2567 ;
  assign n16937 = n5134 & n16936 ;
  assign n16938 = n603 & n16937 ;
  assign n16933 = n12805 ^ n941 ^ 1'b0 ;
  assign n16934 = n16933 ^ n12228 ^ 1'b0 ;
  assign n16935 = n2272 & n16934 ;
  assign n16939 = n16938 ^ n16935 ^ 1'b0 ;
  assign n16940 = n10425 | n16939 ;
  assign n16941 = n15958 ^ n7850 ^ 1'b0 ;
  assign n16942 = n6794 | n16941 ;
  assign n16943 = n16942 ^ n16197 ^ n8815 ;
  assign n16944 = n1529 & n3021 ;
  assign n16945 = n9692 & n16944 ;
  assign n16946 = n4282 ^ n3305 ^ x210 ;
  assign n16947 = n4234 | n16946 ;
  assign n16948 = n1976 & n2688 ;
  assign n16949 = n16697 & n16948 ;
  assign n16950 = n5761 & n16949 ;
  assign n16951 = n16950 ^ n4101 ^ 1'b0 ;
  assign n16952 = n16951 ^ n13764 ^ n3802 ;
  assign n16953 = n16947 | n16952 ;
  assign n16956 = n338 | n2160 ;
  assign n16957 = n10898 & ~n16956 ;
  assign n16954 = x120 & ~n13717 ;
  assign n16955 = ~n14365 & n16954 ;
  assign n16958 = n16957 ^ n16955 ^ 1'b0 ;
  assign n16959 = n5357 & ~n14612 ;
  assign n16960 = n3764 | n7244 ;
  assign n16961 = n16960 ^ n14758 ^ 1'b0 ;
  assign n16962 = ( n3327 & n16959 ) | ( n3327 & ~n16961 ) | ( n16959 & ~n16961 ) ;
  assign n16963 = ~n9642 & n14016 ;
  assign n16964 = ~n808 & n16963 ;
  assign n16965 = n16964 ^ n8253 ^ 1'b0 ;
  assign n16966 = n2133 & ~n16335 ;
  assign n16967 = n14016 | n14870 ;
  assign n16968 = ~n5463 & n16967 ;
  assign n16969 = n1047 | n7144 ;
  assign n16970 = n16969 ^ n10269 ^ n620 ;
  assign n16971 = n2927 & ~n6799 ;
  assign n16972 = ~n14057 & n16971 ;
  assign n16973 = ( n667 & n10636 ) | ( n667 & ~n16972 ) | ( n10636 & ~n16972 ) ;
  assign n16974 = ( n6587 & n10100 ) | ( n6587 & n13499 ) | ( n10100 & n13499 ) ;
  assign n16975 = n16974 ^ n9447 ^ 1'b0 ;
  assign n16976 = n6691 & ~n16975 ;
  assign n16977 = n8653 ^ n3381 ^ 1'b0 ;
  assign n16978 = ( n1413 & ~n14045 ) | ( n1413 & n16977 ) | ( ~n14045 & n16977 ) ;
  assign n16984 = n13972 ^ n1350 ^ 1'b0 ;
  assign n16985 = n6921 | n16984 ;
  assign n16986 = n16911 | n16985 ;
  assign n16979 = n10947 ^ n8075 ^ 1'b0 ;
  assign n16980 = n803 & n1080 ;
  assign n16981 = ~n5760 & n16980 ;
  assign n16982 = ( n2469 & ~n11703 ) | ( n2469 & n16981 ) | ( ~n11703 & n16981 ) ;
  assign n16983 = n16979 & n16982 ;
  assign n16987 = n16986 ^ n16983 ^ 1'b0 ;
  assign n16993 = n1727 | n6005 ;
  assign n16991 = n1284 ^ n545 ^ 1'b0 ;
  assign n16988 = n1055 & n1761 ;
  assign n16989 = ~n1010 & n16988 ;
  assign n16990 = n11581 | n16989 ;
  assign n16992 = n16991 ^ n16990 ^ 1'b0 ;
  assign n16994 = n16993 ^ n16992 ^ n461 ;
  assign n17001 = ( x146 & ~n4047 ) | ( x146 & n5213 ) | ( ~n4047 & n5213 ) ;
  assign n16995 = n1250 | n1626 ;
  assign n16996 = n8722 | n16995 ;
  assign n16997 = n16996 ^ n13645 ^ 1'b0 ;
  assign n16998 = n3555 & ~n10748 ;
  assign n16999 = n16997 & n16998 ;
  assign n17000 = n12663 & n16999 ;
  assign n17002 = n17001 ^ n17000 ^ 1'b0 ;
  assign n17003 = n17002 ^ n7134 ^ 1'b0 ;
  assign n17004 = ~n15835 & n17003 ;
  assign n17005 = n8491 | n9193 ;
  assign n17006 = n17005 ^ n9061 ^ 1'b0 ;
  assign n17007 = n14847 ^ n9321 ^ n1105 ;
  assign n17008 = n12106 & n17007 ;
  assign n17009 = ~n3347 & n17008 ;
  assign n17010 = n17009 ^ n2708 ^ 1'b0 ;
  assign n17011 = n6403 & n17010 ;
  assign n17012 = n10303 ^ n8742 ^ 1'b0 ;
  assign n17013 = ( n1120 & n2473 ) | ( n1120 & ~n12019 ) | ( n2473 & ~n12019 ) ;
  assign n17014 = ( n7800 & n17012 ) | ( n7800 & ~n17013 ) | ( n17012 & ~n17013 ) ;
  assign n17015 = ( ~n320 & n4139 ) | ( ~n320 & n4157 ) | ( n4139 & n4157 ) ;
  assign n17016 = n17015 ^ n5488 ^ 1'b0 ;
  assign n17017 = n2553 | n17016 ;
  assign n17018 = n1693 | n3599 ;
  assign n17019 = n3837 & n10440 ;
  assign n17020 = n17018 & n17019 ;
  assign n17021 = x110 & ~n15335 ;
  assign n17022 = n17021 ^ n9563 ^ 1'b0 ;
  assign n17023 = n11009 & ~n16848 ;
  assign n17024 = n5119 & n5982 ;
  assign n17025 = n17024 ^ n10281 ^ 1'b0 ;
  assign n17026 = n630 | n9873 ;
  assign n17027 = n5408 & ~n17026 ;
  assign n17028 = n8638 & n11087 ;
  assign n17029 = n16523 & n17028 ;
  assign n17032 = n14907 ^ n847 ^ 1'b0 ;
  assign n17033 = n3269 | n17032 ;
  assign n17034 = n804 | n1972 ;
  assign n17035 = n17034 ^ n7915 ^ 1'b0 ;
  assign n17036 = ( n7342 & n17033 ) | ( n7342 & ~n17035 ) | ( n17033 & ~n17035 ) ;
  assign n17037 = n2185 & ~n17036 ;
  assign n17030 = n14274 ^ n10209 ^ n7155 ;
  assign n17031 = n13043 | n17030 ;
  assign n17038 = n17037 ^ n17031 ^ 1'b0 ;
  assign n17041 = n5660 ^ n3040 ^ 1'b0 ;
  assign n17042 = n17041 ^ n11459 ^ n3109 ;
  assign n17039 = n2462 & n3052 ;
  assign n17040 = n13962 & n17039 ;
  assign n17043 = n17042 ^ n17040 ^ 1'b0 ;
  assign n17044 = ~n6385 & n10164 ;
  assign n17045 = n12761 ^ n3410 ^ 1'b0 ;
  assign n17046 = n11231 | n13437 ;
  assign n17047 = n17046 ^ n3937 ^ 1'b0 ;
  assign n17048 = n3039 & ~n6103 ;
  assign n17049 = n6376 & n17048 ;
  assign n17050 = n17049 ^ n5228 ^ n4937 ;
  assign n17051 = n5974 | n9482 ;
  assign n17052 = ~n6836 & n17051 ;
  assign n17053 = ( n10112 & n17050 ) | ( n10112 & n17052 ) | ( n17050 & n17052 ) ;
  assign n17054 = n2948 ^ n1382 ^ 1'b0 ;
  assign n17055 = n16640 & n17054 ;
  assign n17056 = ( n2048 & ~n6968 ) | ( n2048 & n7522 ) | ( ~n6968 & n7522 ) ;
  assign n17057 = n17056 ^ n13399 ^ n8448 ;
  assign n17058 = n2643 & ~n17057 ;
  assign n17059 = n17058 ^ n16757 ^ 1'b0 ;
  assign n17060 = n7774 ^ x97 ^ 1'b0 ;
  assign n17061 = ~n1900 & n17060 ;
  assign n17062 = n6075 & n17061 ;
  assign n17063 = n17062 ^ n8497 ^ 1'b0 ;
  assign n17064 = ( n5468 & n5936 ) | ( n5468 & n8813 ) | ( n5936 & n8813 ) ;
  assign n17065 = ~n9672 & n17064 ;
  assign n17066 = n17065 ^ n6130 ^ 1'b0 ;
  assign n17067 = ( n4565 & n7167 ) | ( n4565 & n15209 ) | ( n7167 & n15209 ) ;
  assign n17068 = n15692 ^ n5595 ^ x169 ;
  assign n17069 = ~n3437 & n7186 ;
  assign n17070 = n10429 | n11462 ;
  assign n17071 = n17070 ^ x82 ^ 1'b0 ;
  assign n17072 = n16312 & ~n17071 ;
  assign n17073 = ( ~n577 & n6124 ) | ( ~n577 & n12693 ) | ( n6124 & n12693 ) ;
  assign n17074 = n17073 ^ n15142 ^ n3624 ;
  assign n17075 = n10009 ^ x160 ^ 1'b0 ;
  assign n17076 = n6179 ^ n1778 ^ n396 ;
  assign n17077 = ( n1882 & n5039 ) | ( n1882 & ~n17076 ) | ( n5039 & ~n17076 ) ;
  assign n17078 = ~n1319 & n17077 ;
  assign n17079 = n7858 & n10820 ;
  assign n17080 = ~n5407 & n17079 ;
  assign n17081 = n6353 ^ n464 ^ 1'b0 ;
  assign n17082 = n499 ^ x1 ^ 1'b0 ;
  assign n17083 = n17082 ^ n8363 ^ n5821 ;
  assign n17084 = n17083 ^ n10863 ^ 1'b0 ;
  assign n17085 = ~n5539 & n6742 ;
  assign n17086 = n1126 & n17085 ;
  assign n17087 = n3300 & ~n17086 ;
  assign n17088 = n17087 ^ n11227 ^ 1'b0 ;
  assign n17093 = ( n5503 & n12109 ) | ( n5503 & ~n12239 ) | ( n12109 & ~n12239 ) ;
  assign n17089 = n363 & ~n3707 ;
  assign n17090 = n11667 & ~n17089 ;
  assign n17091 = n6099 & n17090 ;
  assign n17092 = n4045 & ~n17091 ;
  assign n17094 = n17093 ^ n17092 ^ 1'b0 ;
  assign n17095 = n17094 ^ n5655 ^ 1'b0 ;
  assign n17097 = n14754 ^ n9839 ^ 1'b0 ;
  assign n17098 = ~n3749 & n17097 ;
  assign n17096 = n8319 & ~n12721 ;
  assign n17099 = n17098 ^ n17096 ^ 1'b0 ;
  assign n17100 = n5905 ^ n3133 ^ 1'b0 ;
  assign n17101 = n3591 | n17100 ;
  assign n17105 = n3093 & ~n7536 ;
  assign n17106 = n14527 & n17105 ;
  assign n17103 = ( ~n1201 & n7232 ) | ( ~n1201 & n12498 ) | ( n7232 & n12498 ) ;
  assign n17102 = n2635 ^ n469 ^ n294 ;
  assign n17104 = n17103 ^ n17102 ^ 1'b0 ;
  assign n17107 = n17106 ^ n17104 ^ n5681 ;
  assign n17108 = n4912 ^ n2426 ^ 1'b0 ;
  assign n17116 = n4013 | n7180 ;
  assign n17115 = n2004 ^ n1354 ^ 1'b0 ;
  assign n17110 = n7509 & ~n11007 ;
  assign n17111 = ~n8556 & n17110 ;
  assign n17109 = ~n455 & n6730 ;
  assign n17112 = n17111 ^ n17109 ^ 1'b0 ;
  assign n17113 = n16424 & n17112 ;
  assign n17114 = n750 & n17113 ;
  assign n17117 = n17116 ^ n17115 ^ n17114 ;
  assign n17118 = n6991 | n7611 ;
  assign n17119 = n17118 ^ n4132 ^ 1'b0 ;
  assign n17120 = n10909 & ~n17119 ;
  assign n17121 = n7641 & n17120 ;
  assign n17122 = n17121 ^ n9143 ^ 1'b0 ;
  assign n17123 = ~n9641 & n17122 ;
  assign n17124 = ( n293 & n2648 ) | ( n293 & ~n10067 ) | ( n2648 & ~n10067 ) ;
  assign n17125 = n7549 | n17124 ;
  assign n17126 = n17123 | n17125 ;
  assign n17127 = ~n2671 & n8099 ;
  assign n17128 = n15567 & n17127 ;
  assign n17129 = n16370 ^ n6542 ^ 1'b0 ;
  assign n17130 = n5781 | n17129 ;
  assign n17131 = n17130 ^ n9470 ^ 1'b0 ;
  assign n17132 = n8526 | n12387 ;
  assign n17133 = n3203 & ~n17132 ;
  assign n17134 = ( n3016 & n4720 ) | ( n3016 & ~n16046 ) | ( n4720 & ~n16046 ) ;
  assign n17135 = n17134 ^ n3361 ^ n1690 ;
  assign n17136 = ~n2596 & n17135 ;
  assign n17137 = n17136 ^ n16701 ^ n2713 ;
  assign n17138 = n5209 ^ n3328 ^ 1'b0 ;
  assign n17139 = n5586 | n8688 ;
  assign n17140 = n17139 ^ n12334 ^ 1'b0 ;
  assign n17141 = n10844 ^ n1037 ^ 1'b0 ;
  assign n17142 = n17140 & ~n17141 ;
  assign n17143 = n6829 ^ n5436 ^ 1'b0 ;
  assign n17144 = n2800 ^ n1098 ^ x223 ;
  assign n17145 = n7159 & ~n17144 ;
  assign n17146 = n14634 & n17145 ;
  assign n17147 = ( n9931 & ~n17143 ) | ( n9931 & n17146 ) | ( ~n17143 & n17146 ) ;
  assign n17148 = n13038 ^ n10247 ^ n9201 ;
  assign n17149 = n6437 & n8284 ;
  assign n17150 = ( x88 & n4179 ) | ( x88 & ~n17149 ) | ( n4179 & ~n17149 ) ;
  assign n17151 = n5545 & n12839 ;
  assign n17152 = n17151 ^ n11420 ^ 1'b0 ;
  assign n17153 = n14954 ^ n4132 ^ n3795 ;
  assign n17154 = n4294 & ~n12659 ;
  assign n17155 = n17154 ^ n310 ^ 1'b0 ;
  assign n17156 = ( n2106 & n9634 ) | ( n2106 & n16811 ) | ( n9634 & n16811 ) ;
  assign n17157 = n4187 & n13975 ;
  assign n17158 = ~n8956 & n17157 ;
  assign n17159 = n17158 ^ n8253 ^ n5287 ;
  assign n17160 = n5014 | n11977 ;
  assign n17161 = x225 | n5107 ;
  assign n17162 = n17161 ^ n15515 ^ 1'b0 ;
  assign n17163 = n2886 & n17162 ;
  assign n17164 = n17160 | n17163 ;
  assign n17165 = ( ~n1786 & n6414 ) | ( ~n1786 & n17164 ) | ( n6414 & n17164 ) ;
  assign n17166 = ~n4070 & n6450 ;
  assign n17170 = n2078 | n2251 ;
  assign n17167 = n14023 ^ n6805 ^ 1'b0 ;
  assign n17168 = n8913 ^ n2860 ^ 1'b0 ;
  assign n17169 = ( n6963 & n17167 ) | ( n6963 & n17168 ) | ( n17167 & n17168 ) ;
  assign n17171 = n17170 ^ n17169 ^ n10623 ;
  assign n17172 = ( n3275 & n9857 ) | ( n3275 & ~n12570 ) | ( n9857 & ~n12570 ) ;
  assign n17173 = n4172 ^ n1993 ^ 1'b0 ;
  assign n17174 = ~n8717 & n17173 ;
  assign n17175 = n13391 ^ n8240 ^ 1'b0 ;
  assign n17176 = ~n1022 & n6606 ;
  assign n17177 = n17175 & n17176 ;
  assign n17178 = n17177 ^ n12423 ^ 1'b0 ;
  assign n17179 = n17174 & n17178 ;
  assign n17180 = n8965 & ~n13830 ;
  assign n17181 = n17179 & n17180 ;
  assign n17182 = ~n13886 & n17181 ;
  assign n17183 = n5055 ^ n2819 ^ 1'b0 ;
  assign n17184 = n1359 | n17183 ;
  assign n17185 = ~n7718 & n17184 ;
  assign n17186 = n6868 ^ n1206 ^ 1'b0 ;
  assign n17187 = n17185 & n17186 ;
  assign n17188 = n11557 ^ n10660 ^ n5011 ;
  assign n17189 = ( n6375 & n14116 ) | ( n6375 & ~n17188 ) | ( n14116 & ~n17188 ) ;
  assign n17190 = ~n1836 & n3140 ;
  assign n17191 = n17190 ^ n2236 ^ 1'b0 ;
  assign n17192 = n7543 | n17191 ;
  assign n17193 = n9832 ^ n2515 ^ 1'b0 ;
  assign n17195 = n8021 & n9685 ;
  assign n17194 = n4861 & n13014 ;
  assign n17196 = n17195 ^ n17194 ^ n8145 ;
  assign n17197 = n4321 | n16021 ;
  assign n17198 = n2407 & ~n13017 ;
  assign n17199 = ~n7956 & n17198 ;
  assign n17200 = n14641 ^ n2471 ^ 1'b0 ;
  assign n17201 = n17199 | n17200 ;
  assign n17202 = n17161 ^ n4003 ^ 1'b0 ;
  assign n17203 = n11601 ^ n10748 ^ 1'b0 ;
  assign n17204 = ~n17202 & n17203 ;
  assign n17205 = n2099 ^ n279 ^ 1'b0 ;
  assign n17206 = n2230 & n17205 ;
  assign n17207 = ~n9723 & n17206 ;
  assign n17208 = n2386 & n17207 ;
  assign n17209 = n3932 & n17208 ;
  assign n17210 = n14307 | n17209 ;
  assign n17211 = n17210 ^ n14551 ^ 1'b0 ;
  assign n17212 = n11768 ^ n3750 ^ n3158 ;
  assign n17213 = n966 & ~n17212 ;
  assign n17214 = n17213 ^ n5398 ^ 1'b0 ;
  assign n17215 = n9076 ^ n5186 ^ 1'b0 ;
  assign n17216 = n4422 & ~n4468 ;
  assign n17217 = n4561 & n17216 ;
  assign n17218 = n5066 & ~n17217 ;
  assign n17219 = n17218 ^ n11617 ^ 1'b0 ;
  assign n17220 = n5786 & ~n17219 ;
  assign n17221 = ~n17215 & n17220 ;
  assign n17222 = n3297 ^ n1211 ^ 1'b0 ;
  assign n17223 = n2931 | n17222 ;
  assign n17224 = n17223 ^ n5616 ^ n403 ;
  assign n17225 = n1886 | n7670 ;
  assign n17226 = n9506 ^ n1795 ^ 1'b0 ;
  assign n17227 = ~n12615 & n17226 ;
  assign n17228 = n11048 | n13680 ;
  assign n17229 = n17228 ^ n12912 ^ n9863 ;
  assign n17230 = n6399 ^ n5193 ^ 1'b0 ;
  assign n17231 = n6994 & ~n17230 ;
  assign n17232 = n10145 ^ n8670 ^ 1'b0 ;
  assign n17233 = n13865 & ~n17232 ;
  assign n17234 = n11759 ^ n8524 ^ 1'b0 ;
  assign n17235 = n1182 & ~n13176 ;
  assign n17236 = n17235 ^ n11800 ^ 1'b0 ;
  assign n17237 = n17236 ^ n9640 ^ 1'b0 ;
  assign n17238 = ( n17233 & n17234 ) | ( n17233 & ~n17237 ) | ( n17234 & ~n17237 ) ;
  assign n17239 = n14410 ^ n12068 ^ n428 ;
  assign n17240 = n10884 | n13789 ;
  assign n17241 = n1780 | n17240 ;
  assign n17242 = n17241 ^ n11010 ^ n8497 ;
  assign n17243 = n3902 ^ n976 ^ 1'b0 ;
  assign n17244 = n1079 & n1641 ;
  assign n17245 = n17244 ^ n11703 ^ 1'b0 ;
  assign n17246 = ( n5685 & ~n7144 ) | ( n5685 & n8909 ) | ( ~n7144 & n8909 ) ;
  assign n17247 = n4346 | n17246 ;
  assign n17248 = n17247 ^ n15022 ^ 1'b0 ;
  assign n17249 = n3151 & ~n6428 ;
  assign n17250 = ~n8440 & n17249 ;
  assign n17251 = x51 & n1409 ;
  assign n17252 = n17251 ^ n11758 ^ 1'b0 ;
  assign n17254 = ~n2645 & n7276 ;
  assign n17255 = ~n4001 & n17254 ;
  assign n17256 = n2070 & n17255 ;
  assign n17253 = n3669 & n15879 ;
  assign n17257 = n17256 ^ n17253 ^ 1'b0 ;
  assign n17258 = ~n4287 & n17257 ;
  assign n17259 = ( ~n17250 & n17252 ) | ( ~n17250 & n17258 ) | ( n17252 & n17258 ) ;
  assign n17260 = n3444 & ~n8750 ;
  assign n17261 = n17260 ^ n7342 ^ 1'b0 ;
  assign n17262 = ~n13284 & n16083 ;
  assign n17263 = ( n11474 & n16476 ) | ( n11474 & ~n17262 ) | ( n16476 & ~n17262 ) ;
  assign n17264 = n10341 ^ n7631 ^ 1'b0 ;
  assign n17265 = n3064 | n17264 ;
  assign n17266 = n17265 ^ n9486 ^ 1'b0 ;
  assign n17267 = n7069 | n14365 ;
  assign n17268 = n17267 ^ n2502 ^ 1'b0 ;
  assign n17269 = ~n2967 & n4120 ;
  assign n17270 = n17268 & n17269 ;
  assign n17271 = n12346 ^ n637 ^ 1'b0 ;
  assign n17272 = n5645 ^ n2506 ^ 1'b0 ;
  assign n17273 = ~n1671 & n17272 ;
  assign n17274 = n12036 ^ n1140 ^ 1'b0 ;
  assign n17275 = ~n9068 & n17274 ;
  assign n17276 = n17273 & n17275 ;
  assign n17277 = n3190 ^ n2594 ^ n1754 ;
  assign n17278 = n1962 | n17277 ;
  assign n17279 = ( n3096 & n6270 ) | ( n3096 & ~n17278 ) | ( n6270 & ~n17278 ) ;
  assign n17280 = n11390 & n17279 ;
  assign n17281 = ~n15629 & n17280 ;
  assign n17283 = n12622 ^ n2699 ^ 1'b0 ;
  assign n17284 = n5417 | n17283 ;
  assign n17282 = ( n5676 & n7427 ) | ( n5676 & ~n8903 ) | ( n7427 & ~n8903 ) ;
  assign n17285 = n17284 ^ n17282 ^ n9343 ;
  assign n17286 = ~n13970 & n17285 ;
  assign n17287 = n17286 ^ n9274 ^ n5356 ;
  assign n17288 = n2038 ^ n1105 ^ n639 ;
  assign n17289 = n5330 | n9008 ;
  assign n17292 = n11373 ^ n8293 ^ n2571 ;
  assign n17290 = ( n1773 & ~n7252 ) | ( n1773 & n10524 ) | ( ~n7252 & n10524 ) ;
  assign n17291 = n8309 & ~n17290 ;
  assign n17293 = n17292 ^ n17291 ^ 1'b0 ;
  assign n17295 = ( n879 & n1584 ) | ( n879 & ~n9255 ) | ( n1584 & ~n9255 ) ;
  assign n17294 = n9048 ^ n7088 ^ n2748 ;
  assign n17296 = n17295 ^ n17294 ^ n7420 ;
  assign n17297 = ( n4292 & ~n17293 ) | ( n4292 & n17296 ) | ( ~n17293 & n17296 ) ;
  assign n17300 = n8051 & n9537 ;
  assign n17301 = n15222 ^ n7250 ^ n6713 ;
  assign n17302 = n4063 & n6325 ;
  assign n17303 = n17302 ^ n8058 ^ 1'b0 ;
  assign n17304 = ~n17301 & n17303 ;
  assign n17305 = n17300 & ~n17304 ;
  assign n17298 = n9967 ^ x90 ^ 1'b0 ;
  assign n17299 = n4217 & n17298 ;
  assign n17306 = n17305 ^ n17299 ^ n4592 ;
  assign n17307 = ( n2515 & n8258 ) | ( n2515 & ~n9073 ) | ( n8258 & ~n9073 ) ;
  assign n17308 = n17307 ^ n3476 ^ 1'b0 ;
  assign n17309 = n11923 ^ n11122 ^ 1'b0 ;
  assign n17310 = n5610 & n17309 ;
  assign n17311 = n3996 & n17310 ;
  assign n17312 = n13481 ^ n4756 ^ 1'b0 ;
  assign n17313 = n9872 & n17312 ;
  assign n17314 = n17313 ^ n11575 ^ n5021 ;
  assign n17315 = ( n4517 & ~n10065 ) | ( n4517 & n12106 ) | ( ~n10065 & n12106 ) ;
  assign n17316 = n13800 | n17315 ;
  assign n17317 = n17316 ^ n8422 ^ 1'b0 ;
  assign n17318 = n16334 ^ n447 ^ 1'b0 ;
  assign n17319 = n2048 | n13835 ;
  assign n17320 = ( n1002 & n17318 ) | ( n1002 & ~n17319 ) | ( n17318 & ~n17319 ) ;
  assign n17321 = n3368 ^ x159 ^ 1'b0 ;
  assign n17322 = n17321 ^ n10463 ^ n4600 ;
  assign n17323 = n2606 & n4870 ;
  assign n17324 = n17323 ^ n7743 ^ 1'b0 ;
  assign n17325 = n15919 ^ n1881 ^ 1'b0 ;
  assign n17326 = ( n4546 & ~n5839 ) | ( n4546 & n7135 ) | ( ~n5839 & n7135 ) ;
  assign n17327 = ~n777 & n17326 ;
  assign n17328 = n14628 & n17327 ;
  assign n17329 = n17328 ^ n12861 ^ n3516 ;
  assign n17330 = n7966 | n13275 ;
  assign n17331 = n4223 | n17330 ;
  assign n17332 = n14861 ^ n10459 ^ n5833 ;
  assign n17333 = n3517 & n15320 ;
  assign n17334 = n1863 | n17333 ;
  assign n17335 = n13035 ^ n1010 ^ 1'b0 ;
  assign n17336 = n4086 & n10407 ;
  assign n17337 = ~n17335 & n17336 ;
  assign n17341 = ( n1339 & n1914 ) | ( n1339 & ~n7733 ) | ( n1914 & ~n7733 ) ;
  assign n17338 = n1635 | n3810 ;
  assign n17339 = n16830 & ~n17338 ;
  assign n17340 = n16964 & n17339 ;
  assign n17342 = n17341 ^ n17340 ^ 1'b0 ;
  assign n17343 = ~n10971 & n17342 ;
  assign n17344 = ( n4977 & n10898 ) | ( n4977 & n17343 ) | ( n10898 & n17343 ) ;
  assign n17345 = n1071 & ~n5217 ;
  assign n17346 = n14905 ^ n7088 ^ 1'b0 ;
  assign n17347 = n17346 ^ n3366 ^ 1'b0 ;
  assign n17348 = ~n17345 & n17347 ;
  assign n17349 = n4233 | n17348 ;
  assign n17350 = n13097 ^ n4163 ^ 1'b0 ;
  assign n17351 = n11391 ^ n6626 ^ 1'b0 ;
  assign n17352 = ~n2317 & n17351 ;
  assign n17353 = n496 & n15353 ;
  assign n17354 = n3225 & ~n11084 ;
  assign n17355 = n17354 ^ n1497 ^ 1'b0 ;
  assign n17356 = n17353 & n17355 ;
  assign n17357 = ( ~n4305 & n6764 ) | ( ~n4305 & n12784 ) | ( n6764 & n12784 ) ;
  assign n17358 = ~n325 & n12129 ;
  assign n17359 = n9050 | n15042 ;
  assign n17360 = n9276 & ~n10489 ;
  assign n17361 = n16668 & n17360 ;
  assign n17362 = n12072 | n17361 ;
  assign n17363 = ( n8237 & n10124 ) | ( n8237 & ~n10178 ) | ( n10124 & ~n10178 ) ;
  assign n17364 = n17363 ^ n1536 ^ 1'b0 ;
  assign n17365 = n3722 ^ n2769 ^ 1'b0 ;
  assign n17366 = n17365 ^ n4421 ^ 1'b0 ;
  assign n17367 = n4935 & n17366 ;
  assign n17368 = n17367 ^ n436 ^ x184 ;
  assign n17369 = n14636 | n16434 ;
  assign n17370 = ~n1503 & n2824 ;
  assign n17371 = n4567 | n9845 ;
  assign n17372 = n17371 ^ n16703 ^ 1'b0 ;
  assign n17373 = n12140 ^ n1899 ^ 1'b0 ;
  assign n17374 = n3348 & n13384 ;
  assign n17375 = n17374 ^ n5027 ^ 1'b0 ;
  assign n17376 = n17375 ^ n7841 ^ 1'b0 ;
  assign n17377 = n878 & n9681 ;
  assign n17378 = ~n1487 & n6765 ;
  assign n17379 = n17378 ^ n2836 ^ 1'b0 ;
  assign n17380 = n10652 ^ n5947 ^ 1'b0 ;
  assign n17381 = n17379 & n17380 ;
  assign n17382 = n5838 & n17381 ;
  assign n17383 = n6111 & n17382 ;
  assign n17384 = n4928 & ~n17383 ;
  assign n17385 = n1558 & n17384 ;
  assign n17386 = n5969 & n17385 ;
  assign n17387 = n17345 ^ n12842 ^ n5437 ;
  assign n17388 = ~n9784 & n17387 ;
  assign n17389 = ( n1515 & n11579 ) | ( n1515 & n17388 ) | ( n11579 & n17388 ) ;
  assign n17390 = ~n5230 & n6672 ;
  assign n17391 = ( n13725 & ~n13736 ) | ( n13725 & n17390 ) | ( ~n13736 & n17390 ) ;
  assign n17392 = ~n1682 & n16194 ;
  assign n17393 = n5518 ^ n3328 ^ 1'b0 ;
  assign n17394 = n1197 & n17393 ;
  assign n17395 = n16973 ^ n2985 ^ 1'b0 ;
  assign n17396 = n17394 & n17395 ;
  assign n17398 = n1636 | n1740 ;
  assign n17397 = n4345 | n11371 ;
  assign n17399 = n17398 ^ n17397 ^ 1'b0 ;
  assign n17400 = n1902 & ~n2066 ;
  assign n17401 = n12105 & n17400 ;
  assign n17402 = n12423 ^ n341 ^ 1'b0 ;
  assign n17403 = ~n4567 & n17402 ;
  assign n17404 = n4611 & n17403 ;
  assign n17405 = n277 & n17404 ;
  assign n17406 = n13731 | n17405 ;
  assign n17407 = n17406 ^ n7643 ^ 1'b0 ;
  assign n17408 = n17407 ^ n16862 ^ 1'b0 ;
  assign n17409 = n17401 | n17408 ;
  assign n17412 = ~n4126 & n8737 ;
  assign n17410 = n1970 & ~n8157 ;
  assign n17411 = n17410 ^ n9729 ^ 1'b0 ;
  assign n17413 = n17412 ^ n17411 ^ n13956 ;
  assign n17414 = n4013 ^ n3122 ^ 1'b0 ;
  assign n17415 = ( ~x111 & n5135 ) | ( ~x111 & n17414 ) | ( n5135 & n17414 ) ;
  assign n17416 = ~n2790 & n17415 ;
  assign n17417 = n4067 | n17416 ;
  assign n17418 = n17417 ^ n5085 ^ 1'b0 ;
  assign n17419 = x154 & ~n259 ;
  assign n17420 = n17419 ^ n1995 ^ 1'b0 ;
  assign n17421 = n2907 & ~n13943 ;
  assign n17422 = n17421 ^ n3521 ^ 1'b0 ;
  assign n17423 = n15933 ^ x38 ^ 1'b0 ;
  assign n17424 = n11207 | n17423 ;
  assign n17425 = n4456 ^ n4085 ^ 1'b0 ;
  assign n17426 = n2645 | n7326 ;
  assign n17432 = ~n305 & n725 ;
  assign n17433 = ~x58 & n17432 ;
  assign n17428 = n3165 ^ n1935 ^ x78 ;
  assign n17429 = n17428 ^ n6663 ^ 1'b0 ;
  assign n17430 = ~n8013 & n17429 ;
  assign n17431 = ~n1659 & n17430 ;
  assign n17427 = n5050 ^ n3571 ^ n2149 ;
  assign n17434 = n17433 ^ n17431 ^ n17427 ;
  assign n17435 = n12878 | n17434 ;
  assign n17436 = n17426 & ~n17435 ;
  assign n17437 = ~n341 & n9069 ;
  assign n17438 = ~n8916 & n17437 ;
  assign n17439 = ( n5777 & ~n6329 ) | ( n5777 & n16907 ) | ( ~n6329 & n16907 ) ;
  assign n17440 = ~n2473 & n17439 ;
  assign n17441 = n15239 ^ n11299 ^ n6488 ;
  assign n17442 = n17185 ^ n516 ^ 1'b0 ;
  assign n17443 = n13336 & n17442 ;
  assign n17444 = n4411 & n17443 ;
  assign n17445 = n17444 ^ n9271 ^ 1'b0 ;
  assign n17446 = n12367 ^ n10344 ^ 1'b0 ;
  assign n17447 = ~n17445 & n17446 ;
  assign n17448 = n17441 & ~n17447 ;
  assign n17449 = n5475 & n11062 ;
  assign n17450 = n17449 ^ n14334 ^ 1'b0 ;
  assign n17451 = n11373 | n12875 ;
  assign n17452 = n17451 ^ n10463 ^ 1'b0 ;
  assign n17453 = n17452 ^ n15712 ^ 1'b0 ;
  assign n17454 = n17450 | n17453 ;
  assign n17456 = n1493 | n8447 ;
  assign n17455 = n4020 & ~n4239 ;
  assign n17457 = n17456 ^ n17455 ^ n6073 ;
  assign n17458 = ( n9044 & n11192 ) | ( n9044 & ~n13647 ) | ( n11192 & ~n13647 ) ;
  assign n17459 = n6393 ^ n591 ^ 1'b0 ;
  assign n17460 = n17458 & ~n17459 ;
  assign n17461 = n12133 ^ n9089 ^ 1'b0 ;
  assign n17462 = ~n2616 & n17461 ;
  assign n17463 = n9997 ^ n1659 ^ 1'b0 ;
  assign n17464 = n17463 ^ n4553 ^ n2412 ;
  assign n17465 = ~n6047 & n6080 ;
  assign n17466 = ~n7145 & n17465 ;
  assign n17467 = n1572 | n17466 ;
  assign n17468 = n7325 | n17467 ;
  assign n17469 = ( n5964 & n11128 ) | ( n5964 & ~n17468 ) | ( n11128 & ~n17468 ) ;
  assign n17470 = n13285 & n15656 ;
  assign n17471 = ~n4105 & n4592 ;
  assign n17472 = n8453 | n17471 ;
  assign n17473 = n17472 ^ n12091 ^ 1'b0 ;
  assign n17474 = n9522 & n12828 ;
  assign n17475 = n17474 ^ n12799 ^ 1'b0 ;
  assign n17476 = ~n3269 & n10285 ;
  assign n17477 = ~n12748 & n17476 ;
  assign n17478 = ( n3595 & n13722 ) | ( n3595 & ~n16179 ) | ( n13722 & ~n16179 ) ;
  assign n17479 = n12174 & ~n17478 ;
  assign n17480 = n9952 ^ n1748 ^ 1'b0 ;
  assign n17481 = n4814 & n17480 ;
  assign n17482 = n17481 ^ n13079 ^ 1'b0 ;
  assign n17483 = n9687 & ~n17482 ;
  assign n17484 = ( ~n13189 & n15357 ) | ( ~n13189 & n17483 ) | ( n15357 & n17483 ) ;
  assign n17487 = n12593 ^ n7444 ^ 1'b0 ;
  assign n17485 = n401 | n7803 ;
  assign n17486 = n17485 ^ n11921 ^ 1'b0 ;
  assign n17488 = n17487 ^ n17486 ^ n16867 ;
  assign n17489 = ~n8071 & n12504 ;
  assign n17490 = n6738 ^ n1209 ^ n449 ;
  assign n17491 = n17490 ^ n6688 ^ n2313 ;
  assign n17492 = n17491 ^ n3157 ^ 1'b0 ;
  assign n17493 = n15656 & ~n17492 ;
  assign n17494 = ~n12826 & n17493 ;
  assign n17495 = n5969 & ~n12504 ;
  assign n17496 = ~n6915 & n17495 ;
  assign n17497 = n4623 | n17496 ;
  assign n17498 = ~n17494 & n17497 ;
  assign n17499 = n6675 & n11667 ;
  assign n17500 = n13751 ^ n12165 ^ 1'b0 ;
  assign n17501 = n11105 ^ n3982 ^ 1'b0 ;
  assign n17502 = ~n1272 & n17501 ;
  assign n17503 = ~n17500 & n17502 ;
  assign n17504 = ~n5981 & n7176 ;
  assign n17505 = ( ~n13420 & n13740 ) | ( ~n13420 & n17504 ) | ( n13740 & n17504 ) ;
  assign n17506 = n4361 ^ n3424 ^ 1'b0 ;
  assign n17507 = n1835 | n5393 ;
  assign n17508 = ( ~n9224 & n13668 ) | ( ~n9224 & n17507 ) | ( n13668 & n17507 ) ;
  assign n17509 = n7482 ^ n5557 ^ x173 ;
  assign n17510 = n6807 & n17509 ;
  assign n17511 = ~n476 & n17510 ;
  assign n17512 = n4906 | n5598 ;
  assign n17513 = n368 & ~n17512 ;
  assign n17514 = ( ~n7173 & n8018 ) | ( ~n7173 & n17513 ) | ( n8018 & n17513 ) ;
  assign n17515 = n17514 ^ n13227 ^ n471 ;
  assign n17516 = n7568 ^ n3071 ^ 1'b0 ;
  assign n17517 = ~n16005 & n17516 ;
  assign n17518 = ( n4447 & n9986 ) | ( n4447 & n17517 ) | ( n9986 & n17517 ) ;
  assign n17519 = ~n3108 & n3856 ;
  assign n17520 = n17519 ^ n15787 ^ n4254 ;
  assign n17521 = ( n6318 & n6446 ) | ( n6318 & n17520 ) | ( n6446 & n17520 ) ;
  assign n17522 = n5384 ^ n1394 ^ 1'b0 ;
  assign n17523 = n8168 | n17522 ;
  assign n17526 = ~n4902 & n9607 ;
  assign n17524 = n5339 ^ n5191 ^ 1'b0 ;
  assign n17525 = n17524 ^ n1567 ^ n1024 ;
  assign n17527 = n17526 ^ n17525 ^ 1'b0 ;
  assign n17528 = n718 & n17527 ;
  assign n17529 = ( n12585 & ~n17523 ) | ( n12585 & n17528 ) | ( ~n17523 & n17528 ) ;
  assign n17531 = ( ~n550 & n4155 ) | ( ~n550 & n4625 ) | ( n4155 & n4625 ) ;
  assign n17532 = n17531 ^ n3204 ^ n2365 ;
  assign n17530 = n9662 ^ n3324 ^ n656 ;
  assign n17533 = n17532 ^ n17530 ^ n7353 ;
  assign n17534 = n752 & ~n9025 ;
  assign n17535 = n17534 ^ n970 ^ 1'b0 ;
  assign n17536 = ( n3784 & n6736 ) | ( n3784 & ~n17535 ) | ( n6736 & ~n17535 ) ;
  assign n17537 = n17536 ^ n15922 ^ n8536 ;
  assign n17538 = n16774 & ~n17537 ;
  assign n17539 = ~n9939 & n17538 ;
  assign n17540 = n3347 & ~n5645 ;
  assign n17541 = n3139 & n17540 ;
  assign n17542 = n9485 ^ n6001 ^ x240 ;
  assign n17543 = x39 & ~n8466 ;
  assign n17544 = n17543 ^ n7621 ^ 1'b0 ;
  assign n17545 = n6048 | n17544 ;
  assign n17546 = ( ~n16362 & n17542 ) | ( ~n16362 & n17545 ) | ( n17542 & n17545 ) ;
  assign n17547 = ~n5933 & n17140 ;
  assign n17548 = n4857 | n16172 ;
  assign n17549 = n13911 & ~n17548 ;
  assign n17550 = ( n3261 & ~n7459 ) | ( n3261 & n17549 ) | ( ~n7459 & n17549 ) ;
  assign n17553 = n13551 ^ n8735 ^ n5709 ;
  assign n17551 = ( ~n639 & n2174 ) | ( ~n639 & n9598 ) | ( n2174 & n9598 ) ;
  assign n17552 = n17551 ^ n12353 ^ n3691 ;
  assign n17554 = n17553 ^ n17552 ^ n12540 ;
  assign n17555 = n15807 & n17554 ;
  assign n17556 = n2937 | n5056 ;
  assign n17557 = n13916 & n17556 ;
  assign n17558 = n4692 ^ n3264 ^ 1'b0 ;
  assign n17559 = n13987 ^ n4221 ^ 1'b0 ;
  assign n17560 = n4045 | n17559 ;
  assign n17561 = n727 & n15853 ;
  assign n17562 = n17230 ^ n15710 ^ n6805 ;
  assign n17564 = n7243 ^ n6114 ^ n2619 ;
  assign n17563 = n1835 | n11211 ;
  assign n17565 = n17564 ^ n17563 ^ 1'b0 ;
  assign n17566 = n17565 ^ n14691 ^ 1'b0 ;
  assign n17567 = n17566 ^ n10495 ^ 1'b0 ;
  assign n17568 = n3061 & n17567 ;
  assign n17569 = n2478 | n3172 ;
  assign n17570 = n17569 ^ n5914 ^ 1'b0 ;
  assign n17571 = n2806 ^ x89 ^ 1'b0 ;
  assign n17572 = ( n3798 & n10185 ) | ( n3798 & n17571 ) | ( n10185 & n17571 ) ;
  assign n17573 = n8608 & n17572 ;
  assign n17574 = n17573 ^ n3991 ^ 1'b0 ;
  assign n17575 = n17574 ^ n11458 ^ n4355 ;
  assign n17576 = n17575 ^ n5909 ^ 1'b0 ;
  assign n17578 = x185 & ~n2846 ;
  assign n17579 = n15642 ^ n7155 ^ 1'b0 ;
  assign n17580 = n1814 & ~n17579 ;
  assign n17581 = ~n17578 & n17580 ;
  assign n17577 = n8858 & ~n14929 ;
  assign n17582 = n17581 ^ n17577 ^ 1'b0 ;
  assign n17583 = n10002 & ~n17582 ;
  assign n17584 = n14635 & n14968 ;
  assign n17585 = ( n10495 & n12914 ) | ( n10495 & n17584 ) | ( n12914 & n17584 ) ;
  assign n17586 = n2038 | n5204 ;
  assign n17587 = n17586 ^ n2943 ^ 1'b0 ;
  assign n17588 = n2746 & ~n17256 ;
  assign n17589 = n17587 & n17588 ;
  assign n17590 = n1196 & ~n5988 ;
  assign n17591 = n17589 & n17590 ;
  assign n17592 = n12709 ^ n6513 ^ n737 ;
  assign n17593 = n17592 ^ n3146 ^ 1'b0 ;
  assign n17594 = n11258 & ~n13418 ;
  assign n17596 = n8717 ^ n3585 ^ 1'b0 ;
  assign n17595 = ~n1582 & n17159 ;
  assign n17597 = n17596 ^ n17595 ^ 1'b0 ;
  assign n17598 = ( n2401 & n6626 ) | ( n2401 & ~n7730 ) | ( n6626 & ~n7730 ) ;
  assign n17599 = n16687 & n17598 ;
  assign n17600 = ~n4592 & n17599 ;
  assign n17601 = ~n2865 & n4150 ;
  assign n17602 = n17601 ^ n2496 ^ 1'b0 ;
  assign n17603 = n17602 ^ n12026 ^ 1'b0 ;
  assign n17604 = ( n12594 & n17514 ) | ( n12594 & n17603 ) | ( n17514 & n17603 ) ;
  assign n17605 = n2425 ^ n1120 ^ 1'b0 ;
  assign n17606 = n17605 ^ n1603 ^ 1'b0 ;
  assign n17607 = n8250 ^ n1788 ^ 1'b0 ;
  assign n17608 = ( n1158 & n1880 ) | ( n1158 & n17607 ) | ( n1880 & n17607 ) ;
  assign n17609 = n8018 ^ n6982 ^ n5328 ;
  assign n17610 = n17609 ^ n13821 ^ 1'b0 ;
  assign n17611 = n11140 & ~n17610 ;
  assign n17612 = n8591 & n17611 ;
  assign n17613 = n17612 ^ n15722 ^ 1'b0 ;
  assign n17614 = n12613 ^ n4444 ^ 1'b0 ;
  assign n17615 = n10798 ^ n7250 ^ n5386 ;
  assign n17616 = n15022 & n17615 ;
  assign n17617 = n3956 ^ n915 ^ 1'b0 ;
  assign n17618 = n9741 | n17617 ;
  assign n17619 = n5121 ^ n2106 ^ n1094 ;
  assign n17620 = ~n1024 & n10321 ;
  assign n17621 = ( n14787 & ~n17619 ) | ( n14787 & n17620 ) | ( ~n17619 & n17620 ) ;
  assign n17622 = n8970 & ~n17621 ;
  assign n17623 = n2107 & n17622 ;
  assign n17624 = n5057 ^ n4496 ^ 1'b0 ;
  assign n17625 = n4212 & ~n8670 ;
  assign n17626 = n17624 & ~n17625 ;
  assign n17627 = n5945 & ~n17626 ;
  assign n17628 = n9144 ^ n8902 ^ 1'b0 ;
  assign n17629 = x12 | n3640 ;
  assign n17630 = n17629 ^ n15013 ^ 1'b0 ;
  assign n17631 = n2821 & ~n10298 ;
  assign n17632 = n17631 ^ n16193 ^ n10395 ;
  assign n17633 = ~n3449 & n4896 ;
  assign n17634 = n4825 & n8477 ;
  assign n17635 = n17634 ^ n7916 ^ 1'b0 ;
  assign n17636 = x189 & ~n17635 ;
  assign n17637 = n8799 & ~n13314 ;
  assign n17638 = ~n17636 & n17637 ;
  assign n17639 = n5426 ^ n759 ^ 1'b0 ;
  assign n17640 = ( n11612 & n13797 ) | ( n11612 & ~n17639 ) | ( n13797 & ~n17639 ) ;
  assign n17641 = n16029 & ~n17640 ;
  assign n17642 = n17641 ^ n5761 ^ 1'b0 ;
  assign n17643 = ( n4282 & n9386 ) | ( n4282 & ~n14570 ) | ( n9386 & ~n14570 ) ;
  assign n17644 = n3632 & ~n15610 ;
  assign n17645 = n17644 ^ n9591 ^ 1'b0 ;
  assign n17646 = n12340 ^ n3624 ^ n898 ;
  assign n17648 = n4381 & ~n5398 ;
  assign n17649 = n6491 & n17648 ;
  assign n17650 = n2196 | n17649 ;
  assign n17651 = n5054 & ~n17650 ;
  assign n17652 = n10180 & ~n17651 ;
  assign n17653 = n8415 ^ n5189 ^ n2917 ;
  assign n17654 = ~n17652 & n17653 ;
  assign n17647 = n12394 ^ n11000 ^ 1'b0 ;
  assign n17655 = n17654 ^ n17647 ^ n12138 ;
  assign n17656 = n9824 ^ n1532 ^ 1'b0 ;
  assign n17657 = n1713 & n17656 ;
  assign n17658 = n17655 & n17657 ;
  assign n17659 = n10042 | n10529 ;
  assign n17660 = n17659 ^ n5488 ^ 1'b0 ;
  assign n17661 = n13278 ^ n5839 ^ n4447 ;
  assign n17662 = ( ~n1534 & n1994 ) | ( ~n1534 & n17661 ) | ( n1994 & n17661 ) ;
  assign n17663 = n1933 & n17662 ;
  assign n17664 = n17660 & ~n17663 ;
  assign n17665 = n8043 & ~n17664 ;
  assign n17666 = n15403 ^ n14613 ^ 1'b0 ;
  assign n17669 = n4879 ^ n2199 ^ 1'b0 ;
  assign n17667 = x110 | n1440 ;
  assign n17668 = ( n4767 & n11976 ) | ( n4767 & n17667 ) | ( n11976 & n17667 ) ;
  assign n17670 = n17669 ^ n17668 ^ n2118 ;
  assign n17674 = n8631 ^ x185 ^ 1'b0 ;
  assign n17675 = n3905 & ~n9217 ;
  assign n17676 = n17674 & n17675 ;
  assign n17671 = n8171 ^ n5870 ^ 1'b0 ;
  assign n17672 = n9292 & n17671 ;
  assign n17673 = ( n2348 & n16105 ) | ( n2348 & ~n17672 ) | ( n16105 & ~n17672 ) ;
  assign n17677 = n17676 ^ n17673 ^ 1'b0 ;
  assign n17678 = n16538 & n17677 ;
  assign n17679 = n13352 ^ n7273 ^ 1'b0 ;
  assign n17680 = n11258 & n17679 ;
  assign n17681 = n17680 ^ n15311 ^ x147 ;
  assign n17682 = n2663 | n5878 ;
  assign n17683 = n14442 ^ n13637 ^ 1'b0 ;
  assign n17684 = x23 & ~n2766 ;
  assign n17685 = ~n2469 & n17684 ;
  assign n17686 = n17685 ^ n2588 ^ 1'b0 ;
  assign n17687 = ~n17683 & n17686 ;
  assign n17688 = n15046 & n17687 ;
  assign n17689 = n16755 & n17688 ;
  assign n17690 = n12916 ^ n6182 ^ 1'b0 ;
  assign n17693 = n8609 ^ n4609 ^ 1'b0 ;
  assign n17694 = n968 & n17693 ;
  assign n17691 = ~n522 & n4271 ;
  assign n17692 = n2959 & ~n17691 ;
  assign n17695 = n17694 ^ n17692 ^ 1'b0 ;
  assign n17696 = n9282 | n12664 ;
  assign n17697 = n17696 ^ n8079 ^ 1'b0 ;
  assign n17698 = n6306 ^ x110 ^ 1'b0 ;
  assign n17699 = n16342 & ~n17698 ;
  assign n17700 = ~n7440 & n17699 ;
  assign n17705 = n5063 ^ n2240 ^ n1765 ;
  assign n17706 = n4141 & ~n17705 ;
  assign n17701 = n16624 ^ n3015 ^ 1'b0 ;
  assign n17702 = n1413 & ~n17701 ;
  assign n17703 = n10117 ^ n10108 ^ n4870 ;
  assign n17704 = n17702 & n17703 ;
  assign n17707 = n17706 ^ n17704 ^ 1'b0 ;
  assign n17708 = n12253 ^ n11845 ^ n1559 ;
  assign n17709 = n13452 ^ n8398 ^ 1'b0 ;
  assign n17710 = n17709 ^ n6036 ^ 1'b0 ;
  assign n17711 = n17710 ^ n7995 ^ 1'b0 ;
  assign n17712 = n264 | n13556 ;
  assign n17713 = n17712 ^ n5513 ^ 1'b0 ;
  assign n17717 = ~n4060 & n5821 ;
  assign n17718 = n8748 & n17717 ;
  assign n17714 = n10117 | n14142 ;
  assign n17715 = ~n9539 & n17714 ;
  assign n17716 = ( n1124 & n5739 ) | ( n1124 & ~n17715 ) | ( n5739 & ~n17715 ) ;
  assign n17719 = n17718 ^ n17716 ^ 1'b0 ;
  assign n17720 = n5919 & ~n17719 ;
  assign n17721 = n17720 ^ n14888 ^ n5553 ;
  assign n17722 = n14003 & ~n17721 ;
  assign n17723 = n17713 & n17722 ;
  assign n17724 = n747 | n12469 ;
  assign n17725 = ~n1482 & n17724 ;
  assign n17726 = ~n7386 & n17725 ;
  assign n17727 = ~n1576 & n13433 ;
  assign n17728 = n8486 & ~n17727 ;
  assign n17729 = ( n3052 & n7581 ) | ( n3052 & ~n17728 ) | ( n7581 & ~n17728 ) ;
  assign n17730 = n3764 ^ n1906 ^ 1'b0 ;
  assign n17731 = ~n3324 & n17730 ;
  assign n17732 = ( n369 & n913 ) | ( n369 & ~n4533 ) | ( n913 & ~n4533 ) ;
  assign n17733 = n10388 ^ n8077 ^ 1'b0 ;
  assign n17734 = ~n17732 & n17733 ;
  assign n17735 = ~n17731 & n17734 ;
  assign n17736 = n5437 ^ n3091 ^ n2808 ;
  assign n17737 = ~n8494 & n17736 ;
  assign n17738 = ( n2504 & n2885 ) | ( n2504 & n17737 ) | ( n2885 & n17737 ) ;
  assign n17739 = ( n2049 & n10844 ) | ( n2049 & n17738 ) | ( n10844 & n17738 ) ;
  assign n17740 = n14866 ^ n14110 ^ 1'b0 ;
  assign n17741 = n2554 & n7218 ;
  assign n17742 = n17741 ^ n8839 ^ 1'b0 ;
  assign n17743 = n2908 & n17742 ;
  assign n17744 = ~n16294 & n17743 ;
  assign n17745 = n14016 ^ n3595 ^ 1'b0 ;
  assign n17746 = n1576 | n17745 ;
  assign n17747 = n11737 & ~n17746 ;
  assign n17748 = ~n4498 & n17747 ;
  assign n17749 = n1525 | n6020 ;
  assign n17750 = n17749 ^ n17309 ^ 1'b0 ;
  assign n17752 = n649 | n6567 ;
  assign n17753 = n17752 ^ n981 ^ 1'b0 ;
  assign n17751 = ~n10721 & n12787 ;
  assign n17754 = n17753 ^ n17751 ^ n8622 ;
  assign n17755 = n12360 ^ n9067 ^ n3034 ;
  assign n17756 = ( ~n5475 & n13407 ) | ( ~n5475 & n16334 ) | ( n13407 & n16334 ) ;
  assign n17757 = n7513 ^ n3422 ^ 1'b0 ;
  assign n17758 = ~n1096 & n17757 ;
  assign n17759 = n350 & n659 ;
  assign n17760 = n17759 ^ n3802 ^ 1'b0 ;
  assign n17761 = ( n4904 & n17758 ) | ( n4904 & ~n17760 ) | ( n17758 & ~n17760 ) ;
  assign n17762 = n17118 ^ n14035 ^ 1'b0 ;
  assign n17763 = n1880 | n17762 ;
  assign n17764 = n17761 & ~n17763 ;
  assign n17765 = n1041 | n6189 ;
  assign n17766 = n17765 ^ n4388 ^ 1'b0 ;
  assign n17767 = n17766 ^ n10192 ^ 1'b0 ;
  assign n17768 = n7970 & n13026 ;
  assign n17769 = n2563 & n17768 ;
  assign n17770 = n17769 ^ n10994 ^ 1'b0 ;
  assign n17771 = n13098 ^ n1470 ^ 1'b0 ;
  assign n17772 = ~n4600 & n5362 ;
  assign n17773 = n14003 ^ n12193 ^ n4300 ;
  assign n17774 = ( n17771 & n17772 ) | ( n17771 & n17773 ) | ( n17772 & n17773 ) ;
  assign n17775 = ~n13740 & n17774 ;
  assign n17776 = n17770 & n17775 ;
  assign n17777 = n17767 | n17776 ;
  assign n17778 = n17777 ^ n1149 ^ 1'b0 ;
  assign n17779 = n4679 & ~n14403 ;
  assign n17780 = ~n3953 & n17779 ;
  assign n17781 = n3681 & ~n8012 ;
  assign n17782 = ( n3056 & n11173 ) | ( n3056 & ~n16190 ) | ( n11173 & ~n16190 ) ;
  assign n17783 = n593 & ~n17782 ;
  assign n17784 = ~n17781 & n17783 ;
  assign n17785 = n1154 & ~n17784 ;
  assign n17786 = n17780 & n17785 ;
  assign n17787 = n8043 ^ n7978 ^ n3291 ;
  assign n17788 = ~n5854 & n17787 ;
  assign n17789 = n17788 ^ n9326 ^ 1'b0 ;
  assign n17790 = n2349 | n17789 ;
  assign n17791 = n13494 & ~n17790 ;
  assign n17792 = n8219 & ~n17791 ;
  assign n17793 = n8565 ^ x225 ^ 1'b0 ;
  assign n17794 = n600 & ~n17793 ;
  assign n17795 = ( n4849 & n5179 ) | ( n4849 & ~n17794 ) | ( n5179 & ~n17794 ) ;
  assign n17796 = n17795 ^ n1515 ^ 1'b0 ;
  assign n17797 = n17796 ^ n5370 ^ 1'b0 ;
  assign n17798 = ~n7184 & n17276 ;
  assign n17799 = n15404 ^ n12260 ^ n3977 ;
  assign n17800 = n7562 ^ n2856 ^ 1'b0 ;
  assign n17801 = n17799 & n17800 ;
  assign n17802 = n279 & n4823 ;
  assign n17803 = ~n15426 & n17802 ;
  assign n17809 = n5328 & ~n11597 ;
  assign n17810 = n17809 ^ n9187 ^ 1'b0 ;
  assign n17807 = n2966 & ~n11407 ;
  assign n17808 = n17807 ^ n10421 ^ 1'b0 ;
  assign n17804 = n10848 ^ n1453 ^ 1'b0 ;
  assign n17805 = n2050 | n17804 ;
  assign n17806 = ~n1927 & n17805 ;
  assign n17811 = n17810 ^ n17808 ^ n17806 ;
  assign n17812 = ( n4628 & ~n14621 ) | ( n4628 & n17811 ) | ( ~n14621 & n17811 ) ;
  assign n17813 = n5975 & n15881 ;
  assign n17814 = n17813 ^ n3862 ^ 1'b0 ;
  assign n17817 = n11626 ^ n4561 ^ n3310 ;
  assign n17815 = n2150 & ~n2423 ;
  assign n17816 = n17815 ^ n6487 ^ 1'b0 ;
  assign n17818 = n17817 ^ n17816 ^ 1'b0 ;
  assign n17819 = n17814 & n17818 ;
  assign n17820 = ~n3625 & n10195 ;
  assign n17822 = n13725 ^ n1442 ^ 1'b0 ;
  assign n17821 = ( n8327 & n10094 ) | ( n8327 & ~n11592 ) | ( n10094 & ~n11592 ) ;
  assign n17823 = n17822 ^ n17821 ^ 1'b0 ;
  assign n17824 = n17823 ^ n14850 ^ 1'b0 ;
  assign n17825 = n5060 | n5296 ;
  assign n17826 = n17825 ^ n7731 ^ 1'b0 ;
  assign n17827 = n17826 ^ n10672 ^ n10659 ;
  assign n17828 = n10704 ^ n6905 ^ n1031 ;
  assign n17829 = n2927 & ~n10345 ;
  assign n17830 = ~n10449 & n17829 ;
  assign n17831 = n10092 & ~n12701 ;
  assign n17832 = n7411 ^ n6971 ^ n6847 ;
  assign n17833 = n17832 ^ n9228 ^ n5809 ;
  assign n17834 = n6073 ^ n835 ^ 1'b0 ;
  assign n17835 = ~n17833 & n17834 ;
  assign n17836 = ( n4840 & n4981 ) | ( n4840 & ~n10638 ) | ( n4981 & ~n10638 ) ;
  assign n17837 = n10579 ^ n2661 ^ 1'b0 ;
  assign n17838 = ( ~n14297 & n15610 ) | ( ~n14297 & n17837 ) | ( n15610 & n17837 ) ;
  assign n17839 = n2200 & ~n2846 ;
  assign n17840 = n2948 | n9831 ;
  assign n17841 = ( n4699 & n6612 ) | ( n4699 & n12035 ) | ( n6612 & n12035 ) ;
  assign n17842 = ( n6390 & ~n8066 ) | ( n6390 & n17841 ) | ( ~n8066 & n17841 ) ;
  assign n17843 = n13456 ^ n2225 ^ 1'b0 ;
  assign n17844 = ( n2019 & n8171 ) | ( n2019 & ~n17843 ) | ( n8171 & ~n17843 ) ;
  assign n17845 = ( ~n8021 & n9947 ) | ( ~n8021 & n14906 ) | ( n9947 & n14906 ) ;
  assign n17847 = n7586 ^ n4490 ^ 1'b0 ;
  assign n17846 = n6660 & n10401 ;
  assign n17848 = n17847 ^ n17846 ^ 1'b0 ;
  assign n17849 = n434 | n6406 ;
  assign n17855 = ( ~n339 & n1916 ) | ( ~n339 & n13427 ) | ( n1916 & n13427 ) ;
  assign n17850 = n922 & n2734 ;
  assign n17851 = n17850 ^ n3592 ^ 1'b0 ;
  assign n17852 = n5615 & ~n17851 ;
  assign n17853 = n17852 ^ n11823 ^ 1'b0 ;
  assign n17854 = ~n9699 & n17853 ;
  assign n17856 = n17855 ^ n17854 ^ 1'b0 ;
  assign n17857 = ( n8127 & ~n13735 ) | ( n8127 & n17856 ) | ( ~n13735 & n17856 ) ;
  assign n17858 = ( ~n2275 & n3762 ) | ( ~n2275 & n17574 ) | ( n3762 & n17574 ) ;
  assign n17859 = n17749 ^ n16002 ^ 1'b0 ;
  assign n17860 = n17858 & n17859 ;
  assign n17861 = n9117 ^ n371 ^ 1'b0 ;
  assign n17862 = n17860 & ~n17861 ;
  assign n17863 = ( x94 & n10606 ) | ( x94 & ~n17784 ) | ( n10606 & ~n17784 ) ;
  assign n17864 = n17863 ^ n15255 ^ 1'b0 ;
  assign n17865 = n17862 & n17864 ;
  assign n17866 = ~n1702 & n2448 ;
  assign n17867 = ~n13781 & n15430 ;
  assign n17868 = n17866 & n17867 ;
  assign n17869 = n13878 ^ n3939 ^ 1'b0 ;
  assign n17870 = ~n11200 & n17869 ;
  assign n17871 = n17870 ^ n9411 ^ n5653 ;
  assign n17872 = n17871 ^ n10145 ^ n7589 ;
  assign n17873 = n16177 ^ n7970 ^ 1'b0 ;
  assign n17874 = n12813 & ~n17873 ;
  assign n17875 = ( n1200 & ~n10330 ) | ( n1200 & n17874 ) | ( ~n10330 & n17874 ) ;
  assign n17876 = n6213 & n11620 ;
  assign n17877 = n17876 ^ n3541 ^ 1'b0 ;
  assign n17878 = n6594 & n17877 ;
  assign n17883 = n614 & ~n3073 ;
  assign n17879 = n11449 ^ n2151 ^ 1'b0 ;
  assign n17880 = ~n4185 & n17879 ;
  assign n17881 = n17880 ^ n13866 ^ n5551 ;
  assign n17882 = n14774 | n17881 ;
  assign n17884 = n17883 ^ n17882 ^ 1'b0 ;
  assign n17885 = n9173 & n15971 ;
  assign n17886 = n14894 ^ n4041 ^ 1'b0 ;
  assign n17887 = n3339 & ~n17886 ;
  assign n17888 = ( n14648 & ~n16499 ) | ( n14648 & n17887 ) | ( ~n16499 & n17887 ) ;
  assign n17889 = n17888 ^ n10481 ^ n10465 ;
  assign n17890 = n12511 ^ n12282 ^ 1'b0 ;
  assign n17895 = n3070 | n3459 ;
  assign n17896 = n17895 ^ n3190 ^ 1'b0 ;
  assign n17899 = x240 & n312 ;
  assign n17898 = n9802 ^ n7110 ^ 1'b0 ;
  assign n17900 = n17899 ^ n17898 ^ n2019 ;
  assign n17897 = ~n4495 & n6085 ;
  assign n17901 = n17900 ^ n17897 ^ 1'b0 ;
  assign n17902 = ( n8810 & n17896 ) | ( n8810 & ~n17901 ) | ( n17896 & ~n17901 ) ;
  assign n17903 = ( n347 & ~n3540 ) | ( n347 & n17902 ) | ( ~n3540 & n17902 ) ;
  assign n17891 = n3578 & ~n3919 ;
  assign n17892 = n396 & n17891 ;
  assign n17893 = ( ~n7457 & n12296 ) | ( ~n7457 & n17892 ) | ( n12296 & n17892 ) ;
  assign n17894 = n17893 ^ n1032 ^ 1'b0 ;
  assign n17904 = n17903 ^ n17894 ^ n8639 ;
  assign n17908 = n12933 ^ n2568 ^ 1'b0 ;
  assign n17909 = n595 & n17908 ;
  assign n17905 = ~n848 & n1179 ;
  assign n17906 = n464 & n17905 ;
  assign n17907 = n2394 & ~n17906 ;
  assign n17910 = n17909 ^ n17907 ^ 1'b0 ;
  assign n17911 = n3957 ^ n263 ^ 1'b0 ;
  assign n17912 = n3555 & ~n17911 ;
  assign n17913 = n2904 & n17912 ;
  assign n17914 = n17913 ^ n1906 ^ 1'b0 ;
  assign n17915 = ~n13226 & n17914 ;
  assign n17916 = n17915 ^ n14907 ^ 1'b0 ;
  assign n17917 = ( ~n1061 & n14020 ) | ( ~n1061 & n17916 ) | ( n14020 & n17916 ) ;
  assign n17918 = n2325 & ~n4984 ;
  assign n17919 = n15060 & ~n17918 ;
  assign n17920 = n17919 ^ n3430 ^ 1'b0 ;
  assign n17921 = n16911 ^ n2565 ^ n926 ;
  assign n17922 = n4416 & ~n17921 ;
  assign n17923 = ( n4128 & n17920 ) | ( n4128 & ~n17922 ) | ( n17920 & ~n17922 ) ;
  assign n17924 = n5181 & n17923 ;
  assign n17925 = n13550 ^ n7417 ^ n4734 ;
  assign n17927 = n3285 & n8508 ;
  assign n17926 = ~n7040 & n15590 ;
  assign n17928 = n17927 ^ n17926 ^ 1'b0 ;
  assign n17929 = ~n10919 & n17928 ;
  assign n17930 = ( n277 & n3053 ) | ( n277 & ~n8428 ) | ( n3053 & ~n8428 ) ;
  assign n17931 = n9622 ^ n625 ^ 1'b0 ;
  assign n17932 = n17931 ^ n4960 ^ n4516 ;
  assign n17933 = n17932 ^ n12385 ^ 1'b0 ;
  assign n17934 = ~n4355 & n17933 ;
  assign n17935 = ( n14796 & ~n17930 ) | ( n14796 & n17934 ) | ( ~n17930 & n17934 ) ;
  assign n17936 = n17935 ^ n1335 ^ 1'b0 ;
  assign n17937 = n7163 | n11180 ;
  assign n17938 = n11283 | n17937 ;
  assign n17939 = n8997 | n11588 ;
  assign n17940 = n17939 ^ n12241 ^ 1'b0 ;
  assign n17941 = n17940 ^ n14934 ^ 1'b0 ;
  assign n17942 = n10891 | n14360 ;
  assign n17945 = n15720 ^ n3207 ^ 1'b0 ;
  assign n17946 = n423 & n17945 ;
  assign n17947 = n14470 ^ n2819 ^ 1'b0 ;
  assign n17948 = n17946 & n17947 ;
  assign n17943 = n14273 | n15838 ;
  assign n17944 = x209 | n17943 ;
  assign n17949 = n17948 ^ n17944 ^ n15599 ;
  assign n17950 = ~n5389 & n8171 ;
  assign n17951 = n17950 ^ n5290 ^ 1'b0 ;
  assign n17952 = ~n2727 & n11974 ;
  assign n17953 = ( n7712 & ~n10021 ) | ( n7712 & n17952 ) | ( ~n10021 & n17952 ) ;
  assign n17954 = n17953 ^ n2043 ^ 1'b0 ;
  assign n17955 = n887 & n17954 ;
  assign n17959 = ( n2223 & ~n4050 ) | ( n2223 & n11598 ) | ( ~n4050 & n11598 ) ;
  assign n17957 = n1266 & n7674 ;
  assign n17958 = ~n6569 & n17957 ;
  assign n17960 = n17959 ^ n17958 ^ 1'b0 ;
  assign n17956 = n4662 | n6038 ;
  assign n17961 = n17960 ^ n17956 ^ 1'b0 ;
  assign n17962 = n17961 ^ n3640 ^ 1'b0 ;
  assign n17963 = n3339 & ~n17962 ;
  assign n17964 = n7923 ^ n1160 ^ 1'b0 ;
  assign n17967 = ( n1110 & ~n10780 ) | ( n1110 & n16096 ) | ( ~n10780 & n16096 ) ;
  assign n17965 = n8217 | n15621 ;
  assign n17966 = n3960 & ~n17965 ;
  assign n17968 = n17967 ^ n17966 ^ 1'b0 ;
  assign n17969 = n2106 & ~n5094 ;
  assign n17970 = n17969 ^ n935 ^ 1'b0 ;
  assign n17971 = n14577 & ~n17970 ;
  assign n17972 = n5877 & ~n6118 ;
  assign n17973 = n17972 ^ n9712 ^ 1'b0 ;
  assign n17974 = n17973 ^ n14708 ^ 1'b0 ;
  assign n17975 = n17974 ^ n16358 ^ 1'b0 ;
  assign n17976 = n17971 & ~n17975 ;
  assign n17977 = n1413 & ~n6971 ;
  assign n17978 = n17977 ^ n2645 ^ 1'b0 ;
  assign n17979 = n17921 ^ n14754 ^ 1'b0 ;
  assign n17980 = n13030 ^ n5470 ^ 1'b0 ;
  assign n17981 = ~n11000 & n17980 ;
  assign n17982 = n17981 ^ n2176 ^ 1'b0 ;
  assign n17983 = n17979 & ~n17982 ;
  assign n17984 = ( n9761 & ~n15069 ) | ( n9761 & n17983 ) | ( ~n15069 & n17983 ) ;
  assign n17985 = n7634 ^ n7411 ^ n6609 ;
  assign n17989 = n5133 ^ n3552 ^ 1'b0 ;
  assign n17990 = ~n6545 & n17989 ;
  assign n17986 = ( n9364 & ~n11939 ) | ( n9364 & n17763 ) | ( ~n11939 & n17763 ) ;
  assign n17987 = x66 & n10780 ;
  assign n17988 = n17986 | n17987 ;
  assign n17991 = n17990 ^ n17988 ^ n8177 ;
  assign n17992 = n1852 | n2459 ;
  assign n17993 = n17992 ^ n5277 ^ 1'b0 ;
  assign n17994 = ( n4767 & ~n12589 ) | ( n4767 & n17993 ) | ( ~n12589 & n17993 ) ;
  assign n17995 = n6961 ^ n2778 ^ 1'b0 ;
  assign n17996 = n9919 | n17995 ;
  assign n17997 = n17994 & ~n17996 ;
  assign n18005 = n12804 ^ n4274 ^ 1'b0 ;
  assign n18001 = n5385 ^ n3252 ^ 1'b0 ;
  assign n17998 = n10212 ^ n2399 ^ 1'b0 ;
  assign n17999 = ~n7062 & n17998 ;
  assign n18000 = ~n1182 & n17999 ;
  assign n18002 = n18001 ^ n18000 ^ 1'b0 ;
  assign n18003 = n5608 & n18002 ;
  assign n18004 = n7576 & n18003 ;
  assign n18006 = n18005 ^ n18004 ^ n6472 ;
  assign n18007 = n18006 ^ n13483 ^ 1'b0 ;
  assign n18008 = n7058 | n8632 ;
  assign n18009 = n6596 ^ x34 ^ 1'b0 ;
  assign n18010 = ( n2348 & n18008 ) | ( n2348 & n18009 ) | ( n18008 & n18009 ) ;
  assign n18011 = ( n5106 & ~n5341 ) | ( n5106 & n14578 ) | ( ~n5341 & n14578 ) ;
  assign n18012 = ~n7271 & n18011 ;
  assign n18013 = n8882 ^ n3191 ^ 1'b0 ;
  assign n18014 = n7135 & n9253 ;
  assign n18015 = n18014 ^ n2317 ^ 1'b0 ;
  assign n18016 = n18015 ^ n15799 ^ 1'b0 ;
  assign n18017 = n4824 | n18016 ;
  assign n18018 = n16271 ^ n10009 ^ 1'b0 ;
  assign n18019 = n3945 | n18018 ;
  assign n18020 = n18019 ^ n6843 ^ 1'b0 ;
  assign n18021 = n13004 & n18020 ;
  assign n18022 = n6318 & n16190 ;
  assign n18023 = n18022 ^ n7503 ^ 1'b0 ;
  assign n18024 = n9139 & ~n15665 ;
  assign n18025 = n6874 & ~n18024 ;
  assign n18026 = n4433 & n8345 ;
  assign n18027 = n7169 ^ n6345 ^ 1'b0 ;
  assign n18028 = n18027 ^ n8799 ^ 1'b0 ;
  assign n18029 = ~n18026 & n18028 ;
  assign n18030 = n18029 ^ n10832 ^ n5793 ;
  assign n18031 = ~n5934 & n6661 ;
  assign n18032 = n18031 ^ n7908 ^ n5319 ;
  assign n18033 = n4879 | n18032 ;
  assign n18034 = n18033 ^ n13015 ^ n512 ;
  assign n18035 = n3457 ^ n312 ^ 1'b0 ;
  assign n18036 = ~x240 & n18035 ;
  assign n18037 = n10212 ^ n5266 ^ n868 ;
  assign n18038 = n17279 ^ n9617 ^ 1'b0 ;
  assign n18039 = ~n935 & n18038 ;
  assign n18040 = n12553 ^ n11967 ^ n3213 ;
  assign n18041 = n2136 & ~n6321 ;
  assign n18042 = ~n1939 & n18041 ;
  assign n18043 = n13968 ^ n7730 ^ 1'b0 ;
  assign n18044 = ~n5618 & n11667 ;
  assign n18045 = n18044 ^ x31 ^ 1'b0 ;
  assign n18046 = ( ~n7627 & n9581 ) | ( ~n7627 & n18045 ) | ( n9581 & n18045 ) ;
  assign n18047 = n12486 ^ x166 ^ 1'b0 ;
  assign n18048 = n18046 & n18047 ;
  assign n18049 = n18048 ^ n5840 ^ 1'b0 ;
  assign n18050 = ~n5460 & n18049 ;
  assign n18051 = n18043 & n18050 ;
  assign n18058 = ~n9215 & n17607 ;
  assign n18052 = ~n432 & n14416 ;
  assign n18053 = n18052 ^ n13201 ^ 1'b0 ;
  assign n18054 = n1291 & n18053 ;
  assign n18055 = n18054 ^ n6965 ^ 1'b0 ;
  assign n18056 = n14840 & n18055 ;
  assign n18057 = n11566 & n18056 ;
  assign n18059 = n18058 ^ n18057 ^ n13730 ;
  assign n18060 = n1372 | n3666 ;
  assign n18061 = n3155 | n18060 ;
  assign n18062 = ( n2444 & ~n16159 ) | ( n2444 & n18061 ) | ( ~n16159 & n18061 ) ;
  assign n18063 = n15807 ^ n6715 ^ 1'b0 ;
  assign n18064 = n6992 & ~n9996 ;
  assign n18065 = n1035 & n18064 ;
  assign n18066 = ( n1724 & n3074 ) | ( n1724 & n13216 ) | ( n3074 & n13216 ) ;
  assign n18067 = ( n5729 & n15540 ) | ( n5729 & ~n18066 ) | ( n15540 & ~n18066 ) ;
  assign n18068 = n18007 | n18067 ;
  assign n18069 = n8352 ^ n7285 ^ 1'b0 ;
  assign n18070 = ( n16305 & ~n17887 ) | ( n16305 & n18069 ) | ( ~n17887 & n18069 ) ;
  assign n18071 = n17443 ^ x87 ^ 1'b0 ;
  assign n18072 = n17403 & n18071 ;
  assign n18073 = n5255 | n18072 ;
  assign n18074 = n2220 | n18008 ;
  assign n18075 = n18074 ^ n15480 ^ 1'b0 ;
  assign n18076 = n4081 ^ n706 ^ 1'b0 ;
  assign n18077 = n1251 | n18076 ;
  assign n18078 = ~n856 & n13065 ;
  assign n18079 = n18077 & n18078 ;
  assign n18080 = n2777 ^ n925 ^ 1'b0 ;
  assign n18081 = ~n18079 & n18080 ;
  assign n18082 = n14976 ^ n3136 ^ n797 ;
  assign n18083 = n7100 & n12953 ;
  assign n18084 = ~n18082 & n18083 ;
  assign n18085 = n1374 | n1769 ;
  assign n18086 = n18085 ^ n12911 ^ 1'b0 ;
  assign n18087 = ( n692 & n983 ) | ( n692 & ~n9645 ) | ( n983 & ~n9645 ) ;
  assign n18088 = n18058 | n18087 ;
  assign n18089 = n18086 & ~n18088 ;
  assign n18090 = n18089 ^ n16811 ^ n16148 ;
  assign n18091 = ( n3226 & n5146 ) | ( n3226 & n7070 ) | ( n5146 & n7070 ) ;
  assign n18092 = n3576 & ~n18091 ;
  assign n18093 = ~n11152 & n18092 ;
  assign n18094 = n18093 ^ n9351 ^ 1'b0 ;
  assign n18095 = n18094 ^ n3107 ^ 1'b0 ;
  assign n18096 = n4189 & ~n4980 ;
  assign n18097 = n15008 ^ n1678 ^ n538 ;
  assign n18102 = ( n6547 & n7733 ) | ( n6547 & ~n11550 ) | ( n7733 & ~n11550 ) ;
  assign n18103 = ( n12983 & n16540 ) | ( n12983 & n18102 ) | ( n16540 & n18102 ) ;
  assign n18098 = ~n3069 & n5803 ;
  assign n18099 = n4048 & n18098 ;
  assign n18100 = n3034 | n18099 ;
  assign n18101 = ~n5886 & n18100 ;
  assign n18104 = n18103 ^ n18101 ^ 1'b0 ;
  assign n18105 = n13798 ^ n2701 ^ 1'b0 ;
  assign n18106 = n1091 | n18105 ;
  assign n18107 = n18106 ^ n8253 ^ 1'b0 ;
  assign n18108 = n11076 ^ n10620 ^ 1'b0 ;
  assign n18109 = n5475 & ~n18108 ;
  assign n18110 = n18109 ^ n3789 ^ 1'b0 ;
  assign n18111 = n2991 & n18110 ;
  assign n18113 = ~n2012 & n5077 ;
  assign n18114 = n18113 ^ n3474 ^ 1'b0 ;
  assign n18112 = n16247 ^ n14600 ^ 1'b0 ;
  assign n18115 = n18114 ^ n18112 ^ n9712 ;
  assign n18119 = n2724 & n6776 ;
  assign n18116 = n2814 & ~n16333 ;
  assign n18117 = n12504 | n18116 ;
  assign n18118 = n2490 | n18117 ;
  assign n18120 = n18119 ^ n18118 ^ n15063 ;
  assign n18121 = n5088 ^ n2329 ^ n815 ;
  assign n18122 = n5420 & n18121 ;
  assign n18123 = n18122 ^ n11932 ^ 1'b0 ;
  assign n18124 = n18123 ^ n14299 ^ 1'b0 ;
  assign n18125 = n577 | n7696 ;
  assign n18126 = n16828 ^ n369 ^ 1'b0 ;
  assign n18127 = n6897 | n11159 ;
  assign n18128 = ~n17866 & n18127 ;
  assign n18129 = ~n6177 & n18128 ;
  assign n18130 = n3425 ^ n2283 ^ 1'b0 ;
  assign n18131 = n18130 ^ n16086 ^ 1'b0 ;
  assign n18132 = n17626 | n18131 ;
  assign n18133 = n13884 ^ n1030 ^ 1'b0 ;
  assign n18134 = ~n820 & n18133 ;
  assign n18135 = n18134 ^ n18019 ^ 1'b0 ;
  assign n18136 = n10405 | n18135 ;
  assign n18137 = n2001 & ~n10608 ;
  assign n18141 = n7549 ^ n1452 ^ 1'b0 ;
  assign n18142 = n1240 | n18141 ;
  assign n18138 = n4500 ^ x141 ^ 1'b0 ;
  assign n18139 = n8565 ^ n7086 ^ 1'b0 ;
  assign n18140 = n18138 & ~n18139 ;
  assign n18143 = n18142 ^ n18140 ^ 1'b0 ;
  assign n18144 = n16763 ^ n4373 ^ 1'b0 ;
  assign n18146 = n6675 ^ n847 ^ 1'b0 ;
  assign n18147 = n3654 & n18146 ;
  assign n18145 = n4685 ^ n4659 ^ 1'b0 ;
  assign n18148 = n18147 ^ n18145 ^ n2009 ;
  assign n18149 = n18148 ^ n16828 ^ n15710 ;
  assign n18151 = ( n3557 & n7002 ) | ( n3557 & ~n9058 ) | ( n7002 & ~n9058 ) ;
  assign n18150 = n1516 & ~n8608 ;
  assign n18152 = n18151 ^ n18150 ^ 1'b0 ;
  assign n18153 = ~n1596 & n18152 ;
  assign n18154 = n8679 & ~n11140 ;
  assign n18155 = n5618 ^ n3429 ^ 1'b0 ;
  assign n18156 = n18154 & n18155 ;
  assign n18157 = n12471 & n18156 ;
  assign n18158 = n18157 ^ x209 ^ 1'b0 ;
  assign n18159 = ~n7316 & n13106 ;
  assign n18160 = n18159 ^ n9501 ^ n1672 ;
  assign n18161 = n7921 ^ n3810 ^ 1'b0 ;
  assign n18162 = n13167 ^ x126 ^ 1'b0 ;
  assign n18163 = ~n798 & n11035 ;
  assign n18164 = n18163 ^ n10428 ^ 1'b0 ;
  assign n18165 = n1870 & n11236 ;
  assign n18166 = n18165 ^ n12285 ^ 1'b0 ;
  assign n18167 = n8217 & n13356 ;
  assign n18168 = n14560 & ~n15710 ;
  assign n18169 = n3434 & ~n15013 ;
  assign n18170 = n18169 ^ n12160 ^ 1'b0 ;
  assign n18171 = n15539 & ~n17305 ;
  assign n18172 = ~n7465 & n11801 ;
  assign n18173 = n4090 ^ n1812 ^ 1'b0 ;
  assign n18174 = n6339 & n18173 ;
  assign n18175 = n2055 & n11806 ;
  assign n18176 = n766 & ~n6390 ;
  assign n18177 = ( n15527 & ~n18175 ) | ( n15527 & n18176 ) | ( ~n18175 & n18176 ) ;
  assign n18178 = n8481 ^ x70 ^ 1'b0 ;
  assign n18179 = n7823 & n8579 ;
  assign n18180 = n7016 & n18179 ;
  assign n18181 = n1975 | n3232 ;
  assign n18182 = n7120 ^ n4930 ^ 1'b0 ;
  assign n18183 = n18182 ^ n8346 ^ 1'b0 ;
  assign n18184 = n8927 ^ n398 ^ 1'b0 ;
  assign n18185 = n18183 & ~n18184 ;
  assign n18186 = ~n8159 & n18185 ;
  assign n18187 = n9250 ^ n5992 ^ 1'b0 ;
  assign n18188 = n8102 ^ n3264 ^ 1'b0 ;
  assign n18189 = n6706 & ~n18188 ;
  assign n18190 = n6554 | n18189 ;
  assign n18191 = n1757 & ~n5342 ;
  assign n18192 = n3814 & n5417 ;
  assign n18193 = n2041 & n9571 ;
  assign n18194 = ~n3662 & n18193 ;
  assign n18195 = n18194 ^ n16656 ^ 1'b0 ;
  assign n18196 = n18192 | n18195 ;
  assign n18197 = n3475 | n6549 ;
  assign n18198 = ( n4130 & n6678 ) | ( n4130 & ~n18197 ) | ( n6678 & ~n18197 ) ;
  assign n18199 = n14528 ^ n3557 ^ 1'b0 ;
  assign n18200 = n18199 ^ n12091 ^ 1'b0 ;
  assign n18201 = n9777 ^ n4709 ^ x78 ;
  assign n18202 = ~n8185 & n18201 ;
  assign n18203 = n1524 | n16679 ;
  assign n18204 = n18203 ^ n12709 ^ 1'b0 ;
  assign n18205 = ~n4917 & n11163 ;
  assign n18206 = n15944 & n18205 ;
  assign n18207 = n12968 & ~n16495 ;
  assign n18208 = n5816 & n18207 ;
  assign n18209 = ~n7801 & n18208 ;
  assign n18210 = n12368 & n13206 ;
  assign n18211 = ~n5034 & n18210 ;
  assign n18212 = n8491 ^ n3401 ^ 1'b0 ;
  assign n18213 = n5792 ^ n4955 ^ 1'b0 ;
  assign n18214 = n18212 & ~n18213 ;
  assign n18225 = ( x69 & n4966 ) | ( x69 & n11953 ) | ( n4966 & n11953 ) ;
  assign n18226 = n7003 ^ x184 ^ 1'b0 ;
  assign n18227 = n18225 | n18226 ;
  assign n18221 = n12457 ^ n1423 ^ 1'b0 ;
  assign n18222 = ~n6039 & n18221 ;
  assign n18215 = n4825 & n5739 ;
  assign n18216 = n18215 ^ n5732 ^ 1'b0 ;
  assign n18217 = n1688 & n2259 ;
  assign n18218 = n4347 & n18217 ;
  assign n18219 = n18218 ^ n11886 ^ 1'b0 ;
  assign n18220 = n18216 & ~n18219 ;
  assign n18223 = n18222 ^ n18220 ^ n12539 ;
  assign n18224 = n18223 ^ n12197 ^ n5139 ;
  assign n18228 = n18227 ^ n18224 ^ 1'b0 ;
  assign n18229 = n12919 & ~n18228 ;
  assign n18230 = x120 & ~n5316 ;
  assign n18231 = ( n1285 & n8393 ) | ( n1285 & n18230 ) | ( n8393 & n18230 ) ;
  assign n18232 = n18231 ^ n16830 ^ n13540 ;
  assign n18233 = n9853 | n18232 ;
  assign n18234 = ~n1055 & n1943 ;
  assign n18235 = ~n3090 & n18234 ;
  assign n18236 = n7034 ^ n4391 ^ 1'b0 ;
  assign n18237 = ~n11945 & n12768 ;
  assign n18238 = n18237 ^ n11177 ^ 1'b0 ;
  assign n18239 = n18238 ^ n7512 ^ 1'b0 ;
  assign n18240 = n1814 | n16269 ;
  assign n18241 = n8746 ^ n1661 ^ 1'b0 ;
  assign n18242 = ~n18240 & n18241 ;
  assign n18244 = n1155 | n11451 ;
  assign n18245 = n12615 ^ n5643 ^ 1'b0 ;
  assign n18246 = n18244 & n18245 ;
  assign n18243 = n15139 ^ n10640 ^ 1'b0 ;
  assign n18247 = n18246 ^ n18243 ^ 1'b0 ;
  assign n18248 = n15517 ^ n10063 ^ 1'b0 ;
  assign n18249 = n2584 | n8407 ;
  assign n18250 = n18249 ^ n7457 ^ 1'b0 ;
  assign n18251 = n18250 ^ n17771 ^ 1'b0 ;
  assign n18252 = ~n5018 & n14998 ;
  assign n18253 = n18252 ^ n10261 ^ 1'b0 ;
  assign n18254 = ~n3937 & n5994 ;
  assign n18255 = n8517 & n18254 ;
  assign n18256 = ~n6528 & n18255 ;
  assign n18257 = n18256 ^ n4103 ^ 1'b0 ;
  assign n18258 = n669 & ~n4817 ;
  assign n18259 = ~n895 & n18258 ;
  assign n18260 = n17044 ^ n11103 ^ 1'b0 ;
  assign n18265 = n3231 | n8005 ;
  assign n18266 = n10011 & ~n18265 ;
  assign n18261 = n15188 ^ n4004 ^ 1'b0 ;
  assign n18262 = n9682 & ~n18261 ;
  assign n18263 = ~n15125 & n18262 ;
  assign n18264 = ~n15149 & n18263 ;
  assign n18267 = n18266 ^ n18264 ^ n851 ;
  assign n18268 = n18267 ^ n3532 ^ n1845 ;
  assign n18271 = ( n9537 & n10065 ) | ( n9537 & ~n11531 ) | ( n10065 & ~n11531 ) ;
  assign n18269 = n1209 & ~n9597 ;
  assign n18270 = n1529 & ~n18269 ;
  assign n18272 = n18271 ^ n18270 ^ 1'b0 ;
  assign n18273 = n6422 | n18272 ;
  assign n18274 = ( n9918 & n10048 ) | ( n9918 & n18273 ) | ( n10048 & n18273 ) ;
  assign n18275 = ~n3153 & n6242 ;
  assign n18276 = n7157 & ~n18275 ;
  assign n18277 = ( ~n260 & n15636 ) | ( ~n260 & n18276 ) | ( n15636 & n18276 ) ;
  assign n18278 = n2141 & ~n8157 ;
  assign n18279 = n18278 ^ n4838 ^ 1'b0 ;
  assign n18280 = n5954 | n18279 ;
  assign n18281 = n6817 | n18280 ;
  assign n18282 = x122 | n18281 ;
  assign n18283 = n2354 ^ n809 ^ 1'b0 ;
  assign n18284 = n18282 & n18283 ;
  assign n18285 = ( n300 & n2263 ) | ( n300 & n9653 ) | ( n2263 & n9653 ) ;
  assign n18286 = n18285 ^ n5715 ^ 1'b0 ;
  assign n18287 = ~n6307 & n18286 ;
  assign n18288 = n2498 ^ n843 ^ 1'b0 ;
  assign n18289 = n2493 & n18288 ;
  assign n18290 = n18289 ^ n6912 ^ 1'b0 ;
  assign n18291 = n5813 | n18290 ;
  assign n18292 = ~n1158 & n3819 ;
  assign n18293 = n8346 & ~n18292 ;
  assign n18294 = ( n14008 & n18291 ) | ( n14008 & n18293 ) | ( n18291 & n18293 ) ;
  assign n18295 = n15621 ^ n10728 ^ 1'b0 ;
  assign n18296 = ( ~n3517 & n18294 ) | ( ~n3517 & n18295 ) | ( n18294 & n18295 ) ;
  assign n18297 = n14847 ^ n2628 ^ 1'b0 ;
  assign n18298 = n1241 & ~n6365 ;
  assign n18299 = n18298 ^ n844 ^ 1'b0 ;
  assign n18300 = n3020 & n18139 ;
  assign n18302 = n533 & ~n3532 ;
  assign n18301 = n12014 | n16895 ;
  assign n18303 = n18302 ^ n18301 ^ 1'b0 ;
  assign n18304 = n1896 ^ n699 ^ 1'b0 ;
  assign n18305 = n2867 & ~n18304 ;
  assign n18306 = ( n1203 & n6473 ) | ( n1203 & n7622 ) | ( n6473 & n7622 ) ;
  assign n18307 = ~n18305 & n18306 ;
  assign n18308 = n3514 & ~n17727 ;
  assign n18309 = n11878 & ~n18308 ;
  assign n18310 = ~n18307 & n18309 ;
  assign n18311 = n5719 | n18310 ;
  assign n18312 = n18303 & ~n18311 ;
  assign n18313 = n15800 ^ n6501 ^ 1'b0 ;
  assign n18314 = n2357 | n15936 ;
  assign n18315 = n6519 & ~n18314 ;
  assign n18316 = n7466 | n18315 ;
  assign n18317 = n3063 & ~n18316 ;
  assign n18318 = n943 & ~n15163 ;
  assign n18319 = n6021 & n8041 ;
  assign n18320 = n13652 & ~n18217 ;
  assign n18321 = n12301 & n18320 ;
  assign n18322 = n6290 & ~n18321 ;
  assign n18323 = n18322 ^ n18264 ^ 1'b0 ;
  assign n18324 = ( n2955 & ~n10468 ) | ( n2955 & n17995 ) | ( ~n10468 & n17995 ) ;
  assign n18325 = n18324 ^ n14603 ^ 1'b0 ;
  assign n18326 = n18325 ^ n3229 ^ 1'b0 ;
  assign n18327 = n4148 & ~n14793 ;
  assign n18328 = n18327 ^ n3125 ^ 1'b0 ;
  assign n18329 = n18328 ^ n1759 ^ 1'b0 ;
  assign n18330 = n7580 ^ n3296 ^ 1'b0 ;
  assign n18331 = n2392 & n18330 ;
  assign n18332 = n13597 & n18331 ;
  assign n18333 = n18332 ^ n823 ^ 1'b0 ;
  assign n18335 = n6986 ^ n2912 ^ 1'b0 ;
  assign n18336 = n18335 ^ n7231 ^ 1'b0 ;
  assign n18334 = n8112 ^ n1922 ^ 1'b0 ;
  assign n18337 = n18336 ^ n18334 ^ 1'b0 ;
  assign n18338 = n1650 & n11671 ;
  assign n18339 = n18338 ^ x231 ^ 1'b0 ;
  assign n18340 = n5681 ^ n4614 ^ 1'b0 ;
  assign n18341 = ~n18339 & n18340 ;
  assign n18342 = ~n8259 & n18341 ;
  assign n18343 = n17175 ^ n16710 ^ 1'b0 ;
  assign n18344 = n8325 ^ n1932 ^ 1'b0 ;
  assign n18345 = n5223 & ~n18344 ;
  assign n18346 = ~n4836 & n8424 ;
  assign n18347 = n18346 ^ n9164 ^ 1'b0 ;
  assign n18348 = n18347 ^ n9775 ^ n6626 ;
  assign n18349 = n18348 ^ n13444 ^ 1'b0 ;
  assign n18350 = n5056 ^ n4414 ^ n591 ;
  assign n18351 = n1319 & ~n18350 ;
  assign n18352 = n18351 ^ n2962 ^ 1'b0 ;
  assign n18353 = x196 | n2990 ;
  assign n18354 = ~n5539 & n13743 ;
  assign n18355 = n11767 & n18354 ;
  assign n18356 = n9645 & n18355 ;
  assign n18357 = n13576 ^ n4472 ^ 1'b0 ;
  assign n18358 = n18357 ^ n426 ^ 1'b0 ;
  assign n18359 = n1975 | n18358 ;
  assign n18360 = n2675 ^ x18 ^ 1'b0 ;
  assign n18361 = n9396 | n18360 ;
  assign n18362 = n8755 | n18361 ;
  assign n18363 = ( n2688 & n13873 ) | ( n2688 & ~n18362 ) | ( n13873 & ~n18362 ) ;
  assign n18364 = n7779 ^ n7099 ^ n3431 ;
  assign n18365 = n2042 | n4013 ;
  assign n18366 = ( ~n2272 & n17160 ) | ( ~n2272 & n18365 ) | ( n17160 & n18365 ) ;
  assign n18367 = x174 & n8946 ;
  assign n18368 = ( n18364 & n18366 ) | ( n18364 & n18367 ) | ( n18366 & n18367 ) ;
  assign n18369 = n602 & n5792 ;
  assign n18370 = ~n14866 & n18369 ;
  assign n18371 = n18370 ^ n13321 ^ 1'b0 ;
  assign n18372 = n2820 & ~n8609 ;
  assign n18373 = n18372 ^ n8368 ^ 1'b0 ;
  assign n18374 = n8094 & n18373 ;
  assign n18375 = n7986 | n16191 ;
  assign n18376 = n18374 | n18375 ;
  assign n18377 = n2642 & ~n5248 ;
  assign n18378 = n18377 ^ n3255 ^ 1'b0 ;
  assign n18379 = ~n3079 & n18378 ;
  assign n18380 = n18106 ^ n1182 ^ n633 ;
  assign n18381 = n18380 ^ n7530 ^ 1'b0 ;
  assign n18382 = n18379 & n18381 ;
  assign n18383 = n16887 ^ n9735 ^ 1'b0 ;
  assign n18385 = n7528 ^ n1057 ^ 1'b0 ;
  assign n18386 = n3352 & n18385 ;
  assign n18384 = n3546 & ~n6802 ;
  assign n18387 = n18386 ^ n18384 ^ 1'b0 ;
  assign n18388 = ( ~n9506 & n18223 ) | ( ~n9506 & n18387 ) | ( n18223 & n18387 ) ;
  assign n18389 = n4575 ^ n4209 ^ 1'b0 ;
  assign n18390 = ( n3299 & n9730 ) | ( n3299 & ~n18389 ) | ( n9730 & ~n18389 ) ;
  assign n18393 = ~n389 & n2606 ;
  assign n18394 = ~n12264 & n18393 ;
  assign n18395 = n1000 | n18394 ;
  assign n18391 = n10505 ^ n5410 ^ 1'b0 ;
  assign n18392 = n6549 & n18391 ;
  assign n18396 = n18395 ^ n18392 ^ n15188 ;
  assign n18397 = n14119 ^ n4202 ^ 1'b0 ;
  assign n18398 = n12212 | n18397 ;
  assign n18399 = n1327 & n13439 ;
  assign n18400 = n8215 ^ n3023 ^ n1879 ;
  assign n18401 = n4095 & n17443 ;
  assign n18402 = n17338 & n18401 ;
  assign n18403 = n2299 | n2748 ;
  assign n18404 = x214 & ~n4617 ;
  assign n18405 = n15472 ^ n10044 ^ 1'b0 ;
  assign n18406 = n18404 | n18405 ;
  assign n18407 = n1266 & ~n15228 ;
  assign n18408 = n11355 & n18377 ;
  assign n18409 = ~n4715 & n18408 ;
  assign n18410 = n14193 ^ n6099 ^ 1'b0 ;
  assign n18411 = ~n17649 & n18410 ;
  assign n18412 = n18409 & n18411 ;
  assign n18413 = ( ~n8260 & n11271 ) | ( ~n8260 & n12180 ) | ( n11271 & n12180 ) ;
  assign n18414 = n12480 | n18413 ;
  assign n18415 = n18414 ^ n16269 ^ 1'b0 ;
  assign n18416 = n997 & ~n4989 ;
  assign n18417 = n5873 & n18416 ;
  assign n18418 = n13982 & n18417 ;
  assign n18419 = ( n6114 & ~n7161 ) | ( n6114 & n18418 ) | ( ~n7161 & n18418 ) ;
  assign n18420 = n18419 ^ n1659 ^ n843 ;
  assign n18421 = n11940 ^ n8238 ^ n7404 ;
  assign n18422 = n13583 ^ n4256 ^ 1'b0 ;
  assign n18423 = n18421 | n18422 ;
  assign n18424 = n4285 & n6715 ;
  assign n18425 = n18424 ^ n17592 ^ 1'b0 ;
  assign n18426 = ( ~n3080 & n7220 ) | ( ~n3080 & n15529 ) | ( n7220 & n15529 ) ;
  assign n18427 = x144 & n18426 ;
  assign n18428 = n18427 ^ n1453 ^ 1'b0 ;
  assign n18429 = x185 & n18428 ;
  assign n18431 = ~n3602 & n8317 ;
  assign n18432 = n18431 ^ n4898 ^ 1'b0 ;
  assign n18430 = ( n11085 & ~n11603 ) | ( n11085 & n13860 ) | ( ~n11603 & n13860 ) ;
  assign n18433 = n18432 ^ n18430 ^ 1'b0 ;
  assign n18434 = n1812 & ~n11871 ;
  assign n18435 = n7624 & n18434 ;
  assign n18436 = ~n5698 & n18435 ;
  assign n18437 = n14962 ^ n14130 ^ 1'b0 ;
  assign n18438 = n6306 & ~n18437 ;
  assign n18439 = ~n415 & n7131 ;
  assign n18440 = ( n1927 & ~n6462 ) | ( n1927 & n18439 ) | ( ~n6462 & n18439 ) ;
  assign n18441 = n16811 & n18440 ;
  assign n18442 = ~n476 & n1269 ;
  assign n18443 = n18442 ^ x235 ^ 1'b0 ;
  assign n18444 = n18443 ^ x175 ^ 1'b0 ;
  assign n18447 = n14789 ^ n5904 ^ 1'b0 ;
  assign n18448 = ~n5410 & n18447 ;
  assign n18445 = n868 & ~n1802 ;
  assign n18446 = n1489 & n18445 ;
  assign n18449 = n18448 ^ n18446 ^ 1'b0 ;
  assign n18450 = n18449 ^ n471 ^ 1'b0 ;
  assign n18451 = n12320 & ~n18450 ;
  assign n18452 = n18451 ^ n10643 ^ 1'b0 ;
  assign n18453 = ~n7599 & n11791 ;
  assign n18454 = n1928 ^ n608 ^ 1'b0 ;
  assign n18455 = ~n11998 & n14516 ;
  assign n18456 = ~n18454 & n18455 ;
  assign n18457 = n18453 & ~n18456 ;
  assign n18458 = n5171 & n18457 ;
  assign n18459 = n18458 ^ n5596 ^ 1'b0 ;
  assign n18462 = ~n11661 & n15182 ;
  assign n18460 = n2667 & n5781 ;
  assign n18461 = n7576 | n18460 ;
  assign n18463 = n18462 ^ n18461 ^ 1'b0 ;
  assign n18464 = n6140 ^ n5991 ^ n2046 ;
  assign n18465 = n5377 ^ n3823 ^ 1'b0 ;
  assign n18466 = n1365 & ~n4323 ;
  assign n18467 = n18466 ^ n5763 ^ 1'b0 ;
  assign n18468 = n17554 | n18467 ;
  assign n18469 = ~n286 & n8996 ;
  assign n18470 = n18469 ^ n1816 ^ 1'b0 ;
  assign n18471 = n18470 ^ n11902 ^ 1'b0 ;
  assign n18472 = ~n4364 & n18471 ;
  assign n18473 = n3899 ^ n3220 ^ 1'b0 ;
  assign n18474 = n18472 & n18473 ;
  assign n18475 = n8524 ^ n5264 ^ 1'b0 ;
  assign n18476 = n4878 & ~n6303 ;
  assign n18477 = n18476 ^ n9861 ^ 1'b0 ;
  assign n18478 = n12875 | n15737 ;
  assign n18479 = n18478 ^ n12822 ^ 1'b0 ;
  assign n18480 = n2510 & ~n18479 ;
  assign n18481 = n16347 ^ n9288 ^ n6045 ;
  assign n18482 = n18481 ^ n9643 ^ 1'b0 ;
  assign n18483 = n14124 ^ n13045 ^ n9658 ;
  assign n18484 = ~n5628 & n18483 ;
  assign n18485 = ~n7127 & n18484 ;
  assign n18486 = ~n11698 & n18485 ;
  assign n18487 = ( n15083 & ~n18482 ) | ( n15083 & n18486 ) | ( ~n18482 & n18486 ) ;
  assign n18488 = n6681 ^ n2350 ^ 1'b0 ;
  assign n18489 = n13019 & n18488 ;
  assign n18490 = n9901 & n16695 ;
  assign n18491 = n18490 ^ n3282 ^ 1'b0 ;
  assign n18492 = n17531 ^ n6247 ^ x155 ;
  assign n18493 = ( ~n2769 & n4232 ) | ( ~n2769 & n18492 ) | ( n4232 & n18492 ) ;
  assign n18494 = n18493 ^ n14011 ^ 1'b0 ;
  assign n18500 = n1407 & ~n7216 ;
  assign n18501 = n18500 ^ n1909 ^ 1'b0 ;
  assign n18499 = ~n1597 & n4072 ;
  assign n18502 = n18501 ^ n18499 ^ 1'b0 ;
  assign n18503 = n18502 ^ n3094 ^ 1'b0 ;
  assign n18495 = n9367 & n18481 ;
  assign n18496 = n18495 ^ n14684 ^ 1'b0 ;
  assign n18497 = n10427 & n17185 ;
  assign n18498 = n18496 & ~n18497 ;
  assign n18504 = n18503 ^ n18498 ^ 1'b0 ;
  assign n18505 = n18504 ^ n3891 ^ n1486 ;
  assign n18506 = n15509 ^ x68 ^ 1'b0 ;
  assign n18507 = n7520 ^ n4353 ^ 1'b0 ;
  assign n18508 = ~n4626 & n18507 ;
  assign n18509 = n18508 ^ n5453 ^ 1'b0 ;
  assign n18510 = n16174 ^ n6994 ^ 1'b0 ;
  assign n18511 = n18510 ^ n10257 ^ 1'b0 ;
  assign n18512 = n18509 | n18511 ;
  assign n18513 = n18512 ^ n5611 ^ 1'b0 ;
  assign n18514 = ~n12865 & n18323 ;
  assign n18515 = n18514 ^ n3885 ^ 1'b0 ;
  assign n18516 = n5631 & ~n6527 ;
  assign n18517 = ( ~n1399 & n15267 ) | ( ~n1399 & n18516 ) | ( n15267 & n18516 ) ;
  assign n18518 = n1981 | n18517 ;
  assign n18519 = n2990 & ~n11886 ;
  assign n18520 = ( n18223 & ~n18518 ) | ( n18223 & n18519 ) | ( ~n18518 & n18519 ) ;
  assign n18521 = n7697 & ~n15767 ;
  assign n18522 = n18521 ^ n6344 ^ 1'b0 ;
  assign n18523 = ( n1196 & ~n17379 ) | ( n1196 & n18522 ) | ( ~n17379 & n18522 ) ;
  assign n18524 = n3758 ^ n3064 ^ n2524 ;
  assign n18525 = ~n264 & n18524 ;
  assign n18526 = n18525 ^ n8456 ^ 1'b0 ;
  assign n18527 = n4413 | n11458 ;
  assign n18528 = n18527 ^ n9814 ^ 1'b0 ;
  assign n18529 = n3952 | n17651 ;
  assign n18530 = ~n15913 & n18529 ;
  assign n18531 = n18530 ^ n14663 ^ 1'b0 ;
  assign n18532 = ~n18528 & n18531 ;
  assign n18533 = ~n11372 & n18532 ;
  assign n18534 = ~n6058 & n13450 ;
  assign n18535 = x23 & n9877 ;
  assign n18536 = n12710 & ~n13324 ;
  assign n18537 = n18536 ^ n17304 ^ 1'b0 ;
  assign n18538 = n6930 & ~n17481 ;
  assign n18539 = ( n7447 & n14752 ) | ( n7447 & n18538 ) | ( n14752 & n18538 ) ;
  assign n18540 = n18539 ^ n2978 ^ 1'b0 ;
  assign n18541 = n8970 & ~n18540 ;
  assign n18544 = n5722 & ~n12579 ;
  assign n18545 = n7767 & n18544 ;
  assign n18546 = ( ~n1241 & n10562 ) | ( ~n1241 & n18545 ) | ( n10562 & n18545 ) ;
  assign n18542 = n5135 ^ x62 ^ 1'b0 ;
  assign n18543 = n6267 & n18542 ;
  assign n18547 = n18546 ^ n18543 ^ 1'b0 ;
  assign n18548 = n10016 ^ n8984 ^ 1'b0 ;
  assign n18549 = ~n15448 & n18548 ;
  assign n18550 = n3984 ^ x90 ^ 1'b0 ;
  assign n18551 = n18550 ^ n5926 ^ 1'b0 ;
  assign n18552 = n8622 | n18551 ;
  assign n18553 = ( n4805 & n17188 ) | ( n4805 & ~n18552 ) | ( n17188 & ~n18552 ) ;
  assign n18554 = ~n673 & n7231 ;
  assign n18555 = ( n2645 & ~n15210 ) | ( n2645 & n18554 ) | ( ~n15210 & n18554 ) ;
  assign n18556 = n6999 ^ n1021 ^ 1'b0 ;
  assign n18557 = ~n1609 & n18556 ;
  assign n18558 = n12084 & ~n18557 ;
  assign n18559 = n9346 ^ n7562 ^ 1'b0 ;
  assign n18560 = n7710 & ~n18559 ;
  assign n18561 = ( n7359 & n13606 ) | ( n7359 & n18560 ) | ( n13606 & n18560 ) ;
  assign n18562 = ~n5169 & n18561 ;
  assign n18565 = n16867 ^ n9125 ^ n6207 ;
  assign n18563 = n14304 ^ n5368 ^ 1'b0 ;
  assign n18564 = n7568 & n18563 ;
  assign n18566 = n18565 ^ n18564 ^ n4422 ;
  assign n18567 = n17009 ^ n1062 ^ 1'b0 ;
  assign n18568 = x174 & n9884 ;
  assign n18569 = n18568 ^ n5610 ^ 1'b0 ;
  assign n18570 = n11315 & ~n18569 ;
  assign n18571 = n18570 ^ n5411 ^ 1'b0 ;
  assign n18572 = n3853 & ~n4019 ;
  assign n18573 = n6677 & n18572 ;
  assign n18574 = n1582 | n18573 ;
  assign n18575 = ~n259 & n3184 ;
  assign n18576 = n18575 ^ n9112 ^ 1'b0 ;
  assign n18577 = n18576 ^ n3094 ^ 1'b0 ;
  assign n18578 = n4343 | n14273 ;
  assign n18579 = n2582 | n18578 ;
  assign n18580 = ~n18577 & n18579 ;
  assign n18581 = n18580 ^ n3813 ^ 1'b0 ;
  assign n18582 = n18574 & n18581 ;
  assign n18583 = n11703 ^ n5472 ^ 1'b0 ;
  assign n18584 = n394 & n1476 ;
  assign n18585 = n18584 ^ n10432 ^ 1'b0 ;
  assign n18586 = ( n3672 & n6919 ) | ( n3672 & n7273 ) | ( n6919 & n7273 ) ;
  assign n18587 = n18586 ^ n13645 ^ 1'b0 ;
  assign n18588 = n4612 | n18587 ;
  assign n18589 = n18588 ^ n5641 ^ 1'b0 ;
  assign n18590 = n6010 ^ n3991 ^ 1'b0 ;
  assign n18594 = n4559 & n6094 ;
  assign n18591 = n14870 ^ n12429 ^ 1'b0 ;
  assign n18592 = n7113 | n18591 ;
  assign n18593 = ( n2989 & ~n11501 ) | ( n2989 & n18592 ) | ( ~n11501 & n18592 ) ;
  assign n18595 = n18594 ^ n18593 ^ 1'b0 ;
  assign n18596 = n14134 | n18595 ;
  assign n18597 = n2468 | n9587 ;
  assign n18598 = n1898 & n7187 ;
  assign n18599 = n17317 ^ n15438 ^ 1'b0 ;
  assign n18600 = ~n18598 & n18599 ;
  assign n18601 = ( ~x125 & n18597 ) | ( ~x125 & n18600 ) | ( n18597 & n18600 ) ;
  assign n18605 = n1666 & ~n2954 ;
  assign n18602 = n11234 ^ n8463 ^ 1'b0 ;
  assign n18603 = n5076 | n18602 ;
  assign n18604 = n18603 ^ n2950 ^ 1'b0 ;
  assign n18606 = n18605 ^ n18604 ^ n8066 ;
  assign n18607 = n16242 ^ n13352 ^ n13000 ;
  assign n18608 = n18607 ^ n4033 ^ 1'b0 ;
  assign n18609 = n4355 | n18608 ;
  assign n18610 = n18609 ^ n6406 ^ 1'b0 ;
  assign n18617 = ( ~n1495 & n8278 ) | ( ~n1495 & n8913 ) | ( n8278 & n8913 ) ;
  assign n18618 = n6613 & ~n18617 ;
  assign n18619 = ( n7598 & n13674 ) | ( n7598 & n18618 ) | ( n13674 & n18618 ) ;
  assign n18611 = n13545 ^ n4993 ^ 1'b0 ;
  assign n18612 = n2595 & ~n18611 ;
  assign n18613 = n2064 & ~n12608 ;
  assign n18614 = ~n18612 & n18613 ;
  assign n18615 = n9767 ^ n2103 ^ 1'b0 ;
  assign n18616 = n18614 | n18615 ;
  assign n18620 = n18619 ^ n18616 ^ 1'b0 ;
  assign n18621 = n10968 & ~n17223 ;
  assign n18622 = ~n8145 & n18621 ;
  assign n18623 = n17202 ^ n4776 ^ 1'b0 ;
  assign n18624 = ( n1356 & ~n7980 ) | ( n1356 & n18623 ) | ( ~n7980 & n18623 ) ;
  assign n18625 = ( n6654 & ~n18622 ) | ( n6654 & n18624 ) | ( ~n18622 & n18624 ) ;
  assign n18626 = n7382 & n16025 ;
  assign n18627 = n18626 ^ n16645 ^ 1'b0 ;
  assign n18628 = n10230 & ~n11302 ;
  assign n18629 = n18628 ^ n10121 ^ 1'b0 ;
  assign n18630 = n8391 & ~n16059 ;
  assign n18631 = n4159 & n18630 ;
  assign n18632 = n18631 ^ n1817 ^ 1'b0 ;
  assign n18633 = n11651 & n18632 ;
  assign n18634 = x76 & ~n16663 ;
  assign n18635 = n18634 ^ n11010 ^ 1'b0 ;
  assign n18636 = ( ~n1448 & n1504 ) | ( ~n1448 & n18635 ) | ( n1504 & n18635 ) ;
  assign n18637 = ( n6622 & n15379 ) | ( n6622 & n18636 ) | ( n15379 & n18636 ) ;
  assign n18643 = n6818 & n7550 ;
  assign n18638 = n5190 & ~n5428 ;
  assign n18639 = n7675 & n18638 ;
  assign n18640 = n18639 ^ n7664 ^ 1'b0 ;
  assign n18641 = n5219 | n18640 ;
  assign n18642 = n5920 & ~n18641 ;
  assign n18644 = n18643 ^ n18642 ^ 1'b0 ;
  assign n18645 = n1497 | n1658 ;
  assign n18648 = n5004 | n6848 ;
  assign n18649 = n18648 ^ n10917 ^ 1'b0 ;
  assign n18646 = n5424 & ~n13968 ;
  assign n18647 = n18646 ^ n16108 ^ n4350 ;
  assign n18650 = n18649 ^ n18647 ^ n10828 ;
  assign n18653 = ~n5686 & n14655 ;
  assign n18654 = n18653 ^ n3575 ^ 1'b0 ;
  assign n18655 = n7317 ^ n7169 ^ 1'b0 ;
  assign n18656 = n9447 & ~n18655 ;
  assign n18657 = ( n3525 & n18654 ) | ( n3525 & n18656 ) | ( n18654 & n18656 ) ;
  assign n18651 = n5438 & ~n14790 ;
  assign n18652 = n15154 & ~n18651 ;
  assign n18658 = n18657 ^ n18652 ^ 1'b0 ;
  assign n18659 = n610 & ~n14901 ;
  assign n18660 = n2427 & n9430 ;
  assign n18661 = n18659 & n18660 ;
  assign n18662 = n12672 & ~n18661 ;
  assign n18663 = n5259 & n14811 ;
  assign n18664 = n18663 ^ n1650 ^ 1'b0 ;
  assign n18665 = ~n7004 & n12556 ;
  assign n18666 = n876 & n10705 ;
  assign n18667 = ( ~n8505 & n9851 ) | ( ~n8505 & n18666 ) | ( n9851 & n18666 ) ;
  assign n18668 = n7168 ^ n1600 ^ 1'b0 ;
  assign n18669 = n16194 & ~n18668 ;
  assign n18670 = ~n18667 & n18669 ;
  assign n18674 = n5631 ^ n2692 ^ n2145 ;
  assign n18675 = ( n3842 & n8337 ) | ( n3842 & ~n18674 ) | ( n8337 & ~n18674 ) ;
  assign n18671 = n4756 & n13848 ;
  assign n18672 = n10942 & n18671 ;
  assign n18673 = n13716 & ~n18672 ;
  assign n18676 = n18675 ^ n18673 ^ 1'b0 ;
  assign n18677 = n13006 ^ n9067 ^ 1'b0 ;
  assign n18678 = n18676 & n18677 ;
  assign n18679 = ( n2293 & ~n10162 ) | ( n2293 & n18678 ) | ( ~n10162 & n18678 ) ;
  assign n18680 = n3080 | n16407 ;
  assign n18681 = n18680 ^ n3344 ^ 1'b0 ;
  assign n18682 = n16586 ^ n13704 ^ 1'b0 ;
  assign n18683 = ~n3975 & n18682 ;
  assign n18684 = ( ~n6901 & n8377 ) | ( ~n6901 & n13151 ) | ( n8377 & n13151 ) ;
  assign n18685 = n12427 | n18684 ;
  assign n18686 = n18685 ^ n2841 ^ 1'b0 ;
  assign n18687 = x239 & ~n8239 ;
  assign n18688 = n5763 & ~n18687 ;
  assign n18689 = n7225 & n18688 ;
  assign n18690 = n1659 & ~n11187 ;
  assign n18691 = n18690 ^ n13909 ^ 1'b0 ;
  assign n18692 = n18691 ^ n11143 ^ n10922 ;
  assign n18693 = x226 & n4053 ;
  assign n18694 = n10369 & ~n18693 ;
  assign n18695 = n6991 ^ n750 ^ 1'b0 ;
  assign n18696 = n3067 & n18695 ;
  assign n18697 = n18696 ^ n10642 ^ n6348 ;
  assign n18698 = n18694 & ~n18697 ;
  assign n18699 = n9086 ^ n4939 ^ 1'b0 ;
  assign n18700 = n438 | n18699 ;
  assign n18701 = n5599 & n6866 ;
  assign n18702 = n18701 ^ n4258 ^ 1'b0 ;
  assign n18703 = n680 | n18702 ;
  assign n18704 = ~n6192 & n18703 ;
  assign n18705 = n18704 ^ n6853 ^ 1'b0 ;
  assign n18706 = n18705 ^ n17562 ^ n3902 ;
  assign n18707 = ( n6361 & ~n18700 ) | ( n6361 & n18706 ) | ( ~n18700 & n18706 ) ;
  assign n18708 = n10221 ^ n10127 ^ n9614 ;
  assign n18709 = n1786 & ~n11435 ;
  assign n18710 = n8744 ^ n7976 ^ 1'b0 ;
  assign n18711 = ~n18709 & n18710 ;
  assign n18712 = ~n3644 & n16308 ;
  assign n18713 = ~n18711 & n18712 ;
  assign n18714 = n11363 & ~n18713 ;
  assign n18715 = n18714 ^ x60 ^ 1'b0 ;
  assign n18716 = ~n3525 & n12405 ;
  assign n18717 = n8158 ^ n5420 ^ 1'b0 ;
  assign n18718 = ( ~n468 & n4293 ) | ( ~n468 & n18717 ) | ( n4293 & n18717 ) ;
  assign n18719 = n16085 | n18718 ;
  assign n18720 = n7559 | n18719 ;
  assign n18721 = n11068 & ~n11157 ;
  assign n18722 = ~n4006 & n7716 ;
  assign n18723 = n8424 & n18722 ;
  assign n18724 = n18723 ^ n13362 ^ n12008 ;
  assign n18725 = n18724 ^ n6406 ^ n3126 ;
  assign n18726 = n6190 ^ n659 ^ 1'b0 ;
  assign n18727 = n6626 & ~n18726 ;
  assign n18728 = n1831 & n18727 ;
  assign n18729 = n1460 & ~n18728 ;
  assign n18730 = n3220 | n13645 ;
  assign n18731 = n18729 | n18730 ;
  assign n18732 = ~n7860 & n15473 ;
  assign n18733 = ( n8978 & ~n16350 ) | ( n8978 & n18732 ) | ( ~n16350 & n18732 ) ;
  assign n18734 = n4142 ^ n3472 ^ n2611 ;
  assign n18735 = n18734 ^ n2703 ^ 1'b0 ;
  assign n18736 = n8705 ^ n4278 ^ 1'b0 ;
  assign n18737 = ~n18735 & n18736 ;
  assign n18738 = n2469 & n10296 ;
  assign n18739 = ( n2570 & n13201 ) | ( n2570 & ~n18738 ) | ( n13201 & ~n18738 ) ;
  assign n18740 = n3776 & ~n8954 ;
  assign n18741 = n18740 ^ n3808 ^ n2439 ;
  assign n18742 = n18741 ^ n4305 ^ 1'b0 ;
  assign n18743 = n3109 & ~n18742 ;
  assign n18744 = n18743 ^ n17863 ^ 1'b0 ;
  assign n18745 = n16357 ^ n4717 ^ n1628 ;
  assign n18746 = ( n3613 & n10588 ) | ( n3613 & ~n18745 ) | ( n10588 & ~n18745 ) ;
  assign n18747 = n18746 ^ n6438 ^ 1'b0 ;
  assign n18748 = n12334 & ~n18747 ;
  assign n18749 = ~n9421 & n18748 ;
  assign n18750 = n18749 ^ n6373 ^ 1'b0 ;
  assign n18751 = ~n13680 & n17776 ;
  assign n18752 = n8404 ^ n2859 ^ 1'b0 ;
  assign n18753 = n18631 ^ n7745 ^ n5844 ;
  assign n18754 = n679 & n9258 ;
  assign n18755 = n13894 & n18754 ;
  assign n18756 = n18753 & ~n18755 ;
  assign n18757 = ( n4205 & ~n18752 ) | ( n4205 & n18756 ) | ( ~n18752 & n18756 ) ;
  assign n18758 = n16819 ^ n282 ^ 1'b0 ;
  assign n18759 = n11179 ^ n3254 ^ n976 ;
  assign n18760 = n15546 ^ n12525 ^ n2208 ;
  assign n18761 = n18760 ^ n790 ^ 1'b0 ;
  assign n18762 = ( n2176 & n6927 ) | ( n2176 & n18761 ) | ( n6927 & n18761 ) ;
  assign n18763 = ~n1918 & n8965 ;
  assign n18764 = n18763 ^ n4243 ^ 1'b0 ;
  assign n18765 = x14 | n18764 ;
  assign n18766 = n8000 ^ n2649 ^ 1'b0 ;
  assign n18767 = n13996 & n18766 ;
  assign n18768 = n18767 ^ n4180 ^ 1'b0 ;
  assign n18769 = n18768 ^ n16769 ^ 1'b0 ;
  assign n18770 = n18765 & ~n18769 ;
  assign n18771 = n12285 & ~n18770 ;
  assign n18772 = ~n6782 & n9709 ;
  assign n18773 = n10474 ^ n2634 ^ 1'b0 ;
  assign n18774 = ~n8127 & n18773 ;
  assign n18775 = n11172 & n18774 ;
  assign n18776 = n18775 ^ n9948 ^ 1'b0 ;
  assign n18777 = n9705 & n18776 ;
  assign n18778 = n4224 & n18777 ;
  assign n18779 = n18718 ^ n5696 ^ 1'b0 ;
  assign n18780 = ( n1161 & n11719 ) | ( n1161 & n18779 ) | ( n11719 & n18779 ) ;
  assign n18781 = n12595 ^ n12285 ^ n2349 ;
  assign n18782 = n13004 & n18781 ;
  assign n18783 = n10618 ^ n2439 ^ 1'b0 ;
  assign n18784 = ( n4651 & ~n5105 ) | ( n4651 & n18783 ) | ( ~n5105 & n18783 ) ;
  assign n18785 = ( n2717 & n3437 ) | ( n2717 & ~n12197 ) | ( n3437 & ~n12197 ) ;
  assign n18786 = n11418 & n18785 ;
  assign n18787 = n5492 & ~n6668 ;
  assign n18788 = ~n18786 & n18787 ;
  assign n18789 = ~n13084 & n14930 ;
  assign n18790 = ~n5206 & n18789 ;
  assign n18791 = n11589 ^ n7548 ^ n4006 ;
  assign n18792 = ~n6194 & n18791 ;
  assign n18793 = n18792 ^ n1152 ^ 1'b0 ;
  assign n18794 = n5567 | n18793 ;
  assign n18796 = n8403 | n11093 ;
  assign n18797 = n18796 ^ n5107 ^ 1'b0 ;
  assign n18795 = n8716 | n9287 ;
  assign n18798 = n18797 ^ n18795 ^ 1'b0 ;
  assign n18799 = n18798 ^ n3725 ^ 1'b0 ;
  assign n18800 = n18794 & n18799 ;
  assign n18801 = ~n4153 & n17313 ;
  assign n18802 = ~n929 & n1260 ;
  assign n18803 = n18802 ^ n5172 ^ 1'b0 ;
  assign n18804 = n18803 ^ n11931 ^ 1'b0 ;
  assign n18805 = n15022 & n18804 ;
  assign n18806 = n18805 ^ n18075 ^ n15767 ;
  assign n18807 = n10151 & n13833 ;
  assign n18808 = ( n4498 & n6132 ) | ( n4498 & ~n18807 ) | ( n6132 & ~n18807 ) ;
  assign n18809 = n10507 ^ n4223 ^ 1'b0 ;
  assign n18810 = ( ~n13733 & n18808 ) | ( ~n13733 & n18809 ) | ( n18808 & n18809 ) ;
  assign n18812 = n7721 & ~n14307 ;
  assign n18811 = n12600 | n17209 ;
  assign n18813 = n18812 ^ n18811 ^ 1'b0 ;
  assign n18814 = n15715 ^ n15549 ^ 1'b0 ;
  assign n18815 = n1308 & ~n5437 ;
  assign n18816 = n18814 & n18815 ;
  assign n18817 = ~n2727 & n14946 ;
  assign n18818 = ( x169 & n2953 ) | ( x169 & ~n15219 ) | ( n2953 & ~n15219 ) ;
  assign n18819 = ~n1558 & n18818 ;
  assign n18820 = ~n18817 & n18819 ;
  assign n18821 = ~n1019 & n4719 ;
  assign n18822 = n18820 | n18821 ;
  assign n18823 = n5582 ^ n1685 ^ 1'b0 ;
  assign n18824 = ~n4803 & n18823 ;
  assign n18825 = n10181 | n18824 ;
  assign n18826 = n8620 ^ n5076 ^ 1'b0 ;
  assign n18827 = ~n18825 & n18826 ;
  assign n18828 = n18827 ^ n13253 ^ n5177 ;
  assign n18829 = ~n1661 & n8707 ;
  assign n18830 = n18829 ^ n2348 ^ 1'b0 ;
  assign n18831 = n13448 & n18830 ;
  assign n18832 = n18831 ^ n11655 ^ 1'b0 ;
  assign n18833 = ( n1943 & n7540 ) | ( n1943 & ~n18627 ) | ( n7540 & ~n18627 ) ;
  assign n18835 = n3093 & n5862 ;
  assign n18836 = n1583 & n18835 ;
  assign n18834 = n2852 & n5694 ;
  assign n18837 = n18836 ^ n18834 ^ 1'b0 ;
  assign n18838 = n7712 & n18837 ;
  assign n18839 = n18838 ^ n9630 ^ 1'b0 ;
  assign n18840 = ~n4311 & n5495 ;
  assign n18841 = n18840 ^ n13012 ^ n5627 ;
  assign n18842 = ~n1890 & n16630 ;
  assign n18843 = n4113 & n18842 ;
  assign n18844 = n18843 ^ n11416 ^ 1'b0 ;
  assign n18845 = ( n2133 & n18841 ) | ( n2133 & n18844 ) | ( n18841 & n18844 ) ;
  assign n18846 = n18845 ^ n13619 ^ 1'b0 ;
  assign n18847 = ~n8480 & n14004 ;
  assign n18848 = n12917 & n18847 ;
  assign n18849 = n2229 & ~n18848 ;
  assign n18850 = n8926 & ~n13045 ;
  assign n18851 = n18850 ^ n13626 ^ 1'b0 ;
  assign n18852 = n3147 | n18851 ;
  assign n18853 = n2274 ^ n1155 ^ 1'b0 ;
  assign n18854 = ~n9063 & n15964 ;
  assign n18855 = n6328 ^ n2733 ^ 1'b0 ;
  assign n18856 = n1923 & ~n18855 ;
  assign n18857 = n13352 & ~n18856 ;
  assign n18858 = n18857 ^ n13167 ^ 1'b0 ;
  assign n18859 = n11474 ^ n10416 ^ 1'b0 ;
  assign n18860 = n8752 & n18859 ;
  assign n18861 = ~n4048 & n5114 ;
  assign n18863 = n12906 ^ n1688 ^ 1'b0 ;
  assign n18864 = n7369 | n18863 ;
  assign n18862 = n11367 | n11531 ;
  assign n18865 = n18864 ^ n18862 ^ 1'b0 ;
  assign n18866 = ( ~n13756 & n18861 ) | ( ~n13756 & n18865 ) | ( n18861 & n18865 ) ;
  assign n18867 = n10524 ^ n5183 ^ n4298 ;
  assign n18868 = n18866 | n18867 ;
  assign n18869 = n18868 ^ n6522 ^ 1'b0 ;
  assign n18870 = n10468 & n18869 ;
  assign n18871 = n11758 ^ n7359 ^ 1'b0 ;
  assign n18872 = ( n1158 & n3371 ) | ( n1158 & n18871 ) | ( n3371 & n18871 ) ;
  assign n18873 = n8626 & n17082 ;
  assign n18874 = ( n6103 & n9381 ) | ( n6103 & ~n18873 ) | ( n9381 & ~n18873 ) ;
  assign n18875 = ~n14125 & n18874 ;
  assign n18876 = ~n1009 & n5296 ;
  assign n18877 = n4090 & ~n18876 ;
  assign n18878 = ~n5148 & n6997 ;
  assign n18879 = ~n18683 & n18878 ;
  assign n18880 = n6699 | n8544 ;
  assign n18881 = n8971 ^ n460 ^ 1'b0 ;
  assign n18882 = n12333 | n14177 ;
  assign n18885 = n7525 ^ n4909 ^ 1'b0 ;
  assign n18886 = n4611 & ~n18885 ;
  assign n18883 = n8873 & ~n11075 ;
  assign n18884 = n18883 ^ n1727 ^ 1'b0 ;
  assign n18887 = n18886 ^ n18884 ^ n15681 ;
  assign n18888 = ( n7963 & n12179 ) | ( n7963 & ~n14546 ) | ( n12179 & ~n14546 ) ;
  assign n18889 = ( x136 & n10365 ) | ( x136 & n18888 ) | ( n10365 & n18888 ) ;
  assign n18892 = n6485 ^ n6086 ^ 1'b0 ;
  assign n18890 = ( n3429 & n3593 ) | ( n3429 & n3777 ) | ( n3593 & n3777 ) ;
  assign n18891 = ~n8194 & n18890 ;
  assign n18893 = n18892 ^ n18891 ^ 1'b0 ;
  assign n18894 = ( n11415 & ~n17574 ) | ( n11415 & n18893 ) | ( ~n17574 & n18893 ) ;
  assign n18895 = n9724 ^ n7576 ^ 1'b0 ;
  assign n18896 = n4948 & ~n8218 ;
  assign n18897 = ~n4693 & n12941 ;
  assign n18898 = n18897 ^ n9058 ^ 1'b0 ;
  assign n18899 = n18896 | n18898 ;
  assign n18900 = n15173 ^ n3247 ^ 1'b0 ;
  assign n18901 = n1158 & ~n7813 ;
  assign n18902 = n9635 & ~n18901 ;
  assign n18903 = n3220 & n18902 ;
  assign n18904 = n18903 ^ n15226 ^ 1'b0 ;
  assign n18905 = n13108 & n18904 ;
  assign n18906 = n18355 ^ n11005 ^ n8192 ;
  assign n18907 = ( n3203 & n6207 ) | ( n3203 & ~n18906 ) | ( n6207 & ~n18906 ) ;
  assign n18908 = ~n323 & n8802 ;
  assign n18909 = n14967 & ~n18908 ;
  assign n18910 = n18909 ^ n7426 ^ 1'b0 ;
  assign n18911 = ~n6568 & n18910 ;
  assign n18912 = n8161 & n14577 ;
  assign n18913 = ~n6257 & n18912 ;
  assign n18914 = n2849 | n8626 ;
  assign n18915 = n735 & ~n4203 ;
  assign n18916 = n18915 ^ n7468 ^ 1'b0 ;
  assign n18917 = n18916 ^ n5777 ^ n1160 ;
  assign n18918 = n18917 ^ n10065 ^ 1'b0 ;
  assign n18919 = n6406 & n14739 ;
  assign n18920 = n8702 ^ n736 ^ 1'b0 ;
  assign n18921 = n13673 | n18920 ;
  assign n18922 = n18921 ^ n2616 ^ 1'b0 ;
  assign n18923 = n6192 ^ n597 ^ 1'b0 ;
  assign n18925 = n10298 & ~n11234 ;
  assign n18926 = n18925 ^ n2202 ^ 1'b0 ;
  assign n18924 = n2932 ^ x143 ^ 1'b0 ;
  assign n18927 = n18926 ^ n18924 ^ n14114 ;
  assign n18928 = n16413 ^ n10550 ^ 1'b0 ;
  assign n18929 = n18928 ^ n15356 ^ n11509 ;
  assign n18930 = n15023 ^ n11851 ^ n887 ;
  assign n18931 = ~n4465 & n14887 ;
  assign n18932 = n18931 ^ n13109 ^ n12969 ;
  assign n18933 = ( n5126 & n18930 ) | ( n5126 & ~n18932 ) | ( n18930 & ~n18932 ) ;
  assign n18934 = n11475 ^ n9172 ^ 1'b0 ;
  assign n18935 = ~n7788 & n18934 ;
  assign n18936 = n11035 ^ n8067 ^ n4060 ;
  assign n18937 = n1142 & ~n18936 ;
  assign n18938 = ~n12598 & n18937 ;
  assign n18939 = n4009 & n4941 ;
  assign n18940 = n18939 ^ n7988 ^ 1'b0 ;
  assign n18941 = ~n18938 & n18940 ;
  assign n18942 = n13632 ^ n11584 ^ n9082 ;
  assign n18943 = n2618 | n10416 ;
  assign n18944 = n3694 & ~n18943 ;
  assign n18945 = ( ~n1775 & n15610 ) | ( ~n1775 & n18944 ) | ( n15610 & n18944 ) ;
  assign n18946 = n18033 & ~n18945 ;
  assign n18947 = n17967 ^ n8735 ^ 1'b0 ;
  assign n18948 = n16969 & ~n18947 ;
  assign n18949 = n3926 & n4045 ;
  assign n18950 = n18949 ^ n15733 ^ n15109 ;
  assign n18951 = n18102 & n18950 ;
  assign n18952 = ~n3356 & n18951 ;
  assign n18953 = n11126 ^ n3393 ^ 1'b0 ;
  assign n18954 = n18953 ^ n11232 ^ 1'b0 ;
  assign n18955 = n2488 | n18954 ;
  assign n18956 = ~n3223 & n8381 ;
  assign n18957 = n7873 ^ n7777 ^ 1'b0 ;
  assign n18958 = n11377 | n18957 ;
  assign n18960 = n3440 & n3651 ;
  assign n18959 = n5209 & ~n9263 ;
  assign n18961 = n18960 ^ n18959 ^ 1'b0 ;
  assign n18962 = ( n9764 & n16822 ) | ( n9764 & n18961 ) | ( n16822 & n18961 ) ;
  assign n18963 = n10778 ^ n3862 ^ 1'b0 ;
  assign n18964 = n15088 | n18963 ;
  assign n18965 = n18964 ^ n11425 ^ n275 ;
  assign n18966 = n1479 & ~n11234 ;
  assign n18967 = ~n3207 & n18966 ;
  assign n18968 = n18967 ^ n7739 ^ n6878 ;
  assign n18969 = n9933 ^ n3369 ^ 1'b0 ;
  assign n18970 = n3614 & n16499 ;
  assign n18971 = n10144 & n18970 ;
  assign n18972 = n1357 & ~n4867 ;
  assign n18973 = n8159 & n18972 ;
  assign n18974 = n18973 ^ n10524 ^ 1'b0 ;
  assign n18975 = n2687 & ~n10912 ;
  assign n18976 = n18975 ^ n7647 ^ 1'b0 ;
  assign n18977 = ( ~n7625 & n9047 ) | ( ~n7625 & n18976 ) | ( n9047 & n18976 ) ;
  assign n18978 = ( ~n6828 & n16785 ) | ( ~n6828 & n18977 ) | ( n16785 & n18977 ) ;
  assign n18979 = ( ~n8763 & n9441 ) | ( ~n8763 & n11426 ) | ( n9441 & n11426 ) ;
  assign n18981 = ~n1227 & n1327 ;
  assign n18982 = n18981 ^ n5101 ^ 1'b0 ;
  assign n18980 = n8355 ^ n7872 ^ 1'b0 ;
  assign n18983 = n18982 ^ n18980 ^ 1'b0 ;
  assign n18984 = n12411 | n18983 ;
  assign n18985 = n13298 & n15469 ;
  assign n18986 = n11119 & n18985 ;
  assign n18987 = n18984 & n18986 ;
  assign n18988 = n6332 ^ n3475 ^ 1'b0 ;
  assign n18989 = ~n2865 & n18988 ;
  assign n18990 = n18989 ^ n10919 ^ 1'b0 ;
  assign n18991 = n18990 ^ n13952 ^ n1658 ;
  assign n18992 = ~n1216 & n4074 ;
  assign n18993 = n13048 & n18992 ;
  assign n18994 = n18993 ^ n7589 ^ 1'b0 ;
  assign n18995 = n10334 & n18994 ;
  assign n18996 = n17705 ^ x113 ^ 1'b0 ;
  assign n18997 = n16569 | n18996 ;
  assign n18998 = n2598 & ~n2748 ;
  assign n18999 = ( n9765 & n18997 ) | ( n9765 & ~n18998 ) | ( n18997 & ~n18998 ) ;
  assign n19000 = n7008 ^ n725 ^ 1'b0 ;
  assign n19001 = n11001 | n19000 ;
  assign n19002 = ~n3561 & n10437 ;
  assign n19003 = n2720 & n13092 ;
  assign n19004 = n19003 ^ n4300 ^ 1'b0 ;
  assign n19005 = n19002 | n19004 ;
  assign n19006 = ~n8976 & n12387 ;
  assign n19007 = x254 & n14642 ;
  assign n19008 = n19007 ^ n7622 ^ 1'b0 ;
  assign n19009 = n19006 & n19008 ;
  assign n19010 = n8593 | n12575 ;
  assign n19011 = n19010 ^ n15027 ^ 1'b0 ;
  assign n19012 = n16821 ^ n4592 ^ 1'b0 ;
  assign n19013 = n19011 & ~n19012 ;
  assign n19014 = n4826 | n14583 ;
  assign n19015 = n19013 | n19014 ;
  assign n19016 = n17993 ^ n9579 ^ n8675 ;
  assign n19017 = n5298 ^ n1927 ^ 1'b0 ;
  assign n19018 = n19017 ^ n9244 ^ n8961 ;
  assign n19019 = n16136 & ~n19018 ;
  assign n19020 = n12425 & ~n12976 ;
  assign n19021 = n19020 ^ n8783 ^ 1'b0 ;
  assign n19022 = n17498 ^ n2435 ^ 1'b0 ;
  assign n19023 = x10 & n19022 ;
  assign n19024 = n11248 | n11474 ;
  assign n19025 = n5775 & ~n19024 ;
  assign n19026 = n11187 ^ n5037 ^ 1'b0 ;
  assign n19027 = n14133 ^ n7087 ^ 1'b0 ;
  assign n19028 = n1462 & ~n5090 ;
  assign n19029 = n5059 & n19028 ;
  assign n19030 = n1938 & ~n9378 ;
  assign n19031 = ~n14372 & n19030 ;
  assign n19032 = n14804 & ~n19031 ;
  assign n19033 = ~n19029 & n19032 ;
  assign n19034 = n6678 ^ n317 ^ 1'b0 ;
  assign n19036 = n8584 | n9514 ;
  assign n19037 = n15335 ^ x163 ^ 1'b0 ;
  assign n19038 = n7327 & n19037 ;
  assign n19039 = n3877 & n19038 ;
  assign n19040 = n1689 | n3813 ;
  assign n19041 = n19040 ^ n3907 ^ 1'b0 ;
  assign n19042 = n19041 ^ n11101 ^ n1977 ;
  assign n19043 = ~n3937 & n19042 ;
  assign n19044 = n19043 ^ n12072 ^ 1'b0 ;
  assign n19045 = n2908 & n19044 ;
  assign n19046 = n19045 ^ n16881 ^ n4398 ;
  assign n19047 = n11860 & ~n19046 ;
  assign n19048 = n19047 ^ n8732 ^ 1'b0 ;
  assign n19049 = ( n19036 & ~n19039 ) | ( n19036 & n19048 ) | ( ~n19039 & n19048 ) ;
  assign n19035 = n2332 & n13659 ;
  assign n19050 = n19049 ^ n19035 ^ 1'b0 ;
  assign n19051 = n13227 ^ n4692 ^ 1'b0 ;
  assign n19052 = x230 & ~n19051 ;
  assign n19053 = ~n1022 & n19052 ;
  assign n19054 = n19053 ^ n11173 ^ 1'b0 ;
  assign n19055 = n7529 & ~n14317 ;
  assign n19056 = n3264 & n6502 ;
  assign n19057 = n15112 ^ n1830 ^ 1'b0 ;
  assign n19058 = n9520 & ~n19057 ;
  assign n19059 = ( n12004 & ~n12454 ) | ( n12004 & n18164 ) | ( ~n12454 & n18164 ) ;
  assign n19060 = n2547 & n9754 ;
  assign n19061 = ( n1037 & n18046 ) | ( n1037 & ~n19060 ) | ( n18046 & ~n19060 ) ;
  assign n19062 = n10242 ^ n6915 ^ n6594 ;
  assign n19063 = n5918 | n6005 ;
  assign n19064 = ( ~n4151 & n19062 ) | ( ~n4151 & n19063 ) | ( n19062 & n19063 ) ;
  assign n19065 = ( ~n5779 & n8083 ) | ( ~n5779 & n16206 ) | ( n8083 & n16206 ) ;
  assign n19066 = ( n1324 & ~n4011 ) | ( n1324 & n4210 ) | ( ~n4011 & n4210 ) ;
  assign n19067 = n5329 | n8622 ;
  assign n19068 = n2006 | n19067 ;
  assign n19069 = n19068 ^ n8916 ^ 1'b0 ;
  assign n19070 = ~n2877 & n19069 ;
  assign n19071 = n19070 ^ n15509 ^ 1'b0 ;
  assign n19072 = n5373 & n19071 ;
  assign n19073 = ~n608 & n4738 ;
  assign n19074 = n264 & n19073 ;
  assign n19075 = n19074 ^ n4506 ^ 1'b0 ;
  assign n19076 = ~n1009 & n5610 ;
  assign n19077 = ( n4927 & ~n13116 ) | ( n4927 & n19076 ) | ( ~n13116 & n19076 ) ;
  assign n19078 = n2621 | n19077 ;
  assign n19079 = n19078 ^ n10934 ^ 1'b0 ;
  assign n19080 = n3304 ^ n1476 ^ 1'b0 ;
  assign n19081 = n3434 & ~n19080 ;
  assign n19082 = n4738 & n7629 ;
  assign n19083 = n19082 ^ n10595 ^ 1'b0 ;
  assign n19084 = ~n9308 & n19083 ;
  assign n19085 = ~n19081 & n19084 ;
  assign n19086 = n16014 ^ n15414 ^ n4114 ;
  assign n19087 = n19086 ^ n16558 ^ n4533 ;
  assign n19088 = ( ~n13038 & n15226 ) | ( ~n13038 & n19087 ) | ( n15226 & n19087 ) ;
  assign n19089 = n15686 & n19088 ;
  assign n19090 = ( n992 & n1593 ) | ( n992 & ~n4544 ) | ( n1593 & ~n4544 ) ;
  assign n19091 = n2833 & n8181 ;
  assign n19092 = n19091 ^ n4324 ^ 1'b0 ;
  assign n19093 = n19090 & n19092 ;
  assign n19094 = ~n4769 & n19093 ;
  assign n19095 = ~n906 & n10705 ;
  assign n19096 = n17562 ^ n17089 ^ n12341 ;
  assign n19097 = n3054 & ~n10690 ;
  assign n19098 = n14317 ^ n13068 ^ 1'b0 ;
  assign n19099 = n371 & ~n10075 ;
  assign n19100 = n19099 ^ n16547 ^ n2823 ;
  assign n19101 = ( n1687 & n9048 ) | ( n1687 & n19100 ) | ( n9048 & n19100 ) ;
  assign n19102 = n10942 ^ n783 ^ 1'b0 ;
  assign n19103 = ( x128 & n3788 ) | ( x128 & n6501 ) | ( n3788 & n6501 ) ;
  assign n19104 = n19103 ^ n5800 ^ n5404 ;
  assign n19105 = ( n12401 & n19102 ) | ( n12401 & ~n19104 ) | ( n19102 & ~n19104 ) ;
  assign n19106 = n1206 & ~n4618 ;
  assign n19107 = n17217 ^ n9641 ^ 1'b0 ;
  assign n19108 = ( ~n17714 & n19106 ) | ( ~n17714 & n19107 ) | ( n19106 & n19107 ) ;
  assign n19109 = n2640 & n16926 ;
  assign n19110 = n11334 ^ n3128 ^ 1'b0 ;
  assign n19111 = n9341 ^ x90 ^ 1'b0 ;
  assign n19112 = n3091 & ~n19111 ;
  assign n19113 = n19112 ^ n12206 ^ 1'b0 ;
  assign n19114 = n3123 & ~n19113 ;
  assign n19115 = ( n5069 & n6802 ) | ( n5069 & n19114 ) | ( n6802 & n19114 ) ;
  assign n19116 = n5049 | n19115 ;
  assign n19117 = n19058 | n19116 ;
  assign n19118 = n1935 ^ x4 ^ 1'b0 ;
  assign n19120 = n10428 & ~n16053 ;
  assign n19121 = ~n6375 & n19120 ;
  assign n19122 = ( n389 & ~n2865 ) | ( n389 & n11851 ) | ( ~n2865 & n11851 ) ;
  assign n19123 = n5551 ^ n550 ^ 1'b0 ;
  assign n19124 = n19123 ^ n2228 ^ n1778 ;
  assign n19125 = ~n7816 & n19124 ;
  assign n19126 = n19122 & n19125 ;
  assign n19127 = n19121 | n19126 ;
  assign n19128 = n18890 | n19127 ;
  assign n19119 = n4741 & n14417 ;
  assign n19129 = n19128 ^ n19119 ^ n382 ;
  assign n19130 = n10782 ^ n6442 ^ n6329 ;
  assign n19131 = n19130 ^ n1671 ^ 1'b0 ;
  assign n19132 = ~n7767 & n19131 ;
  assign n19134 = ( n4829 & ~n7334 ) | ( n4829 & n13288 ) | ( ~n7334 & n13288 ) ;
  assign n19133 = n4140 & ~n6328 ;
  assign n19135 = n19134 ^ n19133 ^ 1'b0 ;
  assign n19136 = n4806 & ~n17565 ;
  assign n19137 = n7711 ^ n2867 ^ 1'b0 ;
  assign n19138 = n4604 & ~n5582 ;
  assign n19139 = n16403 & n19138 ;
  assign n19140 = n11019 & n19139 ;
  assign n19141 = n4611 & n10194 ;
  assign n19142 = n1666 & n6295 ;
  assign n19143 = n14988 & n19142 ;
  assign n19144 = n19143 ^ n13072 ^ 1'b0 ;
  assign n19147 = n16690 ^ n10519 ^ n9538 ;
  assign n19145 = n10941 ^ n8001 ^ 1'b0 ;
  assign n19146 = n528 & n19145 ;
  assign n19148 = n19147 ^ n19146 ^ n16674 ;
  assign n19149 = ~n13644 & n18345 ;
  assign n19150 = n11582 & n19149 ;
  assign n19151 = n5441 ^ n729 ^ 1'b0 ;
  assign n19152 = n11715 ^ n1569 ^ 1'b0 ;
  assign n19153 = ~n3587 & n3739 ;
  assign n19154 = n19153 ^ n2064 ^ 1'b0 ;
  assign n19155 = ( n445 & n15493 ) | ( n445 & ~n19154 ) | ( n15493 & ~n19154 ) ;
  assign n19156 = n16709 ^ n4053 ^ x134 ;
  assign n19157 = ~n655 & n19156 ;
  assign n19158 = n19157 ^ n9247 ^ 1'b0 ;
  assign n19159 = n15867 ^ n7812 ^ 1'b0 ;
  assign n19160 = n16397 & n19159 ;
  assign n19161 = n17507 & n19160 ;
  assign n19162 = n6896 ^ n2305 ^ 1'b0 ;
  assign n19163 = n19124 & n19162 ;
  assign n19164 = ( n12100 & n13330 ) | ( n12100 & ~n19163 ) | ( n13330 & ~n19163 ) ;
  assign n19165 = ( n702 & n2649 ) | ( n702 & ~n10346 ) | ( n2649 & ~n10346 ) ;
  assign n19166 = n1940 & n4001 ;
  assign n19167 = ( n2312 & ~n2504 ) | ( n2312 & n14470 ) | ( ~n2504 & n14470 ) ;
  assign n19168 = n6302 & n19167 ;
  assign n19169 = n12906 & n19168 ;
  assign n19173 = n2365 & n6487 ;
  assign n19174 = ~n5681 & n19173 ;
  assign n19170 = n5532 ^ n5408 ^ n1757 ;
  assign n19171 = n7668 ^ n1148 ^ 1'b0 ;
  assign n19172 = ~n19170 & n19171 ;
  assign n19175 = n19174 ^ n19172 ^ 1'b0 ;
  assign n19176 = n16396 ^ n8015 ^ 1'b0 ;
  assign n19177 = n19175 & n19176 ;
  assign n19178 = ~n2025 & n19177 ;
  assign n19179 = n11455 ^ n6093 ^ 1'b0 ;
  assign n19180 = ~n19178 & n19179 ;
  assign n19181 = n19180 ^ n391 ^ 1'b0 ;
  assign n19182 = ~n831 & n13269 ;
  assign n19183 = n3592 & ~n12495 ;
  assign n19184 = ~n19182 & n19183 ;
  assign n19187 = n1658 | n3732 ;
  assign n19188 = n19187 ^ n661 ^ 1'b0 ;
  assign n19189 = ( x153 & x179 ) | ( x153 & ~n1318 ) | ( x179 & ~n1318 ) ;
  assign n19190 = n19188 & ~n19189 ;
  assign n19191 = n1220 | n19190 ;
  assign n19186 = ( ~n3689 & n7439 ) | ( ~n3689 & n16031 ) | ( n7439 & n16031 ) ;
  assign n19185 = n13555 ^ n7373 ^ 1'b0 ;
  assign n19192 = n19191 ^ n19186 ^ n19185 ;
  assign n19193 = ~n12270 & n16580 ;
  assign n19194 = n19193 ^ n3401 ^ 1'b0 ;
  assign n19195 = n11340 ^ n5744 ^ 1'b0 ;
  assign n19196 = n5873 ^ n3631 ^ n1269 ;
  assign n19197 = x203 | n19196 ;
  assign n19198 = n9370 ^ n2266 ^ 1'b0 ;
  assign n19199 = n19197 & n19198 ;
  assign n19200 = n6191 & n19199 ;
  assign n19201 = n18672 ^ n16954 ^ 1'b0 ;
  assign n19202 = n6619 | n19201 ;
  assign n19203 = n12627 ^ n10372 ^ 1'b0 ;
  assign n19204 = n9142 ^ n1151 ^ 1'b0 ;
  assign n19205 = n862 & ~n5591 ;
  assign n19206 = n8520 & n19205 ;
  assign n19207 = n14790 ^ n13354 ^ 1'b0 ;
  assign n19208 = n1804 | n19207 ;
  assign n19209 = n19206 & ~n19208 ;
  assign n19210 = n3273 ^ n1309 ^ 1'b0 ;
  assign n19211 = n5610 & n6960 ;
  assign n19212 = n1256 & n19211 ;
  assign n19213 = n19212 ^ n11363 ^ 1'b0 ;
  assign n19214 = n2313 & n6274 ;
  assign n19215 = n19214 ^ n9172 ^ 1'b0 ;
  assign n19216 = ( n2348 & n9013 ) | ( n2348 & n19215 ) | ( n9013 & n19215 ) ;
  assign n19217 = n7392 | n14031 ;
  assign n19218 = n5289 & n8034 ;
  assign n19219 = n7732 & ~n19218 ;
  assign n19220 = ~n8983 & n19219 ;
  assign n19222 = n2680 ^ n690 ^ 1'b0 ;
  assign n19221 = n4215 | n7589 ;
  assign n19223 = n19222 ^ n19221 ^ 1'b0 ;
  assign n19224 = n19223 ^ n16363 ^ 1'b0 ;
  assign n19225 = ~n19220 & n19224 ;
  assign n19226 = n6748 ^ n5999 ^ 1'b0 ;
  assign n19227 = n6420 & ~n19226 ;
  assign n19228 = n16317 & n16424 ;
  assign n19229 = n19228 ^ n15088 ^ 1'b0 ;
  assign n19230 = n19227 & ~n19229 ;
  assign n19231 = ( n6580 & ~n10445 ) | ( n6580 & n16619 ) | ( ~n10445 & n16619 ) ;
  assign n19232 = n12886 ^ n8042 ^ 1'b0 ;
  assign n19233 = n16413 ^ n10092 ^ 1'b0 ;
  assign n19234 = n13117 ^ n4061 ^ 1'b0 ;
  assign n19235 = n19233 & n19234 ;
  assign n19241 = n12832 ^ n5329 ^ 1'b0 ;
  assign n19240 = n8605 ^ n5524 ^ n4523 ;
  assign n19242 = n19241 ^ n19240 ^ n3104 ;
  assign n19236 = n6444 & ~n9212 ;
  assign n19237 = n2412 & ~n17715 ;
  assign n19238 = n19237 ^ n9685 ^ 1'b0 ;
  assign n19239 = n19236 & n19238 ;
  assign n19243 = n19242 ^ n19239 ^ 1'b0 ;
  assign n19244 = n17450 | n19243 ;
  assign n19245 = n3830 & n12598 ;
  assign n19246 = n12312 | n19245 ;
  assign n19247 = n17944 ^ n1788 ^ x13 ;
  assign n19248 = n8956 & ~n14848 ;
  assign n19249 = n2342 | n3140 ;
  assign n19250 = ~n8593 & n19249 ;
  assign n19251 = n19248 & n19250 ;
  assign n19252 = ~n6891 & n19251 ;
  assign n19253 = n17233 & ~n19252 ;
  assign n19254 = n19247 & n19253 ;
  assign n19256 = n13865 ^ n1838 ^ n983 ;
  assign n19257 = n671 & ~n9755 ;
  assign n19258 = n19257 ^ n14617 ^ x77 ;
  assign n19259 = n19258 ^ n14894 ^ 1'b0 ;
  assign n19260 = n19256 | n19259 ;
  assign n19255 = n1280 & n13385 ;
  assign n19261 = n19260 ^ n19255 ^ 1'b0 ;
  assign n19262 = ~n6941 & n9628 ;
  assign n19263 = n7488 & n17071 ;
  assign n19264 = ~n1452 & n19263 ;
  assign n19265 = n8021 ^ n7561 ^ 1'b0 ;
  assign n19266 = n19265 ^ n5912 ^ 1'b0 ;
  assign n19267 = ( n326 & ~n10202 ) | ( n326 & n10486 ) | ( ~n10202 & n10486 ) ;
  assign n19268 = n19267 ^ n2932 ^ 1'b0 ;
  assign n19269 = n15509 ^ n5201 ^ n3475 ;
  assign n19270 = n1040 & ~n4070 ;
  assign n19271 = n19269 & ~n19270 ;
  assign n19272 = n19271 ^ n15097 ^ n11298 ;
  assign n19273 = ~n629 & n19272 ;
  assign n19275 = n7144 | n12459 ;
  assign n19276 = n5133 | n19275 ;
  assign n19277 = n9853 & n19276 ;
  assign n19278 = n19277 ^ n8066 ^ 1'b0 ;
  assign n19279 = ( ~n4825 & n18280 ) | ( ~n4825 & n19278 ) | ( n18280 & n19278 ) ;
  assign n19274 = n4604 & n10065 ;
  assign n19280 = n19279 ^ n19274 ^ 1'b0 ;
  assign n19281 = n2149 | n15813 ;
  assign n19282 = n19281 ^ n18908 ^ 1'b0 ;
  assign n19283 = n19282 ^ n10683 ^ 1'b0 ;
  assign n19284 = n7086 & n19283 ;
  assign n19285 = n19284 ^ n10231 ^ 1'b0 ;
  assign n19286 = n15901 ^ n10606 ^ n1844 ;
  assign n19287 = n16713 ^ n2406 ^ 1'b0 ;
  assign n19288 = n7325 & ~n14515 ;
  assign n19289 = n19287 & n19288 ;
  assign n19290 = n7517 ^ n4049 ^ 1'b0 ;
  assign n19296 = n1752 ^ n1440 ^ n845 ;
  assign n19295 = n3576 ^ n658 ^ 1'b0 ;
  assign n19293 = ~n2350 & n7836 ;
  assign n19291 = n14407 ^ n5499 ^ 1'b0 ;
  assign n19292 = ~n1624 & n19291 ;
  assign n19294 = n19293 ^ n19292 ^ n5462 ;
  assign n19297 = n19296 ^ n19295 ^ n19294 ;
  assign n19298 = n19297 ^ n17401 ^ 1'b0 ;
  assign n19299 = n19290 | n19298 ;
  assign n19300 = n6612 ^ n3416 ^ 1'b0 ;
  assign n19301 = n3115 & ~n19300 ;
  assign n19302 = n6065 ^ n2476 ^ 1'b0 ;
  assign n19303 = n13901 ^ x61 ^ 1'b0 ;
  assign n19304 = n16954 & ~n19303 ;
  assign n19305 = ~n9226 & n10652 ;
  assign n19306 = n7003 ^ n1250 ^ 1'b0 ;
  assign n19307 = n17531 ^ n2558 ^ 1'b0 ;
  assign n19308 = ~n13680 & n13768 ;
  assign n19309 = ~n17731 & n19308 ;
  assign n19315 = n10654 ^ n2210 ^ 1'b0 ;
  assign n19313 = n10803 ^ n9548 ^ n2711 ;
  assign n19310 = n599 & ~n18983 ;
  assign n19311 = ~n10889 & n19310 ;
  assign n19312 = n9497 & ~n19311 ;
  assign n19314 = n19313 ^ n19312 ^ 1'b0 ;
  assign n19316 = n19315 ^ n19314 ^ 1'b0 ;
  assign n19317 = ~n19309 & n19316 ;
  assign n19318 = ~n11293 & n14528 ;
  assign n19319 = n12188 & n19318 ;
  assign n19320 = n16641 ^ x182 ^ 1'b0 ;
  assign n19321 = n2811 & n19320 ;
  assign n19322 = ~n6205 & n19321 ;
  assign n19323 = ( n1893 & ~n16644 ) | ( n1893 & n19322 ) | ( ~n16644 & n19322 ) ;
  assign n19324 = n19323 ^ n2906 ^ 1'b0 ;
  assign n19325 = ~n9649 & n19324 ;
  assign n19326 = n19325 ^ n18013 ^ 1'b0 ;
  assign n19327 = n19319 | n19326 ;
  assign n19328 = n12090 ^ n8135 ^ 1'b0 ;
  assign n19329 = n1695 | n5437 ;
  assign n19330 = n19329 ^ n3122 ^ 1'b0 ;
  assign n19331 = n18404 & n19330 ;
  assign n19332 = n6031 | n6897 ;
  assign n19333 = n19332 ^ n1690 ^ 1'b0 ;
  assign n19334 = n19333 ^ n5859 ^ 1'b0 ;
  assign n19335 = n9560 & ~n18181 ;
  assign n19336 = ~n9560 & n19335 ;
  assign n19337 = x172 & ~n5337 ;
  assign n19338 = ~n7486 & n19337 ;
  assign n19339 = n19338 ^ n12779 ^ n5197 ;
  assign n19340 = n300 & ~n17603 ;
  assign n19341 = ~n5795 & n8734 ;
  assign n19342 = n19341 ^ n5854 ^ 1'b0 ;
  assign n19343 = n19342 ^ n9614 ^ 1'b0 ;
  assign n19345 = ( n8248 & n12462 ) | ( n8248 & n14820 ) | ( n12462 & n14820 ) ;
  assign n19346 = ( n381 & ~n9891 ) | ( n381 & n19345 ) | ( ~n9891 & n19345 ) ;
  assign n19347 = n515 | n19346 ;
  assign n19344 = ~n5988 & n12722 ;
  assign n19348 = n19347 ^ n19344 ^ 1'b0 ;
  assign n19349 = n559 | n2255 ;
  assign n19350 = n19349 ^ n10385 ^ 1'b0 ;
  assign n19352 = ~n8473 & n13398 ;
  assign n19353 = n1888 & n19352 ;
  assign n19351 = n8642 | n15687 ;
  assign n19354 = n19353 ^ n19351 ^ 1'b0 ;
  assign n19355 = n10753 ^ n567 ^ 1'b0 ;
  assign n19356 = n11802 ^ n282 ^ 1'b0 ;
  assign n19357 = ~n8004 & n19356 ;
  assign n19358 = ~n17286 & n19357 ;
  assign n19359 = n9276 ^ n2009 ^ 1'b0 ;
  assign n19360 = n19358 | n19359 ;
  assign n19361 = n11545 | n19360 ;
  assign n19362 = n10180 ^ n735 ^ 1'b0 ;
  assign n19363 = n3954 & ~n19362 ;
  assign n19364 = ( n1755 & ~n9838 ) | ( n1755 & n19363 ) | ( ~n9838 & n19363 ) ;
  assign n19365 = n14223 ^ n13735 ^ 1'b0 ;
  assign n19366 = n15274 & ~n19365 ;
  assign n19367 = ~n5575 & n19366 ;
  assign n19368 = n19367 ^ n12978 ^ n8386 ;
  assign n19369 = n8447 ^ n1607 ^ 1'b0 ;
  assign n19370 = x156 & n19369 ;
  assign n19371 = n5099 ^ n2702 ^ n1810 ;
  assign n19372 = n19371 ^ n10821 ^ 1'b0 ;
  assign n19373 = ( n9025 & n19285 ) | ( n9025 & ~n19372 ) | ( n19285 & ~n19372 ) ;
  assign n19374 = n5405 ^ n1055 ^ 1'b0 ;
  assign n19375 = n10385 | n19374 ;
  assign n19376 = n19375 ^ n10773 ^ n10474 ;
  assign n19377 = n19376 ^ n16635 ^ n12513 ;
  assign n19378 = n9536 ^ n7171 ^ 1'b0 ;
  assign n19379 = n5377 & n17625 ;
  assign n19380 = n6826 ^ n2699 ^ 1'b0 ;
  assign n19381 = n19380 ^ n4490 ^ 1'b0 ;
  assign n19387 = n16845 ^ n3239 ^ 1'b0 ;
  assign n19388 = n12453 & n19387 ;
  assign n19389 = ~n14314 & n19388 ;
  assign n19390 = n19389 ^ n6030 ^ 1'b0 ;
  assign n19382 = n5320 & n14765 ;
  assign n19383 = ~n3095 & n8991 ;
  assign n19384 = ~n7342 & n19383 ;
  assign n19385 = ( n835 & n19382 ) | ( n835 & n19384 ) | ( n19382 & n19384 ) ;
  assign n19386 = n9664 & n19385 ;
  assign n19391 = n19390 ^ n19386 ^ 1'b0 ;
  assign n19395 = ( n6592 & ~n7222 ) | ( n6592 & n12812 ) | ( ~n7222 & n12812 ) ;
  assign n19392 = n862 & ~n3272 ;
  assign n19393 = n1096 & n19392 ;
  assign n19394 = n19393 ^ n11598 ^ n3369 ;
  assign n19396 = n19395 ^ n19394 ^ n1405 ;
  assign n19397 = ~x53 & n1077 ;
  assign n19399 = n11370 ^ n2986 ^ n1285 ;
  assign n19398 = ~n1382 & n4444 ;
  assign n19400 = n19399 ^ n19398 ^ 1'b0 ;
  assign n19401 = n19397 | n19400 ;
  assign n19402 = n14711 ^ n11372 ^ 1'b0 ;
  assign n19403 = ~n432 & n9094 ;
  assign n19404 = ~n4356 & n19403 ;
  assign n19405 = n19402 & ~n19404 ;
  assign n19406 = n4049 & n16346 ;
  assign n19407 = n19406 ^ n17848 ^ 1'b0 ;
  assign n19408 = n4510 ^ n4369 ^ n2379 ;
  assign n19409 = n19408 ^ n11308 ^ 1'b0 ;
  assign n19410 = n19409 ^ n953 ^ 1'b0 ;
  assign n19411 = ( ~n15428 & n19062 ) | ( ~n15428 & n19410 ) | ( n19062 & n19410 ) ;
  assign n19412 = n14435 | n19411 ;
  assign n19413 = n19412 ^ n2554 ^ 1'b0 ;
  assign n19414 = n17324 ^ n3396 ^ 1'b0 ;
  assign n19415 = n12971 ^ n907 ^ 1'b0 ;
  assign n19416 = n5162 & n19415 ;
  assign n19417 = n6822 ^ n3447 ^ 1'b0 ;
  assign n19418 = n19417 ^ n7525 ^ 1'b0 ;
  assign n19419 = ~n10888 & n19418 ;
  assign n19420 = n19419 ^ n2744 ^ 1'b0 ;
  assign n19421 = n17961 ^ n12232 ^ n12066 ;
  assign n19422 = ( n11147 & n17532 ) | ( n11147 & n19421 ) | ( n17532 & n19421 ) ;
  assign n19423 = n4909 | n5670 ;
  assign n19424 = n19423 ^ n1383 ^ 1'b0 ;
  assign n19425 = n5648 & n19424 ;
  assign n19426 = ~n17488 & n18425 ;
  assign n19427 = ~n402 & n1867 ;
  assign n19428 = n19427 ^ n6064 ^ 1'b0 ;
  assign n19429 = n1856 & n2268 ;
  assign n19430 = n19429 ^ n1266 ^ 1'b0 ;
  assign n19431 = ( ~n8689 & n11445 ) | ( ~n8689 & n19430 ) | ( n11445 & n19430 ) ;
  assign n19432 = n19431 ^ n7300 ^ 1'b0 ;
  assign n19433 = n19428 & ~n19432 ;
  assign n19434 = ~n16555 & n19433 ;
  assign n19435 = ~n8218 & n19434 ;
  assign n19436 = n19435 ^ n5918 ^ 1'b0 ;
  assign n19437 = n580 & n3624 ;
  assign n19438 = ~n2628 & n19437 ;
  assign n19439 = n1734 | n2385 ;
  assign n19440 = n19439 ^ n13252 ^ 1'b0 ;
  assign n19441 = n19440 ^ n9511 ^ n3455 ;
  assign n19444 = x133 | n3894 ;
  assign n19445 = n19444 ^ n12926 ^ n9433 ;
  assign n19446 = n19445 ^ n2427 ^ 1'b0 ;
  assign n19442 = n3982 ^ n3479 ^ n1944 ;
  assign n19443 = ~n6638 & n19442 ;
  assign n19447 = n19446 ^ n19443 ^ 1'b0 ;
  assign n19448 = n8102 | n15139 ;
  assign n19449 = n19448 ^ n7065 ^ 1'b0 ;
  assign n19450 = n11791 & ~n19449 ;
  assign n19451 = n19450 ^ n6636 ^ 1'b0 ;
  assign n19452 = ~n6558 & n19451 ;
  assign n19453 = n19452 ^ n8457 ^ 1'b0 ;
  assign n19454 = n19453 ^ n5609 ^ 1'b0 ;
  assign n19456 = n6425 | n14531 ;
  assign n19457 = n13763 | n19456 ;
  assign n19455 = n15672 | n18449 ;
  assign n19458 = n19457 ^ n19455 ^ 1'b0 ;
  assign n19459 = n11965 ^ n2500 ^ 1'b0 ;
  assign n19460 = ~n2804 & n6767 ;
  assign n19461 = ~n2554 & n19460 ;
  assign n19462 = ~n11357 & n19461 ;
  assign n19463 = n18949 | n19462 ;
  assign n19464 = ~n4168 & n14587 ;
  assign n19465 = n19464 ^ n14108 ^ 1'b0 ;
  assign n19466 = ( n2806 & n3354 ) | ( n2806 & ~n19465 ) | ( n3354 & ~n19465 ) ;
  assign n19467 = n14094 ^ n6829 ^ x232 ;
  assign n19468 = n10626 & ~n12786 ;
  assign n19469 = n19467 & n19468 ;
  assign n19470 = n19469 ^ n12899 ^ n2165 ;
  assign n19471 = n2675 & n17372 ;
  assign n19472 = n15667 ^ n8529 ^ 1'b0 ;
  assign n19473 = n9152 ^ n3514 ^ 1'b0 ;
  assign n19474 = n1682 | n7831 ;
  assign n19475 = n19473 | n19474 ;
  assign n19476 = n729 & n1454 ;
  assign n19477 = n8155 | n14138 ;
  assign n19478 = n19476 | n19477 ;
  assign n19479 = n5342 | n17241 ;
  assign n19480 = n820 & n19479 ;
  assign n19481 = n7075 & n11877 ;
  assign n19482 = n19481 ^ n12289 ^ 1'b0 ;
  assign n19483 = n19482 ^ n13668 ^ 1'b0 ;
  assign n19487 = n10549 ^ x158 ^ 1'b0 ;
  assign n19484 = n19397 ^ n905 ^ 1'b0 ;
  assign n19485 = n13213 & ~n17841 ;
  assign n19486 = n19484 & n19485 ;
  assign n19488 = n19487 ^ n19486 ^ n4472 ;
  assign n19490 = ( n8858 & n10340 ) | ( n8858 & n15125 ) | ( n10340 & n15125 ) ;
  assign n19491 = n17773 & ~n19490 ;
  assign n19489 = ~n10314 & n11013 ;
  assign n19492 = n19491 ^ n19489 ^ 1'b0 ;
  assign n19493 = n19492 ^ n6927 ^ n4631 ;
  assign n19494 = n1937 | n4207 ;
  assign n19495 = n19494 ^ n7044 ^ 1'b0 ;
  assign n19496 = n19495 ^ n18960 ^ n3714 ;
  assign n19497 = n8945 ^ n1257 ^ 1'b0 ;
  assign n19498 = n1385 | n4646 ;
  assign n19499 = n19498 ^ x226 ^ 1'b0 ;
  assign n19500 = n15464 ^ n13667 ^ 1'b0 ;
  assign n19501 = n1374 | n19500 ;
  assign n19502 = n19501 ^ n17233 ^ n13997 ;
  assign n19503 = ~n2901 & n8670 ;
  assign n19504 = ~n7743 & n9704 ;
  assign n19505 = n4277 & ~n14993 ;
  assign n19506 = ~n11578 & n19505 ;
  assign n19507 = ( n8043 & n19504 ) | ( n8043 & n19506 ) | ( n19504 & n19506 ) ;
  assign n19508 = n8418 ^ n7545 ^ n3005 ;
  assign n19509 = ~n5949 & n12059 ;
  assign n19510 = n3791 & n19509 ;
  assign n19511 = ( n5193 & ~n13206 ) | ( n5193 & n13348 ) | ( ~n13206 & n13348 ) ;
  assign n19512 = n4703 & n19511 ;
  assign n19513 = n19510 & n19512 ;
  assign n19514 = n19508 & ~n19513 ;
  assign n19515 = n19514 ^ n9351 ^ 1'b0 ;
  assign n19516 = n11145 ^ n9482 ^ n3458 ;
  assign n19517 = ~n5470 & n13939 ;
  assign n19518 = n13537 & n19517 ;
  assign n19519 = ( n6733 & ~n8981 ) | ( n6733 & n19424 ) | ( ~n8981 & n19424 ) ;
  assign n19520 = ~n604 & n7586 ;
  assign n19521 = n19520 ^ n11161 ^ 1'b0 ;
  assign n19522 = ~n19519 & n19521 ;
  assign n19523 = n19522 ^ n5359 ^ 1'b0 ;
  assign n19524 = n1914 & ~n2985 ;
  assign n19525 = n19524 ^ n16056 ^ n8206 ;
  assign n19526 = ~n19486 & n19525 ;
  assign n19527 = n14548 & n19526 ;
  assign n19528 = n4865 & n18624 ;
  assign n19529 = n3653 ^ n1865 ^ 1'b0 ;
  assign n19530 = n6647 | n19529 ;
  assign n19531 = n19530 ^ n1454 ^ 1'b0 ;
  assign n19532 = ( n11445 & n18864 ) | ( n11445 & n19531 ) | ( n18864 & n19531 ) ;
  assign n19533 = n19532 ^ n2670 ^ 1'b0 ;
  assign n19534 = n15125 ^ n8069 ^ 1'b0 ;
  assign n19535 = n19534 ^ n15550 ^ 1'b0 ;
  assign n19536 = n16756 ^ n9181 ^ 1'b0 ;
  assign n19537 = n12842 & n19536 ;
  assign n19538 = n6536 & n8894 ;
  assign n19539 = n19538 ^ n1930 ^ 1'b0 ;
  assign n19540 = n16927 ^ n13123 ^ n5686 ;
  assign n19541 = ( n1663 & n4411 ) | ( n1663 & ~n17602 ) | ( n4411 & ~n17602 ) ;
  assign n19542 = ( ~n4543 & n11376 ) | ( ~n4543 & n19541 ) | ( n11376 & n19541 ) ;
  assign n19543 = n1661 | n15219 ;
  assign n19544 = n19543 ^ n4851 ^ 1'b0 ;
  assign n19545 = n4448 | n7447 ;
  assign n19546 = n19545 ^ x246 ^ 1'b0 ;
  assign n19547 = n19546 ^ n9662 ^ 1'b0 ;
  assign n19548 = ~n992 & n19547 ;
  assign n19549 = ( ~n3244 & n15325 ) | ( ~n3244 & n19548 ) | ( n15325 & n19548 ) ;
  assign n19550 = n10102 ^ n1983 ^ 1'b0 ;
  assign n19551 = ~n12540 & n19550 ;
  assign n19552 = n5367 | n19551 ;
  assign n19556 = ( n4985 & ~n10618 ) | ( n4985 & n11034 ) | ( ~n10618 & n11034 ) ;
  assign n19553 = ~n1487 & n18027 ;
  assign n19554 = n19553 ^ n6701 ^ 1'b0 ;
  assign n19555 = n1158 & n19554 ;
  assign n19557 = n19556 ^ n19555 ^ n5374 ;
  assign n19558 = n19557 ^ n18723 ^ 1'b0 ;
  assign n19559 = ~n1181 & n7712 ;
  assign n19560 = ~n19558 & n19559 ;
  assign n19561 = n5066 & ~n6654 ;
  assign n19562 = n19561 ^ n8654 ^ 1'b0 ;
  assign n19563 = ( ~n12718 & n14496 ) | ( ~n12718 & n17551 ) | ( n14496 & n17551 ) ;
  assign n19564 = n7197 | n14548 ;
  assign n19565 = n19564 ^ n13348 ^ 1'b0 ;
  assign n19566 = n6260 & n19565 ;
  assign n19568 = n14519 ^ n7242 ^ 1'b0 ;
  assign n19567 = n9259 ^ n9170 ^ n2344 ;
  assign n19569 = n19568 ^ n19567 ^ 1'b0 ;
  assign n19570 = n2401 & ~n8140 ;
  assign n19571 = n19570 ^ n3022 ^ 1'b0 ;
  assign n19572 = n19571 ^ n13423 ^ n6568 ;
  assign n19573 = n19572 ^ n12313 ^ 1'b0 ;
  assign n19574 = ( n12340 & n13501 ) | ( n12340 & ~n15630 ) | ( n13501 & ~n15630 ) ;
  assign n19575 = ~n3274 & n19574 ;
  assign n19576 = ~n814 & n5850 ;
  assign n19577 = n10778 & n19576 ;
  assign n19578 = n1769 & ~n19577 ;
  assign n19579 = n10968 & n17914 ;
  assign n19580 = ~n5904 & n19579 ;
  assign n19581 = n6399 | n19580 ;
  assign n19582 = n19578 & n19581 ;
  assign n19583 = ~n19575 & n19582 ;
  assign n19584 = ~n9100 & n19583 ;
  assign n19592 = ~n4543 & n7225 ;
  assign n19593 = n8859 & ~n11020 ;
  assign n19594 = ~n19592 & n19593 ;
  assign n19585 = n11925 ^ n3767 ^ x161 ;
  assign n19587 = n1955 & n12403 ;
  assign n19586 = n1423 & n6417 ;
  assign n19588 = n19587 ^ n19586 ^ 1'b0 ;
  assign n19589 = n8140 | n8646 ;
  assign n19590 = n19588 & ~n19589 ;
  assign n19591 = ( ~n10422 & n19585 ) | ( ~n10422 & n19590 ) | ( n19585 & n19590 ) ;
  assign n19595 = n19594 ^ n19591 ^ x31 ;
  assign n19597 = ~n8268 & n9314 ;
  assign n19598 = ~n12305 & n19597 ;
  assign n19599 = n19598 ^ n11409 ^ 1'b0 ;
  assign n19600 = ~n14527 & n19599 ;
  assign n19596 = n9518 & ~n15939 ;
  assign n19601 = n19600 ^ n19596 ^ 1'b0 ;
  assign n19603 = n9775 ^ n1853 ^ 1'b0 ;
  assign n19604 = n5548 | n19603 ;
  assign n19602 = n13255 & n15226 ;
  assign n19605 = n19604 ^ n19602 ^ 1'b0 ;
  assign n19606 = n19605 ^ n16781 ^ n1395 ;
  assign n19607 = n19606 ^ n16886 ^ n5592 ;
  assign n19608 = n9752 ^ n4364 ^ n3735 ;
  assign n19609 = n19608 ^ n17104 ^ n12437 ;
  assign n19611 = n3128 | n7411 ;
  assign n19612 = n4767 | n19611 ;
  assign n19613 = ~n7829 & n19612 ;
  assign n19614 = n19613 ^ n2095 ^ 1'b0 ;
  assign n19615 = ( n10493 & n15969 ) | ( n10493 & ~n19614 ) | ( n15969 & ~n19614 ) ;
  assign n19616 = ( ~n3851 & n10557 ) | ( ~n3851 & n19615 ) | ( n10557 & n19615 ) ;
  assign n19610 = ~n3227 & n16887 ;
  assign n19617 = n19616 ^ n19610 ^ n6526 ;
  assign n19618 = n16413 ^ n4699 ^ n1430 ;
  assign n19619 = n5088 & n19618 ;
  assign n19620 = n5077 & n6016 ;
  assign n19621 = n19619 & n19620 ;
  assign n19622 = n9917 | n19621 ;
  assign n19629 = n13090 ^ n10753 ^ n6088 ;
  assign n19625 = n1720 ^ n1425 ^ 1'b0 ;
  assign n19624 = n17191 ^ x136 ^ 1'b0 ;
  assign n19626 = n19625 ^ n19624 ^ 1'b0 ;
  assign n19627 = n15677 | n19626 ;
  assign n19623 = ~n3664 & n12385 ;
  assign n19628 = n19627 ^ n19623 ^ 1'b0 ;
  assign n19630 = n19629 ^ n19628 ^ n1907 ;
  assign n19631 = n16473 ^ n6267 ^ n4156 ;
  assign n19632 = ~n1698 & n9096 ;
  assign n19633 = n10488 | n14807 ;
  assign n19634 = n3269 & n16370 ;
  assign n19635 = n7149 | n19634 ;
  assign n19636 = n19635 ^ n14316 ^ 1'b0 ;
  assign n19637 = n4751 ^ n1006 ^ 1'b0 ;
  assign n19638 = ~n11377 & n19637 ;
  assign n19639 = ~n4982 & n7305 ;
  assign n19640 = n19639 ^ n8603 ^ 1'b0 ;
  assign n19641 = ( n1332 & n13384 ) | ( n1332 & ~n19640 ) | ( n13384 & ~n19640 ) ;
  assign n19642 = n12284 ^ n11945 ^ 1'b0 ;
  assign n19643 = ( n19638 & n19641 ) | ( n19638 & n19642 ) | ( n19641 & n19642 ) ;
  assign n19646 = ~n1309 & n3589 ;
  assign n19647 = n19646 ^ n1257 ^ 1'b0 ;
  assign n19648 = n6725 & ~n19647 ;
  assign n19649 = n2972 | n19648 ;
  assign n19650 = n19649 ^ n16040 ^ 1'b0 ;
  assign n19645 = n18604 ^ n15791 ^ n10838 ;
  assign n19644 = ~n1867 & n16749 ;
  assign n19651 = n19650 ^ n19645 ^ n19644 ;
  assign n19652 = ~n8526 & n18410 ;
  assign n19653 = n19652 ^ n17385 ^ 1'b0 ;
  assign n19654 = n19653 ^ n9320 ^ n5524 ;
  assign n19655 = n6084 ^ n4564 ^ n1145 ;
  assign n19656 = n19655 ^ n9353 ^ n2121 ;
  assign n19657 = n9610 ^ n6517 ^ 1'b0 ;
  assign n19658 = n11388 & ~n19657 ;
  assign n19659 = ~n19656 & n19658 ;
  assign n19660 = n5325 | n19659 ;
  assign n19661 = n19660 ^ n12804 ^ 1'b0 ;
  assign n19662 = ~n1489 & n5481 ;
  assign n19663 = n597 | n1150 ;
  assign n19664 = n19663 ^ n4635 ^ 1'b0 ;
  assign n19665 = n19664 ^ n14954 ^ n8824 ;
  assign n19669 = n5093 & ~n15766 ;
  assign n19667 = n12401 | n16495 ;
  assign n19668 = n3426 & ~n19667 ;
  assign n19666 = ( n1106 & n3389 ) | ( n1106 & n3936 ) | ( n3389 & n3936 ) ;
  assign n19670 = n19669 ^ n19668 ^ n19666 ;
  assign n19671 = n15549 ^ n6807 ^ n417 ;
  assign n19672 = n13399 ^ n5500 ^ 1'b0 ;
  assign n19673 = ( n7976 & ~n19333 ) | ( n7976 & n19672 ) | ( ~n19333 & n19672 ) ;
  assign n19674 = n987 & ~n1530 ;
  assign n19675 = n5749 & n9775 ;
  assign n19676 = n19675 ^ n1393 ^ 1'b0 ;
  assign n19677 = n19674 & ~n19676 ;
  assign n19680 = n13444 ^ n7248 ^ 1'b0 ;
  assign n19678 = n3732 | n8713 ;
  assign n19679 = n19678 ^ n5984 ^ 1'b0 ;
  assign n19681 = n19680 ^ n19679 ^ n4700 ;
  assign n19682 = n19681 ^ n9115 ^ 1'b0 ;
  assign n19683 = n19677 & n19682 ;
  assign n19684 = n7231 & ~n8387 ;
  assign n19685 = ~n2991 & n19684 ;
  assign n19686 = n12903 ^ n10181 ^ n6114 ;
  assign n19687 = n2937 | n18569 ;
  assign n19688 = n19687 ^ n5324 ^ 1'b0 ;
  assign n19689 = ( n10780 & ~n18318 ) | ( n10780 & n19688 ) | ( ~n18318 & n19688 ) ;
  assign n19690 = ( ~n3479 & n8215 ) | ( ~n3479 & n12301 ) | ( n8215 & n12301 ) ;
  assign n19691 = n18780 ^ n14970 ^ n4487 ;
  assign n19692 = n8834 ^ n7005 ^ 1'b0 ;
  assign n19693 = n6411 & n7199 ;
  assign n19694 = n19693 ^ n15290 ^ n1638 ;
  assign n19695 = ( n9937 & ~n19692 ) | ( n9937 & n19694 ) | ( ~n19692 & n19694 ) ;
  assign n19696 = n5404 | n7631 ;
  assign n19697 = ( ~n1326 & n15906 ) | ( ~n1326 & n19696 ) | ( n15906 & n19696 ) ;
  assign n19698 = n2860 & n14922 ;
  assign n19699 = n18008 ^ n4398 ^ 1'b0 ;
  assign n19709 = ~n3983 & n13010 ;
  assign n19710 = n19709 ^ n5417 ^ 1'b0 ;
  assign n19711 = ( n5526 & n9824 ) | ( n5526 & n19710 ) | ( n9824 & n19710 ) ;
  assign n19700 = n5291 & n10016 ;
  assign n19701 = n6472 ^ n3588 ^ n1694 ;
  assign n19702 = ( n6418 & n7550 ) | ( n6418 & n19701 ) | ( n7550 & n19701 ) ;
  assign n19703 = n19702 ^ n7266 ^ 1'b0 ;
  assign n19704 = n19703 ^ n9494 ^ 1'b0 ;
  assign n19705 = n19700 | n19704 ;
  assign n19706 = n8750 & ~n19705 ;
  assign n19707 = ~n10464 & n14201 ;
  assign n19708 = n19706 & n19707 ;
  assign n19712 = n19711 ^ n19708 ^ 1'b0 ;
  assign n19713 = ~n1548 & n19712 ;
  assign n19714 = n18702 | n19713 ;
  assign n19715 = n19714 ^ n3125 ^ 1'b0 ;
  assign n19716 = n11304 & n17427 ;
  assign n19717 = n18661 & n19716 ;
  assign n19718 = n1458 & ~n11437 ;
  assign n19720 = n2567 & ~n10750 ;
  assign n19721 = n338 & ~n7959 ;
  assign n19722 = n19721 ^ n837 ^ 1'b0 ;
  assign n19723 = n8553 & ~n19722 ;
  assign n19724 = ( n4995 & n6275 ) | ( n4995 & n19723 ) | ( n6275 & n19723 ) ;
  assign n19725 = ~n19720 & n19724 ;
  assign n19719 = ( n4693 & n7187 ) | ( n4693 & n8504 ) | ( n7187 & n8504 ) ;
  assign n19726 = n19725 ^ n19719 ^ n10844 ;
  assign n19727 = ( n5042 & n7581 ) | ( n5042 & ~n11472 ) | ( n7581 & ~n11472 ) ;
  assign n19728 = n19058 ^ n16478 ^ 1'b0 ;
  assign n19729 = n6297 | n19728 ;
  assign n19730 = n19729 ^ n5065 ^ 1'b0 ;
  assign n19731 = n445 & n3843 ;
  assign n19732 = n6269 & n19731 ;
  assign n19733 = n19732 ^ n3506 ^ 1'b0 ;
  assign n19734 = n19733 ^ n7586 ^ 1'b0 ;
  assign n19735 = n14819 ^ n13923 ^ n8073 ;
  assign n19736 = n9544 ^ n4031 ^ 1'b0 ;
  assign n19737 = n9840 ^ n7416 ^ 1'b0 ;
  assign n19738 = n19736 & ~n19737 ;
  assign n19739 = n18307 ^ n6167 ^ 1'b0 ;
  assign n19741 = x87 & n7627 ;
  assign n19740 = n12677 ^ n6828 ^ n5527 ;
  assign n19742 = n19741 ^ n19740 ^ 1'b0 ;
  assign n19743 = n19742 ^ n14452 ^ n3943 ;
  assign n19744 = n4150 ^ n1285 ^ 1'b0 ;
  assign n19745 = ~n4889 & n19744 ;
  assign n19746 = n10520 & n19745 ;
  assign n19747 = n19746 ^ n3235 ^ 1'b0 ;
  assign n19748 = ~n16185 & n19747 ;
  assign n19749 = n16328 ^ n13968 ^ 1'b0 ;
  assign n19750 = n2560 | n19749 ;
  assign n19751 = n4305 | n6773 ;
  assign n19752 = n19751 ^ n4258 ^ 1'b0 ;
  assign n19753 = ~n15599 & n19752 ;
  assign n19754 = n18238 ^ n1923 ^ 1'b0 ;
  assign n19755 = n9030 & n19754 ;
  assign n19756 = n15185 ^ n5386 ^ 1'b0 ;
  assign n19757 = n1281 & n19756 ;
  assign n19758 = ~x162 & n19757 ;
  assign n19759 = n4174 & ~n8365 ;
  assign n19761 = n12569 ^ n9340 ^ n2522 ;
  assign n19760 = x158 & ~n17206 ;
  assign n19762 = n19761 ^ n19760 ^ n14943 ;
  assign n19763 = n17246 ^ n15311 ^ n1356 ;
  assign n19764 = n3420 ^ n1850 ^ 1'b0 ;
  assign n19765 = n18304 ^ n2616 ^ 1'b0 ;
  assign n19766 = ( n959 & n8796 ) | ( n959 & ~n11376 ) | ( n8796 & ~n11376 ) ;
  assign n19767 = ~n19765 & n19766 ;
  assign n19768 = n5494 ^ x177 ^ 1'b0 ;
  assign n19769 = n10838 & ~n19768 ;
  assign n19770 = n7049 | n13330 ;
  assign n19771 = n3240 & ~n4033 ;
  assign n19772 = ~n10267 & n19771 ;
  assign n19773 = n19772 ^ n1935 ^ 1'b0 ;
  assign n19774 = n7806 | n14333 ;
  assign n19775 = n19774 ^ x24 ^ 1'b0 ;
  assign n19776 = n5331 & ~n16845 ;
  assign n19777 = ~n19775 & n19776 ;
  assign n19778 = n14835 ^ n1216 ^ 1'b0 ;
  assign n19779 = ~n16004 & n19778 ;
  assign n19780 = n4928 ^ n4230 ^ 1'b0 ;
  assign n19781 = n19780 ^ n18825 ^ n1980 ;
  assign n19782 = n18728 | n19781 ;
  assign n19783 = n701 & ~n17617 ;
  assign n19784 = ~n1958 & n19783 ;
  assign n19785 = n6896 & n12301 ;
  assign n19786 = n16311 ^ n13403 ^ 1'b0 ;
  assign n19787 = n4812 & n19786 ;
  assign n19788 = ~n741 & n5475 ;
  assign n19789 = n19788 ^ n8114 ^ 1'b0 ;
  assign n19790 = n2665 | n7680 ;
  assign n19791 = n19789 | n19790 ;
  assign n19792 = ( n3700 & n11800 ) | ( n3700 & n13850 ) | ( n11800 & n13850 ) ;
  assign n19793 = n15774 ^ n15033 ^ 1'b0 ;
  assign n19794 = ~n4302 & n10326 ;
  assign n19795 = n19794 ^ n8328 ^ 1'b0 ;
  assign n19796 = n19795 ^ n6418 ^ n676 ;
  assign n19797 = n792 | n2534 ;
  assign n19798 = ( n14560 & n18631 ) | ( n14560 & ~n19797 ) | ( n18631 & ~n19797 ) ;
  assign n19799 = n12270 ^ n10111 ^ n5616 ;
  assign n19800 = n10414 & ~n19799 ;
  assign n19801 = n19800 ^ n10521 ^ 1'b0 ;
  assign n19803 = n5989 & n12489 ;
  assign n19804 = n2718 & n19803 ;
  assign n19802 = ~n8302 & n15899 ;
  assign n19805 = n19804 ^ n19802 ^ n8773 ;
  assign n19806 = n9729 | n15222 ;
  assign n19807 = n4034 & n19806 ;
  assign n19808 = ~n12015 & n19807 ;
  assign n19809 = ( n10941 & n15416 ) | ( n10941 & n19808 ) | ( n15416 & n19808 ) ;
  assign n19810 = n5823 ^ n2656 ^ n1007 ;
  assign n19811 = n19810 ^ n5366 ^ n3722 ;
  assign n19812 = ( n6856 & ~n7957 ) | ( n6856 & n8001 ) | ( ~n7957 & n8001 ) ;
  assign n19813 = ~n11988 & n19812 ;
  assign n19814 = n19813 ^ n4916 ^ 1'b0 ;
  assign n19815 = ~n5792 & n19814 ;
  assign n19816 = n19815 ^ n5719 ^ 1'b0 ;
  assign n19817 = n1765 ^ n569 ^ 1'b0 ;
  assign n19818 = n9255 & n19817 ;
  assign n19823 = n9424 & n17212 ;
  assign n19819 = n7851 ^ n3550 ^ 1'b0 ;
  assign n19820 = ~n11595 & n13500 ;
  assign n19821 = n10704 & n19820 ;
  assign n19822 = n19819 & ~n19821 ;
  assign n19824 = n19823 ^ n19822 ^ 1'b0 ;
  assign n19825 = n11913 ^ n9311 ^ 1'b0 ;
  assign n19826 = n7130 & ~n19825 ;
  assign n19827 = n19190 | n19826 ;
  assign n19828 = n8952 ^ n2980 ^ 1'b0 ;
  assign n19829 = n2167 & ~n4085 ;
  assign n19830 = ~n11521 & n19829 ;
  assign n19831 = n14585 ^ n9351 ^ 1'b0 ;
  assign n19832 = n12701 ^ n2473 ^ 1'b0 ;
  assign n19833 = ( n8460 & ~n13308 ) | ( n8460 & n19832 ) | ( ~n13308 & n19832 ) ;
  assign n19834 = n15636 | n19833 ;
  assign n19835 = n16017 | n19834 ;
  assign n19836 = n8183 | n14708 ;
  assign n19837 = n12036 ^ n11338 ^ n2344 ;
  assign n19838 = n7448 & ~n8654 ;
  assign n19839 = n19838 ^ n7044 ^ 1'b0 ;
  assign n19840 = n19839 ^ n17995 ^ n11379 ;
  assign n19841 = n1836 & ~n7011 ;
  assign n19842 = ( ~n7339 & n19840 ) | ( ~n7339 & n19841 ) | ( n19840 & n19841 ) ;
  assign n19843 = ( n6941 & ~n13382 ) | ( n6941 & n14850 ) | ( ~n13382 & n14850 ) ;
  assign n19844 = n19843 ^ n12129 ^ 1'b0 ;
  assign n19845 = n2515 & n3152 ;
  assign n19846 = ~n9632 & n19845 ;
  assign n19847 = n9795 ^ n6262 ^ 1'b0 ;
  assign n19848 = n3269 ^ n2439 ^ 1'b0 ;
  assign n19849 = n1105 ^ n675 ^ 1'b0 ;
  assign n19853 = n13020 ^ n11543 ^ n3302 ;
  assign n19850 = n7790 & ~n14969 ;
  assign n19851 = n19850 ^ n632 ^ 1'b0 ;
  assign n19852 = n2951 & n19851 ;
  assign n19854 = n19853 ^ n19852 ^ 1'b0 ;
  assign n19855 = n19356 & ~n19854 ;
  assign n19856 = ~n13714 & n19855 ;
  assign n19857 = ( n335 & ~n19849 ) | ( n335 & n19856 ) | ( ~n19849 & n19856 ) ;
  assign n19858 = n11076 ^ n7402 ^ n4791 ;
  assign n19859 = n14731 | n19858 ;
  assign n19861 = n5775 ^ n4929 ^ 1'b0 ;
  assign n19862 = n12784 | n19861 ;
  assign n19863 = n3961 | n8500 ;
  assign n19864 = n19862 & ~n19863 ;
  assign n19860 = n17901 | n18686 ;
  assign n19865 = n19864 ^ n19860 ^ 1'b0 ;
  assign n19866 = n7047 & ~n7504 ;
  assign n19867 = ~n16152 & n19866 ;
  assign n19868 = n19867 ^ n8021 ^ 1'b0 ;
  assign n19869 = n14266 & ~n15891 ;
  assign n19870 = n19869 ^ n3625 ^ 1'b0 ;
  assign n19871 = n17129 | n19870 ;
  assign n19872 = ( ~n2223 & n4769 ) | ( ~n2223 & n8149 ) | ( n4769 & n8149 ) ;
  assign n19873 = ~n4555 & n12102 ;
  assign n19874 = n19873 ^ n13505 ^ 1'b0 ;
  assign n19875 = n8393 ^ n5753 ^ n1630 ;
  assign n19876 = n19875 ^ n12812 ^ n10096 ;
  assign n19877 = n19876 ^ n6679 ^ 1'b0 ;
  assign n19878 = ~n3640 & n19877 ;
  assign n19879 = n17553 ^ n4438 ^ 1'b0 ;
  assign n19880 = ~n2921 & n13017 ;
  assign n19881 = ( n498 & ~n1000 ) | ( n498 & n13009 ) | ( ~n1000 & n13009 ) ;
  assign n19882 = n19881 ^ n12539 ^ n2055 ;
  assign n19883 = ~n3080 & n4324 ;
  assign n19884 = n14715 | n19883 ;
  assign n19885 = n5427 & n14416 ;
  assign n19886 = ~n1506 & n14975 ;
  assign n19887 = n4604 & ~n6855 ;
  assign n19888 = n19886 & n19887 ;
  assign n19889 = n13326 ^ n6437 ^ 1'b0 ;
  assign n19890 = n10201 & ~n19889 ;
  assign n19891 = ~n17535 & n19890 ;
  assign n19892 = n8222 | n19891 ;
  assign n19893 = n7741 & n8433 ;
  assign n19894 = n3215 ^ n1476 ^ 1'b0 ;
  assign n19895 = n19894 ^ n6473 ^ 1'b0 ;
  assign n19896 = n19011 ^ n16215 ^ n1463 ;
  assign n19897 = n7776 & n15856 ;
  assign n19898 = n19897 ^ n17184 ^ 1'b0 ;
  assign n19900 = ( n3004 & n10624 ) | ( n3004 & n15969 ) | ( n10624 & n15969 ) ;
  assign n19899 = ~n7708 & n12778 ;
  assign n19901 = n19900 ^ n19899 ^ 1'b0 ;
  assign n19902 = n17129 ^ n13917 ^ 1'b0 ;
  assign n19903 = n18904 & n19902 ;
  assign n19904 = ~n9792 & n18972 ;
  assign n19905 = n19904 ^ n4574 ^ 1'b0 ;
  assign n19906 = n19903 & n19905 ;
  assign n19907 = ( n1940 & ~n2854 ) | ( n1940 & n6395 ) | ( ~n2854 & n6395 ) ;
  assign n19908 = n19907 ^ n12089 ^ n2464 ;
  assign n19909 = ~n13553 & n19908 ;
  assign n19910 = n19305 & n19909 ;
  assign n19911 = n14867 ^ n6603 ^ 1'b0 ;
  assign n19912 = n19911 ^ n333 ^ 1'b0 ;
  assign n19913 = n5580 | n7503 ;
  assign n19914 = ( ~n6447 & n19440 ) | ( ~n6447 & n19913 ) | ( n19440 & n19913 ) ;
  assign n19915 = ( n1294 & n1298 ) | ( n1294 & ~n5791 ) | ( n1298 & ~n5791 ) ;
  assign n19916 = n14032 ^ n7585 ^ n6418 ;
  assign n19917 = n10744 ^ n10488 ^ 1'b0 ;
  assign n19918 = n19917 ^ n16964 ^ 1'b0 ;
  assign n19919 = ~n19916 & n19918 ;
  assign n19920 = ( n14201 & n19915 ) | ( n14201 & ~n19919 ) | ( n19915 & ~n19919 ) ;
  assign n19921 = n15182 ^ n10165 ^ n5528 ;
  assign n19922 = n3192 & ~n13152 ;
  assign n19923 = n16959 & n19922 ;
  assign n19924 = ( ~n16867 & n18748 ) | ( ~n16867 & n19923 ) | ( n18748 & n19923 ) ;
  assign n19925 = n3461 | n7179 ;
  assign n19926 = n19925 ^ n19103 ^ 1'b0 ;
  assign n19927 = n11157 | n19926 ;
  assign n19928 = n13137 | n19927 ;
  assign n19929 = n5305 ^ n2721 ^ n1110 ;
  assign n19930 = n19929 ^ n5897 ^ 1'b0 ;
  assign n19931 = n2645 | n19930 ;
  assign n19933 = ~n11231 & n19656 ;
  assign n19932 = n9590 ^ n5316 ^ n1836 ;
  assign n19934 = n19933 ^ n19932 ^ n5253 ;
  assign n19935 = n7289 & n7613 ;
  assign n19936 = n19935 ^ n1874 ^ 1'b0 ;
  assign n19937 = ~n3104 & n19936 ;
  assign n19938 = n19937 ^ n6137 ^ 1'b0 ;
  assign n19939 = n19938 ^ n2376 ^ 1'b0 ;
  assign n19940 = n19939 ^ n7140 ^ 1'b0 ;
  assign n19941 = n17394 ^ n15715 ^ 1'b0 ;
  assign n19942 = n19940 | n19941 ;
  assign n19943 = n19942 ^ n8217 ^ 1'b0 ;
  assign n19944 = n2331 & n19943 ;
  assign n19945 = n19944 ^ n4653 ^ 1'b0 ;
  assign n19946 = ~n8426 & n17179 ;
  assign n19947 = n18287 ^ n4804 ^ n4133 ;
  assign n19948 = x21 | n6213 ;
  assign n19949 = n2266 & n19948 ;
  assign n19950 = ~n16470 & n19949 ;
  assign n19951 = n19233 ^ n2680 ^ n1181 ;
  assign n19952 = n19951 ^ n6653 ^ 1'b0 ;
  assign n19953 = ~n7791 & n8100 ;
  assign n19954 = n19953 ^ n8310 ^ 1'b0 ;
  assign n19955 = n6227 | n19954 ;
  assign n19956 = ~n5664 & n5809 ;
  assign n19957 = n4091 & n19956 ;
  assign n19958 = ~n18814 & n19957 ;
  assign n19960 = n1937 & ~n18466 ;
  assign n19959 = n2702 & n11926 ;
  assign n19961 = n19960 ^ n19959 ^ 1'b0 ;
  assign n19962 = n8835 ^ n5645 ^ 1'b0 ;
  assign n19963 = n1132 & ~n9123 ;
  assign n19964 = ~n4072 & n19963 ;
  assign n19965 = n14636 ^ n5458 ^ 1'b0 ;
  assign n19966 = n3654 & ~n13336 ;
  assign n19967 = n5775 ^ n947 ^ 1'b0 ;
  assign n19968 = n7172 & n19967 ;
  assign n19969 = n2310 & ~n9035 ;
  assign n19970 = ~n19968 & n19969 ;
  assign n19971 = ( n17922 & ~n19966 ) | ( n17922 & n19970 ) | ( ~n19966 & n19970 ) ;
  assign n19972 = n10602 | n14892 ;
  assign n19973 = n1968 ^ x155 ^ x74 ;
  assign n19974 = n11533 & ~n14081 ;
  assign n19975 = n8315 ^ n5818 ^ 1'b0 ;
  assign n19976 = ( ~n2174 & n11624 ) | ( ~n2174 & n19975 ) | ( n11624 & n19975 ) ;
  assign n19977 = n1416 | n13414 ;
  assign n19978 = ~n7195 & n10002 ;
  assign n19979 = n19978 ^ n15825 ^ n12285 ;
  assign n19980 = ~n9623 & n19979 ;
  assign n19981 = ~n5027 & n6543 ;
  assign n19982 = ~n19980 & n19981 ;
  assign n19983 = n384 ^ x20 ^ 1'b0 ;
  assign n19984 = n2015 & ~n19983 ;
  assign n19985 = n19984 ^ n9375 ^ 1'b0 ;
  assign n19986 = n9845 & n19985 ;
  assign n19987 = n1034 | n19986 ;
  assign n19988 = ~n19982 & n19987 ;
  assign n19989 = n1750 & ~n1979 ;
  assign n19990 = ( n4061 & n10355 ) | ( n4061 & n19257 ) | ( n10355 & n19257 ) ;
  assign n19991 = n3622 | n11313 ;
  assign n19992 = ~n18329 & n19991 ;
  assign n19993 = n6266 ^ n5262 ^ 1'b0 ;
  assign n19994 = n19993 ^ n2828 ^ n1331 ;
  assign n19995 = ( ~n4285 & n10003 ) | ( ~n4285 & n19994 ) | ( n10003 & n19994 ) ;
  assign n19996 = ~n3862 & n5432 ;
  assign n19997 = n19996 ^ n3830 ^ 1'b0 ;
  assign n19998 = n5978 | n10366 ;
  assign n19999 = n12678 ^ n11715 ^ 1'b0 ;
  assign n20000 = ~n18032 & n19999 ;
  assign n20001 = n1500 & ~n6134 ;
  assign n20002 = n2538 & n20001 ;
  assign n20003 = n20002 ^ n10657 ^ 1'b0 ;
  assign n20004 = n13442 | n14138 ;
  assign n20005 = n6071 | n20004 ;
  assign n20007 = n2339 & n5601 ;
  assign n20008 = ~n1910 & n20007 ;
  assign n20009 = ( n615 & ~n675 ) | ( n615 & n20008 ) | ( ~n675 & n20008 ) ;
  assign n20010 = ~n4033 & n20009 ;
  assign n20006 = n7856 & ~n11768 ;
  assign n20011 = n20010 ^ n20006 ^ 1'b0 ;
  assign n20012 = n3402 & ~n8316 ;
  assign n20014 = n5816 & n18035 ;
  assign n20013 = n14030 & ~n18259 ;
  assign n20015 = n20014 ^ n20013 ^ 1'b0 ;
  assign n20016 = n12720 & n16698 ;
  assign n20017 = ~n4150 & n20016 ;
  assign n20018 = ~n1944 & n6885 ;
  assign n20019 = n20018 ^ n428 ^ 1'b0 ;
  assign n20020 = n20017 | n20019 ;
  assign n20021 = n20020 ^ n3086 ^ 1'b0 ;
  assign n20022 = n20021 ^ n16205 ^ n2942 ;
  assign n20023 = n1848 & n6204 ;
  assign n20024 = n18884 & ~n20023 ;
  assign n20025 = n1454 & ~n1675 ;
  assign n20026 = ~n13202 & n20025 ;
  assign n20027 = n20024 & n20026 ;
  assign n20028 = ~n20022 & n20027 ;
  assign n20029 = ~n6310 & n17228 ;
  assign n20033 = n967 | n1345 ;
  assign n20034 = n18302 & ~n20033 ;
  assign n20035 = n20034 ^ n13085 ^ 1'b0 ;
  assign n20030 = n1267 | n2931 ;
  assign n20031 = n20030 ^ n1022 ^ 1'b0 ;
  assign n20032 = n12533 | n20031 ;
  assign n20036 = n20035 ^ n20032 ^ 1'b0 ;
  assign n20037 = n2243 & n11545 ;
  assign n20038 = ~n19798 & n20037 ;
  assign n20039 = n9292 ^ n3317 ^ 1'b0 ;
  assign n20040 = n8507 & n8872 ;
  assign n20041 = n1791 & n19096 ;
  assign n20042 = ~n20040 & n20041 ;
  assign n20043 = n18958 ^ n17106 ^ 1'b0 ;
  assign n20044 = n603 ^ x238 ^ 1'b0 ;
  assign n20045 = n6310 & n20044 ;
  assign n20046 = n6807 & ~n20045 ;
  assign n20048 = n15148 ^ n961 ^ 1'b0 ;
  assign n20049 = n3556 | n20048 ;
  assign n20047 = n10846 & ~n11455 ;
  assign n20050 = n20049 ^ n20047 ^ n13669 ;
  assign n20051 = n20046 & ~n20050 ;
  assign n20052 = n6015 & n20051 ;
  assign n20053 = n6770 & ~n9264 ;
  assign n20054 = n20053 ^ n19632 ^ 1'b0 ;
  assign n20055 = n1051 & ~n7761 ;
  assign n20056 = n11039 & ~n20055 ;
  assign n20057 = n6339 & n9558 ;
  assign n20058 = n2840 | n13409 ;
  assign n20059 = n20058 ^ n11603 ^ 1'b0 ;
  assign n20060 = ( ~n8546 & n11269 ) | ( ~n8546 & n20059 ) | ( n11269 & n20059 ) ;
  assign n20061 = n5658 | n9075 ;
  assign n20062 = n20061 ^ n10247 ^ 1'b0 ;
  assign n20063 = n20062 ^ n6517 ^ 1'b0 ;
  assign n20064 = n14600 ^ n2123 ^ 1'b0 ;
  assign n20065 = n4464 & n20064 ;
  assign n20066 = n20065 ^ n13981 ^ 1'b0 ;
  assign n20067 = n20066 ^ n10811 ^ 1'b0 ;
  assign n20068 = ( n6699 & n7975 ) | ( n6699 & ~n20067 ) | ( n7975 & ~n20067 ) ;
  assign n20069 = n15854 ^ n14164 ^ n1840 ;
  assign n20070 = n1200 & n10923 ;
  assign n20071 = n4832 | n10303 ;
  assign n20072 = n15838 & ~n20071 ;
  assign n20073 = n1145 & ~n20072 ;
  assign n20074 = n20073 ^ n12440 ^ 1'b0 ;
  assign n20075 = n5883 & n14595 ;
  assign n20076 = ( n2275 & ~n10425 ) | ( n2275 & n20075 ) | ( ~n10425 & n20075 ) ;
  assign n20077 = n17123 & n20076 ;
  assign n20078 = ~n20074 & n20077 ;
  assign n20079 = ~n4207 & n19973 ;
  assign n20080 = n18487 & n20079 ;
  assign n20081 = n17778 ^ n17254 ^ 1'b0 ;
  assign n20082 = n19416 ^ n1592 ^ 1'b0 ;
  assign n20083 = n9176 & n20082 ;
  assign n20084 = ( n6087 & ~n14068 ) | ( n6087 & n20083 ) | ( ~n14068 & n20083 ) ;
  assign n20085 = n3259 & n12314 ;
  assign n20086 = n5613 ^ n2408 ^ 1'b0 ;
  assign n20087 = n10757 | n14563 ;
  assign n20088 = n12460 | n20087 ;
  assign n20089 = n20088 ^ n3475 ^ 1'b0 ;
  assign n20090 = n20086 & ~n20089 ;
  assign n20091 = ~n2421 & n2997 ;
  assign n20092 = n7519 | n15112 ;
  assign n20093 = n20091 & ~n20092 ;
  assign n20094 = ( n1713 & n6300 ) | ( n1713 & ~n14226 ) | ( n6300 & ~n14226 ) ;
  assign n20095 = n3873 & ~n4423 ;
  assign n20096 = n20095 ^ n8030 ^ 1'b0 ;
  assign n20097 = n8544 ^ n2900 ^ n559 ;
  assign n20098 = n1870 | n20097 ;
  assign n20099 = n20098 ^ n8403 ^ 1'b0 ;
  assign n20100 = ~n9562 & n20099 ;
  assign n20101 = ~n14793 & n20100 ;
  assign n20102 = ~n6066 & n10982 ;
  assign n20103 = ( n4700 & n6047 ) | ( n4700 & n20102 ) | ( n6047 & n20102 ) ;
  assign n20104 = n3373 ^ n498 ^ 1'b0 ;
  assign n20105 = n20104 ^ n15661 ^ 1'b0 ;
  assign n20106 = x243 & n4100 ;
  assign n20107 = n7408 & n20106 ;
  assign n20108 = n20107 ^ n4544 ^ 1'b0 ;
  assign n20109 = n11942 | n20108 ;
  assign n20110 = n14805 & ~n20109 ;
  assign n20111 = ~n6686 & n17944 ;
  assign n20112 = n5987 & n20111 ;
  assign n20113 = n18588 ^ n8110 ^ 1'b0 ;
  assign n20114 = n13620 & n20113 ;
  assign n20115 = n8590 ^ n1432 ^ 1'b0 ;
  assign n20116 = n20115 ^ n5148 ^ 1'b0 ;
  assign n20120 = n3203 ^ n1450 ^ 1'b0 ;
  assign n20117 = ( n1257 & ~n4228 ) | ( n1257 & n5859 ) | ( ~n4228 & n5859 ) ;
  assign n20118 = n1943 & ~n20117 ;
  assign n20119 = n13099 & n20118 ;
  assign n20121 = n20120 ^ n20119 ^ 1'b0 ;
  assign n20122 = n1446 | n8605 ;
  assign n20123 = n20122 ^ n19363 ^ 1'b0 ;
  assign n20124 = n13261 & n20123 ;
  assign n20125 = ( ~n9799 & n12616 ) | ( ~n9799 & n16516 ) | ( n12616 & n16516 ) ;
  assign n20126 = ~n2263 & n8092 ;
  assign n20127 = ~n20125 & n20126 ;
  assign n20128 = n350 & ~n8456 ;
  assign n20129 = ~n7710 & n20128 ;
  assign n20130 = n20129 ^ n10757 ^ x218 ;
  assign n20131 = n10553 ^ n1149 ^ 1'b0 ;
  assign n20132 = n20131 ^ n7895 ^ n451 ;
  assign n20133 = ~n1168 & n5317 ;
  assign n20134 = n943 & n20133 ;
  assign n20135 = n14357 & n20134 ;
  assign n20136 = n20135 ^ n13597 ^ n9040 ;
  assign n20137 = n17346 ^ n4833 ^ n3949 ;
  assign n20138 = n20137 ^ n2334 ^ n2092 ;
  assign n20139 = n2407 ^ n1374 ^ 1'b0 ;
  assign n20140 = n20139 ^ n16892 ^ 1'b0 ;
  assign n20141 = ( ~n2882 & n4086 ) | ( ~n2882 & n4479 ) | ( n4086 & n4479 ) ;
  assign n20142 = n20141 ^ n1260 ^ 1'b0 ;
  assign n20143 = n12026 & ~n20142 ;
  assign n20144 = n1600 | n6976 ;
  assign n20145 = ~n15107 & n20144 ;
  assign n20146 = n20145 ^ n4212 ^ n2647 ;
  assign n20147 = n5760 & n9676 ;
  assign n20148 = ~n20146 & n20147 ;
  assign n20149 = n20143 & ~n20148 ;
  assign n20150 = n18201 & ~n20149 ;
  assign n20151 = ~n13236 & n20150 ;
  assign n20152 = n14436 ^ n5473 ^ n5242 ;
  assign n20153 = n6387 ^ n1776 ^ 1'b0 ;
  assign n20154 = n18672 ^ n6649 ^ n3100 ;
  assign n20155 = ( n3556 & n5076 ) | ( n3556 & ~n6386 ) | ( n5076 & ~n6386 ) ;
  assign n20156 = n20154 & ~n20155 ;
  assign n20157 = ~n6253 & n10557 ;
  assign n20158 = n7165 | n20157 ;
  assign n20159 = n15382 | n20158 ;
  assign n20160 = n20159 ^ n17680 ^ 1'b0 ;
  assign n20162 = n19853 ^ n3745 ^ n909 ;
  assign n20161 = ~n1286 & n20040 ;
  assign n20163 = n20162 ^ n20161 ^ 1'b0 ;
  assign n20164 = ( n1987 & n2188 ) | ( n1987 & ~n18043 ) | ( n2188 & ~n18043 ) ;
  assign n20168 = n6073 ^ n5816 ^ 1'b0 ;
  assign n20166 = ( n8043 & n16898 ) | ( n8043 & ~n18347 ) | ( n16898 & ~n18347 ) ;
  assign n20165 = n3708 & n7559 ;
  assign n20167 = n20166 ^ n20165 ^ 1'b0 ;
  assign n20169 = n20168 ^ n20167 ^ 1'b0 ;
  assign n20170 = ~n6589 & n20169 ;
  assign n20171 = ( n292 & ~n20164 ) | ( n292 & n20170 ) | ( ~n20164 & n20170 ) ;
  assign n20172 = n3308 ^ n1711 ^ 1'b0 ;
  assign n20173 = ( n1409 & n2626 ) | ( n1409 & n20172 ) | ( n2626 & n20172 ) ;
  assign n20174 = ( x110 & ~n9631 ) | ( x110 & n20173 ) | ( ~n9631 & n20173 ) ;
  assign n20175 = n16422 | n20174 ;
  assign n20176 = n20175 ^ n14768 ^ 1'b0 ;
  assign n20177 = n10034 | n11800 ;
  assign n20178 = n20177 ^ n11045 ^ 1'b0 ;
  assign n20179 = n19618 ^ n10671 ^ 1'b0 ;
  assign n20180 = n10442 & ~n20179 ;
  assign n20181 = n20180 ^ n16899 ^ 1'b0 ;
  assign n20182 = n5994 & ~n20181 ;
  assign n20184 = n4591 ^ n2817 ^ n1103 ;
  assign n20185 = n20184 ^ n13439 ^ n10283 ;
  assign n20186 = ~n7915 & n20185 ;
  assign n20183 = ~n10614 & n11444 ;
  assign n20187 = n20186 ^ n20183 ^ 1'b0 ;
  assign n20188 = n6308 & n20187 ;
  assign n20189 = ~n20182 & n20188 ;
  assign n20190 = n12809 ^ n5263 ^ 1'b0 ;
  assign n20193 = ( ~n7390 & n8624 ) | ( ~n7390 & n10208 ) | ( n8624 & n10208 ) ;
  assign n20191 = n19018 & ~n19873 ;
  assign n20192 = n20191 ^ n16335 ^ 1'b0 ;
  assign n20194 = n20193 ^ n20192 ^ x183 ;
  assign n20195 = n7521 | n15808 ;
  assign n20196 = n20195 ^ n5296 ^ 1'b0 ;
  assign n20197 = ( ~n12032 & n15240 ) | ( ~n12032 & n20196 ) | ( n15240 & n20196 ) ;
  assign n20203 = n2824 & ~n8362 ;
  assign n20204 = ~n14289 & n14951 ;
  assign n20205 = ~n20203 & n20204 ;
  assign n20198 = n688 ^ n356 ^ 1'b0 ;
  assign n20199 = n2001 | n20198 ;
  assign n20200 = n20199 ^ n3047 ^ n841 ;
  assign n20201 = ~n9631 & n20200 ;
  assign n20202 = n17050 & ~n20201 ;
  assign n20206 = n20205 ^ n20202 ^ 1'b0 ;
  assign n20207 = n8424 ^ n7488 ^ 1'b0 ;
  assign n20208 = n14496 & n17946 ;
  assign n20209 = n18629 ^ n5361 ^ 1'b0 ;
  assign n20210 = ~n6728 & n20209 ;
  assign n20211 = n2220 & ~n15250 ;
  assign n20221 = ~n8965 & n11891 ;
  assign n20219 = n4840 ^ x243 ^ 1'b0 ;
  assign n20216 = ~x151 & n17795 ;
  assign n20212 = ( n8223 & n12340 ) | ( n8223 & n16073 ) | ( n12340 & n16073 ) ;
  assign n20213 = n20212 ^ n7740 ^ 1'b0 ;
  assign n20214 = n11197 ^ n1698 ^ 1'b0 ;
  assign n20215 = n20213 & ~n20214 ;
  assign n20217 = n20216 ^ n20215 ^ 1'b0 ;
  assign n20218 = ~n15704 & n20217 ;
  assign n20220 = n20219 ^ n20218 ^ 1'b0 ;
  assign n20222 = n20221 ^ n20220 ^ 1'b0 ;
  assign n20223 = ( n1383 & n9734 ) | ( n1383 & ~n20193 ) | ( n9734 & ~n20193 ) ;
  assign n20224 = ( ~n6371 & n9058 ) | ( ~n6371 & n9785 ) | ( n9058 & n9785 ) ;
  assign n20225 = n4076 & ~n8923 ;
  assign n20226 = n20225 ^ n8693 ^ 1'b0 ;
  assign n20227 = ( n12378 & n20224 ) | ( n12378 & ~n20226 ) | ( n20224 & ~n20226 ) ;
  assign n20228 = n3605 ^ x219 ^ 1'b0 ;
  assign n20229 = n3304 | n20228 ;
  assign n20230 = n20229 ^ n6573 ^ 1'b0 ;
  assign n20232 = ~n3473 & n16603 ;
  assign n20233 = n20232 ^ n4108 ^ 1'b0 ;
  assign n20234 = n20233 ^ n4473 ^ 1'b0 ;
  assign n20235 = n17490 | n20234 ;
  assign n20231 = ~n619 & n3422 ;
  assign n20236 = n20235 ^ n20231 ^ 1'b0 ;
  assign n20237 = n9756 ^ n4698 ^ 1'b0 ;
  assign n20238 = n6483 | n18635 ;
  assign n20239 = ( n5274 & n13003 ) | ( n5274 & n20238 ) | ( n13003 & n20238 ) ;
  assign n20240 = n20239 ^ n3581 ^ 1'b0 ;
  assign n20241 = ( n5440 & ~n20237 ) | ( n5440 & n20240 ) | ( ~n20237 & n20240 ) ;
  assign n20242 = ( n5197 & ~n19414 ) | ( n5197 & n20241 ) | ( ~n19414 & n20241 ) ;
  assign n20243 = ~n15338 & n17112 ;
  assign n20244 = n20243 ^ n6462 ^ 1'b0 ;
  assign n20245 = n8363 & ~n20244 ;
  assign n20246 = n18241 ^ n9564 ^ 1'b0 ;
  assign n20247 = n686 | n4555 ;
  assign n20248 = n20247 ^ n3915 ^ 1'b0 ;
  assign n20249 = n20248 ^ n13301 ^ 1'b0 ;
  assign n20250 = ~n4909 & n20249 ;
  assign n20251 = n16522 ^ n2548 ^ 1'b0 ;
  assign n20252 = ~n2466 & n20251 ;
  assign n20253 = ~n737 & n10041 ;
  assign n20254 = n20253 ^ n8841 ^ 1'b0 ;
  assign n20255 = n20252 & n20254 ;
  assign n20256 = n11493 & n20255 ;
  assign n20257 = ( n17077 & n20250 ) | ( n17077 & ~n20256 ) | ( n20250 & ~n20256 ) ;
  assign n20258 = n7545 | n12094 ;
  assign n20259 = n20257 | n20258 ;
  assign n20260 = n5464 & ~n9802 ;
  assign n20261 = n20260 ^ n2151 ^ 1'b0 ;
  assign n20262 = ~n10780 & n19295 ;
  assign n20263 = n20262 ^ n2967 ^ 1'b0 ;
  assign n20264 = n10856 & ~n20263 ;
  assign n20265 = ~n7611 & n20264 ;
  assign n20266 = n4699 & ~n9921 ;
  assign n20267 = n20265 & n20266 ;
  assign n20268 = ~n464 & n16811 ;
  assign n20269 = n18936 & n20268 ;
  assign n20275 = n16556 ^ n6245 ^ n3050 ;
  assign n20270 = ~n2724 & n2942 ;
  assign n20271 = ~n5057 & n20270 ;
  assign n20272 = n4180 | n20271 ;
  assign n20273 = n20272 ^ n4019 ^ 1'b0 ;
  assign n20274 = n5458 & ~n20273 ;
  assign n20276 = n20275 ^ n20274 ^ 1'b0 ;
  assign n20277 = n3849 & n20276 ;
  assign n20278 = n1071 & n20277 ;
  assign n20279 = n16400 | n20278 ;
  assign n20280 = n5914 & ~n20279 ;
  assign n20281 = n16433 ^ n7448 ^ 1'b0 ;
  assign n20282 = n17486 & n20281 ;
  assign n20283 = n2005 & ~n4752 ;
  assign n20284 = n20283 ^ n10748 ^ n5546 ;
  assign n20285 = n20284 ^ n18762 ^ 1'b0 ;
  assign n20286 = ~n1882 & n4076 ;
  assign n20287 = n935 & n20286 ;
  assign n20288 = n14539 | n19582 ;
  assign n20289 = n741 | n5049 ;
  assign n20290 = n7381 | n20289 ;
  assign n20291 = n20290 ^ n1653 ^ 1'b0 ;
  assign n20292 = n5988 | n20291 ;
  assign n20293 = n20292 ^ n8670 ^ 1'b0 ;
  assign n20294 = n891 & ~n20293 ;
  assign n20295 = n20294 ^ n2908 ^ 1'b0 ;
  assign n20296 = ( n3546 & ~n16003 ) | ( n3546 & n20295 ) | ( ~n16003 & n20295 ) ;
  assign n20297 = x114 & n9172 ;
  assign n20298 = n20297 ^ n6283 ^ 1'b0 ;
  assign n20299 = n20298 ^ n18372 ^ n3269 ;
  assign n20300 = n9398 ^ n6941 ^ n2352 ;
  assign n20301 = ( ~n4061 & n7698 ) | ( ~n4061 & n20300 ) | ( n7698 & n20300 ) ;
  assign n20302 = n14677 | n14912 ;
  assign n20303 = n20301 & ~n20302 ;
  assign n20305 = n3941 & ~n14576 ;
  assign n20304 = n6827 | n13512 ;
  assign n20306 = n20305 ^ n20304 ^ 1'b0 ;
  assign n20307 = n13557 | n20306 ;
  assign n20308 = ( n12234 & n13370 ) | ( n12234 & ~n16488 ) | ( n13370 & ~n16488 ) ;
  assign n20309 = n7145 & ~n13038 ;
  assign n20310 = n2608 & ~n8253 ;
  assign n20311 = n5873 ^ n5179 ^ 1'b0 ;
  assign n20312 = ~n20310 & n20311 ;
  assign n20313 = n6256 ^ n5263 ^ 1'b0 ;
  assign n20314 = n20313 ^ x131 ^ 1'b0 ;
  assign n20315 = n4982 ^ n2651 ^ 1'b0 ;
  assign n20316 = n12463 ^ n10973 ^ n10957 ;
  assign n20317 = n3471 & ~n20316 ;
  assign n20318 = ~n20315 & n20317 ;
  assign n20319 = n17104 ^ n10287 ^ 1'b0 ;
  assign n20320 = n11861 ^ x132 ^ 1'b0 ;
  assign n20321 = n20319 & n20320 ;
  assign n20322 = n5451 ^ n3518 ^ 1'b0 ;
  assign n20323 = ~n1573 & n20322 ;
  assign n20324 = n20323 ^ n18646 ^ 1'b0 ;
  assign n20331 = ~n8903 & n17753 ;
  assign n20332 = n20331 ^ n9936 ^ 1'b0 ;
  assign n20333 = ~n5928 & n20332 ;
  assign n20334 = n20333 ^ n17056 ^ 1'b0 ;
  assign n20326 = n13861 ^ n7384 ^ 1'b0 ;
  assign n20327 = n5466 | n20326 ;
  assign n20325 = n2307 & n6097 ;
  assign n20328 = n20327 ^ n20325 ^ 1'b0 ;
  assign n20329 = n20328 ^ n5723 ^ 1'b0 ;
  assign n20330 = n11771 & n20329 ;
  assign n20335 = n20334 ^ n20330 ^ 1'b0 ;
  assign n20336 = n18200 ^ n9411 ^ n2287 ;
  assign n20337 = n20336 ^ n7791 ^ 1'b0 ;
  assign n20338 = n16817 ^ n6358 ^ 1'b0 ;
  assign n20339 = n14560 & n20338 ;
  assign n20340 = ( n3672 & n11900 ) | ( n3672 & ~n14804 ) | ( n11900 & ~n14804 ) ;
  assign n20341 = n9184 ^ n5509 ^ 1'b0 ;
  assign n20342 = n2840 | n20341 ;
  assign n20343 = n2193 | n20342 ;
  assign n20344 = n4074 & n20343 ;
  assign n20345 = ~n17981 & n20344 ;
  assign n20346 = n2128 & ~n4162 ;
  assign n20347 = n20346 ^ x69 ^ 1'b0 ;
  assign n20348 = ~n2711 & n20347 ;
  assign n20349 = n20305 ^ n9583 ^ 1'b0 ;
  assign n20350 = n11321 ^ n8664 ^ n317 ;
  assign n20351 = ~n1927 & n3434 ;
  assign n20352 = n20351 ^ n16363 ^ 1'b0 ;
  assign n20353 = ( x43 & n20350 ) | ( x43 & n20352 ) | ( n20350 & n20352 ) ;
  assign n20354 = n3125 | n6640 ;
  assign n20355 = n7852 ^ n3535 ^ n1486 ;
  assign n20356 = n20355 ^ n18760 ^ 1'b0 ;
  assign n20357 = n20354 & n20356 ;
  assign n20358 = n5569 | n12597 ;
  assign n20359 = x173 & ~n20358 ;
  assign n20360 = ~n4080 & n20359 ;
  assign n20361 = n20357 & ~n20360 ;
  assign n20362 = n20361 ^ n6296 ^ 1'b0 ;
  assign n20363 = ( ~n7698 & n20353 ) | ( ~n7698 & n20362 ) | ( n20353 & n20362 ) ;
  assign n20364 = n17367 ^ n8525 ^ n7376 ;
  assign n20365 = n9044 & ~n20364 ;
  assign n20366 = ~n15881 & n20365 ;
  assign n20367 = n8812 ^ n2422 ^ 1'b0 ;
  assign n20368 = n16728 ^ n14063 ^ n3510 ;
  assign n20369 = n10348 ^ n7077 ^ n1844 ;
  assign n20370 = n17828 & n20369 ;
  assign n20371 = n20370 ^ n16638 ^ 1'b0 ;
  assign n20372 = n10181 | n14803 ;
  assign n20373 = n20372 ^ n13189 ^ 1'b0 ;
  assign n20374 = n7632 ^ n4783 ^ 1'b0 ;
  assign n20375 = n17000 | n20374 ;
  assign n20376 = ( x139 & ~n1399 ) | ( x139 & n1448 ) | ( ~n1399 & n1448 ) ;
  assign n20377 = n3739 & n3928 ;
  assign n20378 = n20377 ^ n773 ^ 1'b0 ;
  assign n20379 = n20378 ^ n15080 ^ n3169 ;
  assign n20380 = n20379 ^ n1496 ^ 1'b0 ;
  assign n20381 = n11426 & n13249 ;
  assign n20382 = n569 & ~n3904 ;
  assign n20383 = n2157 & ~n5784 ;
  assign n20384 = ~n1194 & n20383 ;
  assign n20385 = ( x187 & n20382 ) | ( x187 & n20384 ) | ( n20382 & n20384 ) ;
  assign n20386 = n7689 & ~n8707 ;
  assign n20387 = n13968 & n20386 ;
  assign n20388 = n9447 ^ n9164 ^ 1'b0 ;
  assign n20389 = n3475 | n20388 ;
  assign n20390 = n19156 ^ n9346 ^ 1'b0 ;
  assign n20391 = ~n20389 & n20390 ;
  assign n20392 = n5674 & ~n13511 ;
  assign n20393 = n20392 ^ n16499 ^ 1'b0 ;
  assign n20394 = n5760 & n16756 ;
  assign n20395 = ~n9189 & n20394 ;
  assign n20396 = n16645 | n17029 ;
  assign n20397 = n9234 | n20396 ;
  assign n20398 = n15547 ^ n8025 ^ 1'b0 ;
  assign n20399 = n780 | n20398 ;
  assign n20400 = n17732 | n20399 ;
  assign n20401 = n20400 ^ n13474 ^ 1'b0 ;
  assign n20403 = n10067 ^ n7634 ^ n3208 ;
  assign n20402 = ( n3309 & ~n8924 ) | ( n3309 & n10124 ) | ( ~n8924 & n10124 ) ;
  assign n20404 = n20403 ^ n20402 ^ 1'b0 ;
  assign n20405 = n14266 | n20404 ;
  assign n20406 = n20405 ^ n10181 ^ 1'b0 ;
  assign n20407 = ~n10317 & n14704 ;
  assign n20408 = n20407 ^ n3621 ^ 1'b0 ;
  assign n20409 = n9581 ^ n1203 ^ 1'b0 ;
  assign n20410 = n11010 & ~n20409 ;
  assign n20411 = n20283 & n20410 ;
  assign n20412 = n20408 & n20411 ;
  assign n20413 = n9173 | n20412 ;
  assign n20414 = n14637 & ~n20413 ;
  assign n20415 = n20414 ^ n2284 ^ 1'b0 ;
  assign n20416 = n7047 & n20415 ;
  assign n20417 = n14328 & n20416 ;
  assign n20418 = n20417 ^ n19612 ^ 1'b0 ;
  assign n20419 = n9346 & ~n9512 ;
  assign n20420 = n11793 & n20419 ;
  assign n20421 = ( n2314 & n10784 ) | ( n2314 & n15202 ) | ( n10784 & n15202 ) ;
  assign n20422 = n20421 ^ n9637 ^ n8231 ;
  assign n20423 = n4308 & n6647 ;
  assign n20424 = n20423 ^ n6119 ^ 1'b0 ;
  assign n20425 = ~n14822 & n20424 ;
  assign n20426 = n13437 ^ n4686 ^ 1'b0 ;
  assign n20427 = ~n7503 & n20426 ;
  assign n20428 = ~n1133 & n20427 ;
  assign n20429 = n13961 & n20428 ;
  assign n20430 = n13869 ^ n10507 ^ n405 ;
  assign n20431 = n7400 & n20430 ;
  assign n20436 = n7252 & ~n11293 ;
  assign n20432 = n18026 ^ n18008 ^ n14147 ;
  assign n20433 = ( n5458 & ~n11998 ) | ( n5458 & n14781 ) | ( ~n11998 & n14781 ) ;
  assign n20434 = n12400 & n20433 ;
  assign n20435 = ~n20432 & n20434 ;
  assign n20437 = n20436 ^ n20435 ^ 1'b0 ;
  assign n20438 = n4158 | n6247 ;
  assign n20439 = n20438 ^ n14938 ^ n2179 ;
  assign n20440 = n13716 ^ n9332 ^ 1'b0 ;
  assign n20441 = n11921 ^ n10194 ^ 1'b0 ;
  assign n20442 = n6113 & n20441 ;
  assign n20443 = n18576 ^ n3110 ^ 1'b0 ;
  assign n20444 = n14481 ^ n4501 ^ 1'b0 ;
  assign n20445 = ( n13648 & n20443 ) | ( n13648 & n20444 ) | ( n20443 & n20444 ) ;
  assign n20446 = n10152 ^ n6562 ^ 1'b0 ;
  assign n20447 = n4280 ^ n1723 ^ 1'b0 ;
  assign n20448 = n20446 & ~n20447 ;
  assign n20449 = n20448 ^ n12902 ^ n7409 ;
  assign n20450 = n20449 ^ n10839 ^ 1'b0 ;
  assign n20451 = n20450 ^ n8492 ^ 1'b0 ;
  assign n20452 = ~n15239 & n20451 ;
  assign n20453 = ( n1322 & n3185 ) | ( n1322 & ~n17082 ) | ( n3185 & ~n17082 ) ;
  assign n20454 = ~n10742 & n20453 ;
  assign n20455 = n20454 ^ n16461 ^ 1'b0 ;
  assign n20456 = ( n1074 & ~n7302 ) | ( n1074 & n20455 ) | ( ~n7302 & n20455 ) ;
  assign n20457 = n20456 ^ n6395 ^ 1'b0 ;
  assign n20458 = n8006 & n20457 ;
  assign n20459 = n7273 ^ n4298 ^ 1'b0 ;
  assign n20460 = ~n7637 & n20459 ;
  assign n20463 = n5195 | n19785 ;
  assign n20464 = n4411 & n20463 ;
  assign n20465 = n20464 ^ n11747 ^ 1'b0 ;
  assign n20461 = n7231 & ~n11691 ;
  assign n20462 = n474 | n20461 ;
  assign n20466 = n20465 ^ n20462 ^ n12370 ;
  assign n20467 = n12670 & n20466 ;
  assign n20468 = n14225 ^ n4940 ^ 1'b0 ;
  assign n20469 = n4426 & n20468 ;
  assign n20470 = n2875 ^ n2816 ^ 1'b0 ;
  assign n20471 = ~n5353 & n20470 ;
  assign n20472 = ~n7912 & n20471 ;
  assign n20473 = ~n3152 & n20472 ;
  assign n20474 = x59 & n20473 ;
  assign n20475 = n12463 ^ n802 ^ n396 ;
  assign n20476 = n9666 ^ n6250 ^ n2912 ;
  assign n20478 = n15219 ^ n1793 ^ 1'b0 ;
  assign n20479 = n743 & ~n20478 ;
  assign n20480 = ( ~n8104 & n15260 ) | ( ~n8104 & n20479 ) | ( n15260 & n20479 ) ;
  assign n20477 = n1651 | n13424 ;
  assign n20481 = n20480 ^ n20477 ^ n20257 ;
  assign n20482 = n3698 & ~n19726 ;
  assign n20483 = ~n1398 & n20482 ;
  assign n20484 = n18661 ^ n5115 ^ n4350 ;
  assign n20485 = ~n13200 & n13273 ;
  assign n20486 = ~n495 & n20485 ;
  assign n20487 = n20486 ^ n7819 ^ n4112 ;
  assign n20488 = n11490 ^ n729 ^ 1'b0 ;
  assign n20489 = n789 & ~n20488 ;
  assign n20490 = ~n2985 & n10342 ;
  assign n20491 = n17420 | n20490 ;
  assign n20492 = n16621 ^ n1962 ^ 1'b0 ;
  assign n20495 = n17602 ^ x124 ^ 1'b0 ;
  assign n20496 = n828 & ~n20495 ;
  assign n20497 = n20496 ^ n2759 ^ 1'b0 ;
  assign n20493 = n4552 | n7553 ;
  assign n20494 = n20493 ^ n10801 ^ n4689 ;
  assign n20498 = n20497 ^ n20494 ^ n17900 ;
  assign n20499 = n13670 ^ n5183 ^ n3256 ;
  assign n20500 = n20499 ^ n5500 ^ 1'b0 ;
  assign n20505 = n14067 ^ n11530 ^ n9538 ;
  assign n20501 = n7530 ^ n1630 ^ 1'b0 ;
  assign n20502 = n20501 ^ n1228 ^ 1'b0 ;
  assign n20503 = n4206 & n20502 ;
  assign n20504 = n20503 ^ n15603 ^ 1'b0 ;
  assign n20506 = n20505 ^ n20504 ^ n11502 ;
  assign n20507 = x141 & n19428 ;
  assign n20508 = n5454 & n20507 ;
  assign n20509 = ( ~n5696 & n15058 ) | ( ~n5696 & n20508 ) | ( n15058 & n20508 ) ;
  assign n20519 = n3543 & ~n17653 ;
  assign n20510 = ~n6471 & n8003 ;
  assign n20512 = n1620 & ~n2824 ;
  assign n20511 = ~n3854 & n3984 ;
  assign n20513 = n20512 ^ n20511 ^ 1'b0 ;
  assign n20514 = n4072 & ~n20513 ;
  assign n20515 = n3989 & n20514 ;
  assign n20516 = n1434 | n20515 ;
  assign n20517 = n5834 | n20516 ;
  assign n20518 = ( n4388 & ~n20510 ) | ( n4388 & n20517 ) | ( ~n20510 & n20517 ) ;
  assign n20520 = n20519 ^ n20518 ^ n10509 ;
  assign n20521 = ( n1415 & n4893 ) | ( n1415 & n11636 ) | ( n4893 & n11636 ) ;
  assign n20522 = n14487 ^ n13359 ^ 1'b0 ;
  assign n20523 = n20521 | n20522 ;
  assign n20524 = n902 ^ n445 ^ 1'b0 ;
  assign n20525 = n1088 ^ x138 ^ 1'b0 ;
  assign n20526 = n20524 | n20525 ;
  assign n20527 = ~n2560 & n4553 ;
  assign n20528 = n20526 & n20527 ;
  assign n20529 = n351 | n8181 ;
  assign n20530 = n2369 | n20529 ;
  assign n20531 = n15893 ^ n8644 ^ 1'b0 ;
  assign n20532 = n20531 ^ n16473 ^ n10757 ;
  assign n20533 = x99 | n14818 ;
  assign n20535 = n4111 & n4385 ;
  assign n20536 = n16051 | n20535 ;
  assign n20537 = n19241 | n20536 ;
  assign n20538 = n20537 ^ n807 ^ 1'b0 ;
  assign n20534 = ~n6001 & n11565 ;
  assign n20539 = n20538 ^ n20534 ^ 1'b0 ;
  assign n20540 = x107 & n1843 ;
  assign n20541 = n20540 ^ n14988 ^ n14125 ;
  assign n20542 = ( n2697 & n5037 ) | ( n2697 & ~n6611 ) | ( n5037 & ~n6611 ) ;
  assign n20543 = n580 & n20542 ;
  assign n20544 = n2068 & ~n8475 ;
  assign n20545 = n8678 & n20544 ;
  assign n20546 = n12059 ^ n11873 ^ n5234 ;
  assign n20547 = n3568 | n20546 ;
  assign n20548 = n10216 | n15385 ;
  assign n20549 = ( ~n6772 & n15750 ) | ( ~n6772 & n20548 ) | ( n15750 & n20548 ) ;
  assign n20550 = n20549 ^ n15630 ^ n1028 ;
  assign n20551 = n12995 ^ n7195 ^ 1'b0 ;
  assign n20552 = n4959 & n20551 ;
  assign n20563 = n7692 ^ n3091 ^ 1'b0 ;
  assign n20564 = n3995 & ~n20563 ;
  assign n20553 = ( n4953 & n10064 ) | ( n4953 & ~n15704 ) | ( n10064 & ~n15704 ) ;
  assign n20554 = n4048 & n8937 ;
  assign n20555 = n20554 ^ n955 ^ 1'b0 ;
  assign n20556 = n5520 | n20555 ;
  assign n20557 = n10816 | n19258 ;
  assign n20558 = n20557 ^ n1389 ^ 1'b0 ;
  assign n20559 = ~n2162 & n20558 ;
  assign n20560 = n20559 ^ n9803 ^ 1'b0 ;
  assign n20561 = n20556 & n20560 ;
  assign n20562 = n20553 & n20561 ;
  assign n20565 = n20564 ^ n20562 ^ 1'b0 ;
  assign n20566 = ( n3409 & n7678 ) | ( n3409 & ~n7927 ) | ( n7678 & ~n7927 ) ;
  assign n20567 = n20566 ^ n10799 ^ 1'b0 ;
  assign n20568 = n13850 | n14951 ;
  assign n20569 = n20568 ^ n12398 ^ n1383 ;
  assign n20570 = ( ~n4093 & n20567 ) | ( ~n4093 & n20569 ) | ( n20567 & n20569 ) ;
  assign n20571 = n13736 ^ n5536 ^ 1'b0 ;
  assign n20572 = n11589 ^ n11293 ^ n2351 ;
  assign n20573 = n9136 & n20572 ;
  assign n20574 = n20573 ^ n9576 ^ 1'b0 ;
  assign n20575 = n19108 & ~n20574 ;
  assign n20576 = ( x183 & ~n4501 ) | ( x183 & n11871 ) | ( ~n4501 & n11871 ) ;
  assign n20577 = n13102 & ~n18292 ;
  assign n20578 = n7136 | n7265 ;
  assign n20579 = n6689 | n18435 ;
  assign n20580 = n20579 ^ n845 ^ 1'b0 ;
  assign n20581 = n13952 | n20580 ;
  assign n20582 = n20581 ^ n368 ^ 1'b0 ;
  assign n20583 = n4157 ^ n1512 ^ 1'b0 ;
  assign n20584 = n3688 & n20583 ;
  assign n20585 = n20584 ^ n7643 ^ n1787 ;
  assign n20586 = n20585 ^ n12483 ^ 1'b0 ;
  assign n20587 = ~n2164 & n20586 ;
  assign n20588 = ~n5104 & n9044 ;
  assign n20589 = n20588 ^ n6725 ^ 1'b0 ;
  assign n20590 = n3244 & n20589 ;
  assign n20591 = n5430 ^ x173 ^ 1'b0 ;
  assign n20592 = n12883 | n20591 ;
  assign n20593 = n11252 & n20592 ;
  assign n20594 = n6612 ^ n580 ^ 1'b0 ;
  assign n20595 = n4604 & ~n13443 ;
  assign n20596 = ( n1851 & ~n3410 ) | ( n1851 & n5795 ) | ( ~n3410 & n5795 ) ;
  assign n20597 = n20596 ^ n8980 ^ 1'b0 ;
  assign n20598 = n20597 ^ n12140 ^ 1'b0 ;
  assign n20600 = n15316 & ~n18876 ;
  assign n20601 = n20600 ^ n12408 ^ 1'b0 ;
  assign n20599 = n2319 & n5793 ;
  assign n20602 = n20601 ^ n20599 ^ 1'b0 ;
  assign n20604 = n13050 ^ n5815 ^ 1'b0 ;
  assign n20605 = ~n2209 & n20604 ;
  assign n20606 = n20605 ^ n11019 ^ 1'b0 ;
  assign n20603 = n12587 ^ n874 ^ 1'b0 ;
  assign n20607 = n20606 ^ n20603 ^ 1'b0 ;
  assign n20608 = n1183 & ~n2680 ;
  assign n20609 = n11409 & n20608 ;
  assign n20610 = ( n12252 & n17047 ) | ( n12252 & n20609 ) | ( n17047 & n20609 ) ;
  assign n20611 = n20610 ^ n7831 ^ 1'b0 ;
  assign n20612 = n6307 ^ n5859 ^ 1'b0 ;
  assign n20613 = n10002 & n20612 ;
  assign n20614 = n20613 ^ n12839 ^ n6917 ;
  assign n20615 = ( ~n4397 & n7840 ) | ( ~n4397 & n20614 ) | ( n7840 & n20614 ) ;
  assign n20616 = n9386 | n12923 ;
  assign n20617 = ( n1031 & n5552 ) | ( n1031 & n20616 ) | ( n5552 & n20616 ) ;
  assign n20618 = ( n1267 & n10119 ) | ( n1267 & ~n16213 ) | ( n10119 & ~n16213 ) ;
  assign n20619 = n1406 | n20618 ;
  assign n20620 = n20617 | n20619 ;
  assign n20621 = n3086 & ~n10584 ;
  assign n20622 = n4874 & ~n19334 ;
  assign n20623 = ~n15635 & n20622 ;
  assign n20624 = n4422 ^ n1751 ^ 1'b0 ;
  assign n20625 = n701 & ~n20624 ;
  assign n20626 = n13830 | n18041 ;
  assign n20627 = ( n7934 & ~n20625 ) | ( n7934 & n20626 ) | ( ~n20625 & n20626 ) ;
  assign n20630 = n16860 ^ n9325 ^ 1'b0 ;
  assign n20628 = n17587 ^ n6757 ^ 1'b0 ;
  assign n20629 = ~n1021 & n20628 ;
  assign n20631 = n20630 ^ n20629 ^ n5020 ;
  assign n20632 = n13922 & n20631 ;
  assign n20640 = n14593 ^ n5737 ^ n2680 ;
  assign n20641 = n20640 ^ n1050 ^ x220 ;
  assign n20633 = ~n8548 & n11068 ;
  assign n20634 = n10636 & n20633 ;
  assign n20635 = n20634 ^ n9751 ^ n4756 ;
  assign n20636 = n1774 | n3575 ;
  assign n20637 = n20636 ^ n12207 ^ n2548 ;
  assign n20638 = n20635 & n20637 ;
  assign n20639 = n20638 ^ n6124 ^ 1'b0 ;
  assign n20642 = n20641 ^ n20639 ^ n9799 ;
  assign n20643 = n16436 ^ n8079 ^ n7850 ;
  assign n20644 = n9143 ^ n8096 ^ 1'b0 ;
  assign n20645 = n14516 & n20644 ;
  assign n20646 = n20645 ^ n11306 ^ 1'b0 ;
  assign n20647 = n11587 | n20646 ;
  assign n20648 = ~n686 & n19688 ;
  assign n20649 = n20648 ^ n19795 ^ n9299 ;
  assign n20650 = n3238 ^ x34 ^ 1'b0 ;
  assign n20651 = n20650 ^ n10105 ^ n6266 ;
  assign n20652 = n20651 ^ n6028 ^ n4700 ;
  assign n20654 = n3945 ^ n507 ^ 1'b0 ;
  assign n20653 = n1941 & n11119 ;
  assign n20655 = n20654 ^ n20653 ^ 1'b0 ;
  assign n20656 = n20655 ^ n4182 ^ n741 ;
  assign n20657 = n6018 ^ n513 ^ 1'b0 ;
  assign n20658 = n17772 & ~n20657 ;
  assign n20663 = n1602 | n9997 ;
  assign n20664 = n5830 & ~n20663 ;
  assign n20665 = ~n16242 & n20664 ;
  assign n20659 = ( ~n5201 & n8148 ) | ( ~n5201 & n14389 ) | ( n8148 & n14389 ) ;
  assign n20660 = n2383 | n5027 ;
  assign n20661 = n20660 ^ n518 ^ 1'b0 ;
  assign n20662 = ~n20659 & n20661 ;
  assign n20666 = n20665 ^ n20662 ^ 1'b0 ;
  assign n20667 = n10847 ^ n6618 ^ 1'b0 ;
  assign n20668 = n2456 & ~n20667 ;
  assign n20670 = n4376 ^ n4059 ^ 1'b0 ;
  assign n20671 = n6563 & n20670 ;
  assign n20669 = n11028 | n13331 ;
  assign n20672 = n20671 ^ n20669 ^ n18134 ;
  assign n20673 = ~n14335 & n20672 ;
  assign n20674 = ~n9874 & n20673 ;
  assign n20675 = n20674 ^ n7566 ^ 1'b0 ;
  assign n20676 = n20668 & ~n20675 ;
  assign n20677 = ~n6130 & n11251 ;
  assign n20678 = n20677 ^ n12977 ^ 1'b0 ;
  assign n20679 = n638 | n20678 ;
  assign n20680 = n20679 ^ n15404 ^ 1'b0 ;
  assign n20681 = n9099 & n20680 ;
  assign n20683 = n2886 & ~n14911 ;
  assign n20682 = n2266 & ~n11913 ;
  assign n20684 = n20683 ^ n20682 ^ 1'b0 ;
  assign n20685 = n8199 | n11020 ;
  assign n20686 = n5077 & ~n20685 ;
  assign n20687 = n14497 | n20686 ;
  assign n20692 = n2321 & ~n18552 ;
  assign n20693 = ~n5123 & n20692 ;
  assign n20694 = n20693 ^ n3674 ^ 1'b0 ;
  assign n20689 = n10075 & ~n15526 ;
  assign n20690 = n20689 ^ n10909 ^ 1'b0 ;
  assign n20688 = n13297 ^ n2340 ^ 1'b0 ;
  assign n20691 = n20690 ^ n20688 ^ n6810 ;
  assign n20695 = n20694 ^ n20691 ^ 1'b0 ;
  assign n20706 = ( n19812 & n20019 ) | ( n19812 & n20097 ) | ( n20019 & n20097 ) ;
  assign n20703 = n6382 ^ x72 ^ 1'b0 ;
  assign n20704 = ~n11190 & n20703 ;
  assign n20705 = n20704 ^ n14940 ^ 1'b0 ;
  assign n20696 = n10432 ^ n5174 ^ n3117 ;
  assign n20697 = n20696 ^ n14789 ^ 1'b0 ;
  assign n20698 = n6430 ^ n5479 ^ 1'b0 ;
  assign n20699 = n10442 & n20698 ;
  assign n20700 = n6050 & n8356 ;
  assign n20701 = n20700 ^ n4214 ^ 1'b0 ;
  assign n20702 = ( n20697 & n20699 ) | ( n20697 & n20701 ) | ( n20699 & n20701 ) ;
  assign n20707 = n20706 ^ n20705 ^ n20702 ;
  assign n20708 = n5975 ^ n4713 ^ 1'b0 ;
  assign n20709 = n2711 & n20708 ;
  assign n20710 = n9030 & ~n11331 ;
  assign n20711 = ~n19857 & n20710 ;
  assign n20712 = n9897 ^ x193 ^ 1'b0 ;
  assign n20713 = n1853 & n20712 ;
  assign n20714 = n20713 ^ n18618 ^ 1'b0 ;
  assign n20715 = ( n4047 & n15348 ) | ( n4047 & n20714 ) | ( n15348 & n20714 ) ;
  assign n20716 = n12483 ^ n12478 ^ 1'b0 ;
  assign n20717 = n20716 ^ n8765 ^ 1'b0 ;
  assign n20718 = ~n12672 & n20717 ;
  assign n20719 = n4881 ^ n3297 ^ 1'b0 ;
  assign n20720 = n19492 ^ n6606 ^ n2567 ;
  assign n20721 = ( n17579 & n20719 ) | ( n17579 & n20720 ) | ( n20719 & n20720 ) ;
  assign n20726 = n1028 & ~n2191 ;
  assign n20722 = n2236 & n11580 ;
  assign n20723 = ( ~n6358 & n10529 ) | ( ~n6358 & n20722 ) | ( n10529 & n20722 ) ;
  assign n20724 = n20723 ^ n9849 ^ n9193 ;
  assign n20725 = n20724 ^ n19916 ^ n8739 ;
  assign n20727 = n20726 ^ n20725 ^ n403 ;
  assign n20728 = n9902 & n20727 ;
  assign n20729 = n20728 ^ n15371 ^ 1'b0 ;
  assign n20730 = ~n5305 & n5877 ;
  assign n20731 = n20730 ^ n515 ^ 1'b0 ;
  assign n20732 = n9408 & n20731 ;
  assign n20733 = n20732 ^ n20645 ^ 1'b0 ;
  assign n20735 = ~n2220 & n4527 ;
  assign n20734 = n4129 & ~n12552 ;
  assign n20736 = n20735 ^ n20734 ^ 1'b0 ;
  assign n20737 = x151 & n2897 ;
  assign n20738 = n4019 | n20737 ;
  assign n20739 = n1538 & ~n20738 ;
  assign n20740 = n20739 ^ n18404 ^ n5245 ;
  assign n20741 = n4670 | n17130 ;
  assign n20742 = n20741 ^ n17118 ^ 1'b0 ;
  assign n20743 = n15912 & ~n20742 ;
  assign n20744 = ~n15959 & n20743 ;
  assign n20745 = n8006 & n12232 ;
  assign n20746 = n15222 & n20745 ;
  assign n20747 = n6376 | n7044 ;
  assign n20748 = n3816 | n17237 ;
  assign n20749 = n20747 | n20748 ;
  assign n20750 = n20749 ^ n1501 ^ x170 ;
  assign n20751 = ( n3961 & n7131 ) | ( n3961 & ~n15893 ) | ( n7131 & ~n15893 ) ;
  assign n20752 = ~n11467 & n20751 ;
  assign n20753 = n4031 | n20752 ;
  assign n20754 = n20753 ^ n394 ^ 1'b0 ;
  assign n20755 = n18842 ^ n3158 ^ n713 ;
  assign n20756 = ~n5446 & n20755 ;
  assign n20757 = n20756 ^ n5318 ^ 1'b0 ;
  assign n20758 = n5860 ^ n3404 ^ 1'b0 ;
  assign n20759 = ~n14694 & n15430 ;
  assign n20760 = n9206 & n20759 ;
  assign n20762 = n12554 ^ n1975 ^ 1'b0 ;
  assign n20763 = n3257 & n20762 ;
  assign n20761 = n4759 | n16874 ;
  assign n20764 = n20763 ^ n20761 ^ 1'b0 ;
  assign n20765 = n6778 | n20556 ;
  assign n20766 = n2727 & ~n20765 ;
  assign n20767 = ~n1090 & n20766 ;
  assign n20768 = n6545 ^ n6256 ^ n2925 ;
  assign n20769 = n2504 ^ n1849 ^ 1'b0 ;
  assign n20770 = n20768 & ~n20769 ;
  assign n20771 = n20770 ^ n9610 ^ 1'b0 ;
  assign n20772 = n1458 & ~n6381 ;
  assign n20773 = ( ~n2005 & n6176 ) | ( ~n2005 & n20772 ) | ( n6176 & n20772 ) ;
  assign n20774 = n20773 ^ n13210 ^ 1'b0 ;
  assign n20775 = n1039 | n20774 ;
  assign n20776 = n20775 ^ n8416 ^ 1'b0 ;
  assign n20777 = n14344 & ~n18963 ;
  assign n20780 = n13261 ^ n9277 ^ 1'b0 ;
  assign n20778 = n2120 ^ x242 ^ 1'b0 ;
  assign n20779 = n13399 & n20778 ;
  assign n20781 = n20780 ^ n20779 ^ 1'b0 ;
  assign n20782 = n17093 | n20781 ;
  assign n20783 = n20782 ^ n13039 ^ 1'b0 ;
  assign n20784 = n2611 ^ n1256 ^ 1'b0 ;
  assign n20785 = n11891 ^ n10036 ^ 1'b0 ;
  assign n20786 = n20785 ^ n4221 ^ 1'b0 ;
  assign n20787 = n10112 ^ n464 ^ 1'b0 ;
  assign n20788 = n14549 | n20787 ;
  assign n20789 = n4849 & ~n20788 ;
  assign n20790 = n14157 & ~n20789 ;
  assign n20791 = n17614 | n20790 ;
  assign n20792 = n20786 & ~n20791 ;
  assign n20797 = n953 | n2287 ;
  assign n20798 = n20797 ^ n8013 ^ 1'b0 ;
  assign n20795 = n1376 & ~n7702 ;
  assign n20796 = n20795 ^ n9115 ^ 1'b0 ;
  assign n20793 = n837 & ~n20159 ;
  assign n20794 = n19031 & n20793 ;
  assign n20799 = n20798 ^ n20796 ^ n20794 ;
  assign n20800 = ( n1389 & n8685 ) | ( n1389 & ~n9967 ) | ( n8685 & ~n9967 ) ;
  assign n20801 = ( n3197 & n14059 ) | ( n3197 & ~n18192 ) | ( n14059 & ~n18192 ) ;
  assign n20802 = n7822 | n20801 ;
  assign n20803 = n1054 & n6794 ;
  assign n20804 = n7599 & n20803 ;
  assign n20807 = n7450 & ~n15519 ;
  assign n20808 = n20807 ^ n11546 ^ 1'b0 ;
  assign n20805 = n1105 | n11422 ;
  assign n20806 = n20805 ^ n5389 ^ 1'b0 ;
  assign n20809 = n20808 ^ n20806 ^ 1'b0 ;
  assign n20810 = n20809 ^ n12469 ^ n2189 ;
  assign n20811 = x125 | n15260 ;
  assign n20812 = n5024 ^ n4277 ^ 1'b0 ;
  assign n20813 = ~n4648 & n20812 ;
  assign n20814 = ~n20495 & n20813 ;
  assign n20815 = ( n8155 & n12115 ) | ( n8155 & n20814 ) | ( n12115 & n20814 ) ;
  assign n20816 = n7075 ^ n5916 ^ 1'b0 ;
  assign n20817 = ~n4809 & n19793 ;
  assign n20818 = ~n716 & n20817 ;
  assign n20819 = n3851 & ~n13668 ;
  assign n20820 = n5662 & n20819 ;
  assign n20821 = n14235 & n20820 ;
  assign n20822 = n1695 ^ n887 ^ 1'b0 ;
  assign n20823 = ~n20821 & n20822 ;
  assign n20824 = n7577 | n8453 ;
  assign n20825 = n20824 ^ n4784 ^ 1'b0 ;
  assign n20826 = n20825 ^ n9598 ^ 1'b0 ;
  assign n20827 = ~n16075 & n20826 ;
  assign n20828 = ~n2463 & n14655 ;
  assign n20829 = n20828 ^ n2317 ^ 1'b0 ;
  assign n20830 = n1741 & n20829 ;
  assign n20831 = n20830 ^ n19244 ^ 1'b0 ;
  assign n20832 = ~n6043 & n20831 ;
  assign n20833 = ~n3459 & n5253 ;
  assign n20834 = ~n14822 & n20833 ;
  assign n20835 = n20834 ^ n11871 ^ 1'b0 ;
  assign n20836 = ( ~n15420 & n17811 ) | ( ~n15420 & n20835 ) | ( n17811 & n20835 ) ;
  assign n20837 = n4959 & n7957 ;
  assign n20838 = n6540 ^ n3877 ^ 1'b0 ;
  assign n20839 = n6543 & n20838 ;
  assign n20840 = n20839 ^ n8264 ^ n6745 ;
  assign n20841 = n16919 ^ n8689 ^ n5419 ;
  assign n20842 = n20840 & ~n20841 ;
  assign n20843 = n20842 ^ n10709 ^ 1'b0 ;
  assign n20844 = ( n10261 & ~n15919 ) | ( n10261 & n20843 ) | ( ~n15919 & n20843 ) ;
  assign n20845 = n20837 & ~n20844 ;
  assign n20846 = ( n2553 & n5751 ) | ( n2553 & ~n17874 ) | ( n5751 & ~n17874 ) ;
  assign n20847 = ( n4203 & ~n10642 ) | ( n4203 & n20846 ) | ( ~n10642 & n20846 ) ;
  assign n20854 = n3950 ^ n3469 ^ 1'b0 ;
  assign n20855 = n14300 | n20854 ;
  assign n20851 = n2733 & n3965 ;
  assign n20852 = n20851 ^ n5648 ^ 1'b0 ;
  assign n20848 = n3700 & ~n4761 ;
  assign n20849 = n20848 ^ n761 ^ 1'b0 ;
  assign n20850 = n20849 ^ n9131 ^ n7552 ;
  assign n20853 = n20852 ^ n20850 ^ n9168 ;
  assign n20856 = n20855 ^ n20853 ^ n19883 ;
  assign n20857 = n658 & ~n2106 ;
  assign n20858 = ~n14158 & n17494 ;
  assign n20859 = ( ~n2607 & n20857 ) | ( ~n2607 & n20858 ) | ( n20857 & n20858 ) ;
  assign n20860 = n12622 ^ n2039 ^ 1'b0 ;
  assign n20861 = n6471 & ~n20860 ;
  assign n20862 = n1341 & ~n20861 ;
  assign n20863 = ~n8258 & n17582 ;
  assign n20872 = ~n8588 & n9520 ;
  assign n20869 = ~n10333 & n15785 ;
  assign n20870 = n20869 ^ n16858 ^ 1'b0 ;
  assign n20868 = n3286 | n20139 ;
  assign n20871 = n20870 ^ n20868 ^ 1'b0 ;
  assign n20873 = n20872 ^ n20871 ^ 1'b0 ;
  assign n20874 = n7347 & ~n20873 ;
  assign n20866 = n15710 ^ n10285 ^ n6080 ;
  assign n20864 = n17513 ^ n10095 ^ 1'b0 ;
  assign n20865 = n20864 ^ n18768 ^ 1'b0 ;
  assign n20867 = n20866 ^ n20865 ^ n18216 ;
  assign n20875 = n20874 ^ n20867 ^ 1'b0 ;
  assign n20876 = ( n2272 & n11300 ) | ( n2272 & n20875 ) | ( n11300 & n20875 ) ;
  assign n20879 = ~n4210 & n11926 ;
  assign n20877 = n10281 & n14241 ;
  assign n20878 = n6127 & n20877 ;
  assign n20880 = n20879 ^ n20878 ^ 1'b0 ;
  assign n20881 = ~n20876 & n20880 ;
  assign n20882 = n17389 & ~n17866 ;
  assign n20883 = n20882 ^ n10681 ^ 1'b0 ;
  assign n20884 = ( n7208 & n12110 ) | ( n7208 & ~n18841 ) | ( n12110 & ~n18841 ) ;
  assign n20885 = n6350 | n7076 ;
  assign n20886 = n7823 | n20885 ;
  assign n20890 = n10832 ^ n5175 ^ 1'b0 ;
  assign n20887 = n3182 & ~n11599 ;
  assign n20888 = n20887 ^ n14974 ^ 1'b0 ;
  assign n20889 = ~n2425 & n20888 ;
  assign n20891 = n20890 ^ n20889 ^ n5509 ;
  assign n20892 = x18 & n9078 ;
  assign n20893 = n14749 & n20892 ;
  assign n20894 = n19415 ^ n16437 ^ 1'b0 ;
  assign n20895 = ( n5978 & ~n11554 ) | ( n5978 & n15910 ) | ( ~n11554 & n15910 ) ;
  assign n20896 = ~n18443 & n20895 ;
  assign n20897 = n20896 ^ n5162 ^ 1'b0 ;
  assign n20898 = n814 | n5139 ;
  assign n20899 = n3245 & n20898 ;
  assign n20900 = n2760 & n10532 ;
  assign n20901 = n589 | n1145 ;
  assign n20902 = ~n2790 & n20901 ;
  assign n20903 = ~n20900 & n20902 ;
  assign n20904 = ( n5099 & n20899 ) | ( n5099 & ~n20903 ) | ( n20899 & ~n20903 ) ;
  assign n20905 = n13714 ^ n9033 ^ 1'b0 ;
  assign n20906 = n20905 ^ n19062 ^ 1'b0 ;
  assign n20907 = n16370 ^ n5213 ^ n4485 ;
  assign n20908 = ( n460 & ~n6783 ) | ( n460 & n12439 ) | ( ~n6783 & n12439 ) ;
  assign n20909 = n17516 ^ n11775 ^ n5162 ;
  assign n20910 = n9630 | n20909 ;
  assign n20911 = n20908 & ~n20910 ;
  assign n20912 = n20911 ^ n931 ^ 1'b0 ;
  assign n20913 = n2363 | n20912 ;
  assign n20914 = n11353 ^ n2671 ^ 1'b0 ;
  assign n20915 = ~n1434 & n20914 ;
  assign n20916 = x94 & ~n8435 ;
  assign n20917 = n20916 ^ n18786 ^ n12929 ;
  assign n20918 = ( n5266 & n9797 ) | ( n5266 & ~n20917 ) | ( n9797 & ~n20917 ) ;
  assign n20919 = ~n5377 & n20918 ;
  assign n20920 = ( n495 & ~n8310 ) | ( n495 & n14334 ) | ( ~n8310 & n14334 ) ;
  assign n20921 = n20920 ^ n6396 ^ 1'b0 ;
  assign n20922 = n20921 ^ n8446 ^ 1'b0 ;
  assign n20923 = ~n6296 & n11759 ;
  assign n20924 = n9664 ^ n4084 ^ n513 ;
  assign n20925 = n20924 ^ n5081 ^ 1'b0 ;
  assign n20926 = n4065 & n15977 ;
  assign n20927 = ( n16930 & n20029 ) | ( n16930 & ~n20926 ) | ( n20029 & ~n20926 ) ;
  assign n20928 = n3540 & n20802 ;
  assign n20929 = n20928 ^ n18045 ^ 1'b0 ;
  assign n20930 = ~n1935 & n2760 ;
  assign n20931 = ~n12671 & n15116 ;
  assign n20932 = n20931 ^ n9122 ^ 1'b0 ;
  assign n20933 = n20158 ^ n15101 ^ 1'b0 ;
  assign n20934 = ( n13998 & ~n17928 ) | ( n13998 & n20933 ) | ( ~n17928 & n20933 ) ;
  assign n20935 = n15415 ^ n7132 ^ 1'b0 ;
  assign n20938 = n17892 ^ n630 ^ 1'b0 ;
  assign n20939 = ( n5513 & n5855 ) | ( n5513 & n20938 ) | ( n5855 & n20938 ) ;
  assign n20936 = ( n11149 & n19731 ) | ( n11149 & n19936 ) | ( n19731 & n19936 ) ;
  assign n20937 = n7769 | n20936 ;
  assign n20940 = n20939 ^ n20937 ^ 1'b0 ;
  assign n20941 = n4197 ^ n2919 ^ 1'b0 ;
  assign n20942 = n20941 ^ n11089 ^ n3549 ;
  assign n20943 = n10753 ^ n7359 ^ 1'b0 ;
  assign n20944 = n7275 ^ n576 ^ 1'b0 ;
  assign n20945 = ~n12648 & n20944 ;
  assign n20946 = n2509 | n20945 ;
  assign n20948 = n15931 ^ x129 ^ 1'b0 ;
  assign n20947 = n9201 & ~n10142 ;
  assign n20949 = n20948 ^ n20947 ^ 1'b0 ;
  assign n20951 = ~n12231 & n19250 ;
  assign n20952 = n20951 ^ n9680 ^ 1'b0 ;
  assign n20950 = n4676 | n9996 ;
  assign n20953 = n20952 ^ n20950 ^ n13396 ;
  assign n20954 = n9210 | n19577 ;
  assign n20955 = n13378 | n20954 ;
  assign n20956 = n4669 & n9068 ;
  assign n20957 = n20956 ^ n9827 ^ 1'b0 ;
  assign n20958 = ~n7120 & n20957 ;
  assign n20959 = n20731 ^ n13545 ^ 1'b0 ;
  assign n20960 = ( n20955 & n20958 ) | ( n20955 & n20959 ) | ( n20958 & n20959 ) ;
  assign n20961 = n6010 | n9238 ;
  assign n20962 = ~n20199 & n20961 ;
  assign n20963 = n20962 ^ n12868 ^ 1'b0 ;
  assign n20967 = n6797 | n16767 ;
  assign n20966 = n13662 ^ n3724 ^ n2189 ;
  assign n20964 = n16845 ^ n3675 ^ 1'b0 ;
  assign n20965 = n11410 & n20964 ;
  assign n20968 = n20967 ^ n20966 ^ n20965 ;
  assign n20969 = n6720 ^ n2151 ^ 1'b0 ;
  assign n20970 = n15429 & n20969 ;
  assign n20971 = ~n2903 & n20970 ;
  assign n20972 = n17888 ^ n3791 ^ 1'b0 ;
  assign n20973 = ~n20971 & n20972 ;
  assign n20974 = ~n3790 & n20973 ;
  assign n20975 = n12008 & ~n18066 ;
  assign n20976 = n20575 ^ n5377 ^ 1'b0 ;
  assign n20977 = n16474 & n20976 ;
  assign n20978 = n2884 & ~n5491 ;
  assign n20979 = n6652 & n20978 ;
  assign n20980 = n20979 ^ n669 ^ 1'b0 ;
  assign n20981 = n6623 & n20980 ;
  assign n20982 = n7399 ^ n1969 ^ 1'b0 ;
  assign n20983 = n20982 ^ n4179 ^ 1'b0 ;
  assign n20984 = n20146 ^ n19797 ^ 1'b0 ;
  assign n20985 = n17786 | n20984 ;
  assign n20986 = n5472 ^ n4916 ^ n2644 ;
  assign n20987 = n12298 & ~n20986 ;
  assign n20988 = n20987 ^ n15275 ^ 1'b0 ;
  assign n20989 = n314 | n18109 ;
  assign n20990 = n20989 ^ n19491 ^ 1'b0 ;
  assign n20991 = n1980 & ~n2662 ;
  assign n20992 = n12303 ^ n9185 ^ n6827 ;
  assign n20993 = n20992 ^ n6927 ^ n6435 ;
  assign n20996 = n7257 ^ n6948 ^ n2633 ;
  assign n20994 = ( n4517 & ~n5226 ) | ( n4517 & n11347 ) | ( ~n5226 & n11347 ) ;
  assign n20995 = n20994 ^ n2103 ^ 1'b0 ;
  assign n20997 = n20996 ^ n20995 ^ 1'b0 ;
  assign n20998 = n7545 | n20997 ;
  assign n20999 = n13512 ^ n2155 ^ 1'b0 ;
  assign n21000 = n3316 & ~n20999 ;
  assign n21001 = ~n11880 & n21000 ;
  assign n21002 = n21001 ^ n20980 ^ 1'b0 ;
  assign n21003 = ( ~n6855 & n14079 ) | ( ~n6855 & n21002 ) | ( n14079 & n21002 ) ;
  assign n21004 = ( n3725 & n13603 ) | ( n3725 & n21003 ) | ( n13603 & n21003 ) ;
  assign n21005 = n21004 ^ n12837 ^ 1'b0 ;
  assign n21006 = n20998 | n21005 ;
  assign n21007 = n15449 & n17488 ;
  assign n21008 = ~n11186 & n21007 ;
  assign n21009 = n7115 ^ n4514 ^ 1'b0 ;
  assign n21010 = x37 & ~n21009 ;
  assign n21011 = n3551 & n21010 ;
  assign n21012 = n5041 & n21011 ;
  assign n21013 = n19871 ^ n11276 ^ 1'b0 ;
  assign n21014 = n15897 & ~n21013 ;
  assign n21015 = n21014 ^ n17654 ^ 1'b0 ;
  assign n21016 = n17880 ^ n16168 ^ n2192 ;
  assign n21017 = ( ~n5065 & n15835 ) | ( ~n5065 & n21016 ) | ( n15835 & n21016 ) ;
  assign n21018 = n16244 ^ n410 ^ 1'b0 ;
  assign n21019 = n18672 ^ n6650 ^ 1'b0 ;
  assign n21020 = n3210 & n8063 ;
  assign n21021 = n8127 | n21020 ;
  assign n21022 = n5386 & ~n21021 ;
  assign n21023 = n21022 ^ n2660 ^ 1'b0 ;
  assign n21024 = ~n12005 & n21023 ;
  assign n21025 = n14774 & n21024 ;
  assign n21026 = n9820 ^ n7590 ^ n5034 ;
  assign n21027 = ( n1486 & n9304 ) | ( n1486 & ~n21026 ) | ( n9304 & ~n21026 ) ;
  assign n21028 = n1741 & ~n21027 ;
  assign n21029 = n21028 ^ n16817 ^ 1'b0 ;
  assign n21030 = ( n2244 & n9772 ) | ( n2244 & n21029 ) | ( n9772 & n21029 ) ;
  assign n21031 = n5159 | n13587 ;
  assign n21032 = n5426 ^ n2755 ^ 1'b0 ;
  assign n21033 = n11757 & ~n21032 ;
  assign n21034 = n3100 | n8600 ;
  assign n21035 = n21034 ^ n19041 ^ 1'b0 ;
  assign n21036 = n19897 | n21035 ;
  assign n21037 = n21033 | n21036 ;
  assign n21038 = n1265 & n9963 ;
  assign n21039 = n6298 & ~n12964 ;
  assign n21040 = ~n18516 & n21039 ;
  assign n21041 = ~n4313 & n6393 ;
  assign n21042 = n19598 & n21041 ;
  assign n21043 = ( n16445 & ~n17309 ) | ( n16445 & n21042 ) | ( ~n17309 & n21042 ) ;
  assign n21044 = ~n2836 & n3150 ;
  assign n21045 = n2722 & n21044 ;
  assign n21046 = n21045 ^ n19719 ^ n9864 ;
  assign n21047 = n10239 | n20379 ;
  assign n21048 = n21047 ^ n4531 ^ 1'b0 ;
  assign n21049 = n4510 | n21048 ;
  assign n21050 = ( n12060 & n18305 ) | ( n12060 & ~n19957 ) | ( n18305 & ~n19957 ) ;
  assign n21051 = ( ~n3067 & n8251 ) | ( ~n3067 & n21050 ) | ( n8251 & n21050 ) ;
  assign n21052 = n9266 ^ n5485 ^ 1'b0 ;
  assign n21053 = n15133 & ~n21052 ;
  assign n21054 = n9740 ^ n9025 ^ 1'b0 ;
  assign n21055 = n3315 & ~n21054 ;
  assign n21056 = n21055 ^ n9850 ^ n6437 ;
  assign n21057 = n21056 ^ x156 ^ 1'b0 ;
  assign n21058 = n12439 ^ n9874 ^ n6325 ;
  assign n21059 = n21058 ^ n4917 ^ 1'b0 ;
  assign n21060 = n5106 & ~n11538 ;
  assign n21061 = n914 & ~n5775 ;
  assign n21062 = ~n21060 & n21061 ;
  assign n21063 = n21059 & ~n21062 ;
  assign n21064 = n21063 ^ n14900 ^ n10157 ;
  assign n21065 = n11234 | n14244 ;
  assign n21066 = ~n11743 & n21065 ;
  assign n21067 = n21066 ^ n18856 ^ 1'b0 ;
  assign n21068 = ( n11173 & n11889 ) | ( n11173 & ~n21067 ) | ( n11889 & ~n21067 ) ;
  assign n21069 = n4884 | n5502 ;
  assign n21070 = n4911 | n21069 ;
  assign n21071 = n21070 ^ n14344 ^ n407 ;
  assign n21072 = n3962 & ~n21071 ;
  assign n21073 = n21072 ^ x124 ^ 1'b0 ;
  assign n21074 = n4754 ^ n3420 ^ 1'b0 ;
  assign n21075 = n21074 ^ n7252 ^ n1178 ;
  assign n21076 = n21075 ^ n5677 ^ 1'b0 ;
  assign n21077 = n4974 | n18569 ;
  assign n21078 = n1054 ^ x17 ^ 1'b0 ;
  assign n21079 = n8941 ^ n4039 ^ 1'b0 ;
  assign n21080 = n21078 & ~n21079 ;
  assign n21081 = n11649 | n15267 ;
  assign n21082 = n11845 | n21081 ;
  assign n21083 = n6204 ^ n4052 ^ 1'b0 ;
  assign n21084 = ~n11449 & n21083 ;
  assign n21085 = n19849 ^ n3995 ^ 1'b0 ;
  assign n21086 = n2680 & ~n16887 ;
  assign n21087 = n21085 & n21086 ;
  assign n21088 = n21084 & ~n21087 ;
  assign n21089 = n17888 & n21088 ;
  assign n21093 = ( n3085 & n13685 ) | ( n3085 & ~n20104 ) | ( n13685 & ~n20104 ) ;
  assign n21090 = n20157 ^ n5840 ^ 1'b0 ;
  assign n21091 = n3059 & n21090 ;
  assign n21092 = ~n1578 & n21091 ;
  assign n21094 = n21093 ^ n21092 ^ 1'b0 ;
  assign n21095 = n13521 & ~n14751 ;
  assign n21096 = n5386 & n6186 ;
  assign n21097 = n10317 & ~n10634 ;
  assign n21098 = ~n9360 & n21097 ;
  assign n21099 = n2819 ^ n1142 ^ x146 ;
  assign n21100 = n12090 ^ n3376 ^ 1'b0 ;
  assign n21101 = n21100 ^ n7345 ^ n2986 ;
  assign n21102 = x23 | n21101 ;
  assign n21105 = ( n2859 & n3637 ) | ( n2859 & n4310 ) | ( n3637 & n4310 ) ;
  assign n21104 = n6342 & n10439 ;
  assign n21106 = n21105 ^ n21104 ^ 1'b0 ;
  assign n21103 = n1179 & ~n15891 ;
  assign n21107 = n21106 ^ n21103 ^ x144 ;
  assign n21108 = ( ~x161 & n5133 ) | ( ~x161 & n6781 ) | ( n5133 & n6781 ) ;
  assign n21109 = n8572 & n21108 ;
  assign n21110 = n10606 ^ n4090 ^ n471 ;
  assign n21111 = ( n9033 & ~n15149 ) | ( n9033 & n21110 ) | ( ~n15149 & n21110 ) ;
  assign n21112 = ~n14473 & n21111 ;
  assign n21113 = n1479 & ~n8337 ;
  assign n21114 = n757 & ~n11567 ;
  assign n21115 = n21114 ^ n2541 ^ 1'b0 ;
  assign n21116 = ~x143 & n21115 ;
  assign n21117 = n12137 ^ n4664 ^ n424 ;
  assign n21118 = n823 & ~n1687 ;
  assign n21119 = n21118 ^ n3510 ^ 1'b0 ;
  assign n21120 = n13798 ^ n12535 ^ 1'b0 ;
  assign n21121 = n21119 & n21120 ;
  assign n21122 = ~n14968 & n15979 ;
  assign n21123 = ( ~n21117 & n21121 ) | ( ~n21117 & n21122 ) | ( n21121 & n21122 ) ;
  assign n21124 = n21123 ^ n18924 ^ 1'b0 ;
  assign n21125 = n15356 ^ n6321 ^ 1'b0 ;
  assign n21126 = n12904 & ~n21125 ;
  assign n21127 = x170 & n21126 ;
  assign n21128 = n21127 ^ n12704 ^ 1'b0 ;
  assign n21129 = n8305 ^ n7190 ^ n485 ;
  assign n21130 = ~n13124 & n21129 ;
  assign n21131 = ( n4763 & ~n8193 ) | ( n4763 & n17489 ) | ( ~n8193 & n17489 ) ;
  assign n21132 = n20503 ^ n15356 ^ n9795 ;
  assign n21133 = ~n7196 & n14877 ;
  assign n21135 = n20097 ^ n9280 ^ 1'b0 ;
  assign n21134 = n11017 & n14239 ;
  assign n21136 = n21135 ^ n21134 ^ 1'b0 ;
  assign n21137 = n11073 | n21136 ;
  assign n21138 = n6194 & ~n21137 ;
  assign n21139 = n10852 & n11809 ;
  assign n21140 = n21139 ^ n12762 ^ n9345 ;
  assign n21141 = n11463 | n21140 ;
  assign n21142 = n21138 & ~n21141 ;
  assign n21143 = n1326 & ~n15334 ;
  assign n21144 = n21143 ^ n7493 ^ 1'b0 ;
  assign n21145 = n5037 & n6695 ;
  assign n21146 = ~n15795 & n21145 ;
  assign n21147 = n21146 ^ n18392 ^ 1'b0 ;
  assign n21148 = n1405 & n15550 ;
  assign n21149 = n21148 ^ n4214 ^ 1'b0 ;
  assign n21150 = n15346 | n21149 ;
  assign n21151 = n4700 | n21150 ;
  assign n21152 = n2244 & n10426 ;
  assign n21153 = ~n21151 & n21152 ;
  assign n21154 = n15051 ^ n8627 ^ 1'b0 ;
  assign n21155 = ( n19655 & n21153 ) | ( n19655 & n21154 ) | ( n21153 & n21154 ) ;
  assign n21156 = n4740 & n6335 ;
  assign n21157 = n1931 & n4154 ;
  assign n21158 = n20191 & n21157 ;
  assign n21159 = ~n21156 & n21158 ;
  assign n21160 = n19138 ^ n15964 ^ n2831 ;
  assign n21161 = n18610 & n21160 ;
  assign n21162 = n4118 & ~n6000 ;
  assign n21163 = ( n472 & n3589 ) | ( n472 & ~n20640 ) | ( n3589 & ~n20640 ) ;
  assign n21164 = n21163 ^ n3339 ^ x98 ;
  assign n21165 = n21164 ^ n14319 ^ 1'b0 ;
  assign n21166 = n11951 & ~n21165 ;
  assign n21167 = n21166 ^ n18623 ^ 1'b0 ;
  assign n21168 = ~n17301 & n21167 ;
  assign n21169 = n5090 ^ n3866 ^ 1'b0 ;
  assign n21170 = n7037 ^ n5259 ^ 1'b0 ;
  assign n21171 = ( n6879 & n7753 ) | ( n6879 & ~n21170 ) | ( n7753 & ~n21170 ) ;
  assign n21172 = n3436 | n9276 ;
  assign n21173 = n21172 ^ n18305 ^ 1'b0 ;
  assign n21174 = n10980 & ~n18349 ;
  assign n21175 = n3436 | n12587 ;
  assign n21176 = n6364 & ~n21175 ;
  assign n21177 = n21176 ^ n19520 ^ n300 ;
  assign n21178 = n21177 ^ n13423 ^ n9174 ;
  assign n21181 = n16668 ^ n13717 ^ n513 ;
  assign n21179 = n9203 ^ n5420 ^ n1145 ;
  assign n21180 = ( n5186 & n12122 ) | ( n5186 & ~n21179 ) | ( n12122 & ~n21179 ) ;
  assign n21182 = n21181 ^ n21180 ^ n10365 ;
  assign n21183 = ( ~n6448 & n8546 ) | ( ~n6448 & n9102 ) | ( n8546 & n9102 ) ;
  assign n21184 = n3065 & ~n21183 ;
  assign n21185 = n14091 & n21184 ;
  assign n21186 = n10401 & ~n17551 ;
  assign n21187 = n21186 ^ n7508 ^ 1'b0 ;
  assign n21188 = n16677 & n21187 ;
  assign n21189 = n12196 ^ n7698 ^ 1'b0 ;
  assign n21190 = ~n5004 & n21189 ;
  assign n21191 = n21190 ^ n20269 ^ 1'b0 ;
  assign n21192 = n21188 | n21191 ;
  assign n21194 = n6124 & n19363 ;
  assign n21193 = ~n3764 & n10811 ;
  assign n21195 = n21194 ^ n21193 ^ 1'b0 ;
  assign n21202 = n5428 ^ n1463 ^ 1'b0 ;
  assign n21203 = ~n1617 & n21202 ;
  assign n21204 = n21203 ^ n7812 ^ 1'b0 ;
  assign n21198 = n4540 ^ n2376 ^ 1'b0 ;
  assign n21199 = n9112 & ~n13039 ;
  assign n21200 = n21198 & n21199 ;
  assign n21201 = ( n2859 & ~n7591 ) | ( n2859 & n21200 ) | ( ~n7591 & n21200 ) ;
  assign n21205 = n21204 ^ n21201 ^ n14791 ;
  assign n21206 = n9206 | n21205 ;
  assign n21196 = n8573 ^ n6008 ^ 1'b0 ;
  assign n21197 = ~n13021 & n21196 ;
  assign n21207 = n21206 ^ n21197 ^ 1'b0 ;
  assign n21208 = n2721 | n9822 ;
  assign n21209 = n15981 & ~n21208 ;
  assign n21210 = n21095 ^ n9155 ^ 1'b0 ;
  assign n21211 = n5367 | n21210 ;
  assign n21212 = ( n5456 & n8930 ) | ( n5456 & n10529 ) | ( n8930 & n10529 ) ;
  assign n21213 = n9588 ^ n852 ^ 1'b0 ;
  assign n21214 = n21213 ^ n8043 ^ 1'b0 ;
  assign n21215 = n21214 ^ n16848 ^ 1'b0 ;
  assign n21216 = n12654 ^ n3970 ^ 1'b0 ;
  assign n21217 = n20796 & ~n21216 ;
  assign n21218 = n18737 & n21217 ;
  assign n21219 = n21218 ^ n20187 ^ 1'b0 ;
  assign n21220 = x53 & ~n6509 ;
  assign n21221 = ( x116 & n12925 ) | ( x116 & ~n21220 ) | ( n12925 & ~n21220 ) ;
  assign n21222 = ~n8093 & n21221 ;
  assign n21223 = ( n1090 & n4611 ) | ( n1090 & ~n9719 ) | ( n4611 & ~n9719 ) ;
  assign n21224 = n895 & n21223 ;
  assign n21225 = n19282 ^ n19250 ^ 1'b0 ;
  assign n21226 = ~n18370 & n21225 ;
  assign n21227 = n21226 ^ n9276 ^ 1'b0 ;
  assign n21228 = n18830 ^ n3232 ^ 1'b0 ;
  assign n21229 = n5860 & ~n21228 ;
  assign n21230 = n21229 ^ n10072 ^ 1'b0 ;
  assign n21231 = n21230 ^ n2733 ^ n1051 ;
  assign n21232 = n21231 ^ n14011 ^ 1'b0 ;
  assign n21233 = n17664 & ~n21232 ;
  assign n21241 = n3688 & ~n15780 ;
  assign n21242 = n3791 & n21241 ;
  assign n21237 = ~n3487 & n19037 ;
  assign n21238 = n10485 & n21237 ;
  assign n21234 = n1521 ^ n932 ^ 1'b0 ;
  assign n21235 = ~n4867 & n21234 ;
  assign n21236 = n2828 & n21235 ;
  assign n21239 = n21238 ^ n21236 ^ 1'b0 ;
  assign n21240 = ~n5094 & n21239 ;
  assign n21243 = n21242 ^ n21240 ^ 1'b0 ;
  assign n21244 = n11667 ^ n6078 ^ n4867 ;
  assign n21245 = n15391 ^ n14636 ^ n3585 ;
  assign n21246 = n10099 | n12682 ;
  assign n21247 = n7668 | n21246 ;
  assign n21248 = ~n13414 & n20723 ;
  assign n21249 = n14017 & n21248 ;
  assign n21250 = n4760 & n10742 ;
  assign n21251 = n9921 | n16621 ;
  assign n21252 = n21251 ^ n15825 ^ 1'b0 ;
  assign n21253 = ( n1022 & ~n17639 ) | ( n1022 & n21252 ) | ( ~n17639 & n21252 ) ;
  assign n21254 = n5362 ^ n3304 ^ 1'b0 ;
  assign n21255 = n12718 ^ n2711 ^ 1'b0 ;
  assign n21256 = ( n12418 & ~n21254 ) | ( n12418 & n21255 ) | ( ~n21254 & n21255 ) ;
  assign n21257 = n10735 | n21256 ;
  assign n21258 = n21257 ^ n20888 ^ 1'b0 ;
  assign n21259 = n16131 ^ n5685 ^ n2832 ;
  assign n21260 = ( n2128 & n3795 ) | ( n2128 & n5556 ) | ( n3795 & n5556 ) ;
  assign n21261 = n21260 ^ n10517 ^ n10125 ;
  assign n21262 = n15229 ^ n13616 ^ 1'b0 ;
  assign n21263 = ~n2202 & n9662 ;
  assign n21264 = ~n4411 & n21263 ;
  assign n21265 = n21262 | n21264 ;
  assign n21266 = n21261 & ~n21265 ;
  assign n21267 = n17616 & ~n21266 ;
  assign n21268 = ~n21259 & n21267 ;
  assign n21269 = n1664 & ~n5815 ;
  assign n21270 = n21269 ^ n13127 ^ n10659 ;
  assign n21271 = n10190 ^ n9515 ^ 1'b0 ;
  assign n21272 = ~n2131 & n21271 ;
  assign n21273 = n21272 ^ n7302 ^ 1'b0 ;
  assign n21274 = ~n21270 & n21273 ;
  assign n21275 = ~n18715 & n21274 ;
  assign n21276 = ~n8853 & n12367 ;
  assign n21277 = n21276 ^ n11341 ^ 1'b0 ;
  assign n21278 = n5898 ^ x19 ^ 1'b0 ;
  assign n21279 = n21277 & ~n21278 ;
  assign n21280 = x129 & n21279 ;
  assign n21281 = ~n16824 & n21280 ;
  assign n21282 = n9345 ^ n759 ^ 1'b0 ;
  assign n21283 = n6742 & n21282 ;
  assign n21284 = x0 & n14004 ;
  assign n21285 = ~n19066 & n21284 ;
  assign n21286 = n580 | n15759 ;
  assign n21287 = n21286 ^ n16512 ^ n7177 ;
  assign n21288 = ( n4224 & ~n6719 ) | ( n4224 & n10845 ) | ( ~n6719 & n10845 ) ;
  assign n21289 = n17983 & ~n20120 ;
  assign n21290 = n10182 | n21289 ;
  assign n21291 = n16841 & ~n21290 ;
  assign n21292 = ( n2064 & n4020 ) | ( n2064 & ~n12804 ) | ( n4020 & ~n12804 ) ;
  assign n21293 = n5134 & ~n6491 ;
  assign n21294 = ~n21292 & n21293 ;
  assign n21295 = n17341 ^ n11315 ^ n9837 ;
  assign n21296 = n17530 | n21295 ;
  assign n21297 = n7936 ^ n2019 ^ 1'b0 ;
  assign n21298 = x19 & ~n17587 ;
  assign n21299 = ~n6645 & n21298 ;
  assign n21300 = n9906 & ~n12963 ;
  assign n21301 = n21299 & n21300 ;
  assign n21302 = n6555 & ~n17357 ;
  assign n21303 = n21302 ^ n20164 ^ 1'b0 ;
  assign n21304 = n14206 ^ n12499 ^ 1'b0 ;
  assign n21305 = n6376 & ~n21304 ;
  assign n21306 = ~n2071 & n21305 ;
  assign n21307 = n21306 ^ n12495 ^ 1'b0 ;
  assign n21308 = ~n8613 & n21307 ;
  assign n21309 = n4493 | n13388 ;
  assign n21310 = n13086 ^ n4426 ^ 1'b0 ;
  assign n21311 = x80 & ~n3724 ;
  assign n21312 = n12265 & ~n21311 ;
  assign n21313 = n1271 & ~n2937 ;
  assign n21314 = n21313 ^ n8357 ^ 1'b0 ;
  assign n21315 = n21314 ^ n7464 ^ n6606 ;
  assign n21317 = n952 & ~n3040 ;
  assign n21318 = n21317 ^ n15686 ^ 1'b0 ;
  assign n21319 = n21318 ^ n3692 ^ 1'b0 ;
  assign n21316 = ( n1168 & n10902 ) | ( n1168 & ~n20224 ) | ( n10902 & ~n20224 ) ;
  assign n21320 = n21319 ^ n21316 ^ n8760 ;
  assign n21321 = n21320 ^ n8151 ^ 1'b0 ;
  assign n21322 = n8731 | n21321 ;
  assign n21323 = n21315 & ~n21322 ;
  assign n21324 = ( n4097 & ~n6182 ) | ( n4097 & n11045 ) | ( ~n6182 & n11045 ) ;
  assign n21326 = n5060 & ~n9172 ;
  assign n21325 = n2399 | n4372 ;
  assign n21327 = n21326 ^ n21325 ^ n15096 ;
  assign n21328 = n2811 & n13150 ;
  assign n21329 = n21328 ^ n7542 ^ 1'b0 ;
  assign n21330 = n17428 ^ n10755 ^ n8762 ;
  assign n21331 = n21330 ^ n13858 ^ n4303 ;
  assign n21332 = n21329 | n21331 ;
  assign n21333 = ~n12720 & n20470 ;
  assign n21334 = n21333 ^ n4992 ^ 1'b0 ;
  assign n21335 = n10654 ^ n2005 ^ 1'b0 ;
  assign n21336 = ~n11118 & n21335 ;
  assign n21337 = n19915 ^ n8775 ^ n5539 ;
  assign n21338 = n21337 ^ n7244 ^ 1'b0 ;
  assign n21339 = n21336 & n21338 ;
  assign n21340 = n19780 ^ n2843 ^ 1'b0 ;
  assign n21341 = n17883 ^ n11802 ^ n595 ;
  assign n21345 = n2688 | n6206 ;
  assign n21342 = n1709 ^ x136 ^ 1'b0 ;
  assign n21343 = n11791 & ~n21342 ;
  assign n21344 = n21343 ^ n20952 ^ n335 ;
  assign n21346 = n21345 ^ n21344 ^ 1'b0 ;
  assign n21347 = n21341 | n21346 ;
  assign n21348 = n18004 & ~n21347 ;
  assign n21349 = n2836 | n7378 ;
  assign n21350 = n11966 | n21349 ;
  assign n21351 = ( n7478 & ~n9506 ) | ( n7478 & n21350 ) | ( ~n9506 & n21350 ) ;
  assign n21352 = n21351 ^ n19220 ^ n11391 ;
  assign n21353 = n7315 ^ n5320 ^ 1'b0 ;
  assign n21354 = ~n7677 & n21353 ;
  assign n21355 = n20460 ^ n4220 ^ 1'b0 ;
  assign n21356 = n21354 & ~n21355 ;
  assign n21357 = ( ~n1390 & n4527 ) | ( ~n1390 & n12936 ) | ( n4527 & n12936 ) ;
  assign n21358 = n7740 & n21357 ;
  assign n21359 = n11256 & ~n20481 ;
  assign n21363 = n1752 & ~n5500 ;
  assign n21362 = ~n6952 & n10437 ;
  assign n21360 = n4652 ^ n669 ^ 1'b0 ;
  assign n21361 = n21360 ^ n6927 ^ n5325 ;
  assign n21364 = n21363 ^ n21362 ^ n21361 ;
  assign n21368 = n6385 | n10922 ;
  assign n21369 = n21368 ^ n10543 ^ 1'b0 ;
  assign n21365 = n9732 | n15027 ;
  assign n21366 = n12731 | n21365 ;
  assign n21367 = n3664 | n21366 ;
  assign n21370 = n21369 ^ n21367 ^ 1'b0 ;
  assign n21372 = ~n4019 & n7517 ;
  assign n21371 = n4239 ^ n794 ^ 1'b0 ;
  assign n21373 = n21372 ^ n21371 ^ 1'b0 ;
  assign n21374 = n11454 & ~n11626 ;
  assign n21375 = n21374 ^ n11593 ^ 1'b0 ;
  assign n21376 = n21357 & ~n21375 ;
  assign n21377 = n3211 & n21376 ;
  assign n21378 = n18429 ^ n14096 ^ 1'b0 ;
  assign n21379 = n9426 & n21378 ;
  assign n21384 = ( n1403 & n7723 ) | ( n1403 & n11031 ) | ( n7723 & n11031 ) ;
  assign n21385 = ( n3795 & ~n5385 ) | ( n3795 & n21384 ) | ( ~n5385 & n21384 ) ;
  assign n21386 = n21385 ^ n6649 ^ n2225 ;
  assign n21380 = n9184 ^ n8361 ^ n4600 ;
  assign n21381 = n21380 ^ n10906 ^ n1933 ;
  assign n21382 = n21381 ^ n3474 ^ 1'b0 ;
  assign n21383 = ~n8536 & n21382 ;
  assign n21387 = n21386 ^ n21383 ^ 1'b0 ;
  assign n21388 = n21387 ^ n857 ^ 1'b0 ;
  assign n21389 = n2679 & n15950 ;
  assign n21390 = n21389 ^ n3475 ^ 1'b0 ;
  assign n21391 = n2394 & ~n5228 ;
  assign n21392 = n21391 ^ n9421 ^ 1'b0 ;
  assign n21393 = n11753 & n19285 ;
  assign n21394 = ~n11100 & n21393 ;
  assign n21399 = n20693 ^ n844 ^ 1'b0 ;
  assign n21400 = ~n4453 & n21399 ;
  assign n21397 = n13798 ^ n2539 ^ 1'b0 ;
  assign n21395 = n16842 ^ n9102 ^ 1'b0 ;
  assign n21396 = n17264 | n21395 ;
  assign n21398 = n21397 ^ n21396 ^ n13086 ;
  assign n21401 = n21400 ^ n21398 ^ 1'b0 ;
  assign n21402 = n1657 & ~n21401 ;
  assign n21403 = n19619 ^ n8613 ^ n2120 ;
  assign n21404 = n13649 & n21403 ;
  assign n21405 = x154 & ~n21404 ;
  assign n21406 = ( ~n2504 & n3068 ) | ( ~n2504 & n19648 ) | ( n3068 & n19648 ) ;
  assign n21407 = n6188 & n8494 ;
  assign n21408 = n21407 ^ x215 ^ 1'b0 ;
  assign n21409 = n4013 & ~n10904 ;
  assign n21410 = n21409 ^ x117 ^ 1'b0 ;
  assign n21411 = n18888 ^ n18130 ^ 1'b0 ;
  assign n21412 = n15987 & n21411 ;
  assign n21413 = n11659 ^ n8214 ^ 1'b0 ;
  assign n21414 = n976 | n8774 ;
  assign n21415 = n6129 & n21414 ;
  assign n21416 = n2824 & n12907 ;
  assign n21417 = n21416 ^ n450 ^ 1'b0 ;
  assign n21420 = ( n8137 & n13659 ) | ( n8137 & n21260 ) | ( n13659 & n21260 ) ;
  assign n21421 = ( n8163 & n8754 ) | ( n8163 & ~n21420 ) | ( n8754 & ~n21420 ) ;
  assign n21418 = x155 | n733 ;
  assign n21419 = n21418 ^ n21319 ^ n18779 ;
  assign n21422 = n21421 ^ n21419 ^ 1'b0 ;
  assign n21423 = ~n8928 & n21422 ;
  assign n21424 = ~n17566 & n21423 ;
  assign n21425 = n20660 ^ n6835 ^ 1'b0 ;
  assign n21426 = n15799 ^ n12794 ^ n8496 ;
  assign n21427 = ( n3152 & n11045 ) | ( n3152 & ~n21426 ) | ( n11045 & ~n21426 ) ;
  assign n21428 = ~n6458 & n21427 ;
  assign n21429 = n21428 ^ n6710 ^ 1'b0 ;
  assign n21430 = n15694 ^ n8458 ^ n4569 ;
  assign n21431 = ~n5712 & n21430 ;
  assign n21432 = x104 & n21431 ;
  assign n21433 = n21432 ^ n4979 ^ 1'b0 ;
  assign n21434 = ( n2531 & n14954 ) | ( n2531 & n21433 ) | ( n14954 & n21433 ) ;
  assign n21435 = n10064 ^ n6533 ^ n4694 ;
  assign n21436 = n20889 ^ n16375 ^ 1'b0 ;
  assign n21437 = n21436 ^ n8818 ^ n1158 ;
  assign n21438 = ~n10046 & n12457 ;
  assign n21439 = ~n7223 & n21438 ;
  assign n21440 = n21439 ^ n10830 ^ 1'b0 ;
  assign n21441 = n11252 & n21440 ;
  assign n21442 = n21437 & n21441 ;
  assign n21443 = n6915 & n8641 ;
  assign n21444 = n21443 ^ n8013 ^ 1'b0 ;
  assign n21445 = ~n15677 & n21444 ;
  assign n21446 = n16341 & n21445 ;
  assign n21447 = ~n4579 & n9044 ;
  assign n21448 = ~n9336 & n21447 ;
  assign n21455 = n5830 | n11880 ;
  assign n21456 = n5521 & ~n21455 ;
  assign n21457 = n21456 ^ n10388 ^ n2296 ;
  assign n21449 = n2727 | n5103 ;
  assign n21450 = n21449 ^ n4725 ^ 1'b0 ;
  assign n21451 = n16167 ^ n9100 ^ 1'b0 ;
  assign n21452 = n6643 | n21451 ;
  assign n21453 = n21452 ^ n18231 ^ n14976 ;
  assign n21454 = ~n21450 & n21453 ;
  assign n21458 = n21457 ^ n21454 ^ n11806 ;
  assign n21459 = n8261 ^ n3173 ^ 1'b0 ;
  assign n21460 = n11571 | n17102 ;
  assign n21461 = ( n2665 & n21459 ) | ( n2665 & n21460 ) | ( n21459 & n21460 ) ;
  assign n21462 = n4695 ^ n584 ^ 1'b0 ;
  assign n21464 = n1820 | n3322 ;
  assign n21463 = ( n3017 & n9418 ) | ( n3017 & n13278 ) | ( n9418 & n13278 ) ;
  assign n21465 = n21464 ^ n21463 ^ n3592 ;
  assign n21466 = ~n4141 & n21465 ;
  assign n21467 = n21466 ^ n15710 ^ 1'b0 ;
  assign n21468 = ~n21462 & n21467 ;
  assign n21469 = n10703 & ~n11264 ;
  assign n21470 = n18127 | n21469 ;
  assign n21471 = n4563 ^ n2648 ^ 1'b0 ;
  assign n21472 = n21471 ^ n2313 ^ 1'b0 ;
  assign n21473 = ( n808 & n4306 ) | ( n808 & ~n10412 ) | ( n4306 & ~n10412 ) ;
  assign n21474 = ~n18774 & n21473 ;
  assign n21475 = n3675 ^ n3393 ^ 1'b0 ;
  assign n21476 = n21475 ^ n11420 ^ 1'b0 ;
  assign n21477 = n2507 & ~n10643 ;
  assign n21478 = n21477 ^ n13850 ^ 1'b0 ;
  assign n21479 = n21478 ^ n15901 ^ n6357 ;
  assign n21480 = n12592 | n13278 ;
  assign n21481 = n21480 ^ n7366 ^ 1'b0 ;
  assign n21482 = ( ~n12808 & n15282 ) | ( ~n12808 & n21481 ) | ( n15282 & n21481 ) ;
  assign n21485 = n2347 ^ n911 ^ 1'b0 ;
  assign n21484 = n2680 | n3390 ;
  assign n21486 = n21485 ^ n21484 ^ 1'b0 ;
  assign n21483 = n12382 ^ n884 ^ 1'b0 ;
  assign n21487 = n21486 ^ n21483 ^ n4479 ;
  assign n21488 = n21487 ^ n6189 ^ 1'b0 ;
  assign n21489 = n19688 ^ n13994 ^ n7808 ;
  assign n21490 = ( n15451 & n18770 ) | ( n15451 & ~n21489 ) | ( n18770 & ~n21489 ) ;
  assign n21491 = ~n1076 & n2110 ;
  assign n21492 = n3950 & n21491 ;
  assign n21493 = n6788 | n21492 ;
  assign n21494 = n6952 | n10068 ;
  assign n21495 = n21494 ^ n1227 ^ 1'b0 ;
  assign n21496 = ( n3825 & ~n10214 ) | ( n3825 & n15428 ) | ( ~n10214 & n15428 ) ;
  assign n21497 = n7917 & ~n21496 ;
  assign n21498 = n21495 & n21497 ;
  assign n21499 = n5639 & n18874 ;
  assign n21500 = ( n5925 & ~n7049 ) | ( n5925 & n17654 ) | ( ~n7049 & n17654 ) ;
  assign n21501 = ( n8015 & n16443 ) | ( n8015 & n21500 ) | ( n16443 & n21500 ) ;
  assign n21502 = n2035 & ~n21122 ;
  assign n21503 = n3393 & n21502 ;
  assign n21507 = n7448 & ~n10912 ;
  assign n21508 = n21507 ^ n12648 ^ 1'b0 ;
  assign n21509 = ~n15969 & n21508 ;
  assign n21510 = n15969 & n21509 ;
  assign n21511 = n16997 & ~n21510 ;
  assign n21512 = n21510 & n21511 ;
  assign n21513 = n7324 | n21512 ;
  assign n21514 = n21512 & ~n21513 ;
  assign n21515 = n13029 | n21514 ;
  assign n21516 = n21514 & ~n21515 ;
  assign n21504 = n4827 | n12087 ;
  assign n21505 = n21504 ^ n10440 ^ 1'b0 ;
  assign n21506 = ( n15864 & n17159 ) | ( n15864 & n21505 ) | ( n17159 & n21505 ) ;
  assign n21517 = n21516 ^ n21506 ^ n16400 ;
  assign n21518 = n1932 & ~n8545 ;
  assign n21519 = ~n1932 & n21518 ;
  assign n21520 = ( n4247 & n9815 ) | ( n4247 & n19079 ) | ( n9815 & n19079 ) ;
  assign n21521 = n14521 ^ n5857 ^ 1'b0 ;
  assign n21522 = ( n2046 & n18297 ) | ( n2046 & n21521 ) | ( n18297 & n21521 ) ;
  assign n21523 = n7442 ^ n6602 ^ 1'b0 ;
  assign n21524 = n7012 & n8989 ;
  assign n21525 = n21524 ^ n4048 ^ 1'b0 ;
  assign n21526 = ( n3363 & n8805 ) | ( n3363 & n15081 ) | ( n8805 & n15081 ) ;
  assign n21527 = n15316 ^ n7480 ^ 1'b0 ;
  assign n21529 = ~n6922 & n10923 ;
  assign n21530 = n21529 ^ n517 ^ 1'b0 ;
  assign n21528 = n17620 & ~n20566 ;
  assign n21531 = n21530 ^ n21528 ^ 1'b0 ;
  assign n21532 = ~n538 & n21531 ;
  assign n21533 = n21532 ^ n8563 ^ 1'b0 ;
  assign n21534 = n21533 ^ n18509 ^ 1'b0 ;
  assign n21535 = n21527 & ~n21534 ;
  assign n21536 = n12493 & n14632 ;
  assign n21537 = n21536 ^ x160 ^ 1'b0 ;
  assign n21538 = ( n1943 & n3605 ) | ( n1943 & ~n11746 ) | ( n3605 & ~n11746 ) ;
  assign n21539 = n9925 & n21538 ;
  assign n21540 = n5762 & n21539 ;
  assign n21541 = n19276 & ~n21540 ;
  assign n21542 = n15736 ^ n827 ^ 1'b0 ;
  assign n21543 = ( n1084 & ~n2726 ) | ( n1084 & n5475 ) | ( ~n2726 & n5475 ) ;
  assign n21544 = n7517 | n21543 ;
  assign n21545 = n18266 ^ n6756 ^ 1'b0 ;
  assign n21546 = n21545 ^ n12581 ^ n9897 ;
  assign n21547 = ( n9607 & n15431 ) | ( n9607 & n21546 ) | ( n15431 & n21546 ) ;
  assign n21548 = ~n3005 & n10838 ;
  assign n21549 = n21548 ^ n5011 ^ 1'b0 ;
  assign n21550 = ( n8962 & n15307 ) | ( n8962 & ~n21549 ) | ( n15307 & ~n21549 ) ;
  assign n21551 = n3449 | n19138 ;
  assign n21552 = n21551 ^ n15429 ^ 1'b0 ;
  assign n21553 = n15793 ^ n13519 ^ 1'b0 ;
  assign n21556 = n3150 ^ n1265 ^ 1'b0 ;
  assign n21557 = n14980 & n21556 ;
  assign n21554 = n7069 ^ n5262 ^ 1'b0 ;
  assign n21555 = ( ~n12715 & n14487 ) | ( ~n12715 & n21554 ) | ( n14487 & n21554 ) ;
  assign n21558 = n21557 ^ n21555 ^ 1'b0 ;
  assign n21559 = n7581 & ~n16965 ;
  assign n21564 = n3687 | n9723 ;
  assign n21565 = n21564 ^ n4098 ^ 1'b0 ;
  assign n21566 = n8221 ^ n545 ^ 1'b0 ;
  assign n21567 = ~n21565 & n21566 ;
  assign n21563 = ( x37 & n8094 ) | ( x37 & n12488 ) | ( n8094 & n12488 ) ;
  assign n21560 = n2657 ^ x102 ^ 1'b0 ;
  assign n21561 = n21560 ^ n11355 ^ n7459 ;
  assign n21562 = ( n2836 & n3445 ) | ( n2836 & ~n21561 ) | ( n3445 & ~n21561 ) ;
  assign n21568 = n21567 ^ n21563 ^ n21562 ;
  assign n21569 = n3042 & ~n11841 ;
  assign n21570 = n21569 ^ n5502 ^ n4026 ;
  assign n21572 = n2468 & ~n9587 ;
  assign n21573 = n12219 & n21572 ;
  assign n21571 = n1948 | n9670 ;
  assign n21574 = n21573 ^ n21571 ^ n14563 ;
  assign n21575 = n21574 ^ n20845 ^ n10355 ;
  assign n21576 = n17317 ^ n13326 ^ 1'b0 ;
  assign n21580 = ~n3739 & n5662 ;
  assign n21577 = n17661 ^ n17301 ^ 1'b0 ;
  assign n21578 = ~n8061 & n21577 ;
  assign n21579 = n21578 ^ n19936 ^ n19680 ;
  assign n21581 = n21580 ^ n21579 ^ 1'b0 ;
  assign n21582 = n21299 ^ n7309 ^ n4928 ;
  assign n21583 = ~n19213 & n21582 ;
  assign n21584 = ~n16060 & n21583 ;
  assign n21585 = n5334 & n8018 ;
  assign n21586 = ( ~n711 & n17223 ) | ( ~n711 & n21585 ) | ( n17223 & n21585 ) ;
  assign n21587 = n13874 ^ n11027 ^ 1'b0 ;
  assign n21588 = n6172 & ~n21587 ;
  assign n21589 = n10408 ^ n478 ^ 1'b0 ;
  assign n21590 = n2554 ^ n1280 ^ 1'b0 ;
  assign n21591 = n12549 & n21590 ;
  assign n21592 = n21591 ^ n17428 ^ n6514 ;
  assign n21593 = n15221 ^ n6621 ^ 1'b0 ;
  assign n21595 = n14349 ^ n13625 ^ n6129 ;
  assign n21594 = n20316 ^ n20024 ^ n12481 ;
  assign n21596 = n21595 ^ n21594 ^ 1'b0 ;
  assign n21597 = n21593 & ~n21596 ;
  assign n21598 = n6581 ^ n5502 ^ 1'b0 ;
  assign n21599 = n21598 ^ n9318 ^ 1'b0 ;
  assign n21600 = n854 | n21599 ;
  assign n21601 = n17163 & ~n21600 ;
  assign n21602 = n4585 & n21601 ;
  assign n21603 = n3169 & ~n5027 ;
  assign n21604 = ( n3758 & n6549 ) | ( n3758 & n21603 ) | ( n6549 & n21603 ) ;
  assign n21605 = n13288 & ~n21604 ;
  assign n21606 = n8629 & ~n14847 ;
  assign n21607 = ~n21605 & n21606 ;
  assign n21608 = ~n10837 & n19577 ;
  assign n21609 = n8616 ^ n2662 ^ 1'b0 ;
  assign n21612 = ~n8606 & n9073 ;
  assign n21610 = n7716 & ~n10852 ;
  assign n21611 = n21610 ^ n4592 ^ 1'b0 ;
  assign n21613 = n21612 ^ n21611 ^ n16406 ;
  assign n21614 = n6332 | n14978 ;
  assign n21615 = n9784 | n21614 ;
  assign n21616 = n21615 ^ n15969 ^ n9463 ;
  assign n21617 = n7545 | n19692 ;
  assign n21618 = n21617 ^ n14091 ^ 1'b0 ;
  assign n21619 = n7790 & n18371 ;
  assign n21620 = n10758 & n21619 ;
  assign n21624 = n1406 | n9018 ;
  assign n21625 = n6032 ^ n5117 ^ n3753 ;
  assign n21626 = n21625 ^ n7390 ^ 1'b0 ;
  assign n21627 = n21624 & ~n21626 ;
  assign n21621 = n4439 & n6684 ;
  assign n21622 = n4078 & n21621 ;
  assign n21623 = ~n8403 & n21622 ;
  assign n21628 = n21627 ^ n21623 ^ n5042 ;
  assign n21629 = n21628 ^ n15766 ^ 1'b0 ;
  assign n21630 = n21354 & n21629 ;
  assign n21631 = n9976 & n18156 ;
  assign n21632 = n21631 ^ n16385 ^ 1'b0 ;
  assign n21633 = n13678 ^ n5365 ^ 1'b0 ;
  assign n21634 = n21633 ^ n843 ^ 1'b0 ;
  assign n21635 = n5860 & ~n21634 ;
  assign n21639 = ~n410 & n6646 ;
  assign n21640 = n8130 & n21639 ;
  assign n21636 = n7879 ^ n2445 ^ n2290 ;
  assign n21637 = ( n3831 & ~n12070 ) | ( n3831 & n21636 ) | ( ~n12070 & n21636 ) ;
  assign n21638 = n21637 ^ n5186 ^ 1'b0 ;
  assign n21641 = n21640 ^ n21638 ^ 1'b0 ;
  assign n21642 = ~n6218 & n9059 ;
  assign n21643 = n21642 ^ n9312 ^ 1'b0 ;
  assign n21644 = n10598 | n21643 ;
  assign n21645 = ( n7361 & ~n10501 ) | ( n7361 & n21644 ) | ( ~n10501 & n21644 ) ;
  assign n21646 = n1702 & n2970 ;
  assign n21647 = n2819 & n21646 ;
  assign n21648 = ( n3029 & n12188 ) | ( n3029 & ~n21647 ) | ( n12188 & ~n21647 ) ;
  assign n21649 = ( n7012 & ~n12861 ) | ( n7012 & n21648 ) | ( ~n12861 & n21648 ) ;
  assign n21650 = ( n7263 & ~n17445 ) | ( n7263 & n21570 ) | ( ~n17445 & n21570 ) ;
  assign n21651 = n16663 ^ n12939 ^ n9314 ;
  assign n21652 = n21651 ^ n7912 ^ 1'b0 ;
  assign n21653 = n6087 & n21652 ;
  assign n21654 = ~n5601 & n21653 ;
  assign n21656 = ( n932 & n6156 ) | ( n932 & ~n6901 ) | ( n6156 & ~n6901 ) ;
  assign n21657 = n21656 ^ n21202 ^ 1'b0 ;
  assign n21658 = n17167 & n21657 ;
  assign n21655 = ( ~n5754 & n6389 ) | ( ~n5754 & n13092 ) | ( n6389 & n13092 ) ;
  assign n21659 = n21658 ^ n21655 ^ 1'b0 ;
  assign n21660 = n3998 & ~n21659 ;
  assign n21661 = ~n312 & n8295 ;
  assign n21662 = n21661 ^ n17952 ^ n11023 ;
  assign n21663 = n8698 | n14765 ;
  assign n21664 = ~n9012 & n21663 ;
  assign n21665 = n1098 & n21664 ;
  assign n21666 = ~n4572 & n6747 ;
  assign n21667 = ( n10661 & ~n20950 ) | ( n10661 & n21666 ) | ( ~n20950 & n21666 ) ;
  assign n21668 = n5576 & n9498 ;
  assign n21669 = n21668 ^ n2634 ^ 1'b0 ;
  assign n21670 = ~n7466 & n21669 ;
  assign n21671 = n21670 ^ n14185 ^ 1'b0 ;
  assign n21672 = ~n12374 & n21671 ;
  assign n21673 = n13997 & ~n20399 ;
  assign n21674 = ~x229 & n6506 ;
  assign n21675 = n21674 ^ n18766 ^ n1465 ;
  assign n21676 = n18302 ^ n3731 ^ 1'b0 ;
  assign n21677 = n5515 ^ n2901 ^ 1'b0 ;
  assign n21678 = ~n1996 & n21677 ;
  assign n21679 = n21678 ^ n8145 ^ 1'b0 ;
  assign n21680 = n16315 & n20805 ;
  assign n21681 = n6453 & n9721 ;
  assign n21682 = ~n4338 & n4446 ;
  assign n21683 = n21682 ^ n1374 ^ 1'b0 ;
  assign n21684 = n10365 & n12407 ;
  assign n21685 = ~n21683 & n21684 ;
  assign n21686 = n6913 & ~n21685 ;
  assign n21687 = n12116 & ~n19744 ;
  assign n21688 = n7905 | n9702 ;
  assign n21689 = n5767 | n21688 ;
  assign n21693 = n8198 ^ n1063 ^ 1'b0 ;
  assign n21694 = n6287 & ~n21693 ;
  assign n21695 = n7872 & n21694 ;
  assign n21690 = n619 & ~n5480 ;
  assign n21691 = ( n7117 & n19766 ) | ( n7117 & n21690 ) | ( n19766 & n21690 ) ;
  assign n21692 = n21691 ^ n8343 ^ 1'b0 ;
  assign n21696 = n21695 ^ n21692 ^ 1'b0 ;
  assign n21697 = x137 & ~n21696 ;
  assign n21698 = n1123 ^ n421 ^ 1'b0 ;
  assign n21699 = n3015 & n21698 ;
  assign n21700 = n9736 & ~n12094 ;
  assign n21701 = ~n21699 & n21700 ;
  assign n21702 = n14827 | n21701 ;
  assign n21703 = n21702 ^ n9694 ^ 1'b0 ;
  assign n21704 = n8618 & n21703 ;
  assign n21705 = n9705 & n12374 ;
  assign n21707 = n11061 | n13862 ;
  assign n21708 = n21707 ^ n5254 ^ 1'b0 ;
  assign n21706 = ~n2263 & n8343 ;
  assign n21709 = n21708 ^ n21706 ^ 1'b0 ;
  assign n21710 = n16929 ^ n5153 ^ 1'b0 ;
  assign n21711 = n21709 & ~n21710 ;
  assign n21712 = n9453 ^ n7416 ^ 1'b0 ;
  assign n21713 = n20655 ^ n15502 ^ 1'b0 ;
  assign n21714 = x23 & n1746 ;
  assign n21715 = n21714 ^ n15959 ^ n10324 ;
  assign n21716 = n21715 ^ n12868 ^ 1'b0 ;
  assign n21717 = n12207 & ~n21716 ;
  assign n21718 = ( n14529 & n16042 ) | ( n14529 & ~n21717 ) | ( n16042 & ~n21717 ) ;
  assign n21719 = ~n9277 & n18488 ;
  assign n21720 = n21718 & n21719 ;
  assign n21721 = n13109 ^ n10793 ^ 1'b0 ;
  assign n21722 = n21720 | n21721 ;
  assign n21724 = n5710 & n6046 ;
  assign n21725 = n14107 | n21724 ;
  assign n21723 = n9718 ^ n3145 ^ 1'b0 ;
  assign n21726 = n21725 ^ n21723 ^ n20569 ;
  assign n21727 = n5712 ^ n5245 ^ n2756 ;
  assign n21728 = n1702 & ~n11953 ;
  assign n21729 = ~n7637 & n21728 ;
  assign n21730 = n21729 ^ n17295 ^ n9367 ;
  assign n21731 = n10034 | n21730 ;
  assign n21732 = n14874 ^ n6385 ^ 1'b0 ;
  assign n21733 = n8916 ^ n3688 ^ 1'b0 ;
  assign n21734 = ( ~x144 & n12352 ) | ( ~x144 & n19017 ) | ( n12352 & n19017 ) ;
  assign n21735 = n18668 ^ n14299 ^ 1'b0 ;
  assign n21736 = ( n1629 & n14700 ) | ( n1629 & ~n21735 ) | ( n14700 & ~n21735 ) ;
  assign n21737 = n16830 & n18398 ;
  assign n21738 = n10592 & ~n18897 ;
  assign n21739 = ~n10531 & n21738 ;
  assign n21740 = x246 & n4481 ;
  assign n21741 = ~n13104 & n21740 ;
  assign n21742 = n3180 | n4840 ;
  assign n21743 = n21741 & ~n21742 ;
  assign n21744 = n21743 ^ n17452 ^ n4865 ;
  assign n21745 = ( ~n3056 & n4103 ) | ( ~n3056 & n19689 ) | ( n4103 & n19689 ) ;
  assign n21746 = ~n8263 & n8295 ;
  assign n21747 = n19063 ^ n2453 ^ 1'b0 ;
  assign n21748 = n21746 | n21747 ;
  assign n21749 = n8083 & ~n8858 ;
  assign n21750 = n16424 & n21749 ;
  assign n21751 = n13301 & n21750 ;
  assign n21752 = n2607 & n11419 ;
  assign n21753 = n21752 ^ n6824 ^ 1'b0 ;
  assign n21754 = n8281 & ~n21753 ;
  assign n21755 = n21754 ^ n6479 ^ 1'b0 ;
  assign n21756 = n9721 & n14348 ;
  assign n21757 = n21756 ^ n10162 ^ n5067 ;
  assign n21758 = n21757 ^ n16718 ^ n10102 ;
  assign n21759 = ( ~n580 & n5857 ) | ( ~n580 & n20980 ) | ( n5857 & n20980 ) ;
  assign n21760 = n21759 ^ n8246 ^ n8160 ;
  assign n21761 = n21760 ^ n13267 ^ 1'b0 ;
  assign n21762 = ~n1337 & n2133 ;
  assign n21763 = n21762 ^ n19092 ^ 1'b0 ;
  assign n21764 = n21763 ^ n1709 ^ 1'b0 ;
  assign n21765 = ~n5419 & n21764 ;
  assign n21766 = ( ~n8001 & n10034 ) | ( ~n8001 & n21765 ) | ( n10034 & n21765 ) ;
  assign n21767 = ~n6776 & n7948 ;
  assign n21768 = n11972 & ~n12110 ;
  assign n21769 = n5104 ^ n3742 ^ 1'b0 ;
  assign n21770 = ~n21768 & n21769 ;
  assign n21771 = n6812 & n21770 ;
  assign n21772 = ( n15813 & n21767 ) | ( n15813 & ~n21771 ) | ( n21767 & ~n21771 ) ;
  assign n21773 = n3455 & n10081 ;
  assign n21774 = n21773 ^ n6946 ^ n2106 ;
  assign n21775 = ( ~n21713 & n21772 ) | ( ~n21713 & n21774 ) | ( n21772 & n21774 ) ;
  assign n21777 = n9546 ^ n4943 ^ x175 ;
  assign n21776 = n3732 | n19524 ;
  assign n21778 = n21777 ^ n21776 ^ 1'b0 ;
  assign n21779 = x158 & ~n6415 ;
  assign n21780 = n21779 ^ n3624 ^ 1'b0 ;
  assign n21781 = n11504 | n21780 ;
  assign n21782 = n8448 & n19076 ;
  assign n21783 = n21782 ^ n953 ^ 1'b0 ;
  assign n21784 = n818 | n21783 ;
  assign n21785 = n21784 ^ n12029 ^ n371 ;
  assign n21786 = n11296 ^ n8075 ^ n2453 ;
  assign n21787 = ~n13297 & n21786 ;
  assign n21788 = n21787 ^ n9721 ^ 1'b0 ;
  assign n21789 = n11584 ^ n7380 ^ n3316 ;
  assign n21790 = n21789 ^ n10498 ^ n9875 ;
  assign n21791 = ( n2196 & ~n20334 ) | ( n2196 & n21790 ) | ( ~n20334 & n21790 ) ;
  assign n21792 = x238 & n7022 ;
  assign n21793 = n5179 ^ n1525 ^ n655 ;
  assign n21794 = n21793 ^ n5225 ^ 1'b0 ;
  assign n21795 = n21794 ^ n17175 ^ n4939 ;
  assign n21796 = ( n2787 & n17496 ) | ( n2787 & ~n21795 ) | ( n17496 & ~n21795 ) ;
  assign n21797 = n21792 | n21796 ;
  assign n21798 = n14353 | n21797 ;
  assign n21799 = n16344 & ~n21798 ;
  assign n21800 = ( n16502 & n20785 ) | ( n16502 & ~n21799 ) | ( n20785 & ~n21799 ) ;
  assign n21801 = n12999 & ~n19518 ;
  assign n21802 = n10370 & n21801 ;
  assign n21803 = n3073 ^ n1510 ^ 1'b0 ;
  assign n21804 = n7757 & n21803 ;
  assign n21805 = n21804 ^ n5440 ^ n2674 ;
  assign n21806 = n19483 ^ n12553 ^ 1'b0 ;
  assign n21807 = n21805 & n21806 ;
  assign n21808 = n2392 & ~n5979 ;
  assign n21809 = ~n2392 & n21808 ;
  assign n21810 = n6509 & ~n21809 ;
  assign n21811 = ~n6509 & n21810 ;
  assign n21812 = n21661 | n21811 ;
  assign n21813 = n21661 & ~n21812 ;
  assign n21814 = n1118 | n9743 ;
  assign n21815 = n21813 & ~n21814 ;
  assign n21816 = ~n584 & n5188 ;
  assign n21817 = ~n21815 & n21816 ;
  assign n21818 = n21817 ^ n11035 ^ 1'b0 ;
  assign n21823 = n7039 ^ n4615 ^ x202 ;
  assign n21821 = n7296 & ~n8538 ;
  assign n21822 = ~n17794 & n21821 ;
  assign n21819 = n800 | n16058 ;
  assign n21820 = n14370 & ~n21819 ;
  assign n21824 = n21823 ^ n21822 ^ n21820 ;
  assign n21825 = ( n5206 & n9745 ) | ( n5206 & n16917 ) | ( n9745 & n16917 ) ;
  assign n21826 = ~n6992 & n12443 ;
  assign n21827 = n6024 ^ n5263 ^ 1'b0 ;
  assign n21828 = n21827 ^ n663 ^ 1'b0 ;
  assign n21829 = n4699 & ~n21828 ;
  assign n21830 = n21829 ^ n16512 ^ n14366 ;
  assign n21831 = n21830 ^ n4302 ^ 1'b0 ;
  assign n21832 = n8028 ^ n4369 ^ 1'b0 ;
  assign n21833 = n9424 ^ n8356 ^ 1'b0 ;
  assign n21834 = n21833 ^ n4991 ^ 1'b0 ;
  assign n21835 = n21834 ^ n20233 ^ 1'b0 ;
  assign n21836 = n9241 | n14759 ;
  assign n21837 = n21836 ^ n7326 ^ 1'b0 ;
  assign n21838 = n21837 ^ n14044 ^ n11764 ;
  assign n21839 = n21835 | n21838 ;
  assign n21840 = n4485 & n11471 ;
  assign n21841 = n8143 & ~n21840 ;
  assign n21842 = ~n4661 & n21841 ;
  assign n21843 = n21842 ^ n15724 ^ 1'b0 ;
  assign n21844 = n922 & n18675 ;
  assign n21845 = n11140 & ~n21844 ;
  assign n21846 = n21845 ^ n20963 ^ 1'b0 ;
  assign n21847 = n964 | n20980 ;
  assign n21848 = n19077 | n21847 ;
  assign n21849 = ( n6772 & n9997 ) | ( n6772 & ~n21848 ) | ( n9997 & ~n21848 ) ;
  assign n21850 = n13721 | n16502 ;
  assign n21851 = n13279 & ~n14381 ;
  assign n21852 = n21851 ^ n8863 ^ 1'b0 ;
  assign n21853 = n21850 & n21852 ;
  assign n21854 = n8276 ^ n528 ^ 1'b0 ;
  assign n21855 = n1452 & n21854 ;
  assign n21856 = n21855 ^ n5325 ^ n2547 ;
  assign n21857 = ( n15562 & ~n18102 ) | ( n15562 & n21856 ) | ( ~n18102 & n21856 ) ;
  assign n21858 = n19503 & ~n21857 ;
  assign n21859 = n21858 ^ n6547 ^ 1'b0 ;
  assign n21860 = ( n8865 & n10181 ) | ( n8865 & ~n20043 ) | ( n10181 & ~n20043 ) ;
  assign n21861 = ~n2911 & n5463 ;
  assign n21862 = n21861 ^ n16123 ^ 1'b0 ;
  assign n21863 = n21862 ^ n5413 ^ 1'b0 ;
  assign n21864 = n10551 ^ n9399 ^ n6786 ;
  assign n21865 = n19004 ^ n3105 ^ 1'b0 ;
  assign n21866 = n13043 | n21865 ;
  assign n21867 = n15062 ^ n2709 ^ 1'b0 ;
  assign n21868 = n12874 ^ n4402 ^ 1'b0 ;
  assign n21869 = ( n1586 & n12358 ) | ( n1586 & n21868 ) | ( n12358 & n21868 ) ;
  assign n21870 = n1994 & ~n21869 ;
  assign n21871 = n21870 ^ n14204 ^ 1'b0 ;
  assign n21872 = n7305 & n21871 ;
  assign n21874 = n4506 & ~n9257 ;
  assign n21875 = n21874 ^ n4838 ^ 1'b0 ;
  assign n21873 = ~n19709 & n20448 ;
  assign n21876 = n21875 ^ n21873 ^ 1'b0 ;
  assign n21877 = n21876 ^ n20571 ^ 1'b0 ;
  assign n21878 = n12378 ^ n7745 ^ n4991 ;
  assign n21879 = n20965 ^ n18700 ^ 1'b0 ;
  assign n21880 = ~n1757 & n8632 ;
  assign n21881 = n15397 & n21880 ;
  assign n21882 = n1253 & n3074 ;
  assign n21883 = n3113 & n21882 ;
  assign n21884 = n8834 ^ n3204 ^ n3011 ;
  assign n21885 = n11891 ^ n1630 ^ 1'b0 ;
  assign n21886 = ~n21884 & n21885 ;
  assign n21887 = n21886 ^ n18091 ^ n2573 ;
  assign n21888 = n21887 ^ n6329 ^ n2972 ;
  assign n21889 = n3900 ^ x213 ^ 1'b0 ;
  assign n21890 = n21888 | n21889 ;
  assign n21891 = n15057 | n21890 ;
  assign n21892 = n13104 | n14318 ;
  assign n21895 = n349 | n11010 ;
  assign n21896 = n354 & ~n21895 ;
  assign n21893 = ~n3281 & n5146 ;
  assign n21894 = ~n290 & n21893 ;
  assign n21897 = n21896 ^ n21894 ^ 1'b0 ;
  assign n21898 = n21897 ^ n4997 ^ n4760 ;
  assign n21899 = n21898 ^ n10804 ^ 1'b0 ;
  assign n21900 = ~n21892 & n21899 ;
  assign n21901 = n21900 ^ n5449 ^ 1'b0 ;
  assign n21902 = ~n15288 & n21901 ;
  assign n21903 = n20355 ^ n9513 ^ 1'b0 ;
  assign n21904 = n19044 | n21903 ;
  assign n21905 = n9525 ^ n522 ^ 1'b0 ;
  assign n21906 = n21905 ^ n928 ^ 1'b0 ;
  assign n21907 = n2236 & ~n11659 ;
  assign n21908 = ( n1037 & n3403 ) | ( n1037 & n10500 ) | ( n3403 & n10500 ) ;
  assign n21909 = n16880 | n21908 ;
  assign n21913 = n1351 & ~n10941 ;
  assign n21910 = ~n4890 & n6154 ;
  assign n21911 = n13970 & n21910 ;
  assign n21912 = n20501 & ~n21911 ;
  assign n21914 = n21913 ^ n21912 ^ 1'b0 ;
  assign n21915 = n16441 ^ n14409 ^ n709 ;
  assign n21916 = n957 | n9300 ;
  assign n21917 = n10892 | n21916 ;
  assign n21918 = ( n5867 & n17030 ) | ( n5867 & ~n21917 ) | ( n17030 & ~n21917 ) ;
  assign n21919 = n11680 & ~n18279 ;
  assign n21920 = n21919 ^ n5798 ^ 1'b0 ;
  assign n21921 = n11676 ^ n539 ^ 1'b0 ;
  assign n21922 = n21920 | n21921 ;
  assign n21923 = ( n7836 & n15414 ) | ( n7836 & ~n21922 ) | ( n15414 & ~n21922 ) ;
  assign n21925 = n7847 | n13521 ;
  assign n21926 = n3305 | n21925 ;
  assign n21924 = n9794 | n14145 ;
  assign n21927 = n21926 ^ n21924 ^ 1'b0 ;
  assign n21928 = n7740 ^ n520 ^ 1'b0 ;
  assign n21929 = ~n2945 & n7327 ;
  assign n21930 = ( n19841 & n21928 ) | ( n19841 & n21929 ) | ( n21928 & n21929 ) ;
  assign n21931 = n2628 | n8593 ;
  assign n21932 = n21931 ^ n750 ^ 1'b0 ;
  assign n21933 = n9890 & n12155 ;
  assign n21934 = n21933 ^ n11652 ^ 1'b0 ;
  assign n21935 = ~n21932 & n21934 ;
  assign n21936 = n18268 ^ n3905 ^ 1'b0 ;
  assign n21937 = n6611 ^ n4374 ^ 1'b0 ;
  assign n21938 = n16885 & ~n20634 ;
  assign n21939 = ( n9864 & ~n18445 ) | ( n9864 & n19042 ) | ( ~n18445 & n19042 ) ;
  assign n21940 = n3072 & ~n4173 ;
  assign n21941 = n21940 ^ n20463 ^ 1'b0 ;
  assign n21942 = n6968 & n21941 ;
  assign n21943 = n19063 ^ n16518 ^ n10886 ;
  assign n21944 = ( n550 & n7029 ) | ( n550 & n7210 ) | ( n7029 & n7210 ) ;
  assign n21945 = n21944 ^ n3795 ^ 1'b0 ;
  assign n21946 = ~n21943 & n21945 ;
  assign n21947 = n18421 ^ n14970 ^ 1'b0 ;
  assign n21948 = ~n4471 & n20895 ;
  assign n21949 = ~n4999 & n21948 ;
  assign n21950 = n16644 | n18310 ;
  assign n21951 = n15997 & ~n21950 ;
  assign n21952 = ( n5923 & n21949 ) | ( n5923 & n21951 ) | ( n21949 & n21951 ) ;
  assign n21953 = n8942 ^ n2871 ^ n2742 ;
  assign n21954 = ~n6468 & n21953 ;
  assign n21955 = ~n7289 & n21954 ;
  assign n21956 = n425 & ~n1366 ;
  assign n21957 = ( n2942 & n7380 ) | ( n2942 & n21956 ) | ( n7380 & n21956 ) ;
  assign n21958 = n10116 ^ n9121 ^ 1'b0 ;
  assign n21959 = n21957 & ~n21958 ;
  assign n21960 = ( n1088 & ~n9562 ) | ( n1088 & n14874 ) | ( ~n9562 & n14874 ) ;
  assign n21961 = ~n1688 & n6645 ;
  assign n21963 = n785 | n21956 ;
  assign n21962 = ~n4264 & n11909 ;
  assign n21964 = n21963 ^ n21962 ^ n3252 ;
  assign n21965 = n8093 ^ n6992 ^ n5582 ;
  assign n21966 = n8296 ^ n5106 ^ n2147 ;
  assign n21967 = n15737 ^ n14451 ^ 1'b0 ;
  assign n21968 = ( n9875 & n21963 ) | ( n9875 & ~n21967 ) | ( n21963 & ~n21967 ) ;
  assign n21969 = n21968 ^ n13949 ^ 1'b0 ;
  assign n21970 = n3605 & n21969 ;
  assign n21971 = n13892 ^ n9182 ^ 1'b0 ;
  assign n21972 = n5313 & n21971 ;
  assign n21973 = n21972 ^ n15572 ^ 1'b0 ;
  assign n21974 = ( n21966 & n21970 ) | ( n21966 & ~n21973 ) | ( n21970 & ~n21973 ) ;
  assign n21975 = ~n2064 & n13886 ;
  assign n21976 = ~n11445 & n18721 ;
  assign n21977 = n21976 ^ n19709 ^ 1'b0 ;
  assign n21978 = ( ~x157 & n1713 ) | ( ~x157 & n7520 ) | ( n1713 & n7520 ) ;
  assign n21979 = n20162 & n21978 ;
  assign n21980 = n21979 ^ n3329 ^ 1'b0 ;
  assign n21981 = n21980 ^ n13895 ^ 1'b0 ;
  assign n21982 = x77 & ~n12385 ;
  assign n21983 = ~n6717 & n17823 ;
  assign n21984 = ( n6356 & n21982 ) | ( n6356 & n21983 ) | ( n21982 & n21983 ) ;
  assign n21985 = ~n7545 & n9258 ;
  assign n21986 = n8106 ^ n578 ^ 1'b0 ;
  assign n21987 = ~n15936 & n21986 ;
  assign n21988 = n709 & n5612 ;
  assign n21989 = ~n4736 & n21988 ;
  assign n21990 = n358 | n9295 ;
  assign n21991 = n21989 & ~n21990 ;
  assign n21992 = n21991 ^ n19381 ^ 1'b0 ;
  assign n21993 = ~n14863 & n15879 ;
  assign n21994 = n21993 ^ n14230 ^ 1'b0 ;
  assign n21995 = n15451 & n21994 ;
  assign n21996 = n7388 ^ n522 ^ 1'b0 ;
  assign n21997 = n1379 & ~n21996 ;
  assign n21998 = ( n1941 & n17346 ) | ( n1941 & ~n21997 ) | ( n17346 & ~n21997 ) ;
  assign n21999 = n21998 ^ n5897 ^ 1'b0 ;
  assign n22000 = ~n2948 & n7001 ;
  assign n22001 = n22000 ^ n17519 ^ 1'b0 ;
  assign n22002 = ( n7471 & ~n8717 ) | ( n7471 & n22001 ) | ( ~n8717 & n22001 ) ;
  assign n22003 = n22002 ^ n7959 ^ 1'b0 ;
  assign n22004 = ( ~n2435 & n15107 ) | ( ~n2435 & n18217 ) | ( n15107 & n18217 ) ;
  assign n22005 = n4198 & n22004 ;
  assign n22006 = n22005 ^ n9672 ^ 1'b0 ;
  assign n22007 = n20878 | n22006 ;
  assign n22008 = n718 & ~n21506 ;
  assign n22009 = n18643 ^ n860 ^ 1'b0 ;
  assign n22010 = n2970 & ~n16735 ;
  assign n22011 = n9468 | n15890 ;
  assign n22012 = n22011 ^ n7942 ^ 1'b0 ;
  assign n22013 = n6071 & ~n22012 ;
  assign n22014 = n22013 ^ n18084 ^ 1'b0 ;
  assign n22015 = n14133 | n21331 ;
  assign n22016 = n14840 & n16380 ;
  assign n22017 = n7448 & ~n11908 ;
  assign n22018 = n17389 & n22017 ;
  assign n22019 = n8815 & n22018 ;
  assign n22020 = n22016 & ~n22019 ;
  assign n22021 = n15856 ^ n3580 ^ 1'b0 ;
  assign n22022 = n5432 & n6776 ;
  assign n22023 = n4493 & ~n21656 ;
  assign n22024 = n21574 ^ n11023 ^ n9321 ;
  assign n22025 = n11495 ^ n6253 ^ 1'b0 ;
  assign n22026 = n21607 ^ n18086 ^ 1'b0 ;
  assign n22027 = n19744 & n22026 ;
  assign n22028 = n6256 | n11747 ;
  assign n22029 = n562 | n22028 ;
  assign n22030 = ( ~n968 & n8106 ) | ( ~n968 & n22029 ) | ( n8106 & n22029 ) ;
  assign n22031 = n13170 ^ n5996 ^ 1'b0 ;
  assign n22032 = n21275 ^ n15562 ^ 1'b0 ;
  assign n22033 = ( n10055 & n15988 ) | ( n10055 & n20958 ) | ( n15988 & n20958 ) ;
  assign n22042 = n10918 & n12429 ;
  assign n22043 = n22042 ^ n4650 ^ 1'b0 ;
  assign n22044 = ( n5451 & n7293 ) | ( n5451 & ~n22043 ) | ( n7293 & ~n22043 ) ;
  assign n22036 = n5582 ^ n256 ^ 1'b0 ;
  assign n22037 = n680 & n22036 ;
  assign n22038 = ~n16812 & n22037 ;
  assign n22034 = ~n696 & n6127 ;
  assign n22035 = n22034 ^ n3924 ^ 1'b0 ;
  assign n22039 = n22038 ^ n22035 ^ 1'b0 ;
  assign n22040 = ~n20271 & n22039 ;
  assign n22041 = n7442 & n22040 ;
  assign n22045 = n22044 ^ n22041 ^ 1'b0 ;
  assign n22046 = n19087 ^ n13940 ^ 1'b0 ;
  assign n22047 = n14397 & ~n22046 ;
  assign n22050 = n10763 ^ n6275 ^ n6075 ;
  assign n22051 = ( ~n3255 & n6465 ) | ( ~n3255 & n22050 ) | ( n6465 & n22050 ) ;
  assign n22048 = n21085 ^ n14235 ^ n2782 ;
  assign n22049 = n14886 | n22048 ;
  assign n22052 = n22051 ^ n22049 ^ 1'b0 ;
  assign n22053 = n717 & n20271 ;
  assign n22054 = n22053 ^ n18262 ^ n7863 ;
  assign n22055 = n339 & ~n16860 ;
  assign n22056 = n22055 ^ n14416 ^ 1'b0 ;
  assign n22057 = n6681 & ~n22056 ;
  assign n22058 = ~n21359 & n22057 ;
  assign n22059 = n860 | n2052 ;
  assign n22060 = n22059 ^ n13295 ^ 1'b0 ;
  assign n22061 = n455 | n22060 ;
  assign n22062 = ~n1898 & n8697 ;
  assign n22063 = n22061 | n22062 ;
  assign n22064 = n22063 ^ n10990 ^ 1'b0 ;
  assign n22065 = n2035 & n4258 ;
  assign n22066 = n8321 | n22065 ;
  assign n22067 = n20470 ^ n18525 ^ 1'b0 ;
  assign n22068 = n13454 ^ n8440 ^ 1'b0 ;
  assign n22069 = n8941 & ~n22068 ;
  assign n22070 = n8538 & ~n13862 ;
  assign n22071 = n10472 | n18836 ;
  assign n22072 = n22070 & ~n22071 ;
  assign n22073 = n22072 ^ n13320 ^ 1'b0 ;
  assign n22074 = ~n6994 & n22073 ;
  assign n22075 = n7880 ^ n2036 ^ 1'b0 ;
  assign n22076 = ~n7378 & n22075 ;
  assign n22077 = n22076 ^ n7803 ^ n6461 ;
  assign n22078 = n9892 & ~n12041 ;
  assign n22079 = n7434 ^ n704 ^ 1'b0 ;
  assign n22080 = ~n5882 & n16967 ;
  assign n22081 = n866 & ~n11635 ;
  assign n22082 = n22081 ^ n11860 ^ 1'b0 ;
  assign n22083 = n20723 ^ n10388 ^ 1'b0 ;
  assign n22084 = ~n12023 & n22083 ;
  assign n22085 = n22084 ^ n16991 ^ n14906 ;
  assign n22086 = n10600 ^ n9020 ^ n5226 ;
  assign n22087 = n18531 ^ n3024 ^ 1'b0 ;
  assign n22088 = n4578 ^ n1976 ^ n295 ;
  assign n22089 = n6172 & ~n22088 ;
  assign n22090 = n22089 ^ n15379 ^ 1'b0 ;
  assign n22091 = n9276 | n15710 ;
  assign n22092 = n1173 | n22091 ;
  assign n22093 = n22090 & n22092 ;
  assign n22094 = n20967 & n22093 ;
  assign n22095 = n10924 ^ n5285 ^ 1'b0 ;
  assign n22096 = ~n3909 & n22095 ;
  assign n22097 = n8639 | n13857 ;
  assign n22098 = n3904 & ~n19668 ;
  assign n22099 = ( n5296 & n9664 ) | ( n5296 & n22098 ) | ( n9664 & n22098 ) ;
  assign n22100 = n22099 ^ n1711 ^ 1'b0 ;
  assign n22101 = n3679 | n22100 ;
  assign n22102 = ( n6091 & n6515 ) | ( n6091 & ~n7066 ) | ( n6515 & ~n7066 ) ;
  assign n22103 = x57 & ~n4947 ;
  assign n22104 = n22103 ^ n16979 ^ 1'b0 ;
  assign n22105 = n22104 ^ n1217 ^ 1'b0 ;
  assign n22106 = n22102 & ~n22105 ;
  assign n22107 = n1368 | n9439 ;
  assign n22108 = ( n13041 & ~n15230 ) | ( n13041 & n22107 ) | ( ~n15230 & n22107 ) ;
  assign n22109 = n22108 ^ n20648 ^ 1'b0 ;
  assign n22110 = x221 & n22109 ;
  assign n22111 = ~n2701 & n6771 ;
  assign n22112 = n22111 ^ n3110 ^ 1'b0 ;
  assign n22113 = ~n7395 & n22112 ;
  assign n22114 = n12615 ^ n8294 ^ 1'b0 ;
  assign n22115 = n16358 ^ n12423 ^ n4879 ;
  assign n22126 = n7373 | n14223 ;
  assign n22127 = n22126 ^ n9803 ^ 1'b0 ;
  assign n22116 = ~n5257 & n7657 ;
  assign n22117 = n22116 ^ n6773 ^ 1'b0 ;
  assign n22118 = ~n19736 & n22117 ;
  assign n22119 = n4664 & n22118 ;
  assign n22120 = n22119 ^ n13588 ^ 1'b0 ;
  assign n22121 = n8553 & ~n11112 ;
  assign n22122 = ~n21782 & n22121 ;
  assign n22123 = n8606 & n22122 ;
  assign n22124 = n22123 ^ n14805 ^ 1'b0 ;
  assign n22125 = n22120 | n22124 ;
  assign n22128 = n22127 ^ n22125 ^ 1'b0 ;
  assign n22130 = n7540 ^ n3836 ^ 1'b0 ;
  assign n22131 = n1749 & n22130 ;
  assign n22129 = n5698 | n15246 ;
  assign n22132 = n22131 ^ n22129 ^ 1'b0 ;
  assign n22133 = n22132 ^ n21289 ^ n1944 ;
  assign n22134 = n10426 ^ n5655 ^ 1'b0 ;
  assign n22135 = n7537 & n22134 ;
  assign n22136 = n18948 ^ n3666 ^ 1'b0 ;
  assign n22137 = ~n21492 & n22136 ;
  assign n22138 = n7159 & n12839 ;
  assign n22139 = n22138 ^ n2001 ^ 1'b0 ;
  assign n22140 = n11982 ^ n9431 ^ n4265 ;
  assign n22141 = n22140 ^ n16422 ^ n7051 ;
  assign n22142 = x10 | n5679 ;
  assign n22143 = n8186 ^ n4130 ^ 1'b0 ;
  assign n22144 = ~n2504 & n22143 ;
  assign n22145 = n6558 & n22144 ;
  assign n22146 = n2637 & n3868 ;
  assign n22147 = ( n8900 & n17667 ) | ( n8900 & ~n22146 ) | ( n17667 & ~n22146 ) ;
  assign n22148 = ( n7854 & n11240 ) | ( n7854 & n22147 ) | ( n11240 & n22147 ) ;
  assign n22149 = n22148 ^ n8460 ^ 1'b0 ;
  assign n22155 = n19511 ^ n17553 ^ n5768 ;
  assign n22150 = n4829 ^ x123 ^ 1'b0 ;
  assign n22151 = n11712 | n22150 ;
  assign n22152 = n22151 ^ n1055 ^ 1'b0 ;
  assign n22153 = n2325 & n8756 ;
  assign n22154 = ~n22152 & n22153 ;
  assign n22156 = n22155 ^ n22154 ^ 1'b0 ;
  assign n22157 = n1778 & ~n22156 ;
  assign n22158 = n5203 & ~n7848 ;
  assign n22159 = ~n18960 & n22158 ;
  assign n22160 = n282 & ~n22159 ;
  assign n22161 = n22160 ^ n19921 ^ 1'b0 ;
  assign n22162 = n10775 & n22161 ;
  assign n22163 = ( ~n3628 & n5460 ) | ( ~n3628 & n5792 ) | ( n5460 & n5792 ) ;
  assign n22164 = ( n4696 & n7488 ) | ( n4696 & n22163 ) | ( n7488 & n22163 ) ;
  assign n22165 = ~n13592 & n19685 ;
  assign n22166 = n22165 ^ n14478 ^ n5014 ;
  assign n22169 = n9928 & n19163 ;
  assign n22170 = ~n6878 & n22169 ;
  assign n22167 = n6436 ^ n2478 ^ n637 ;
  assign n22168 = n22167 ^ n19124 ^ 1'b0 ;
  assign n22171 = n22170 ^ n22168 ^ n5824 ;
  assign n22172 = n15154 ^ n10108 ^ 1'b0 ;
  assign n22175 = n12284 ^ n600 ^ 1'b0 ;
  assign n22173 = n20399 ^ n12193 ^ n1288 ;
  assign n22174 = ~n11692 & n22173 ;
  assign n22176 = n22175 ^ n22174 ^ 1'b0 ;
  assign n22177 = n22172 & ~n22176 ;
  assign n22183 = n1482 ^ n1479 ^ 1'b0 ;
  assign n22184 = n5155 | n22183 ;
  assign n22178 = n16635 ^ n9643 ^ 1'b0 ;
  assign n22179 = ( n2349 & n10764 ) | ( n2349 & ~n13215 ) | ( n10764 & ~n13215 ) ;
  assign n22180 = n16898 & ~n22179 ;
  assign n22181 = n22180 ^ n15068 ^ 1'b0 ;
  assign n22182 = n22178 | n22181 ;
  assign n22185 = n22184 ^ n22182 ^ 1'b0 ;
  assign n22186 = n4694 ^ n3274 ^ 1'b0 ;
  assign n22187 = ~n4882 & n20012 ;
  assign n22188 = n22187 ^ n15953 ^ 1'b0 ;
  assign n22189 = ( n4257 & ~n13881 ) | ( n4257 & n15165 ) | ( ~n13881 & n15165 ) ;
  assign n22190 = n6167 ^ n4195 ^ n314 ;
  assign n22191 = ~n2680 & n6433 ;
  assign n22192 = n22190 & n22191 ;
  assign n22193 = n6034 & n22192 ;
  assign n22194 = x136 & n9174 ;
  assign n22195 = n22194 ^ n2538 ^ 1'b0 ;
  assign n22196 = n18166 ^ n11909 ^ 1'b0 ;
  assign n22197 = n19677 & n22196 ;
  assign n22198 = ~n6769 & n19558 ;
  assign n22199 = ( n4055 & n11426 ) | ( n4055 & ~n17771 ) | ( n11426 & ~n17771 ) ;
  assign n22203 = ~n1262 & n11426 ;
  assign n22200 = n2372 & ~n3238 ;
  assign n22201 = n22200 ^ n4103 ^ 1'b0 ;
  assign n22202 = n7361 & n22201 ;
  assign n22204 = n22203 ^ n22202 ^ 1'b0 ;
  assign n22205 = ( n879 & ~n16031 ) | ( n879 & n19862 ) | ( ~n16031 & n19862 ) ;
  assign n22206 = n14997 ^ n1940 ^ 1'b0 ;
  assign n22207 = n8124 | n22206 ;
  assign n22208 = n8261 | n10135 ;
  assign n22209 = n2471 & ~n6306 ;
  assign n22210 = n22208 | n22209 ;
  assign n22211 = n22210 ^ n21074 ^ 1'b0 ;
  assign n22212 = n16234 & ~n22211 ;
  assign n22213 = n21983 ^ n2267 ^ n1538 ;
  assign n22217 = n12720 & ~n15402 ;
  assign n22218 = ~n1253 & n22217 ;
  assign n22216 = n7140 ^ x149 ^ x131 ;
  assign n22214 = n15704 ^ n7586 ^ 1'b0 ;
  assign n22215 = n1458 & ~n22214 ;
  assign n22219 = n22218 ^ n22216 ^ n22215 ;
  assign n22220 = n1285 & n10369 ;
  assign n22221 = n15575 & n22220 ;
  assign n22222 = n16083 ^ n629 ^ 1'b0 ;
  assign n22223 = n10220 & n22222 ;
  assign n22224 = x51 & n22223 ;
  assign n22225 = n22221 & n22224 ;
  assign n22226 = ( n4869 & n8252 ) | ( n4869 & n14128 ) | ( n8252 & n14128 ) ;
  assign n22227 = n22226 ^ n8762 ^ n6870 ;
  assign n22228 = n15083 & n22227 ;
  assign n22229 = n22228 ^ n3628 ^ 1'b0 ;
  assign n22230 = ( ~n1607 & n7758 ) | ( ~n1607 & n8958 ) | ( n7758 & n8958 ) ;
  assign n22231 = n22230 ^ n18049 ^ 1'b0 ;
  assign n22232 = ~n2845 & n4891 ;
  assign n22233 = n8748 & n22232 ;
  assign n22234 = ( ~n9058 & n15040 ) | ( ~n9058 & n18776 ) | ( n15040 & n18776 ) ;
  assign n22235 = n19325 ^ n13501 ^ n10646 ;
  assign n22236 = n7447 ^ n6534 ^ n2852 ;
  assign n22237 = n12565 & ~n22236 ;
  assign n22238 = n22237 ^ n2389 ^ 1'b0 ;
  assign n22239 = n15512 ^ n15482 ^ 1'b0 ;
  assign n22240 = n1264 & n22239 ;
  assign n22241 = ~n3835 & n13341 ;
  assign n22242 = n22241 ^ n16415 ^ 1'b0 ;
  assign n22243 = n17845 ^ n12676 ^ 1'b0 ;
  assign n22244 = ~n2261 & n22243 ;
  assign n22245 = n16638 ^ n11733 ^ 1'b0 ;
  assign n22246 = n1716 & n22245 ;
  assign n22247 = n2260 & n19115 ;
  assign n22250 = n10002 & n12358 ;
  assign n22248 = ~n2874 & n16340 ;
  assign n22249 = n6522 & n22248 ;
  assign n22251 = n22250 ^ n22249 ^ 1'b0 ;
  assign n22252 = n3736 & n8419 ;
  assign n22253 = n22252 ^ n469 ^ 1'b0 ;
  assign n22257 = x77 & ~n7691 ;
  assign n22258 = ( n2882 & n3540 ) | ( n2882 & n16580 ) | ( n3540 & n16580 ) ;
  assign n22259 = n9656 & ~n22258 ;
  assign n22260 = n19176 ^ n7591 ^ 1'b0 ;
  assign n22261 = ~n22259 & n22260 ;
  assign n22262 = ~n22257 & n22261 ;
  assign n22254 = n3540 & ~n4013 ;
  assign n22255 = n4405 ^ n783 ^ 1'b0 ;
  assign n22256 = n22254 & ~n22255 ;
  assign n22263 = n22262 ^ n22256 ^ n9230 ;
  assign n22264 = n13357 ^ n5244 ^ n2071 ;
  assign n22265 = n22264 ^ n5815 ^ 1'b0 ;
  assign n22266 = n17549 ^ n3517 ^ 1'b0 ;
  assign n22268 = n3593 & n20630 ;
  assign n22269 = ~n4825 & n22268 ;
  assign n22267 = n15050 ^ n8204 ^ n4458 ;
  assign n22270 = n22269 ^ n22267 ^ n14238 ;
  assign n22271 = ( n6580 & n8765 ) | ( n6580 & n21205 ) | ( n8765 & n21205 ) ;
  assign n22272 = n5844 & ~n18371 ;
  assign n22273 = ( n13391 & ~n18057 ) | ( n13391 & n18482 ) | ( ~n18057 & n18482 ) ;
  assign n22274 = n6129 ^ n4487 ^ 1'b0 ;
  assign n22275 = n8732 ^ n1285 ^ 1'b0 ;
  assign n22276 = n19580 & n22275 ;
  assign n22280 = n9037 & ~n14998 ;
  assign n22277 = n14648 ^ n6705 ^ 1'b0 ;
  assign n22278 = n1356 | n22277 ;
  assign n22279 = n2200 | n22278 ;
  assign n22281 = n22280 ^ n22279 ^ 1'b0 ;
  assign n22283 = ~n8783 & n14191 ;
  assign n22284 = n8155 & n22283 ;
  assign n22282 = ( n5665 & n8461 ) | ( n5665 & ~n17041 ) | ( n8461 & ~n17041 ) ;
  assign n22285 = n22284 ^ n22282 ^ n13030 ;
  assign n22286 = ~n501 & n6447 ;
  assign n22287 = n5058 & n22286 ;
  assign n22288 = n22287 ^ n8409 ^ n2152 ;
  assign n22289 = ( n4273 & n9422 ) | ( n4273 & n10463 ) | ( n9422 & n10463 ) ;
  assign n22294 = n735 ^ n665 ^ 1'b0 ;
  assign n22290 = ~n1501 & n4938 ;
  assign n22291 = ~n6373 & n22290 ;
  assign n22292 = n7584 ^ n7070 ^ 1'b0 ;
  assign n22293 = ( n2565 & n22291 ) | ( n2565 & n22292 ) | ( n22291 & n22292 ) ;
  assign n22295 = n22294 ^ n22293 ^ 1'b0 ;
  assign n22296 = ~n22289 & n22295 ;
  assign n22297 = n22288 & ~n22296 ;
  assign n22298 = n22297 ^ n3157 ^ 1'b0 ;
  assign n22299 = ( ~n282 & n8496 ) | ( ~n282 & n8664 ) | ( n8496 & n8664 ) ;
  assign n22300 = ( ~n7676 & n15604 ) | ( ~n7676 & n22299 ) | ( n15604 & n22299 ) ;
  assign n22301 = n6071 & n15153 ;
  assign n22302 = n22301 ^ n17705 ^ 1'b0 ;
  assign n22303 = ~n12348 & n13295 ;
  assign n22304 = ~n12449 & n22303 ;
  assign n22305 = n22304 ^ n10836 ^ n7127 ;
  assign n22306 = ( ~n5660 & n7168 ) | ( ~n5660 & n12222 ) | ( n7168 & n12222 ) ;
  assign n22307 = n22306 ^ n16099 ^ 1'b0 ;
  assign n22308 = n9638 | n22307 ;
  assign n22309 = n6149 ^ n5901 ^ n5265 ;
  assign n22310 = ( n2459 & n8705 ) | ( n2459 & ~n13619 ) | ( n8705 & ~n13619 ) ;
  assign n22311 = n22310 ^ n20275 ^ n3977 ;
  assign n22312 = n6742 & ~n22311 ;
  assign n22313 = ~n22309 & n22312 ;
  assign n22314 = ~n5515 & n14618 ;
  assign n22315 = n11336 & n22314 ;
  assign n22316 = n22315 ^ n15440 ^ 1'b0 ;
  assign n22317 = n18993 | n22316 ;
  assign n22318 = n8762 ^ n5302 ^ n1164 ;
  assign n22319 = n15449 ^ n6652 ^ n6111 ;
  assign n22320 = n17989 ^ n4155 ^ 1'b0 ;
  assign n22321 = ( n1064 & ~n10896 ) | ( n1064 & n22320 ) | ( ~n10896 & n22320 ) ;
  assign n22322 = ~n294 & n22321 ;
  assign n22323 = ~x148 & n1787 ;
  assign n22324 = n22322 & ~n22323 ;
  assign n22325 = n4454 | n8466 ;
  assign n22326 = n22325 ^ n16221 ^ n6170 ;
  assign n22327 = n22326 ^ n13715 ^ 1'b0 ;
  assign n22328 = ~n13370 & n22327 ;
  assign n22329 = ~n3742 & n12912 ;
  assign n22330 = n22329 ^ n4701 ^ 1'b0 ;
  assign n22331 = n5815 | n14058 ;
  assign n22332 = n22330 & ~n22331 ;
  assign n22334 = n15370 ^ n9336 ^ 1'b0 ;
  assign n22335 = ( n10801 & ~n17912 ) | ( n10801 & n22334 ) | ( ~n17912 & n22334 ) ;
  assign n22333 = ~n1740 & n10480 ;
  assign n22336 = n22335 ^ n22333 ^ 1'b0 ;
  assign n22337 = n15493 ^ n1162 ^ n327 ;
  assign n22338 = n20992 ^ n6001 ^ n4679 ;
  assign n22339 = n22338 ^ n3999 ^ 1'b0 ;
  assign n22340 = n22337 | n22339 ;
  assign n22341 = n22340 ^ n6515 ^ 1'b0 ;
  assign n22342 = n20284 | n22341 ;
  assign n22343 = ~n3730 & n6457 ;
  assign n22344 = n20381 ^ n16413 ^ n6894 ;
  assign n22345 = ( n9148 & n19590 ) | ( n9148 & n20879 ) | ( n19590 & n20879 ) ;
  assign n22346 = ( n3974 & ~n5426 ) | ( n3974 & n5466 ) | ( ~n5426 & n5466 ) ;
  assign n22347 = n423 & ~n22346 ;
  assign n22348 = n22347 ^ n17840 ^ n1938 ;
  assign n22349 = n1392 & n1856 ;
  assign n22350 = ~n4628 & n22349 ;
  assign n22351 = n22350 ^ n2433 ^ 1'b0 ;
  assign n22352 = n22351 ^ n15677 ^ n11620 ;
  assign n22353 = n13798 ^ n7821 ^ 1'b0 ;
  assign n22354 = n12079 & ~n22353 ;
  assign n22355 = n2052 | n11842 ;
  assign n22356 = ~n9022 & n22355 ;
  assign n22357 = ~n22354 & n22356 ;
  assign n22358 = n18072 ^ n12140 ^ n10757 ;
  assign n22359 = n11967 & n22358 ;
  assign n22360 = n16218 ^ n15677 ^ 1'b0 ;
  assign n22361 = ~n933 & n22360 ;
  assign n22362 = ~n10032 & n22361 ;
  assign n22363 = n14050 | n20924 ;
  assign n22364 = n21283 ^ n13057 ^ 1'b0 ;
  assign n22365 = n8858 ^ n5405 ^ 1'b0 ;
  assign n22366 = n20248 ^ n3546 ^ 1'b0 ;
  assign n22367 = ~n22365 & n22366 ;
  assign n22368 = n9331 & ~n17505 ;
  assign n22369 = n22368 ^ n9702 ^ 1'b0 ;
  assign n22370 = n12983 ^ n1022 ^ 1'b0 ;
  assign n22371 = n3572 & n10304 ;
  assign n22372 = n22371 ^ n12404 ^ n3476 ;
  assign n22373 = n22372 ^ n21580 ^ n20433 ;
  assign n22374 = ( n20479 & n21635 ) | ( n20479 & ~n22373 ) | ( n21635 & ~n22373 ) ;
  assign n22375 = n3576 & ~n15511 ;
  assign n22376 = n22375 ^ n17827 ^ 1'b0 ;
  assign n22377 = ( n9015 & n12272 ) | ( n9015 & n16128 ) | ( n12272 & n16128 ) ;
  assign n22378 = n8177 | n22377 ;
  assign n22379 = n1118 & ~n22378 ;
  assign n22381 = ( n2670 & n2989 ) | ( n2670 & n12585 ) | ( n2989 & n12585 ) ;
  assign n22380 = n6944 & ~n8521 ;
  assign n22382 = n22381 ^ n22380 ^ 1'b0 ;
  assign n22383 = n19445 ^ n4260 ^ 1'b0 ;
  assign n22384 = x183 & n22383 ;
  assign n22385 = n22384 ^ n22296 ^ n12722 ;
  assign n22389 = n13511 ^ n7395 ^ 1'b0 ;
  assign n22386 = ( n2357 & ~n5211 ) | ( n2357 & n7288 ) | ( ~n5211 & n7288 ) ;
  assign n22387 = n22386 ^ n615 ^ 1'b0 ;
  assign n22388 = n2606 & ~n22387 ;
  assign n22390 = n22389 ^ n22388 ^ 1'b0 ;
  assign n22391 = ( x210 & ~n9834 ) | ( x210 & n22390 ) | ( ~n9834 & n22390 ) ;
  assign n22392 = n10998 & ~n13949 ;
  assign n22393 = ~n5365 & n22392 ;
  assign n22394 = n22393 ^ n3742 ^ 1'b0 ;
  assign n22395 = ~n12579 & n22394 ;
  assign n22396 = n6608 & n21831 ;
  assign n22397 = n2504 | n17607 ;
  assign n22398 = n8934 | n22397 ;
  assign n22399 = ~n4448 & n22398 ;
  assign n22400 = n14711 & n22399 ;
  assign n22401 = ~n12885 & n14178 ;
  assign n22402 = ~n6149 & n22401 ;
  assign n22403 = n520 | n974 ;
  assign n22404 = n22403 ^ n5744 ^ 1'b0 ;
  assign n22405 = n6908 | n22404 ;
  assign n22406 = n17921 | n22405 ;
  assign n22407 = n8623 & n22406 ;
  assign n22408 = n14791 & n22407 ;
  assign n22409 = ( n20226 & n20262 ) | ( n20226 & n22408 ) | ( n20262 & n22408 ) ;
  assign n22410 = n7547 ^ n6105 ^ 1'b0 ;
  assign n22411 = n10130 & ~n22410 ;
  assign n22412 = n22411 ^ n14543 ^ 1'b0 ;
  assign n22413 = ~n1707 & n4857 ;
  assign n22414 = n4416 & n22413 ;
  assign n22415 = n22414 ^ n1829 ^ 1'b0 ;
  assign n22416 = ~n16250 & n22415 ;
  assign n22417 = n22412 & n22416 ;
  assign n22418 = n21033 | n22417 ;
  assign n22419 = n22418 ^ n16468 ^ 1'b0 ;
  assign n22420 = n21202 ^ n7465 ^ n5798 ;
  assign n22421 = n18082 & n22420 ;
  assign n22422 = n6065 & n22421 ;
  assign n22423 = n8394 ^ n2490 ^ 1'b0 ;
  assign n22424 = n10086 & ~n11583 ;
  assign n22425 = x169 & n22424 ;
  assign n22426 = n22425 ^ n11883 ^ 1'b0 ;
  assign n22427 = n22423 | n22426 ;
  assign n22428 = n17471 ^ n14519 ^ 1'b0 ;
  assign n22429 = n654 & ~n1661 ;
  assign n22430 = n3910 & n22429 ;
  assign n22431 = n2574 | n6485 ;
  assign n22432 = ~n22430 & n22431 ;
  assign n22433 = ~n1369 & n4140 ;
  assign n22434 = n5588 & n22433 ;
  assign n22435 = n22434 ^ n17365 ^ n5377 ;
  assign n22436 = ( n20852 & ~n22432 ) | ( n20852 & n22435 ) | ( ~n22432 & n22435 ) ;
  assign n22437 = n5740 | n11318 ;
  assign n22438 = n14651 & ~n22437 ;
  assign n22439 = n18550 & ~n22438 ;
  assign n22440 = n13923 & ~n18041 ;
  assign n22441 = n22440 ^ n4104 ^ 1'b0 ;
  assign n22442 = ~n12382 & n22441 ;
  assign n22443 = n22442 ^ n5933 ^ 1'b0 ;
  assign n22444 = n22439 | n22443 ;
  assign n22445 = n8280 ^ n6820 ^ 1'b0 ;
  assign n22446 = n20805 ^ n391 ^ 1'b0 ;
  assign n22447 = n1489 & ~n22446 ;
  assign n22448 = n10636 ^ n1459 ^ 1'b0 ;
  assign n22449 = n18285 | n22448 ;
  assign n22450 = ~n1022 & n4724 ;
  assign n22451 = n22450 ^ n6913 ^ 1'b0 ;
  assign n22452 = n1613 | n10157 ;
  assign n22453 = ~n21050 & n22452 ;
  assign n22454 = n22453 ^ n19696 ^ 1'b0 ;
  assign n22455 = n13754 | n22454 ;
  assign n22456 = ( n4592 & n22451 ) | ( n4592 & n22455 ) | ( n22451 & n22455 ) ;
  assign n22457 = n19175 ^ n8752 ^ 1'b0 ;
  assign n22458 = ~n20248 & n22457 ;
  assign n22459 = n6191 ^ n542 ^ 1'b0 ;
  assign n22460 = n18008 | n22459 ;
  assign n22461 = n22460 ^ n20921 ^ n8323 ;
  assign n22462 = n14041 ^ n10401 ^ 1'b0 ;
  assign n22463 = ( n7806 & n19628 ) | ( n7806 & n22462 ) | ( n19628 & n22462 ) ;
  assign n22464 = n18094 ^ n13524 ^ 1'b0 ;
  assign n22465 = n21508 & ~n22464 ;
  assign n22466 = ~n13073 & n22465 ;
  assign n22467 = n13363 ^ n4673 ^ n4091 ;
  assign n22468 = n17566 & ~n22467 ;
  assign n22469 = n15759 ^ x24 ^ 1'b0 ;
  assign n22470 = n22469 ^ n13618 ^ n2840 ;
  assign n22471 = n22470 ^ n22216 ^ 1'b0 ;
  assign n22472 = n9516 ^ n6312 ^ 1'b0 ;
  assign n22473 = n8422 & ~n9070 ;
  assign n22474 = n22472 & n22473 ;
  assign n22479 = ( x197 & ~n11187 ) | ( x197 & n16413 ) | ( ~n11187 & n16413 ) ;
  assign n22475 = n2476 & ~n11291 ;
  assign n22476 = n2183 & n22475 ;
  assign n22477 = ~n11807 & n12870 ;
  assign n22478 = n22476 & n22477 ;
  assign n22480 = n22479 ^ n22478 ^ 1'b0 ;
  assign n22481 = n17537 | n22480 ;
  assign n22482 = n8027 ^ n1586 ^ 1'b0 ;
  assign n22483 = n5043 | n22482 ;
  assign n22484 = n5734 & ~n16907 ;
  assign n22485 = n12721 ^ n12514 ^ n517 ;
  assign n22486 = n1884 & ~n7910 ;
  assign n22487 = ( n6784 & ~n16512 ) | ( n6784 & n22486 ) | ( ~n16512 & n22486 ) ;
  assign n22488 = n22487 ^ n12875 ^ n5492 ;
  assign n22489 = ( ~n16898 & n22485 ) | ( ~n16898 & n22488 ) | ( n22485 & n22488 ) ;
  assign n22490 = n4592 & n13896 ;
  assign n22491 = n14232 ^ n672 ^ 1'b0 ;
  assign n22492 = ( n7936 & ~n22490 ) | ( n7936 & n22491 ) | ( ~n22490 & n22491 ) ;
  assign n22493 = n16508 ^ n8858 ^ 1'b0 ;
  assign n22494 = n9426 & ~n22493 ;
  assign n22495 = x172 & ~n13844 ;
  assign n22496 = n8263 & n22495 ;
  assign n22497 = n12775 & n22496 ;
  assign n22498 = ~n12478 & n22497 ;
  assign n22499 = ( n2342 & n5793 ) | ( n2342 & n6618 ) | ( n5793 & n6618 ) ;
  assign n22500 = n14660 ^ n4891 ^ 1'b0 ;
  assign n22501 = n22499 & n22500 ;
  assign n22502 = n22501 ^ n1063 ^ 1'b0 ;
  assign n22503 = n14136 ^ n7873 ^ 1'b0 ;
  assign n22504 = n4464 & n22503 ;
  assign n22505 = n13420 | n14058 ;
  assign n22506 = n22505 ^ n14164 ^ n13837 ;
  assign n22507 = n16197 ^ n1651 ^ 1'b0 ;
  assign n22508 = ( n9717 & n11455 ) | ( n9717 & n22507 ) | ( n11455 & n22507 ) ;
  assign n22509 = n12505 ^ n8616 ^ n8387 ;
  assign n22510 = n22509 ^ n18661 ^ n4619 ;
  assign n22511 = ( ~n917 & n11077 ) | ( ~n917 & n22510 ) | ( n11077 & n22510 ) ;
  assign n22512 = x143 & n2992 ;
  assign n22513 = n22512 ^ n16066 ^ 1'b0 ;
  assign n22520 = n7087 ^ n6673 ^ 1'b0 ;
  assign n22521 = ~n1870 & n6434 ;
  assign n22522 = n22521 ^ n5215 ^ 1'b0 ;
  assign n22523 = n22520 | n22522 ;
  assign n22514 = n8094 & ~n16201 ;
  assign n22515 = ~n8065 & n22514 ;
  assign n22516 = n18977 & ~n22515 ;
  assign n22517 = n9575 & n22516 ;
  assign n22518 = n22517 ^ n3722 ^ 1'b0 ;
  assign n22519 = n18626 & ~n22518 ;
  assign n22524 = n22523 ^ n22519 ^ 1'b0 ;
  assign n22525 = n15879 & ~n22524 ;
  assign n22526 = n5972 & n16711 ;
  assign n22527 = n22526 ^ n8858 ^ 1'b0 ;
  assign n22528 = n22527 ^ n17774 ^ 1'b0 ;
  assign n22529 = n9782 & n17082 ;
  assign n22530 = n22529 ^ n9872 ^ 1'b0 ;
  assign n22531 = n4439 & ~n22530 ;
  assign n22534 = ~n8300 & n8979 ;
  assign n22532 = ~n10199 & n11659 ;
  assign n22533 = ~n4931 & n22532 ;
  assign n22535 = n22534 ^ n22533 ^ n4069 ;
  assign n22536 = n11007 ^ n10230 ^ 1'b0 ;
  assign n22537 = n15478 | n22536 ;
  assign n22538 = n7311 ^ n4416 ^ 1'b0 ;
  assign n22539 = n7471 | n22538 ;
  assign n22542 = ~n7488 & n11410 ;
  assign n22540 = n12256 ^ n1928 ^ 1'b0 ;
  assign n22541 = n3796 | n22540 ;
  assign n22543 = n22542 ^ n22541 ^ n5263 ;
  assign n22550 = n21065 ^ n10703 ^ 1'b0 ;
  assign n22544 = n841 | n3866 ;
  assign n22545 = n7142 & n10764 ;
  assign n22546 = ~n2189 & n22545 ;
  assign n22547 = n1015 & n22546 ;
  assign n22548 = ~n22544 & n22547 ;
  assign n22549 = n10333 & n22548 ;
  assign n22551 = n22550 ^ n22549 ^ n22033 ;
  assign n22556 = n7335 & n10909 ;
  assign n22552 = n6769 ^ n6427 ^ 1'b0 ;
  assign n22553 = n11331 & n22552 ;
  assign n22554 = ~n5330 & n22553 ;
  assign n22555 = ~n9802 & n22554 ;
  assign n22557 = n22556 ^ n22555 ^ 1'b0 ;
  assign n22558 = ~n12335 & n19444 ;
  assign n22559 = n16083 | n22558 ;
  assign n22560 = n22557 | n22559 ;
  assign n22561 = n2878 & ~n12700 ;
  assign n22562 = n22561 ^ n17940 ^ 1'b0 ;
  assign n22563 = n16568 ^ n537 ^ 1'b0 ;
  assign n22564 = n5728 ^ x161 ^ 1'b0 ;
  assign n22565 = ( n19510 & n22098 ) | ( n19510 & ~n22564 ) | ( n22098 & ~n22564 ) ;
  assign n22566 = n4945 & ~n12998 ;
  assign n22567 = ( n7066 & n15112 ) | ( n7066 & n16542 ) | ( n15112 & n16542 ) ;
  assign n22568 = n12495 & ~n22567 ;
  assign n22570 = n7028 & n8508 ;
  assign n22571 = n22570 ^ n12227 ^ 1'b0 ;
  assign n22569 = n5003 | n21369 ;
  assign n22572 = n22571 ^ n22569 ^ 1'b0 ;
  assign n22573 = ( n11491 & n11965 ) | ( n11491 & ~n22572 ) | ( n11965 & ~n22572 ) ;
  assign n22574 = x227 | n7235 ;
  assign n22575 = n17931 ^ n13725 ^ 1'b0 ;
  assign n22576 = n14442 & n22575 ;
  assign n22577 = ~n22574 & n22576 ;
  assign n22578 = n5877 ^ n5710 ^ 1'b0 ;
  assign n22579 = n17396 & n22578 ;
  assign n22580 = n18748 ^ n3872 ^ 1'b0 ;
  assign n22581 = n18251 ^ n16846 ^ 1'b0 ;
  assign n22582 = n1239 & n22581 ;
  assign n22583 = n17264 ^ n12760 ^ n10018 ;
  assign n22584 = n12587 | n22583 ;
  assign n22585 = ( n8406 & ~n8624 ) | ( n8406 & n12624 ) | ( ~n8624 & n12624 ) ;
  assign n22586 = n15601 ^ n14398 ^ n2885 ;
  assign n22587 = n22586 ^ n7260 ^ 1'b0 ;
  assign n22588 = n5181 & n5752 ;
  assign n22589 = n4126 & n22588 ;
  assign n22590 = n10016 & ~n16529 ;
  assign n22591 = n11441 & ~n22590 ;
  assign n22592 = n4242 & ~n7465 ;
  assign n22593 = n13561 & n22592 ;
  assign n22594 = n6310 & ~n22593 ;
  assign n22595 = ~n9600 & n22594 ;
  assign n22596 = n22595 ^ n8991 ^ 1'b0 ;
  assign n22597 = n20382 ^ n540 ^ 1'b0 ;
  assign n22598 = n2889 & ~n22597 ;
  assign n22599 = n22598 ^ n15909 ^ 1'b0 ;
  assign n22600 = ( n14259 & n18197 ) | ( n14259 & ~n22599 ) | ( n18197 & ~n22599 ) ;
  assign n22601 = n11736 ^ n11381 ^ 1'b0 ;
  assign n22602 = n15418 & n20406 ;
  assign n22605 = n7399 & n12445 ;
  assign n22606 = n22605 ^ n7672 ^ 1'b0 ;
  assign n22604 = n3900 & n11412 ;
  assign n22607 = n22606 ^ n22604 ^ 1'b0 ;
  assign n22603 = ~n17825 & n21651 ;
  assign n22608 = n22607 ^ n22603 ^ 1'b0 ;
  assign n22609 = n4422 | n12700 ;
  assign n22614 = n7152 & n15078 ;
  assign n22615 = n22614 ^ n4280 ^ 1'b0 ;
  assign n22616 = n22615 ^ n1564 ^ 1'b0 ;
  assign n22617 = n1567 & ~n22616 ;
  assign n22618 = n412 & n3277 ;
  assign n22619 = n22618 ^ n10696 ^ 1'b0 ;
  assign n22620 = n22619 ^ n7649 ^ 1'b0 ;
  assign n22621 = ~n5261 & n22620 ;
  assign n22622 = ( n866 & n12476 ) | ( n866 & n22621 ) | ( n12476 & n22621 ) ;
  assign n22623 = n22622 ^ n4355 ^ 1'b0 ;
  assign n22624 = n22617 | n22623 ;
  assign n22610 = n12437 ^ n7404 ^ 1'b0 ;
  assign n22611 = ( n8043 & ~n16502 ) | ( n8043 & n22610 ) | ( ~n16502 & n22610 ) ;
  assign n22612 = n22611 ^ n19533 ^ 1'b0 ;
  assign n22613 = n3589 & ~n22612 ;
  assign n22625 = n22624 ^ n22613 ^ 1'b0 ;
  assign n22626 = n19218 | n22625 ;
  assign n22627 = n3955 & n9061 ;
  assign n22628 = n3188 & ~n22627 ;
  assign n22629 = n22628 ^ n7127 ^ 1'b0 ;
  assign n22630 = x73 & ~n22629 ;
  assign n22631 = n22630 ^ n9906 ^ 1'b0 ;
  assign n22632 = n17412 & ~n22631 ;
  assign n22633 = ( x27 & n815 ) | ( x27 & ~n12081 ) | ( n815 & ~n12081 ) ;
  assign n22634 = n22633 ^ n20055 ^ 1'b0 ;
  assign n22635 = n13921 ^ n3049 ^ 1'b0 ;
  assign n22636 = n7215 | n22635 ;
  assign n22637 = n6858 ^ n6453 ^ 1'b0 ;
  assign n22638 = n9682 | n18365 ;
  assign n22639 = n3541 ^ n3017 ^ n1385 ;
  assign n22640 = n22639 ^ n4190 ^ 1'b0 ;
  assign n22641 = n6627 & n12168 ;
  assign n22642 = ~n18223 & n22641 ;
  assign n22643 = n7223 & n11531 ;
  assign n22644 = n22643 ^ n7553 ^ 1'b0 ;
  assign n22645 = ~n9687 & n22644 ;
  assign n22646 = n22645 ^ n8533 ^ 1'b0 ;
  assign n22647 = n18939 ^ n5131 ^ 1'b0 ;
  assign n22648 = n1659 & ~n22647 ;
  assign n22649 = ( ~n12059 & n14038 ) | ( ~n12059 & n19089 ) | ( n14038 & n19089 ) ;
  assign n22650 = n22649 ^ n15756 ^ 1'b0 ;
  assign n22651 = n3545 ^ n1890 ^ 1'b0 ;
  assign n22652 = n22651 ^ n5912 ^ 1'b0 ;
  assign n22653 = x53 | n7658 ;
  assign n22654 = x224 & ~n1853 ;
  assign n22655 = ~n3344 & n22654 ;
  assign n22656 = n22655 ^ n16907 ^ n16493 ;
  assign n22657 = n22653 & ~n22656 ;
  assign n22658 = n22558 & n22657 ;
  assign n22659 = n20115 ^ n16385 ^ 1'b0 ;
  assign n22660 = n16109 & n16573 ;
  assign n22661 = n4446 & ~n13100 ;
  assign n22662 = n6708 & ~n16917 ;
  assign n22663 = n22662 ^ n6068 ^ 1'b0 ;
  assign n22664 = n3477 & ~n15703 ;
  assign n22665 = n15210 & n22664 ;
  assign n22666 = n7236 & ~n11373 ;
  assign n22667 = ~n3688 & n22666 ;
  assign n22668 = n9874 & n22667 ;
  assign n22669 = n16042 ^ n13356 ^ n3847 ;
  assign n22670 = n3738 & n18525 ;
  assign n22671 = n22670 ^ n13682 ^ 1'b0 ;
  assign n22672 = ( n6822 & ~n7788 ) | ( n6822 & n9002 ) | ( ~n7788 & n9002 ) ;
  assign n22673 = n8631 ^ n7430 ^ 1'b0 ;
  assign n22674 = n18768 & ~n22673 ;
  assign n22675 = n6463 | n8215 ;
  assign n22676 = n19780 & ~n22675 ;
  assign n22678 = ~n4322 & n13035 ;
  assign n22679 = n18134 ^ n4302 ^ 1'b0 ;
  assign n22680 = n22679 ^ n9872 ^ n5195 ;
  assign n22681 = ( n19178 & n22678 ) | ( n19178 & n22680 ) | ( n22678 & n22680 ) ;
  assign n22677 = ~n10436 & n17946 ;
  assign n22682 = n22681 ^ n22677 ^ 1'b0 ;
  assign n22683 = n22682 ^ n11409 ^ 1'b0 ;
  assign n22684 = n18394 | n22683 ;
  assign n22685 = n22676 & ~n22684 ;
  assign n22690 = n3379 | n5385 ;
  assign n22691 = n22690 ^ n305 ^ 1'b0 ;
  assign n22686 = ~n1688 & n6623 ;
  assign n22687 = n22686 ^ n6355 ^ 1'b0 ;
  assign n22688 = n4759 | n22687 ;
  assign n22689 = n22688 ^ n6271 ^ 1'b0 ;
  assign n22692 = n22691 ^ n22689 ^ 1'b0 ;
  assign n22693 = ( ~n11469 & n16005 ) | ( ~n11469 & n22692 ) | ( n16005 & n22692 ) ;
  assign n22694 = n6629 | n15746 ;
  assign n22695 = n22693 | n22694 ;
  assign n22696 = n22695 ^ n1778 ^ 1'b0 ;
  assign n22697 = n11028 & ~n22696 ;
  assign n22698 = ( n756 & n1374 ) | ( n756 & ~n22697 ) | ( n1374 & ~n22697 ) ;
  assign n22699 = n7262 ^ n6829 ^ 1'b0 ;
  assign n22700 = n12155 & n22699 ;
  assign n22701 = n5011 ^ n1885 ^ 1'b0 ;
  assign n22702 = n22701 ^ n10626 ^ 1'b0 ;
  assign n22703 = n1637 & n6660 ;
  assign n22704 = n11200 ^ n2885 ^ 1'b0 ;
  assign n22705 = n22703 | n22704 ;
  assign n22706 = n8278 & n10780 ;
  assign n22707 = n12954 & ~n14180 ;
  assign n22708 = n22706 & n22707 ;
  assign n22715 = ( ~n1361 & n2026 ) | ( ~n1361 & n17526 ) | ( n2026 & n17526 ) ;
  assign n22711 = n3381 & n8036 ;
  assign n22712 = n8650 & n22711 ;
  assign n22713 = n22712 ^ n3986 ^ n1733 ;
  assign n22714 = n10565 & n22713 ;
  assign n22716 = n22715 ^ n22714 ^ 1'b0 ;
  assign n22709 = n22653 ^ n3974 ^ 1'b0 ;
  assign n22710 = n4205 | n22709 ;
  assign n22717 = n22716 ^ n22710 ^ 1'b0 ;
  assign n22718 = n14391 ^ n13604 ^ 1'b0 ;
  assign n22719 = n13757 & n22718 ;
  assign n22720 = n21661 ^ x74 ^ 1'b0 ;
  assign n22721 = ( n19359 & n19700 ) | ( n19359 & ~n22720 ) | ( n19700 & ~n22720 ) ;
  assign n22723 = n885 | n1640 ;
  assign n22724 = n22723 ^ n18825 ^ 1'b0 ;
  assign n22725 = n15436 & n22724 ;
  assign n22722 = ~n5577 & n10468 ;
  assign n22726 = n22725 ^ n22722 ^ 1'b0 ;
  assign n22727 = ( n20865 & n21875 ) | ( n20865 & ~n22726 ) | ( n21875 & ~n22726 ) ;
  assign n22728 = ( n1519 & ~n1874 ) | ( n1519 & n7553 ) | ( ~n1874 & n7553 ) ;
  assign n22729 = n22728 ^ x151 ^ 1'b0 ;
  assign n22730 = n19379 | n22729 ;
  assign n22731 = n7952 | n10129 ;
  assign n22732 = n22731 ^ n18325 ^ 1'b0 ;
  assign n22733 = n1814 & n8531 ;
  assign n22734 = n1966 ^ n472 ^ x170 ;
  assign n22735 = n11875 | n22734 ;
  assign n22736 = n22733 | n22735 ;
  assign n22737 = n5269 ^ n2908 ^ n1174 ;
  assign n22738 = n10961 & ~n22737 ;
  assign n22739 = ~n22736 & n22738 ;
  assign n22740 = n7899 | n9521 ;
  assign n22741 = n22739 & ~n22740 ;
  assign n22742 = ~n9726 & n22741 ;
  assign n22743 = n14270 & n18502 ;
  assign n22744 = n22743 ^ n15401 ^ n6748 ;
  assign n22746 = n3768 & ~n16495 ;
  assign n22747 = ~n10998 & n22746 ;
  assign n22748 = n22747 ^ n12514 ^ 1'b0 ;
  assign n22745 = ~n2826 & n6106 ;
  assign n22749 = n22748 ^ n22745 ^ 1'b0 ;
  assign n22750 = n5839 | n19848 ;
  assign n22751 = n19157 & ~n22750 ;
  assign n22752 = n3967 | n7765 ;
  assign n22753 = n13438 ^ n7353 ^ 1'b0 ;
  assign n22758 = n1327 | n19252 ;
  assign n22759 = n22758 ^ n8439 ^ 1'b0 ;
  assign n22757 = ~n9775 & n16558 ;
  assign n22754 = n8158 & n8454 ;
  assign n22755 = n22754 ^ n8081 ^ 1'b0 ;
  assign n22756 = n1590 & n22755 ;
  assign n22760 = n22759 ^ n22757 ^ n22756 ;
  assign n22761 = n13513 ^ n3471 ^ 1'b0 ;
  assign n22762 = n9919 ^ n5713 ^ 1'b0 ;
  assign n22763 = n6931 | n14692 ;
  assign n22770 = ( ~n1634 & n7250 ) | ( ~n1634 & n11848 ) | ( n7250 & n11848 ) ;
  assign n22764 = n13121 ^ n2362 ^ 1'b0 ;
  assign n22765 = n21560 | n22764 ;
  assign n22766 = n22765 ^ n2275 ^ 1'b0 ;
  assign n22767 = n15684 ^ x112 ^ 1'b0 ;
  assign n22768 = ~n22766 & n22767 ;
  assign n22769 = n22768 ^ n6223 ^ 1'b0 ;
  assign n22771 = n22770 ^ n22769 ^ n1476 ;
  assign n22781 = n12718 ^ n11430 ^ 1'b0 ;
  assign n22782 = n7102 & ~n22781 ;
  assign n22783 = n22782 ^ n620 ^ 1'b0 ;
  assign n22780 = n816 | n5355 ;
  assign n22784 = n22783 ^ n22780 ^ 1'b0 ;
  assign n22777 = n5515 | n6667 ;
  assign n22778 = ( n10907 & n20835 ) | ( n10907 & ~n22777 ) | ( n20835 & ~n22777 ) ;
  assign n22772 = n1939 & ~n7101 ;
  assign n22773 = n22772 ^ n3723 ^ 1'b0 ;
  assign n22774 = n13359 & ~n22773 ;
  assign n22775 = n22774 ^ n16051 ^ 1'b0 ;
  assign n22776 = ~n1399 & n22775 ;
  assign n22779 = n22778 ^ n22776 ^ 1'b0 ;
  assign n22785 = n22784 ^ n22779 ^ n16556 ;
  assign n22786 = n17865 & n22785 ;
  assign n22787 = n22786 ^ n8072 ^ 1'b0 ;
  assign n22788 = ( n1413 & n6474 ) | ( n1413 & n7921 ) | ( n6474 & n7921 ) ;
  assign n22789 = n22788 ^ x35 ^ 1'b0 ;
  assign n22790 = n1831 | n22789 ;
  assign n22791 = n22790 ^ n20301 ^ 1'b0 ;
  assign n22792 = ~n8919 & n12553 ;
  assign n22793 = n17301 | n17631 ;
  assign n22794 = n6915 ^ n1653 ^ 1'b0 ;
  assign n22797 = ( ~n3990 & n8340 ) | ( ~n3990 & n22183 ) | ( n8340 & n22183 ) ;
  assign n22795 = n8732 | n17217 ;
  assign n22796 = n13219 & n22795 ;
  assign n22798 = n22797 ^ n22796 ^ n7324 ;
  assign n22799 = n22798 ^ n16885 ^ n4361 ;
  assign n22800 = n5131 & n22799 ;
  assign n22801 = ~n22794 & n22800 ;
  assign n22802 = ( ~n1938 & n7358 ) | ( ~n1938 & n10950 ) | ( n7358 & n10950 ) ;
  assign n22803 = ( n9659 & ~n16206 ) | ( n9659 & n22802 ) | ( ~n16206 & n22802 ) ;
  assign n22804 = n22803 ^ n5391 ^ 1'b0 ;
  assign n22805 = n10560 ^ n6713 ^ n5376 ;
  assign n22806 = n22805 ^ n15672 ^ n8345 ;
  assign n22807 = n8143 ^ n2624 ^ 1'b0 ;
  assign n22808 = n8919 ^ n3158 ^ 1'b0 ;
  assign n22810 = n4122 & n8847 ;
  assign n22809 = n17039 & n17185 ;
  assign n22811 = n22810 ^ n22809 ^ 1'b0 ;
  assign n22812 = n13067 ^ n7236 ^ 1'b0 ;
  assign n22813 = n22811 & n22812 ;
  assign n22814 = n15973 ^ n6518 ^ n4715 ;
  assign n22815 = n14157 ^ n6219 ^ 1'b0 ;
  assign n22816 = x78 & n22815 ;
  assign n22817 = n9156 ^ n3907 ^ 1'b0 ;
  assign n22818 = n22816 & n22817 ;
  assign n22819 = n256 & n22818 ;
  assign n22822 = n831 & n8507 ;
  assign n22823 = n8365 | n12331 ;
  assign n22824 = n22822 & ~n22823 ;
  assign n22820 = n9048 | n13721 ;
  assign n22821 = n22820 ^ n17142 ^ n10660 ;
  assign n22825 = n22824 ^ n22821 ^ 1'b0 ;
  assign n22826 = ~n12074 & n22825 ;
  assign n22827 = ( n872 & ~n1229 ) | ( n872 & n10272 ) | ( ~n1229 & n10272 ) ;
  assign n22828 = n22827 ^ n6850 ^ n1154 ;
  assign n22832 = n3254 | n4067 ;
  assign n22830 = n7774 ^ n6053 ^ n2167 ;
  assign n22831 = ( n1605 & ~n3599 ) | ( n1605 & n22830 ) | ( ~n3599 & n22830 ) ;
  assign n22829 = n13275 ^ n10584 ^ n4264 ;
  assign n22833 = n22832 ^ n22831 ^ n22829 ;
  assign n22834 = n22828 & ~n22833 ;
  assign n22835 = n16927 ^ n1228 ^ 1'b0 ;
  assign n22836 = ( n5803 & n5823 ) | ( n5803 & n22835 ) | ( n5823 & n22835 ) ;
  assign n22837 = n22836 ^ n17984 ^ n10755 ;
  assign n22838 = n326 & n10164 ;
  assign n22842 = ~n5233 & n8047 ;
  assign n22839 = n2513 ^ n1609 ^ 1'b0 ;
  assign n22840 = n18602 ^ n6560 ^ 1'b0 ;
  assign n22841 = n22839 & ~n22840 ;
  assign n22843 = n22842 ^ n22841 ^ 1'b0 ;
  assign n22844 = n14694 ^ x49 ^ 1'b0 ;
  assign n22845 = n1214 | n22844 ;
  assign n22846 = n10152 ^ n9396 ^ n5089 ;
  assign n22847 = n22845 | n22846 ;
  assign n22848 = ( n2396 & ~n7569 ) | ( n2396 & n22847 ) | ( ~n7569 & n22847 ) ;
  assign n22849 = n10487 ^ n7096 ^ n2086 ;
  assign n22850 = n22849 ^ n1673 ^ 1'b0 ;
  assign n22851 = n22850 ^ n22447 ^ x25 ;
  assign n22854 = ( n3191 & ~n5153 ) | ( n3191 & n6287 ) | ( ~n5153 & n6287 ) ;
  assign n22855 = n1389 & n13877 ;
  assign n22856 = ~n22854 & n22855 ;
  assign n22852 = n3972 ^ n2048 ^ 1'b0 ;
  assign n22853 = n22852 ^ x158 ^ 1'b0 ;
  assign n22857 = n22856 ^ n22853 ^ n22190 ;
  assign n22858 = n12457 & n22857 ;
  assign n22859 = n22858 ^ n11019 ^ 1'b0 ;
  assign n22860 = ~n8538 & n19947 ;
  assign n22861 = n20959 ^ n6358 ^ 1'b0 ;
  assign n22862 = n22861 ^ n18602 ^ n12247 ;
  assign n22863 = ( ~n5408 & n10757 ) | ( ~n5408 & n22862 ) | ( n10757 & n22862 ) ;
  assign n22864 = ~n1853 & n19592 ;
  assign n22865 = n11795 & n22864 ;
  assign n22866 = n2144 & ~n4886 ;
  assign n22867 = n5166 & n8531 ;
  assign n22868 = n3996 & n22867 ;
  assign n22869 = n22868 ^ n13397 ^ n4498 ;
  assign n22875 = n5782 & ~n9300 ;
  assign n22876 = ~n2430 & n22875 ;
  assign n22870 = n15760 ^ n15568 ^ 1'b0 ;
  assign n22871 = n12818 ^ n9781 ^ 1'b0 ;
  assign n22872 = n22870 | n22871 ;
  assign n22873 = ~n3510 & n22872 ;
  assign n22874 = n13172 & ~n22873 ;
  assign n22877 = n22876 ^ n22874 ^ 1'b0 ;
  assign n22880 = n15114 ^ n9757 ^ 1'b0 ;
  assign n22878 = n1379 & ~n12197 ;
  assign n22879 = n379 & n22878 ;
  assign n22881 = n22880 ^ n22879 ^ n459 ;
  assign n22882 = n2548 & n9539 ;
  assign n22883 = n12772 & n22882 ;
  assign n22884 = ( ~x197 & n407 ) | ( ~x197 & n22883 ) | ( n407 & n22883 ) ;
  assign n22885 = ~n9583 & n10753 ;
  assign n22886 = n22885 ^ n18960 ^ n9121 ;
  assign n22887 = n13155 ^ n3674 ^ 1'b0 ;
  assign n22888 = n22886 | n22887 ;
  assign n22889 = n1118 | n22888 ;
  assign n22890 = n22889 ^ n21380 ^ 1'b0 ;
  assign n22891 = n1691 & ~n5079 ;
  assign n22892 = n22891 ^ n9176 ^ 1'b0 ;
  assign n22893 = n11306 | n22892 ;
  assign n22894 = n12556 | n16581 ;
  assign n22895 = n1309 | n3389 ;
  assign n22896 = n3712 | n22895 ;
  assign n22897 = n15261 & n22896 ;
  assign n22898 = n12418 ^ n11601 ^ n10526 ;
  assign n22899 = ~n17106 & n22898 ;
  assign n22900 = ~n22897 & n22899 ;
  assign n22901 = n21185 ^ n9187 ^ n8876 ;
  assign n22902 = n485 & ~n22901 ;
  assign n22903 = n10186 ^ n2974 ^ 1'b0 ;
  assign n22904 = n2125 & n7488 ;
  assign n22905 = ~n15576 & n22904 ;
  assign n22906 = n22905 ^ n13346 ^ 1'b0 ;
  assign n22907 = ( n983 & n22903 ) | ( n983 & n22906 ) | ( n22903 & n22906 ) ;
  assign n22908 = n22907 ^ n16121 ^ n294 ;
  assign n22909 = n22908 ^ n20659 ^ 1'b0 ;
  assign n22910 = n1150 | n21543 ;
  assign n22911 = n1129 | n22910 ;
  assign n22912 = ( n953 & n11973 ) | ( n953 & n18842 ) | ( n11973 & n18842 ) ;
  assign n22913 = n10977 ^ n993 ^ 1'b0 ;
  assign n22914 = n11562 | n22913 ;
  assign n22916 = n12263 ^ n10062 ^ 1'b0 ;
  assign n22917 = n13729 & n22916 ;
  assign n22915 = ~n11965 & n19649 ;
  assign n22918 = n22917 ^ n22915 ^ 1'b0 ;
  assign n22919 = n3743 & ~n5270 ;
  assign n22920 = n9436 ^ n4499 ^ 1'b0 ;
  assign n22921 = n22919 & ~n22920 ;
  assign n22922 = ~n9701 & n17412 ;
  assign n22923 = ~n18082 & n22922 ;
  assign n22924 = ( n10032 & n12723 ) | ( n10032 & n22923 ) | ( n12723 & n22923 ) ;
  assign n22925 = ( n5191 & ~n8465 ) | ( n5191 & n22924 ) | ( ~n8465 & n22924 ) ;
  assign n22926 = n22925 ^ n3279 ^ 1'b0 ;
  assign n22929 = n11682 ^ n9631 ^ n4011 ;
  assign n22930 = n22929 ^ n7425 ^ n2950 ;
  assign n22927 = ( n957 & n8122 ) | ( n957 & n16094 ) | ( n8122 & n16094 ) ;
  assign n22928 = n1795 & ~n22927 ;
  assign n22931 = n22930 ^ n22928 ^ 1'b0 ;
  assign n22932 = n8682 ^ n4735 ^ 1'b0 ;
  assign n22933 = n1168 & n22932 ;
  assign n22934 = ( ~n4072 & n10873 ) | ( ~n4072 & n22933 ) | ( n10873 & n22933 ) ;
  assign n22935 = n15884 ^ n12351 ^ 1'b0 ;
  assign n22936 = n12341 ^ n8559 ^ 1'b0 ;
  assign n22937 = n22935 | n22936 ;
  assign n22938 = n11135 & ~n15054 ;
  assign n22939 = n7245 & n22938 ;
  assign n22940 = ~n1576 & n3891 ;
  assign n22941 = n11709 & ~n22940 ;
  assign n22942 = n5003 | n7034 ;
  assign n22943 = n14364 | n22942 ;
  assign n22944 = ~n17093 & n22943 ;
  assign n22945 = n1005 & n22944 ;
  assign n22946 = n1328 & n6693 ;
  assign n22947 = n15085 | n22946 ;
  assign n22948 = ( n1281 & n1446 ) | ( n1281 & ~n14023 ) | ( n1446 & ~n14023 ) ;
  assign n22949 = n22948 ^ n9074 ^ 1'b0 ;
  assign n22950 = n8821 ^ n3794 ^ n2245 ;
  assign n22951 = ( n1306 & n2730 ) | ( n1306 & n22950 ) | ( n2730 & n22950 ) ;
  assign n22952 = n9054 & ~n10255 ;
  assign n22953 = n22952 ^ n5328 ^ n3029 ;
  assign n22959 = ~n7180 & n7386 ;
  assign n22958 = ~n4255 & n6420 ;
  assign n22954 = ~n6296 & n17578 ;
  assign n22955 = n7646 & n22954 ;
  assign n22956 = n16485 | n22955 ;
  assign n22957 = n22956 ^ n16970 ^ 1'b0 ;
  assign n22960 = n22959 ^ n22958 ^ n22957 ;
  assign n22962 = n8351 & n20254 ;
  assign n22961 = ( n13089 & n17372 ) | ( n13089 & n20995 ) | ( n17372 & n20995 ) ;
  assign n22963 = n22962 ^ n22961 ^ 1'b0 ;
  assign n22964 = n3299 & ~n6919 ;
  assign n22965 = n3992 & n12811 ;
  assign n22966 = n10669 & n22965 ;
  assign n22967 = n8698 ^ n1164 ^ 1'b0 ;
  assign n22968 = ( x98 & n8420 ) | ( x98 & ~n22967 ) | ( n8420 & ~n22967 ) ;
  assign n22969 = n16640 ^ n12526 ^ 1'b0 ;
  assign n22970 = n11087 ^ n10682 ^ 1'b0 ;
  assign n22971 = n20334 ^ n13163 ^ 1'b0 ;
  assign n22972 = n6607 ^ n4619 ^ 1'b0 ;
  assign n22973 = n6450 & ~n14440 ;
  assign n22974 = ~n22940 & n22973 ;
  assign n22975 = ( n1787 & n3746 ) | ( n1787 & ~n17464 ) | ( n3746 & ~n17464 ) ;
  assign n22976 = n22975 ^ n16397 ^ 1'b0 ;
  assign n22977 = n7840 & n22976 ;
  assign n22978 = n6132 ^ n428 ^ 1'b0 ;
  assign n22979 = ~n6474 & n22978 ;
  assign n22980 = x67 & n9250 ;
  assign n22981 = n16154 ^ n1768 ^ 1'b0 ;
  assign n22982 = ~n22980 & n22981 ;
  assign n22983 = ( n6526 & n11886 ) | ( n6526 & n22982 ) | ( n11886 & n22982 ) ;
  assign n22984 = ( n13587 & n13685 ) | ( n13587 & n17159 ) | ( n13685 & n17159 ) ;
  assign n22985 = n998 | n16823 ;
  assign n22986 = n22985 ^ n1869 ^ 1'b0 ;
  assign n22987 = n2452 | n13108 ;
  assign n22988 = n22987 ^ n3213 ^ 1'b0 ;
  assign n22989 = n21299 ^ n13454 ^ n9431 ;
  assign n22990 = n3791 ^ n717 ^ 1'b0 ;
  assign n22991 = ~n4236 & n22990 ;
  assign n22992 = n22991 ^ n21213 ^ 1'b0 ;
  assign n22993 = n22748 | n22992 ;
  assign n22994 = n20280 & ~n22993 ;
  assign n22995 = n4291 ^ n682 ^ 1'b0 ;
  assign n22996 = ~n22994 & n22995 ;
  assign n22997 = n22472 ^ n20660 ^ 1'b0 ;
  assign n22998 = ~n4153 & n22997 ;
  assign n23000 = n12460 & n13550 ;
  assign n22999 = n13035 ^ n2756 ^ n2600 ;
  assign n23001 = n23000 ^ n22999 ^ 1'b0 ;
  assign n23002 = n4243 & ~n14378 ;
  assign n23003 = n20723 ^ n16860 ^ 1'b0 ;
  assign n23004 = n1800 | n23003 ;
  assign n23005 = n23004 ^ n5525 ^ 1'b0 ;
  assign n23006 = ~n19721 & n23005 ;
  assign n23007 = ~n23002 & n23006 ;
  assign n23008 = n11584 ^ n1848 ^ 1'b0 ;
  assign n23009 = n15071 & n23008 ;
  assign n23010 = n23009 ^ n16837 ^ 1'b0 ;
  assign n23011 = ~n7282 & n7478 ;
  assign n23012 = n23011 ^ n1963 ^ 1'b0 ;
  assign n23013 = n945 & n7375 ;
  assign n23014 = n17731 & ~n23013 ;
  assign n23015 = n23012 | n23014 ;
  assign n23016 = n1649 & ~n7577 ;
  assign n23017 = n2169 | n9783 ;
  assign n23018 = n23016 | n23017 ;
  assign n23019 = ( n12959 & n13450 ) | ( n12959 & ~n16195 ) | ( n13450 & ~n16195 ) ;
  assign n23020 = n23019 ^ n18125 ^ 1'b0 ;
  assign n23021 = n402 & ~n6292 ;
  assign n23022 = n6608 & ~n23021 ;
  assign n23023 = n23022 ^ n21570 ^ 1'b0 ;
  assign n23024 = n7125 ^ n2565 ^ 1'b0 ;
  assign n23025 = n23024 ^ n21003 ^ n14665 ;
  assign n23026 = n1275 & n4019 ;
  assign n23027 = n1835 | n9146 ;
  assign n23028 = n4192 & ~n23027 ;
  assign n23029 = n23028 ^ n10926 ^ 1'b0 ;
  assign n23030 = ~n19294 & n23029 ;
  assign n23031 = n23026 & n23030 ;
  assign n23032 = n12124 & n23031 ;
  assign n23033 = n1249 | n23032 ;
  assign n23034 = x121 & n11589 ;
  assign n23035 = n23034 ^ n6247 ^ 1'b0 ;
  assign n23036 = n2199 | n23035 ;
  assign n23037 = n4004 | n23036 ;
  assign n23038 = n23037 ^ n18702 ^ 1'b0 ;
  assign n23039 = n10629 & ~n23038 ;
  assign n23040 = n11951 & n23039 ;
  assign n23041 = ~n21834 & n23040 ;
  assign n23042 = n5475 & n19138 ;
  assign n23043 = ~n20899 & n23042 ;
  assign n23044 = n15461 & ~n23043 ;
  assign n23045 = n1850 & n23044 ;
  assign n23046 = ( n329 & n11211 ) | ( n329 & ~n15719 ) | ( n11211 & ~n15719 ) ;
  assign n23047 = n23046 ^ n21454 ^ n8548 ;
  assign n23048 = ~n1258 & n2720 ;
  assign n23049 = n8345 | n23048 ;
  assign n23050 = n13283 & n23049 ;
  assign n23051 = ~n8828 & n23050 ;
  assign n23052 = n14490 ^ n10861 ^ 1'b0 ;
  assign n23053 = n1523 & n5397 ;
  assign n23054 = n23053 ^ n14490 ^ 1'b0 ;
  assign n23055 = n9030 & ~n23054 ;
  assign n23056 = n805 & n23055 ;
  assign n23057 = n15906 & n23056 ;
  assign n23058 = n15436 & ~n16004 ;
  assign n23059 = n14281 & n23058 ;
  assign n23060 = ( n12189 & ~n23057 ) | ( n12189 & n23059 ) | ( ~n23057 & n23059 ) ;
  assign n23061 = n1481 & n14183 ;
  assign n23063 = n10111 ^ n387 ^ 1'b0 ;
  assign n23064 = n961 & n23063 ;
  assign n23062 = n2077 | n16497 ;
  assign n23065 = n23064 ^ n23062 ^ 1'b0 ;
  assign n23066 = n23065 ^ n15963 ^ n13331 ;
  assign n23068 = ( n8251 & n10339 ) | ( n8251 & n11238 ) | ( n10339 & n11238 ) ;
  assign n23067 = n11044 & ~n15246 ;
  assign n23069 = n23068 ^ n23067 ^ n15719 ;
  assign n23070 = ~n12666 & n23069 ;
  assign n23071 = n23070 ^ n6062 ^ 1'b0 ;
  assign n23072 = n1331 & ~n10450 ;
  assign n23073 = n4988 & n10877 ;
  assign n23074 = n18833 ^ n18240 ^ n17974 ;
  assign n23075 = n23073 & ~n23074 ;
  assign n23076 = n23072 & n23075 ;
  assign n23077 = n20772 ^ n3727 ^ 1'b0 ;
  assign n23078 = ( n8627 & n11590 ) | ( n8627 & n16356 ) | ( n11590 & n16356 ) ;
  assign n23079 = n13420 & n21235 ;
  assign n23080 = ~x149 & n23079 ;
  assign n23081 = n20248 ^ n7375 ^ 1'b0 ;
  assign n23082 = ~n15969 & n23081 ;
  assign n23083 = ~n15387 & n23082 ;
  assign n23084 = n23083 ^ n1476 ^ 1'b0 ;
  assign n23085 = ( ~n6232 & n10617 ) | ( ~n6232 & n21886 ) | ( n10617 & n21886 ) ;
  assign n23086 = n23085 ^ n9757 ^ n8996 ;
  assign n23087 = n23084 & n23086 ;
  assign n23088 = n23087 ^ n1971 ^ 1'b0 ;
  assign n23089 = n9731 ^ n1937 ^ n1918 ;
  assign n23090 = ~n3154 & n18158 ;
  assign n23091 = ~n5328 & n23090 ;
  assign n23092 = n23091 ^ n5967 ^ 1'b0 ;
  assign n23093 = ~n1523 & n23092 ;
  assign n23094 = n6485 & ~n23093 ;
  assign n23095 = ~n23089 & n23094 ;
  assign n23096 = ( n403 & n2200 ) | ( n403 & n2310 ) | ( n2200 & n2310 ) ;
  assign n23097 = n11168 ^ n7789 ^ 1'b0 ;
  assign n23098 = ( n10112 & n15760 ) | ( n10112 & n23097 ) | ( n15760 & n23097 ) ;
  assign n23099 = n16345 & ~n23098 ;
  assign n23100 = n16919 | n23099 ;
  assign n23101 = n18892 ^ n2348 ^ 1'b0 ;
  assign n23102 = n4520 & n20336 ;
  assign n23103 = n23102 ^ n3900 ^ 1'b0 ;
  assign n23104 = n23101 & n23103 ;
  assign n23106 = n7096 ^ n6218 ^ 1'b0 ;
  assign n23105 = n8634 ^ n7364 ^ 1'b0 ;
  assign n23107 = n23106 ^ n23105 ^ n1916 ;
  assign n23108 = n18575 & n23107 ;
  assign n23109 = n7080 & n23108 ;
  assign n23110 = n23109 ^ n13493 ^ n13215 ;
  assign n23111 = n2883 & ~n7420 ;
  assign n23112 = n23111 ^ n18684 ^ n3755 ;
  assign n23113 = n1763 & n14093 ;
  assign n23114 = n12700 ^ n10734 ^ 1'b0 ;
  assign n23115 = n6118 ^ n2900 ^ 1'b0 ;
  assign n23116 = ( n7500 & n21822 ) | ( n7500 & ~n23115 ) | ( n21822 & ~n23115 ) ;
  assign n23117 = n23116 ^ n7899 ^ n5913 ;
  assign n23118 = n3314 ^ x200 ^ 1'b0 ;
  assign n23119 = n2830 & n23118 ;
  assign n23120 = ~n23117 & n23119 ;
  assign n23123 = n7240 & ~n20305 ;
  assign n23121 = ~n6024 & n16699 ;
  assign n23122 = n23121 ^ n6979 ^ 1'b0 ;
  assign n23124 = n23123 ^ n23122 ^ 1'b0 ;
  assign n23125 = ~n573 & n4580 ;
  assign n23126 = ( n16569 & n23089 ) | ( n16569 & ~n23125 ) | ( n23089 & ~n23125 ) ;
  assign n23127 = n2106 & ~n5878 ;
  assign n23128 = ~n8934 & n23127 ;
  assign n23129 = n23128 ^ n10405 ^ n6352 ;
  assign n23130 = n18266 ^ n6186 ^ 1'b0 ;
  assign n23131 = n23130 ^ n3132 ^ 1'b0 ;
  assign n23132 = n23029 ^ n7284 ^ 1'b0 ;
  assign n23133 = n23132 ^ n19966 ^ n6062 ;
  assign n23134 = ~n6503 & n14938 ;
  assign n23135 = n5872 & ~n16965 ;
  assign n23136 = n10713 & n23135 ;
  assign n23137 = ~n2061 & n2323 ;
  assign n23138 = n13182 & ~n23137 ;
  assign n23139 = n2500 & ~n23138 ;
  assign n23140 = n943 ^ n690 ^ 1'b0 ;
  assign n23141 = ~n14449 & n23140 ;
  assign n23142 = n23141 ^ n11009 ^ 1'b0 ;
  assign n23143 = x76 & ~n21459 ;
  assign n23144 = n16599 ^ n7213 ^ n6124 ;
  assign n23145 = n23143 | n23144 ;
  assign n23146 = n18420 ^ n11062 ^ 1'b0 ;
  assign n23147 = n17542 ^ n10528 ^ 1'b0 ;
  assign n23148 = ~n11008 & n23147 ;
  assign n23149 = n18896 ^ n18493 ^ 1'b0 ;
  assign n23150 = n23149 ^ n22350 ^ n14628 ;
  assign n23151 = n22236 ^ n10355 ^ 1'b0 ;
  assign n23152 = n15398 ^ n10794 ^ n4074 ;
  assign n23153 = n23152 ^ n1976 ^ 1'b0 ;
  assign n23154 = n4448 ^ n1909 ^ n898 ;
  assign n23155 = ~n8800 & n23154 ;
  assign n23156 = n1999 & ~n6367 ;
  assign n23157 = n5967 & n23156 ;
  assign n23158 = n23157 ^ n19138 ^ n12024 ;
  assign n23159 = n8161 & n11300 ;
  assign n23160 = ~n5535 & n23159 ;
  assign n23161 = n23160 ^ n682 ^ 1'b0 ;
  assign n23162 = n16407 & ~n19309 ;
  assign n23168 = n4242 & ~n15950 ;
  assign n23163 = ~n14126 & n20131 ;
  assign n23164 = n2506 | n23163 ;
  assign n23165 = n11174 & ~n23164 ;
  assign n23166 = n11358 & ~n23165 ;
  assign n23167 = ~x47 & n23166 ;
  assign n23169 = n23168 ^ n23167 ^ 1'b0 ;
  assign n23170 = n15770 & n23169 ;
  assign n23171 = n4646 | n23170 ;
  assign n23173 = n12849 ^ n3639 ^ 1'b0 ;
  assign n23172 = ( n974 & ~n5662 ) | ( n974 & n7068 ) | ( ~n5662 & n7068 ) ;
  assign n23174 = n23173 ^ n23172 ^ x59 ;
  assign n23175 = n12455 & ~n23174 ;
  assign n23176 = ( n2665 & n3440 ) | ( n2665 & ~n8466 ) | ( n3440 & ~n8466 ) ;
  assign n23177 = x250 & n23176 ;
  assign n23178 = ~n13035 & n23177 ;
  assign n23179 = n7971 ^ n2266 ^ 1'b0 ;
  assign n23180 = n8132 & n23179 ;
  assign n23181 = n8328 ^ n6558 ^ 1'b0 ;
  assign n23182 = ~n256 & n23181 ;
  assign n23183 = ~n13756 & n23182 ;
  assign n23184 = n23183 ^ n2144 ^ 1'b0 ;
  assign n23185 = ( n11022 & n23180 ) | ( n11022 & ~n23184 ) | ( n23180 & ~n23184 ) ;
  assign n23186 = n23185 ^ n5195 ^ 1'b0 ;
  assign n23187 = n16817 ^ n7197 ^ 1'b0 ;
  assign n23188 = n17355 | n22554 ;
  assign n23189 = n20255 ^ x204 ^ 1'b0 ;
  assign n23190 = ~n1216 & n23189 ;
  assign n23191 = n3408 & ~n10010 ;
  assign n23192 = n23191 ^ n7290 ^ n6736 ;
  assign n23193 = x110 & n5351 ;
  assign n23194 = n23192 & n23193 ;
  assign n23195 = n1201 & ~n9231 ;
  assign n23196 = ~n2687 & n23195 ;
  assign n23197 = n5055 ^ n3984 ^ 1'b0 ;
  assign n23198 = n7957 ^ n1963 ^ 1'b0 ;
  assign n23199 = ( n23196 & ~n23197 ) | ( n23196 & n23198 ) | ( ~n23197 & n23198 ) ;
  assign n23200 = n23199 ^ n21714 ^ n16640 ;
  assign n23201 = n8430 ^ n1795 ^ 1'b0 ;
  assign n23202 = n23201 ^ n6435 ^ 1'b0 ;
  assign n23203 = x21 & ~n23202 ;
  assign n23204 = n16753 & n17682 ;
  assign n23205 = n23204 ^ n16866 ^ 1'b0 ;
  assign n23206 = ( n10793 & ~n17018 ) | ( n10793 & n20683 ) | ( ~n17018 & n20683 ) ;
  assign n23207 = n17338 | n23206 ;
  assign n23208 = ( n4767 & n19313 ) | ( n4767 & ~n19977 ) | ( n19313 & ~n19977 ) ;
  assign n23209 = n12214 & ~n22349 ;
  assign n23210 = n20005 ^ n4020 ^ 1'b0 ;
  assign n23212 = ( n1291 & ~n1347 ) | ( n1291 & n2352 ) | ( ~n1347 & n2352 ) ;
  assign n23211 = n3561 | n5524 ;
  assign n23213 = n23212 ^ n23211 ^ n2802 ;
  assign n23214 = ( n8426 & n10212 ) | ( n8426 & n18121 ) | ( n10212 & n18121 ) ;
  assign n23216 = ~n2616 & n6728 ;
  assign n23217 = n23216 ^ n2961 ^ 1'b0 ;
  assign n23215 = n968 & ~n13502 ;
  assign n23218 = n23217 ^ n23215 ^ 1'b0 ;
  assign n23220 = n15311 ^ n3957 ^ 1'b0 ;
  assign n23219 = ( n1598 & n2183 ) | ( n1598 & ~n4817 ) | ( n2183 & ~n4817 ) ;
  assign n23221 = n23220 ^ n23219 ^ 1'b0 ;
  assign n23223 = n20781 ^ n13701 ^ 1'b0 ;
  assign n23222 = n6816 | n14478 ;
  assign n23224 = n23223 ^ n23222 ^ n19270 ;
  assign n23225 = n23224 ^ n7736 ^ 1'b0 ;
  assign n23226 = x227 & n8862 ;
  assign n23227 = n23226 ^ n4896 ^ 1'b0 ;
  assign n23229 = n519 | n9281 ;
  assign n23230 = n18292 & ~n23229 ;
  assign n23231 = ~n1063 & n2775 ;
  assign n23232 = ~n2775 & n23231 ;
  assign n23233 = n23230 | n23232 ;
  assign n23234 = n23230 & ~n23233 ;
  assign n23228 = n8588 | n18186 ;
  assign n23235 = n23234 ^ n23228 ^ 1'b0 ;
  assign n23236 = n3240 & ~n9165 ;
  assign n23237 = n19869 ^ n9840 ^ n5544 ;
  assign n23238 = ( n8671 & n23236 ) | ( n8671 & ~n23237 ) | ( n23236 & ~n23237 ) ;
  assign n23239 = n12800 ^ n6870 ^ n2313 ;
  assign n23240 = n17544 | n23239 ;
  assign n23241 = ~n1285 & n23240 ;
  assign n23242 = n8327 ^ n2850 ^ n2071 ;
  assign n23243 = ~n5004 & n16599 ;
  assign n23244 = ~n805 & n23243 ;
  assign n23245 = ( n1664 & ~n4423 ) | ( n1664 & n7854 ) | ( ~n4423 & n7854 ) ;
  assign n23246 = ( n8964 & n23244 ) | ( n8964 & n23245 ) | ( n23244 & n23245 ) ;
  assign n23247 = ~n5009 & n23246 ;
  assign n23248 = ~n13346 & n23247 ;
  assign n23249 = n2248 | n19962 ;
  assign n23250 = n6213 & n23249 ;
  assign n23251 = ~n16609 & n23250 ;
  assign n23252 = n9993 | n18324 ;
  assign n23253 = n23252 ^ n15902 ^ 1'b0 ;
  assign n23254 = ~n1806 & n4458 ;
  assign n23255 = n7231 | n23254 ;
  assign n23256 = x73 & n3056 ;
  assign n23257 = n23256 ^ n6996 ^ 1'b0 ;
  assign n23258 = ~n8247 & n23257 ;
  assign n23259 = n23258 ^ n9656 ^ 1'b0 ;
  assign n23260 = n18589 ^ n16514 ^ 1'b0 ;
  assign n23261 = n17714 ^ n17194 ^ n14651 ;
  assign n23264 = n16525 ^ n9794 ^ n639 ;
  assign n23265 = n21085 ^ n12622 ^ 1'b0 ;
  assign n23266 = n23264 & n23265 ;
  assign n23262 = n6506 | n9090 ;
  assign n23263 = n11062 | n23262 ;
  assign n23267 = n23266 ^ n23263 ^ n6795 ;
  assign n23268 = n14217 ^ n5102 ^ n2998 ;
  assign n23269 = n771 & n23268 ;
  assign n23270 = n16423 ^ n15346 ^ 1'b0 ;
  assign n23271 = n2782 & n23270 ;
  assign n23272 = ~n12107 & n23271 ;
  assign n23274 = n16080 ^ n3652 ^ n1543 ;
  assign n23273 = n7818 & ~n10563 ;
  assign n23275 = n23274 ^ n23273 ^ 1'b0 ;
  assign n23276 = ( ~x76 & n7901 ) | ( ~x76 & n8830 ) | ( n7901 & n8830 ) ;
  assign n23277 = n23276 ^ n10941 ^ 1'b0 ;
  assign n23278 = n976 | n23277 ;
  assign n23279 = ( n1904 & n12375 ) | ( n1904 & ~n14850 ) | ( n12375 & ~n14850 ) ;
  assign n23280 = ( n15248 & ~n20768 ) | ( n15248 & n23279 ) | ( ~n20768 & n23279 ) ;
  assign n23281 = n23280 ^ n22258 ^ 1'b0 ;
  assign n23282 = n11072 ^ n5965 ^ 1'b0 ;
  assign n23283 = n5933 & ~n23282 ;
  assign n23284 = ~n1667 & n23283 ;
  assign n23285 = n23284 ^ n21100 ^ n4205 ;
  assign n23286 = n10288 ^ n6674 ^ 1'b0 ;
  assign n23287 = n21271 & n23286 ;
  assign n23288 = n5470 & ~n23287 ;
  assign n23289 = n10322 & ~n22490 ;
  assign n23290 = n3046 & n23289 ;
  assign n23291 = n4327 & n9141 ;
  assign n23292 = n23291 ^ n4282 ^ 1'b0 ;
  assign n23293 = n23292 ^ n4307 ^ 1'b0 ;
  assign n23294 = n6967 ^ n3917 ^ n1185 ;
  assign n23295 = n13698 & n23294 ;
  assign n23296 = n9632 & n13704 ;
  assign n23297 = n905 | n9919 ;
  assign n23298 = n2577 & ~n23297 ;
  assign n23299 = n20012 ^ n12180 ^ 1'b0 ;
  assign n23300 = n23298 | n23299 ;
  assign n23301 = n23300 ^ n14531 ^ n7616 ;
  assign n23302 = ( n12273 & ~n23296 ) | ( n12273 & n23301 ) | ( ~n23296 & n23301 ) ;
  assign n23304 = n15703 ^ n2257 ^ 1'b0 ;
  assign n23303 = n2942 & ~n9377 ;
  assign n23305 = n23304 ^ n23303 ^ 1'b0 ;
  assign n23306 = n14125 & ~n18100 ;
  assign n23307 = n12439 & n23306 ;
  assign n23308 = ~n10498 & n12288 ;
  assign n23309 = n14040 & n15402 ;
  assign n23310 = n14779 ^ n13630 ^ n807 ;
  assign n23311 = ~n5839 & n23310 ;
  assign n23312 = n17172 & n23311 ;
  assign n23313 = n20751 ^ n15382 ^ n6250 ;
  assign n23314 = n4695 & ~n7425 ;
  assign n23315 = ~n4695 & n23314 ;
  assign n23316 = n7127 & ~n23315 ;
  assign n23317 = ~n7127 & n23316 ;
  assign n23318 = n4592 | n23317 ;
  assign n23319 = n4592 & ~n23318 ;
  assign n23320 = n12290 | n23319 ;
  assign n23321 = n23319 & ~n23320 ;
  assign n23322 = n23321 ^ n5671 ^ 1'b0 ;
  assign n23323 = n20969 & ~n23322 ;
  assign n23324 = n18604 ^ n16108 ^ 1'b0 ;
  assign n23325 = n23324 ^ n21194 ^ n9266 ;
  assign n23326 = ~n12118 & n21414 ;
  assign n23327 = n23326 ^ x126 ^ 1'b0 ;
  assign n23328 = n2879 | n6800 ;
  assign n23329 = n5632 & ~n23328 ;
  assign n23330 = n1500 & n9792 ;
  assign n23331 = n23330 ^ n2431 ^ 1'b0 ;
  assign n23332 = ( n3357 & ~n8180 ) | ( n3357 & n17961 ) | ( ~n8180 & n17961 ) ;
  assign n23333 = n12575 ^ n8626 ^ n1037 ;
  assign n23334 = n23333 ^ n23265 ^ 1'b0 ;
  assign n23335 = ~n12282 & n18271 ;
  assign n23336 = ~n12644 & n23335 ;
  assign n23337 = n23336 ^ n13461 ^ 1'b0 ;
  assign n23338 = ( n1890 & n4699 ) | ( n1890 & n9113 ) | ( n4699 & n9113 ) ;
  assign n23339 = n23338 ^ n13499 ^ 1'b0 ;
  assign n23340 = n9647 & ~n23339 ;
  assign n23341 = n8958 & n23340 ;
  assign n23342 = n18462 ^ n15300 ^ n13821 ;
  assign n23343 = ~n925 & n5365 ;
  assign n23344 = ( n1025 & ~n18256 ) | ( n1025 & n23343 ) | ( ~n18256 & n23343 ) ;
  assign n23345 = ( n15877 & n23342 ) | ( n15877 & ~n23344 ) | ( n23342 & ~n23344 ) ;
  assign n23350 = n479 & n7157 ;
  assign n23351 = n5524 & n23350 ;
  assign n23346 = n7439 & ~n11357 ;
  assign n23347 = n23346 ^ n738 ^ 1'b0 ;
  assign n23348 = n21894 | n23347 ;
  assign n23349 = n2867 | n23348 ;
  assign n23352 = n23351 ^ n23349 ^ n5704 ;
  assign n23353 = n2157 ^ n1975 ^ 1'b0 ;
  assign n23354 = n23353 ^ n14271 ^ n2695 ;
  assign n23355 = n18597 ^ n7971 ^ 1'b0 ;
  assign n23356 = n10125 & n23355 ;
  assign n23357 = ( n7830 & n12750 ) | ( n7830 & n23356 ) | ( n12750 & n23356 ) ;
  assign n23358 = n13043 ^ n7236 ^ 1'b0 ;
  assign n23359 = ( n2405 & n14618 ) | ( n2405 & ~n23358 ) | ( n14618 & ~n23358 ) ;
  assign n23360 = n2970 & ~n9472 ;
  assign n23361 = n14986 ^ n2818 ^ 1'b0 ;
  assign n23362 = x4 & ~n10566 ;
  assign n23363 = ~n17050 & n23362 ;
  assign n23364 = n23361 | n23363 ;
  assign n23365 = ( n3203 & ~n12121 ) | ( n3203 & n15378 ) | ( ~n12121 & n15378 ) ;
  assign n23366 = n12228 & n19848 ;
  assign n23367 = ~n13842 & n15996 ;
  assign n23368 = n22860 ^ n4303 ^ 1'b0 ;
  assign n23369 = n13818 ^ n3391 ^ 1'b0 ;
  assign n23370 = n21888 ^ n11723 ^ 1'b0 ;
  assign n23371 = n23370 ^ n14968 ^ n264 ;
  assign n23372 = n10655 & n23371 ;
  assign n23373 = n6093 & ~n20332 ;
  assign n23374 = ~n11145 & n23373 ;
  assign n23375 = n735 & ~n13897 ;
  assign n23376 = n23374 & n23375 ;
  assign n23377 = ( n4730 & n11225 ) | ( n4730 & n21928 ) | ( n11225 & n21928 ) ;
  assign n23378 = ( n11385 & n23376 ) | ( n11385 & n23377 ) | ( n23376 & n23377 ) ;
  assign n23379 = ~n1176 & n10028 ;
  assign n23380 = n7725 | n20221 ;
  assign n23381 = n23380 ^ x129 ^ 1'b0 ;
  assign n23382 = n13089 ^ n10194 ^ n9530 ;
  assign n23383 = ~n6406 & n23382 ;
  assign n23384 = n939 | n23383 ;
  assign n23385 = n20343 | n23384 ;
  assign n23386 = ~n1671 & n3892 ;
  assign n23387 = n1711 & n23386 ;
  assign n23388 = ( n1385 & ~n1533 ) | ( n1385 & n23387 ) | ( ~n1533 & n23387 ) ;
  assign n23389 = ( n6137 & ~n11262 ) | ( n6137 & n23388 ) | ( ~n11262 & n23388 ) ;
  assign n23390 = n7630 & n23389 ;
  assign n23393 = ~n1733 & n4703 ;
  assign n23394 = ~n14847 & n23393 ;
  assign n23391 = n5030 & ~n8632 ;
  assign n23392 = n2991 & ~n23391 ;
  assign n23395 = n23394 ^ n23392 ^ n2201 ;
  assign n23396 = n18661 | n23395 ;
  assign n23397 = n18746 ^ n4101 ^ 1'b0 ;
  assign n23398 = ( n1034 & n11873 ) | ( n1034 & n23397 ) | ( n11873 & n23397 ) ;
  assign n23399 = n11861 ^ n8790 ^ 1'b0 ;
  assign n23400 = n14391 & ~n23399 ;
  assign n23401 = n23400 ^ n7206 ^ 1'b0 ;
  assign n23402 = n23401 ^ n20591 ^ n2090 ;
  assign n23405 = n7526 ^ n4038 ^ 1'b0 ;
  assign n23406 = n6646 & ~n23405 ;
  assign n23403 = n5245 | n12027 ;
  assign n23404 = n2908 & ~n23403 ;
  assign n23407 = n23406 ^ n23404 ^ n19738 ;
  assign n23408 = n7019 & ~n17587 ;
  assign n23409 = n23408 ^ n801 ^ 1'b0 ;
  assign n23410 = n7165 & ~n23409 ;
  assign n23411 = ~n3724 & n23410 ;
  assign n23412 = n22627 ^ n7070 ^ 1'b0 ;
  assign n23413 = ( n7665 & n17880 ) | ( n7665 & ~n23412 ) | ( n17880 & ~n23412 ) ;
  assign n23415 = n7291 & n11055 ;
  assign n23416 = ~n682 & n23415 ;
  assign n23414 = n10671 | n23253 ;
  assign n23417 = n23416 ^ n23414 ^ 1'b0 ;
  assign n23418 = n7060 ^ n3982 ^ n1989 ;
  assign n23419 = n23418 ^ n22782 ^ 1'b0 ;
  assign n23420 = n7885 & n23419 ;
  assign n23421 = n8777 ^ n5059 ^ n3344 ;
  assign n23422 = n19939 | n23421 ;
  assign n23423 = n13267 ^ n5464 ^ n3079 ;
  assign n23424 = n8828 & n10440 ;
  assign n23425 = n10543 & n23424 ;
  assign n23426 = n15912 & n17254 ;
  assign n23427 = ~n5185 & n18568 ;
  assign n23428 = n2236 & n23427 ;
  assign n23429 = ~n8907 & n23428 ;
  assign n23430 = n5797 & ~n15736 ;
  assign n23431 = n23430 ^ n15982 ^ 1'b0 ;
  assign n23432 = n21052 & n23431 ;
  assign n23433 = ~n9341 & n18055 ;
  assign n23434 = n20430 & n23433 ;
  assign n23435 = n9073 | n23434 ;
  assign n23436 = ~n5557 & n22447 ;
  assign n23437 = n23436 ^ n347 ^ 1'b0 ;
  assign n23438 = ( n11495 & n14948 ) | ( n11495 & ~n17052 ) | ( n14948 & ~n17052 ) ;
  assign n23439 = ~n18729 & n23438 ;
  assign n23440 = n4258 | n10898 ;
  assign n23441 = ( ~n17617 & n23439 ) | ( ~n17617 & n23440 ) | ( n23439 & n23440 ) ;
  assign n23442 = ( ~n4090 & n9363 ) | ( ~n4090 & n20955 ) | ( n9363 & n20955 ) ;
  assign n23443 = n10492 & n12812 ;
  assign n23444 = n2456 & n23443 ;
  assign n23445 = n6759 & n23444 ;
  assign n23447 = n8985 ^ n6164 ^ n5836 ;
  assign n23446 = n6793 & n9122 ;
  assign n23448 = n23447 ^ n23446 ^ 1'b0 ;
  assign n23449 = n4695 ^ n4652 ^ 1'b0 ;
  assign n23450 = ( ~n4271 & n23448 ) | ( ~n4271 & n23449 ) | ( n23448 & n23449 ) ;
  assign n23451 = ~n1164 & n4715 ;
  assign n23452 = ~n8339 & n23451 ;
  assign n23453 = n23452 ^ n8918 ^ 1'b0 ;
  assign n23454 = ~n5419 & n23453 ;
  assign n23455 = n8800 | n11723 ;
  assign n23456 = n23455 ^ n8815 ^ 1'b0 ;
  assign n23457 = n2270 & ~n23456 ;
  assign n23458 = n23457 ^ n9936 ^ 1'b0 ;
  assign n23459 = n8058 & ~n23458 ;
  assign n23460 = ~n1334 & n3085 ;
  assign n23461 = ~n3085 & n23460 ;
  assign n23462 = x2 & n16183 ;
  assign n23463 = ~n23461 & n23462 ;
  assign n23464 = ~n23048 & n23463 ;
  assign n23465 = n20481 ^ n13587 ^ 1'b0 ;
  assign n23466 = n3288 & n11822 ;
  assign n23467 = n5166 ^ n4996 ^ 1'b0 ;
  assign n23469 = n11897 ^ n1361 ^ 1'b0 ;
  assign n23470 = n763 & n23469 ;
  assign n23468 = n7661 ^ n7016 ^ n2783 ;
  assign n23471 = n23470 ^ n23468 ^ 1'b0 ;
  assign n23472 = ( n17685 & n23467 ) | ( n17685 & ~n23471 ) | ( n23467 & ~n23471 ) ;
  assign n23473 = n16485 ^ n483 ^ 1'b0 ;
  assign n23474 = n21460 & ~n23473 ;
  assign n23475 = n22877 ^ n9607 ^ 1'b0 ;
  assign n23476 = n13026 ^ n5002 ^ n427 ;
  assign n23477 = n23476 ^ n20739 ^ n11502 ;
  assign n23478 = n4997 ^ n729 ^ 1'b0 ;
  assign n23479 = n23477 | n23478 ;
  assign n23482 = n1441 ^ x84 ^ 1'b0 ;
  assign n23483 = n907 & ~n23482 ;
  assign n23480 = n4013 | n21919 ;
  assign n23481 = n8993 & ~n23480 ;
  assign n23484 = n23483 ^ n23481 ^ n16663 ;
  assign n23486 = n4731 & n19189 ;
  assign n23487 = n21894 & n23486 ;
  assign n23488 = n23487 ^ n10505 ^ n7100 ;
  assign n23485 = n4232 & n8045 ;
  assign n23489 = n23488 ^ n23485 ^ 1'b0 ;
  assign n23490 = n13418 & n13907 ;
  assign n23491 = ~n13418 & n23490 ;
  assign n23492 = ~n3481 & n7086 ;
  assign n23493 = n14454 & n23492 ;
  assign n23494 = n13869 & n19692 ;
  assign n23495 = ~n15157 & n23494 ;
  assign n23496 = n23495 ^ n16386 ^ 1'b0 ;
  assign n23497 = n949 | n17041 ;
  assign n23498 = n13058 ^ n9983 ^ 1'b0 ;
  assign n23499 = ( n3788 & n23497 ) | ( n3788 & ~n23498 ) | ( n23497 & ~n23498 ) ;
  assign n23500 = n11548 & n23499 ;
  assign n23504 = n20073 ^ n3322 ^ 1'b0 ;
  assign n23505 = n12065 & ~n23504 ;
  assign n23506 = n11010 & n23505 ;
  assign n23503 = ( n1069 & n4439 ) | ( n1069 & n12334 ) | ( n4439 & n12334 ) ;
  assign n23501 = n9707 | n14464 ;
  assign n23502 = n23501 ^ n13113 ^ 1'b0 ;
  assign n23507 = n23506 ^ n23503 ^ n23502 ;
  assign n23508 = ~n7829 & n7900 ;
  assign n23509 = n23508 ^ n15859 ^ 1'b0 ;
  assign n23510 = n6578 & n23509 ;
  assign n23512 = n8365 ^ n1980 ^ 1'b0 ;
  assign n23513 = n1966 | n6417 ;
  assign n23514 = n23513 ^ n13129 ^ 1'b0 ;
  assign n23515 = ~n5067 & n23514 ;
  assign n23516 = ~n23512 & n23515 ;
  assign n23511 = x216 & ~n391 ;
  assign n23517 = n23516 ^ n23511 ^ 1'b0 ;
  assign n23518 = ~n5311 & n14262 ;
  assign n23519 = ~n23517 & n23518 ;
  assign n23520 = n23510 & n23519 ;
  assign n23521 = n15836 ^ n14833 ^ n7517 ;
  assign n23522 = n16344 ^ n2649 ^ 1'b0 ;
  assign n23523 = n23522 ^ n8376 ^ 1'b0 ;
  assign n23524 = n15524 ^ n3235 ^ 1'b0 ;
  assign n23525 = n1916 | n23524 ;
  assign n23526 = n16715 & ~n23525 ;
  assign n23527 = ( n11873 & n12065 ) | ( n11873 & n12520 ) | ( n12065 & n12520 ) ;
  assign n23528 = ~n23526 & n23527 ;
  assign n23529 = n8578 & n21826 ;
  assign n23530 = n10072 & n23529 ;
  assign n23531 = n4875 ^ n958 ^ 1'b0 ;
  assign n23532 = ~n4807 & n23531 ;
  assign n23533 = ~n22839 & n23532 ;
  assign n23534 = n6518 ^ n1326 ^ n1307 ;
  assign n23535 = ( n2061 & n2770 ) | ( n2061 & n3640 ) | ( n2770 & n3640 ) ;
  assign n23536 = n23534 & ~n23535 ;
  assign n23537 = n23536 ^ n5419 ^ n3909 ;
  assign n23538 = n2183 | n7639 ;
  assign n23539 = n23538 ^ n4699 ^ 1'b0 ;
  assign n23540 = n8009 & n10002 ;
  assign n23541 = ~n23539 & n23540 ;
  assign n23542 = n23541 ^ x242 ^ 1'b0 ;
  assign n23543 = n1162 & ~n23542 ;
  assign n23544 = n13397 ^ n5485 ^ 1'b0 ;
  assign n23545 = n23544 ^ n16691 ^ n15410 ;
  assign n23546 = n23545 ^ n12329 ^ n768 ;
  assign n23547 = n12748 & ~n23546 ;
  assign n23548 = n23547 ^ n17001 ^ 1'b0 ;
  assign n23549 = ~n2541 & n13427 ;
  assign n23550 = n23549 ^ n16148 ^ 1'b0 ;
  assign n23551 = n23550 ^ n3192 ^ 1'b0 ;
  assign n23552 = n12314 ^ n6186 ^ 1'b0 ;
  assign n23553 = n23551 | n23552 ;
  assign n23555 = ( n4094 & ~n5196 ) | ( n4094 & n10470 ) | ( ~n5196 & n10470 ) ;
  assign n23556 = n23555 ^ n13861 ^ n8922 ;
  assign n23554 = n1160 & ~n5496 ;
  assign n23557 = n23556 ^ n23554 ^ 1'b0 ;
  assign n23558 = n23557 ^ n13254 ^ n10663 ;
  assign n23559 = n1053 & ~n6708 ;
  assign n23560 = n23559 ^ n16407 ^ 1'b0 ;
  assign n23561 = n18723 & n23560 ;
  assign n23564 = n13162 & ~n15225 ;
  assign n23565 = n23564 ^ n3508 ^ 1'b0 ;
  assign n23566 = n23565 ^ n10357 ^ 1'b0 ;
  assign n23567 = n7601 | n23566 ;
  assign n23563 = n4604 & ~n5879 ;
  assign n23562 = n19736 ^ n9599 ^ n3237 ;
  assign n23568 = n23567 ^ n23563 ^ n23562 ;
  assign n23569 = n21656 ^ n11156 ^ n3274 ;
  assign n23570 = n23569 ^ n17655 ^ 1'b0 ;
  assign n23571 = n12758 ^ n4986 ^ n4411 ;
  assign n23572 = n23571 ^ n18202 ^ 1'b0 ;
  assign n23573 = ~n1086 & n23572 ;
  assign n23574 = ( ~n3153 & n3157 ) | ( ~n3153 & n12617 ) | ( n3157 & n12617 ) ;
  assign n23575 = n22044 ^ n759 ^ 1'b0 ;
  assign n23576 = n14424 ^ n6406 ^ 1'b0 ;
  assign n23577 = n5065 & n23576 ;
  assign n23578 = n23577 ^ n8439 ^ 1'b0 ;
  assign n23579 = ~n11844 & n23578 ;
  assign n23580 = n17789 ^ n6910 ^ 1'b0 ;
  assign n23581 = ( n3437 & n18873 ) | ( n3437 & ~n23580 ) | ( n18873 & ~n23580 ) ;
  assign n23582 = n12813 ^ n2319 ^ 1'b0 ;
  assign n23583 = ~n638 & n7096 ;
  assign n23584 = n23583 ^ n22150 ^ 1'b0 ;
  assign n23585 = ~n12392 & n23584 ;
  assign n23586 = ~n8575 & n15044 ;
  assign n23587 = ~n11258 & n23586 ;
  assign n23588 = n16603 & ~n23587 ;
  assign n23589 = n1424 & n13030 ;
  assign n23590 = ~n23588 & n23589 ;
  assign n23591 = n23590 ^ n8276 ^ 1'b0 ;
  assign n23592 = n2275 | n23591 ;
  assign n23593 = n7950 | n11575 ;
  assign n23594 = n2808 & ~n23593 ;
  assign n23595 = n23592 & n23594 ;
  assign n23596 = n11368 | n11764 ;
  assign n23597 = n6494 ^ n1678 ^ 1'b0 ;
  assign n23598 = ~n16788 & n23597 ;
  assign n23599 = n22179 ^ n19499 ^ 1'b0 ;
  assign n23600 = ~n18387 & n23599 ;
  assign n23601 = n9754 & n22127 ;
  assign n23602 = ~n14252 & n23601 ;
  assign n23603 = n11875 | n23602 ;
  assign n23604 = n22386 ^ n21266 ^ n18037 ;
  assign n23605 = n23604 ^ n4041 ^ 1'b0 ;
  assign n23606 = n10080 & n23605 ;
  assign n23607 = n23606 ^ n11054 ^ n6328 ;
  assign n23609 = n10875 ^ n2937 ^ 1'b0 ;
  assign n23608 = ( n339 & ~n8164 ) | ( n339 & n11555 ) | ( ~n8164 & n11555 ) ;
  assign n23610 = n23609 ^ n23608 ^ 1'b0 ;
  assign n23611 = ~n3312 & n23610 ;
  assign n23612 = n18459 & ~n22930 ;
  assign n23613 = n23612 ^ n559 ^ 1'b0 ;
  assign n23614 = n5825 ^ n4342 ^ 1'b0 ;
  assign n23615 = n23614 ^ n17817 ^ 1'b0 ;
  assign n23616 = n4723 ^ n4606 ^ n2784 ;
  assign n23617 = n23616 ^ n10862 ^ n2997 ;
  assign n23618 = n19190 | n23617 ;
  assign n23619 = n23618 ^ n18119 ^ 1'b0 ;
  assign n23620 = n10068 & n18824 ;
  assign n23621 = n23619 & n23620 ;
  assign n23622 = n3539 | n4056 ;
  assign n23623 = n23622 ^ n3538 ^ 1'b0 ;
  assign n23624 = n9076 & ~n15687 ;
  assign n23625 = ~n5034 & n23624 ;
  assign n23626 = n23625 ^ n13484 ^ 1'b0 ;
  assign n23627 = n23623 | n23626 ;
  assign n23629 = n1364 | n21669 ;
  assign n23630 = x76 | n23629 ;
  assign n23634 = n19417 ^ n18598 ^ 1'b0 ;
  assign n23631 = n6936 ^ n1583 ^ n462 ;
  assign n23632 = n23631 ^ n20497 ^ 1'b0 ;
  assign n23633 = ~n12343 & n23632 ;
  assign n23635 = n23634 ^ n23633 ^ x100 ;
  assign n23636 = n7085 | n23635 ;
  assign n23637 = n23636 ^ n6919 ^ 1'b0 ;
  assign n23638 = n23630 & n23637 ;
  assign n23628 = ~n12635 & n23049 ;
  assign n23639 = n23638 ^ n23628 ^ 1'b0 ;
  assign n23640 = n17974 ^ n13207 ^ 1'b0 ;
  assign n23641 = n334 | n23640 ;
  assign n23642 = n4008 & n15812 ;
  assign n23643 = n10025 & n23642 ;
  assign n23644 = ( n19810 & ~n23641 ) | ( n19810 & n23643 ) | ( ~n23641 & n23643 ) ;
  assign n23645 = ( n6430 & n10109 ) | ( n6430 & n11173 ) | ( n10109 & n11173 ) ;
  assign n23646 = ( ~n6606 & n9948 ) | ( ~n6606 & n15010 ) | ( n9948 & n15010 ) ;
  assign n23647 = ( n4016 & n4414 ) | ( n4016 & n9745 ) | ( n4414 & n9745 ) ;
  assign n23648 = n3559 & n23647 ;
  assign n23649 = n23648 ^ n10050 ^ 1'b0 ;
  assign n23650 = ~n5001 & n23649 ;
  assign n23651 = n23650 ^ n8112 ^ 1'b0 ;
  assign n23652 = n20680 & n23651 ;
  assign n23653 = n11108 & n23652 ;
  assign n23654 = ~n14454 & n20613 ;
  assign n23655 = n22681 & n23654 ;
  assign n23656 = n7254 & ~n20019 ;
  assign n23657 = n13604 ^ n5526 ^ 1'b0 ;
  assign n23658 = n8529 | n23657 ;
  assign n23659 = ~n4323 & n18636 ;
  assign n23660 = n2940 & n16136 ;
  assign n23661 = n2401 | n23660 ;
  assign n23662 = n17995 & ~n19869 ;
  assign n23663 = n11555 ^ n6149 ^ 1'b0 ;
  assign n23664 = n14551 | n23663 ;
  assign n23665 = ( n8218 & ~n11437 ) | ( n8218 & n12828 ) | ( ~n11437 & n12828 ) ;
  assign n23666 = ( ~n9751 & n10941 ) | ( ~n9751 & n23665 ) | ( n10941 & n23665 ) ;
  assign n23667 = n15069 ^ n12147 ^ 1'b0 ;
  assign n23668 = n23666 & n23667 ;
  assign n23669 = n1797 & ~n3817 ;
  assign n23670 = ( n5519 & n10164 ) | ( n5519 & ~n19677 ) | ( n10164 & ~n19677 ) ;
  assign n23671 = n23670 ^ n13584 ^ 1'b0 ;
  assign n23672 = n23669 & ~n23671 ;
  assign n23673 = n8181 ^ n7590 ^ 1'b0 ;
  assign n23675 = ( n3791 & ~n6534 ) | ( n3791 & n7447 ) | ( ~n6534 & n7447 ) ;
  assign n23676 = ~n825 & n23675 ;
  assign n23677 = n23676 ^ n19329 ^ n12334 ;
  assign n23674 = ( n11031 & n13343 ) | ( n11031 & ~n23184 ) | ( n13343 & ~n23184 ) ;
  assign n23678 = n23677 ^ n23674 ^ x223 ;
  assign n23679 = n11722 ^ n10050 ^ n5311 ;
  assign n23682 = x108 & ~n2494 ;
  assign n23683 = n8913 & n23682 ;
  assign n23684 = ~n2124 & n2683 ;
  assign n23685 = n23684 ^ n2140 ^ 1'b0 ;
  assign n23686 = n2644 & ~n23685 ;
  assign n23687 = ( n22951 & n23683 ) | ( n22951 & ~n23686 ) | ( n23683 & ~n23686 ) ;
  assign n23680 = n16899 ^ n5351 ^ 1'b0 ;
  assign n23681 = n3960 | n23680 ;
  assign n23688 = n23687 ^ n23681 ^ 1'b0 ;
  assign n23689 = n6865 | n16972 ;
  assign n23690 = ( ~n516 & n4392 ) | ( ~n516 & n5655 ) | ( n4392 & n5655 ) ;
  assign n23691 = n23690 ^ n1267 ^ n1141 ;
  assign n23692 = ~n10500 & n11258 ;
  assign n23693 = n23692 ^ n544 ^ 1'b0 ;
  assign n23694 = n9402 ^ n1172 ^ 1'b0 ;
  assign n23695 = n4396 & ~n19926 ;
  assign n23696 = n23694 & n23695 ;
  assign n23697 = n7206 | n23696 ;
  assign n23698 = ( x136 & n6189 ) | ( x136 & ~n13738 ) | ( n6189 & ~n13738 ) ;
  assign n23699 = n11348 ^ n6522 ^ n877 ;
  assign n23703 = n8473 | n11531 ;
  assign n23704 = ~n3064 & n12129 ;
  assign n23705 = n23703 & n23704 ;
  assign n23700 = n8025 | n11028 ;
  assign n23701 = x158 & ~n2489 ;
  assign n23702 = n23700 & n23701 ;
  assign n23706 = n23705 ^ n23702 ^ n15239 ;
  assign n23707 = ~n17214 & n23706 ;
  assign n23708 = ~n23699 & n23707 ;
  assign n23709 = n23708 ^ n12914 ^ 1'b0 ;
  assign n23710 = x243 & ~n23709 ;
  assign n23711 = n4752 ^ n4321 ^ 1'b0 ;
  assign n23712 = ~n8465 & n23711 ;
  assign n23713 = n23712 ^ n6626 ^ n2977 ;
  assign n23714 = n6994 ^ n3905 ^ 1'b0 ;
  assign n23715 = n1533 | n23714 ;
  assign n23716 = n16769 ^ n14636 ^ 1'b0 ;
  assign n23717 = n461 & ~n23716 ;
  assign n23718 = n6499 & ~n9932 ;
  assign n23719 = n3079 | n23718 ;
  assign n23720 = n23719 ^ n11995 ^ 1'b0 ;
  assign n23721 = n10145 ^ n3654 ^ n2296 ;
  assign n23722 = n2551 & n23721 ;
  assign n23723 = n18033 & n23722 ;
  assign n23724 = n2585 & ~n20275 ;
  assign n23725 = n3531 ^ n3057 ^ 1'b0 ;
  assign n23726 = n3868 & ~n23725 ;
  assign n23727 = n1970 & n2312 ;
  assign n23728 = ~n15373 & n23727 ;
  assign n23729 = ( ~n4136 & n9247 ) | ( ~n4136 & n12493 ) | ( n9247 & n12493 ) ;
  assign n23730 = n16947 & n23729 ;
  assign n23731 = n5636 | n15568 ;
  assign n23732 = n22619 ^ n16140 ^ 1'b0 ;
  assign n23733 = n3104 & ~n18939 ;
  assign n23735 = n9858 & ~n13942 ;
  assign n23734 = n16476 | n22831 ;
  assign n23736 = n23735 ^ n23734 ^ 1'b0 ;
  assign n23744 = n10521 ^ n1288 ^ 1'b0 ;
  assign n23742 = n2227 | n15468 ;
  assign n23743 = n23742 ^ n2562 ^ 1'b0 ;
  assign n23740 = x128 & ~n5072 ;
  assign n23741 = n23740 ^ n11351 ^ 1'b0 ;
  assign n23745 = n23744 ^ n23743 ^ n23741 ;
  assign n23737 = n1843 ^ n1061 ^ 1'b0 ;
  assign n23738 = n3572 & ~n23737 ;
  assign n23739 = n3090 & n23738 ;
  assign n23746 = n23745 ^ n23739 ^ 1'b0 ;
  assign n23747 = ~n1582 & n4141 ;
  assign n23748 = ~n1969 & n23747 ;
  assign n23749 = ( n8587 & n17294 ) | ( n8587 & n23748 ) | ( n17294 & n23748 ) ;
  assign n23750 = n23057 | n23749 ;
  assign n23751 = n23750 ^ n18732 ^ 1'b0 ;
  assign n23752 = n16148 ^ n15526 ^ 1'b0 ;
  assign n23753 = n15838 | n23752 ;
  assign n23754 = n23753 ^ n5795 ^ 1'b0 ;
  assign n23761 = x82 & ~n1327 ;
  assign n23755 = n369 | n3144 ;
  assign n23756 = n9493 | n23755 ;
  assign n23757 = n11113 ^ n9327 ^ n5762 ;
  assign n23758 = n23757 ^ n9123 ^ n460 ;
  assign n23759 = n23758 ^ n11342 ^ 1'b0 ;
  assign n23760 = n23756 & n23759 ;
  assign n23762 = n23761 ^ n23760 ^ 1'b0 ;
  assign n23764 = n1439 & n7963 ;
  assign n23763 = n14319 | n22564 ;
  assign n23765 = n23764 ^ n23763 ^ 1'b0 ;
  assign n23766 = ( n3115 & ~n7392 ) | ( n3115 & n9761 ) | ( ~n7392 & n9761 ) ;
  assign n23767 = n21956 ^ n17521 ^ 1'b0 ;
  assign n23768 = n8457 & ~n23767 ;
  assign n23771 = n18529 ^ n14870 ^ 1'b0 ;
  assign n23772 = n16561 ^ n5196 ^ 1'b0 ;
  assign n23773 = n23771 & n23772 ;
  assign n23774 = ( ~n10172 & n22990 ) | ( ~n10172 & n23773 ) | ( n22990 & n23773 ) ;
  assign n23769 = n4845 ^ n4729 ^ 1'b0 ;
  assign n23770 = n20070 & ~n23769 ;
  assign n23775 = n23774 ^ n23770 ^ 1'b0 ;
  assign n23776 = ( n5006 & n6100 ) | ( n5006 & ~n11782 ) | ( n6100 & ~n11782 ) ;
  assign n23777 = n5453 ^ n1015 ^ 1'b0 ;
  assign n23778 = n23777 ^ n10626 ^ 1'b0 ;
  assign n23779 = n17761 ^ n17700 ^ 1'b0 ;
  assign n23780 = n4763 & ~n23779 ;
  assign n23781 = n11819 & n18944 ;
  assign n23782 = n23781 ^ n11100 ^ x70 ;
  assign n23784 = n982 & n10875 ;
  assign n23783 = n8181 & ~n11583 ;
  assign n23785 = n23784 ^ n23783 ^ n16800 ;
  assign n23786 = n4240 & ~n15552 ;
  assign n23787 = ~n9430 & n23786 ;
  assign n23788 = n11112 ^ n5111 ^ 1'b0 ;
  assign n23789 = n10470 & ~n23788 ;
  assign n23790 = n23789 ^ n3024 ^ 1'b0 ;
  assign n23792 = n22430 ^ n3100 ^ 1'b0 ;
  assign n23791 = n4572 & n9749 ;
  assign n23793 = n23792 ^ n23791 ^ 1'b0 ;
  assign n23794 = ~n4270 & n6944 ;
  assign n23795 = n5237 ^ n5060 ^ n3343 ;
  assign n23796 = n4538 | n23795 ;
  assign n23797 = n23796 ^ n4298 ^ 1'b0 ;
  assign n23798 = n9963 ^ n7058 ^ 1'b0 ;
  assign n23799 = n23798 ^ n11142 ^ 1'b0 ;
  assign n23800 = n23799 ^ n11009 ^ 1'b0 ;
  assign n23801 = n23797 & ~n23800 ;
  assign n23802 = n8678 ^ n7553 ^ 1'b0 ;
  assign n23803 = n22478 | n23802 ;
  assign n23804 = n13220 ^ n9344 ^ 1'b0 ;
  assign n23805 = n20693 ^ n10262 ^ 1'b0 ;
  assign n23806 = ~n3333 & n20474 ;
  assign n23807 = n14208 ^ n7154 ^ n4878 ;
  assign n23808 = n7727 & ~n23807 ;
  assign n23809 = n21834 ^ n6297 ^ 1'b0 ;
  assign n23810 = ~n3957 & n23809 ;
  assign n23811 = ( n13439 & ~n23808 ) | ( n13439 & n23810 ) | ( ~n23808 & n23810 ) ;
  assign n23812 = n8929 & n13657 ;
  assign n23813 = n6358 & n23812 ;
  assign n23814 = n22403 ^ n2001 ^ 1'b0 ;
  assign n23815 = n21188 & n23814 ;
  assign n23816 = n18376 | n22278 ;
  assign n23817 = n16431 & n23816 ;
  assign n23818 = n23817 ^ n11805 ^ 1'b0 ;
  assign n23819 = n5518 & ~n9327 ;
  assign n23820 = n23819 ^ n6137 ^ 1'b0 ;
  assign n23821 = n10174 ^ x15 ^ 1'b0 ;
  assign n23822 = n14137 & ~n23821 ;
  assign n23823 = ( n11152 & ~n23820 ) | ( n11152 & n23822 ) | ( ~n23820 & n23822 ) ;
  assign n23824 = ( n1154 & ~n10568 ) | ( n1154 & n16366 ) | ( ~n10568 & n16366 ) ;
  assign n23825 = x223 & ~n2885 ;
  assign n23826 = ( n4799 & ~n11501 ) | ( n4799 & n23825 ) | ( ~n11501 & n23825 ) ;
  assign n23827 = n6253 | n10835 ;
  assign n23828 = n5892 | n15875 ;
  assign n23829 = n7457 & ~n7867 ;
  assign n23830 = n23829 ^ n4288 ^ 1'b0 ;
  assign n23831 = n5360 ^ n4130 ^ n1875 ;
  assign n23832 = n8821 ^ n3296 ^ 1'b0 ;
  assign n23833 = ~n23831 & n23832 ;
  assign n23834 = n4277 & n7260 ;
  assign n23835 = n23834 ^ n6769 ^ 1'b0 ;
  assign n23836 = n15202 | n23835 ;
  assign n23837 = n1474 | n23836 ;
  assign n23838 = n5199 & n13629 ;
  assign n23839 = ~n23837 & n23838 ;
  assign n23840 = n10073 ^ n4217 ^ 1'b0 ;
  assign n23841 = n23840 ^ n11791 ^ 1'b0 ;
  assign n23842 = n4615 & n23841 ;
  assign n23846 = x224 & n3474 ;
  assign n23847 = n3172 & n23846 ;
  assign n23843 = ~n8387 & n8916 ;
  assign n23844 = n23843 ^ n1932 ^ 1'b0 ;
  assign n23845 = n23844 ^ n3286 ^ 1'b0 ;
  assign n23848 = n23847 ^ n23845 ^ n20129 ;
  assign n23849 = n16413 ^ n7196 ^ 1'b0 ;
  assign n23850 = n17860 & n23849 ;
  assign n23851 = n6549 | n6689 ;
  assign n23856 = ~n8172 & n15010 ;
  assign n23857 = n9634 & n23856 ;
  assign n23858 = n23857 ^ n12941 ^ n1773 ;
  assign n23852 = n2843 & ~n7163 ;
  assign n23853 = ( n3656 & ~n8757 ) | ( n3656 & n23852 ) | ( ~n8757 & n23852 ) ;
  assign n23854 = n23853 ^ n15435 ^ 1'b0 ;
  assign n23855 = n22854 & ~n23854 ;
  assign n23859 = n23858 ^ n23855 ^ 1'b0 ;
  assign n23860 = n13218 ^ n3312 ^ 1'b0 ;
  assign n23861 = n23860 ^ n17647 ^ n3932 ;
  assign n23862 = n2970 & n4258 ;
  assign n23863 = n12933 & n23862 ;
  assign n23864 = n2399 & n23863 ;
  assign n23865 = n23864 ^ n23513 ^ n9386 ;
  assign n23867 = n4888 | n7655 ;
  assign n23866 = ~n5662 & n8323 ;
  assign n23868 = n23867 ^ n23866 ^ 1'b0 ;
  assign n23869 = n23868 ^ n21941 ^ 1'b0 ;
  assign n23870 = n6642 | n17562 ;
  assign n23871 = n23870 ^ n4451 ^ 1'b0 ;
  assign n23876 = n17952 ^ n17175 ^ n13155 ;
  assign n23874 = n3414 ^ n3401 ^ 1'b0 ;
  assign n23872 = n2226 | n2674 ;
  assign n23873 = n23872 ^ n18479 ^ 1'b0 ;
  assign n23875 = n23874 ^ n23873 ^ n16471 ;
  assign n23877 = n23876 ^ n23875 ^ n17416 ;
  assign n23878 = n2804 | n10348 ;
  assign n23879 = n4743 | n23878 ;
  assign n23880 = n23879 ^ n4112 ^ 1'b0 ;
  assign n23881 = ~n12341 & n23880 ;
  assign n23882 = n10640 & n23881 ;
  assign n23883 = n23882 ^ n8454 ^ 1'b0 ;
  assign n23884 = n20924 ^ n7483 ^ n4482 ;
  assign n23885 = n23884 ^ n9464 ^ 1'b0 ;
  assign n23886 = n23885 ^ n4847 ^ 1'b0 ;
  assign n23887 = x143 & n8076 ;
  assign n23888 = n10116 & n14700 ;
  assign n23889 = n23887 | n23888 ;
  assign n23890 = n23889 ^ n15074 ^ 1'b0 ;
  assign n23891 = n16416 ^ n3197 ^ 1'b0 ;
  assign n23892 = n23306 ^ n17443 ^ 1'b0 ;
  assign n23893 = n23892 ^ n18805 ^ 1'b0 ;
  assign n23894 = n15477 & ~n19164 ;
  assign n23895 = n23894 ^ n8826 ^ 1'b0 ;
  assign n23898 = n12039 & n14382 ;
  assign n23899 = n1677 | n23898 ;
  assign n23900 = n23899 ^ n1079 ^ 1'b0 ;
  assign n23896 = n3677 | n11795 ;
  assign n23897 = n23896 ^ n5913 ^ n884 ;
  assign n23901 = n23900 ^ n23897 ^ 1'b0 ;
  assign n23902 = n23901 ^ n17808 ^ 1'b0 ;
  assign n23903 = n21398 ^ n7039 ^ 1'b0 ;
  assign n23904 = n7002 & n23903 ;
  assign n23905 = n10839 & n23904 ;
  assign n23906 = n9852 ^ n9779 ^ 1'b0 ;
  assign n23907 = ( n10383 & n14487 ) | ( n10383 & ~n23906 ) | ( n14487 & ~n23906 ) ;
  assign n23908 = n3755 & ~n5077 ;
  assign n23909 = n23908 ^ n1016 ^ 1'b0 ;
  assign n23910 = n17170 & ~n23909 ;
  assign n23911 = n715 & ~n21914 ;
  assign n23912 = n23911 ^ n3376 ^ 1'b0 ;
  assign n23913 = n2099 ^ n1895 ^ 1'b0 ;
  assign n23914 = n3688 & n23913 ;
  assign n23915 = n23914 ^ n6102 ^ 1'b0 ;
  assign n23916 = n17599 & n23915 ;
  assign n23917 = n23916 ^ n10201 ^ 1'b0 ;
  assign n23918 = ( ~n17715 & n19513 ) | ( ~n17715 & n23917 ) | ( n19513 & n23917 ) ;
  assign n23919 = n22534 ^ n15325 ^ n6879 ;
  assign n23920 = n23294 ^ n17334 ^ n16020 ;
  assign n23921 = n18715 | n23920 ;
  assign n23922 = n9402 ^ n1455 ^ 1'b0 ;
  assign n23924 = x35 & n2418 ;
  assign n23925 = n23924 ^ n17995 ^ 1'b0 ;
  assign n23926 = n23925 ^ n15476 ^ 1'b0 ;
  assign n23927 = n23926 ^ n12265 ^ n9764 ;
  assign n23923 = n5186 & n14428 ;
  assign n23928 = n23927 ^ n23923 ^ 1'b0 ;
  assign n23929 = n19408 ^ n6498 ^ 1'b0 ;
  assign n23930 = n15955 ^ x126 ^ 1'b0 ;
  assign n23931 = n11259 & ~n11907 ;
  assign n23932 = n10016 & n23931 ;
  assign n23933 = n23932 ^ n15877 ^ 1'b0 ;
  assign n23934 = n12071 & n12656 ;
  assign n23935 = n23933 & n23934 ;
  assign n23936 = n3730 & ~n9118 ;
  assign n23937 = n23936 ^ x102 ^ 1'b0 ;
  assign n23938 = n15086 ^ n8957 ^ 1'b0 ;
  assign n23939 = n19810 ^ n14572 ^ 1'b0 ;
  assign n23940 = n4592 | n6018 ;
  assign n23941 = n23940 ^ n14498 ^ 1'b0 ;
  assign n23942 = n23941 ^ n17307 ^ n13436 ;
  assign n23943 = n6463 ^ n4373 ^ 1'b0 ;
  assign n23944 = n23943 ^ n11750 ^ n1265 ;
  assign n23945 = n23944 ^ n12023 ^ 1'b0 ;
  assign n23946 = n8999 ^ n3619 ^ 1'b0 ;
  assign n23947 = n16817 & n23946 ;
  assign n23948 = n12256 ^ n1035 ^ 1'b0 ;
  assign n23949 = x80 & ~n23948 ;
  assign n23950 = ~n5618 & n12700 ;
  assign n23951 = n23950 ^ n9611 ^ 1'b0 ;
  assign n23952 = x158 | n13994 ;
  assign n23953 = n6706 ^ n5156 ^ 1'b0 ;
  assign n23954 = n13896 ^ n8842 ^ 1'b0 ;
  assign n23955 = n23953 | n23954 ;
  assign n23956 = ~n8806 & n23955 ;
  assign n23957 = n17455 ^ n10891 ^ n6318 ;
  assign n23958 = n9281 | n21884 ;
  assign n23959 = n23958 ^ n12883 ^ 1'b0 ;
  assign n23962 = n323 & ~n7842 ;
  assign n23963 = n884 & n23962 ;
  assign n23967 = ~x56 & n7858 ;
  assign n23968 = n610 & n1993 ;
  assign n23969 = n14605 & ~n23968 ;
  assign n23970 = n23967 & n23969 ;
  assign n23965 = n7161 ^ n3710 ^ 1'b0 ;
  assign n23964 = n996 & n5792 ;
  assign n23966 = n23965 ^ n23964 ^ 1'b0 ;
  assign n23971 = n23970 ^ n23966 ^ 1'b0 ;
  assign n23972 = ~n9146 & n23971 ;
  assign n23973 = n11587 & n23972 ;
  assign n23974 = ( n2403 & ~n23963 ) | ( n2403 & n23973 ) | ( ~n23963 & n23973 ) ;
  assign n23960 = n8960 ^ n3338 ^ 1'b0 ;
  assign n23961 = n13791 & n23960 ;
  assign n23975 = n23974 ^ n23961 ^ n8774 ;
  assign n23976 = ( n2401 & ~n23118 ) | ( n2401 & n23664 ) | ( ~n23118 & n23664 ) ;
  assign n23977 = n4932 & ~n21132 ;
  assign n23978 = n12947 ^ n12710 ^ 1'b0 ;
  assign n23979 = n2899 & ~n6225 ;
  assign n23980 = ~n23978 & n23979 ;
  assign n23981 = n13546 ^ n2692 ^ n632 ;
  assign n23982 = n23981 ^ n18954 ^ n16908 ;
  assign n23983 = n10267 & ~n22852 ;
  assign n23984 = n5437 & n23983 ;
  assign n23985 = n23984 ^ n12521 ^ 1'b0 ;
  assign n23986 = n6310 & n7963 ;
  assign n23987 = n23986 ^ n8967 ^ 1'b0 ;
  assign n23988 = ( n317 & n10856 ) | ( n317 & ~n20634 ) | ( n10856 & ~n20634 ) ;
  assign n23989 = n23988 ^ n1553 ^ 1'b0 ;
  assign n23990 = n16270 & n23989 ;
  assign n23991 = n21545 ^ n2551 ^ 1'b0 ;
  assign n23992 = n17458 & ~n23991 ;
  assign n23993 = ( ~n6160 & n22387 ) | ( ~n6160 & n23992 ) | ( n22387 & n23992 ) ;
  assign n23994 = n20925 ^ n7525 ^ 1'b0 ;
  assign n23995 = n22715 & n23994 ;
  assign n23996 = n18849 ^ n1862 ^ 1'b0 ;
  assign n23997 = n3091 & ~n13200 ;
  assign n23998 = n23997 ^ n9283 ^ 1'b0 ;
  assign n23999 = n358 | n4263 ;
  assign n24000 = n4950 | n23999 ;
  assign n24002 = n5934 ^ n2386 ^ 1'b0 ;
  assign n24001 = n3161 | n18045 ;
  assign n24003 = n24002 ^ n24001 ^ 1'b0 ;
  assign n24004 = n24003 ^ n16109 ^ 1'b0 ;
  assign n24005 = ~n8230 & n11860 ;
  assign n24006 = n19670 & ~n24005 ;
  assign n24007 = n24006 ^ n5592 ^ 1'b0 ;
  assign n24008 = ( n24000 & ~n24004 ) | ( n24000 & n24007 ) | ( ~n24004 & n24007 ) ;
  assign n24009 = ~n9286 & n13605 ;
  assign n24010 = n24009 ^ n3357 ^ 1'b0 ;
  assign n24011 = ~n3502 & n12889 ;
  assign n24012 = n24011 ^ n11500 ^ 1'b0 ;
  assign n24013 = n24012 ^ n5264 ^ n268 ;
  assign n24014 = ~n10459 & n24013 ;
  assign n24015 = n24014 ^ n3087 ^ 1'b0 ;
  assign n24016 = n24015 ^ n12679 ^ 1'b0 ;
  assign n24017 = n10044 & ~n12520 ;
  assign n24018 = n5500 & n9278 ;
  assign n24019 = n24018 ^ n7589 ^ 1'b0 ;
  assign n24020 = n24019 ^ n17300 ^ n17111 ;
  assign n24021 = n3634 & ~n22865 ;
  assign n24022 = n24021 ^ n21274 ^ 1'b0 ;
  assign n24023 = n3776 & ~n11031 ;
  assign n24024 = n24023 ^ n1494 ^ 1'b0 ;
  assign n24025 = n24024 ^ n7864 ^ 1'b0 ;
  assign n24026 = n22990 ^ n13587 ^ 1'b0 ;
  assign n24027 = n24025 & n24026 ;
  assign n24028 = n3345 & n23992 ;
  assign n24029 = n24028 ^ n18706 ^ 1'b0 ;
  assign n24030 = ( n4690 & n5543 ) | ( n4690 & ~n20952 ) | ( n5543 & ~n20952 ) ;
  assign n24033 = n8208 & n19866 ;
  assign n24031 = n485 & n19499 ;
  assign n24032 = n24031 ^ n18462 ^ 1'b0 ;
  assign n24034 = n24033 ^ n24032 ^ 1'b0 ;
  assign n24035 = ( n2247 & ~n2760 ) | ( n2247 & n9232 ) | ( ~n2760 & n9232 ) ;
  assign n24036 = n8100 & ~n17661 ;
  assign n24037 = ~n24035 & n24036 ;
  assign n24038 = n11805 | n24037 ;
  assign n24039 = n7503 ^ n7152 ^ 1'b0 ;
  assign n24040 = n5557 | n5564 ;
  assign n24041 = n24039 & ~n24040 ;
  assign n24042 = n3356 & ~n11230 ;
  assign n24043 = n24042 ^ n14099 ^ 1'b0 ;
  assign n24044 = ~n6792 & n8084 ;
  assign n24045 = ( ~x244 & n12506 ) | ( ~x244 & n23064 ) | ( n12506 & n23064 ) ;
  assign n24047 = n402 & ~n5721 ;
  assign n24046 = n3855 | n20306 ;
  assign n24048 = n24047 ^ n24046 ^ 1'b0 ;
  assign n24049 = n21329 ^ n9174 ^ 1'b0 ;
  assign n24050 = n10866 | n24049 ;
  assign n24051 = ( n3252 & n12487 ) | ( n3252 & n14907 ) | ( n12487 & n14907 ) ;
  assign n24052 = n24051 ^ n7232 ^ 1'b0 ;
  assign n24053 = n2339 & ~n24052 ;
  assign n24054 = n931 & n24053 ;
  assign n24055 = n15965 & n24054 ;
  assign n24060 = n19408 ^ n12027 ^ 1'b0 ;
  assign n24061 = ~n15936 & n24060 ;
  assign n24062 = n24061 ^ n4422 ^ 1'b0 ;
  assign n24056 = n7795 & n8613 ;
  assign n24057 = n24056 ^ n9068 ^ 1'b0 ;
  assign n24058 = n24057 ^ n13029 ^ x31 ;
  assign n24059 = n22292 & n24058 ;
  assign n24063 = n24062 ^ n24059 ^ 1'b0 ;
  assign n24066 = n2145 & ~n2791 ;
  assign n24067 = n17513 & n24066 ;
  assign n24064 = n19868 | n19883 ;
  assign n24065 = n11472 & ~n24064 ;
  assign n24068 = n24067 ^ n24065 ^ n16478 ;
  assign n24069 = n14048 ^ n1998 ^ 1'b0 ;
  assign n24070 = n14489 & n24069 ;
  assign n24071 = n1175 & n11185 ;
  assign n24072 = n24070 & ~n24071 ;
  assign n24073 = ~n2598 & n18771 ;
  assign n24074 = ~n24072 & n24073 ;
  assign n24075 = n16458 ^ n10573 ^ 1'b0 ;
  assign n24076 = n16081 ^ n12553 ^ 1'b0 ;
  assign n24078 = n2228 | n6316 ;
  assign n24077 = n2394 & n8969 ;
  assign n24079 = n24078 ^ n24077 ^ n22940 ;
  assign n24080 = n24076 & n24079 ;
  assign n24081 = n24080 ^ n4987 ^ 1'b0 ;
  assign n24082 = ~n262 & n1194 ;
  assign n24083 = n24082 ^ n12679 ^ 1'b0 ;
  assign n24089 = n4743 ^ n752 ^ 1'b0 ;
  assign n24084 = n1566 & ~n2453 ;
  assign n24085 = n6249 & n24084 ;
  assign n24086 = n24085 ^ n6663 ^ n6130 ;
  assign n24087 = n24086 ^ n23455 ^ 1'b0 ;
  assign n24088 = n18458 | n24087 ;
  assign n24090 = n24089 ^ n24088 ^ 1'b0 ;
  assign n24092 = ~n7200 & n12519 ;
  assign n24091 = ~n7758 & n8084 ;
  assign n24093 = n24092 ^ n24091 ^ 1'b0 ;
  assign n24097 = n5973 | n18552 ;
  assign n24096 = n4793 & n14114 ;
  assign n24094 = n5112 ^ n1044 ^ 1'b0 ;
  assign n24095 = ( n6276 & n17148 ) | ( n6276 & ~n24094 ) | ( n17148 & ~n24094 ) ;
  assign n24098 = n24097 ^ n24096 ^ n24095 ;
  assign n24099 = n13735 & n21033 ;
  assign n24100 = n24099 ^ n958 ^ 1'b0 ;
  assign n24101 = n19784 ^ n2917 ^ 1'b0 ;
  assign n24103 = ( ~n1409 & n1729 ) | ( ~n1409 & n17082 ) | ( n1729 & n17082 ) ;
  assign n24104 = ~n12300 & n24103 ;
  assign n24105 = n9296 ^ n8420 ^ 1'b0 ;
  assign n24106 = n24104 & n24105 ;
  assign n24102 = n996 & ~n4357 ;
  assign n24107 = n24106 ^ n24102 ^ 1'b0 ;
  assign n24108 = n8332 | n15821 ;
  assign n24109 = n15851 & ~n24108 ;
  assign n24110 = n4993 ^ n3980 ^ 1'b0 ;
  assign n24111 = n3153 & n24110 ;
  assign n24112 = ~n7450 & n24111 ;
  assign n24113 = ( ~n1407 & n2645 ) | ( ~n1407 & n7929 ) | ( n2645 & n7929 ) ;
  assign n24114 = ( n12544 & ~n15106 ) | ( n12544 & n24113 ) | ( ~n15106 & n24113 ) ;
  assign n24115 = n1409 | n24114 ;
  assign n24116 = n24115 ^ n22870 ^ 1'b0 ;
  assign n24117 = x250 & ~n4822 ;
  assign n24118 = n24116 & n24117 ;
  assign n24119 = ( n15035 & n20876 ) | ( n15035 & ~n24118 ) | ( n20876 & ~n24118 ) ;
  assign n24120 = n5818 | n16130 ;
  assign n24121 = n14980 ^ n3327 ^ 1'b0 ;
  assign n24122 = n10770 & n24121 ;
  assign n24123 = ( n1602 & ~n24120 ) | ( n1602 & n24122 ) | ( ~n24120 & n24122 ) ;
  assign n24124 = n15014 ^ x218 ^ 1'b0 ;
  assign n24125 = n12841 & ~n21600 ;
  assign n24126 = ~n9755 & n24125 ;
  assign n24127 = ( n4542 & n21221 ) | ( n4542 & n24126 ) | ( n21221 & n24126 ) ;
  assign n24128 = ( n2516 & n3291 ) | ( n2516 & ~n3845 ) | ( n3291 & ~n3845 ) ;
  assign n24129 = n1320 & n19342 ;
  assign n24130 = n15986 ^ n11692 ^ 1'b0 ;
  assign n24131 = ~n24129 & n24130 ;
  assign n24132 = n24131 ^ n14264 ^ 1'b0 ;
  assign n24133 = ~n4893 & n24132 ;
  assign n24134 = n4995 ^ n2216 ^ 1'b0 ;
  assign n24135 = n9214 & n24134 ;
  assign n24136 = ~n2151 & n18848 ;
  assign n24137 = n15148 ^ n10691 ^ n2551 ;
  assign n24138 = n19772 ^ n16301 ^ n15944 ;
  assign n24139 = n4696 ^ n1248 ^ 1'b0 ;
  assign n24140 = n7940 ^ n6744 ^ 1'b0 ;
  assign n24141 = n8309 & ~n24140 ;
  assign n24142 = n1420 | n4253 ;
  assign n24143 = n24142 ^ n10976 ^ 1'b0 ;
  assign n24144 = n24141 & ~n24143 ;
  assign n24145 = n14405 & n24144 ;
  assign n24146 = n9478 ^ n5816 ^ 1'b0 ;
  assign n24149 = n22802 ^ n3776 ^ 1'b0 ;
  assign n24150 = n8559 & ~n24149 ;
  assign n24147 = n3317 | n6846 ;
  assign n24148 = n24147 ^ n10998 ^ 1'b0 ;
  assign n24151 = n24150 ^ n24148 ^ 1'b0 ;
  assign n24152 = n24146 & n24151 ;
  assign n24153 = n24060 ^ n9044 ^ 1'b0 ;
  assign n24154 = n24153 ^ n16867 ^ 1'b0 ;
  assign n24155 = n22838 | n24154 ;
  assign n24156 = n24155 ^ n14107 ^ 1'b0 ;
  assign n24157 = n375 | n5676 ;
  assign n24158 = n24157 ^ n2823 ^ 1'b0 ;
  assign n24159 = ~n13074 & n24158 ;
  assign n24160 = n24159 ^ n5228 ^ 1'b0 ;
  assign n24161 = n20668 ^ n13291 ^ n9676 ;
  assign n24162 = n13407 ^ n2178 ^ 1'b0 ;
  assign n24163 = n11046 ^ n6674 ^ 1'b0 ;
  assign n24164 = n8949 & n24163 ;
  assign n24165 = ( n4109 & n21520 ) | ( n4109 & n24164 ) | ( n21520 & n24164 ) ;
  assign n24166 = n6293 ^ n1321 ^ x128 ;
  assign n24167 = n1018 & n13348 ;
  assign n24168 = n7819 & n24167 ;
  assign n24169 = ~n3168 & n24168 ;
  assign n24170 = n24166 | n24169 ;
  assign n24171 = ( n1261 & n2927 ) | ( n1261 & ~n4845 ) | ( n2927 & ~n4845 ) ;
  assign n24172 = n24171 ^ n10853 ^ 1'b0 ;
  assign n24173 = n2580 & n5258 ;
  assign n24174 = n24173 ^ n14379 ^ 1'b0 ;
  assign n24175 = n24172 & ~n24174 ;
  assign n24176 = ( n777 & ~n2874 ) | ( n777 & n14874 ) | ( ~n2874 & n14874 ) ;
  assign n24177 = n460 & ~n22141 ;
  assign n24178 = ~n24176 & n24177 ;
  assign n24179 = ( n3408 & n9101 ) | ( n3408 & ~n9592 ) | ( n9101 & ~n9592 ) ;
  assign n24180 = n24179 ^ n8013 ^ 1'b0 ;
  assign n24181 = ~n17270 & n24180 ;
  assign n24188 = n7715 ^ n3310 ^ 1'b0 ;
  assign n24189 = n24188 ^ n1550 ^ 1'b0 ;
  assign n24190 = n2448 & ~n24189 ;
  assign n24184 = ~n8027 & n11321 ;
  assign n24182 = n9740 ^ n8894 ^ n1447 ;
  assign n24183 = n9558 | n24182 ;
  assign n24185 = n24184 ^ n24183 ^ 1'b0 ;
  assign n24186 = n16605 & n24185 ;
  assign n24187 = ~n6441 & n24186 ;
  assign n24191 = n24190 ^ n24187 ^ 1'b0 ;
  assign n24195 = n8305 & ~n10553 ;
  assign n24196 = n24195 ^ n5311 ^ 1'b0 ;
  assign n24197 = n5144 & ~n6750 ;
  assign n24198 = n24196 & n24197 ;
  assign n24192 = ~n10221 & n14356 ;
  assign n24193 = n5406 & n24192 ;
  assign n24194 = n16977 & ~n24193 ;
  assign n24199 = n24198 ^ n24194 ^ 1'b0 ;
  assign n24200 = n16652 ^ n5912 ^ 1'b0 ;
  assign n24201 = n24200 ^ n5936 ^ 1'b0 ;
  assign n24202 = n11279 ^ n4416 ^ 1'b0 ;
  assign n24203 = n24201 & ~n24202 ;
  assign n24204 = n2517 & n9011 ;
  assign n24205 = n3770 & n24204 ;
  assign n24206 = n327 & ~n19616 ;
  assign n24207 = n12292 ^ n8643 ^ 1'b0 ;
  assign n24208 = ( n19425 & n24206 ) | ( n19425 & ~n24207 ) | ( n24206 & ~n24207 ) ;
  assign n24209 = n9077 ^ n9004 ^ 1'b0 ;
  assign n24210 = n17427 & n24209 ;
  assign n24211 = n6063 ^ n1715 ^ x161 ;
  assign n24212 = n6445 ^ n1251 ^ 1'b0 ;
  assign n24213 = n24211 & ~n24212 ;
  assign n24214 = n11457 ^ n10129 ^ 1'b0 ;
  assign n24215 = n17293 ^ n941 ^ 1'b0 ;
  assign n24216 = n24214 & n24215 ;
  assign n24217 = n22778 & n24216 ;
  assign n24218 = ~n24213 & n24217 ;
  assign n24219 = ( ~n4245 & n24210 ) | ( ~n4245 & n24218 ) | ( n24210 & n24218 ) ;
  assign n24220 = n3585 & ~n12771 ;
  assign n24221 = ~n9532 & n11342 ;
  assign n24222 = n24221 ^ n3081 ^ n1164 ;
  assign n24223 = n4402 ^ n1517 ^ n936 ;
  assign n24224 = n24223 ^ n6981 ^ n3123 ;
  assign n24225 = n15162 ^ n10512 ^ 1'b0 ;
  assign n24226 = n20138 & n24225 ;
  assign n24227 = ~n12206 & n24226 ;
  assign n24228 = n24227 ^ x48 ^ 1'b0 ;
  assign n24229 = n13213 ^ n12445 ^ 1'b0 ;
  assign n24230 = n2077 | n24229 ;
  assign n24231 = n24230 ^ n9562 ^ n8475 ;
  assign n24232 = ( n1611 & n5996 ) | ( n1611 & ~n18443 ) | ( n5996 & ~n18443 ) ;
  assign n24233 = n24231 & ~n24232 ;
  assign n24234 = ~n1432 & n24233 ;
  assign n24235 = ( n3693 & ~n11668 ) | ( n3693 & n20755 ) | ( ~n11668 & n20755 ) ;
  assign n24236 = n9711 & ~n16062 ;
  assign n24237 = ~n1739 & n24236 ;
  assign n24238 = n9836 ^ n5867 ^ 1'b0 ;
  assign n24239 = n24237 | n24238 ;
  assign n24240 = ( n11392 & ~n20200 ) | ( n11392 & n24239 ) | ( ~n20200 & n24239 ) ;
  assign n24241 = n2903 & ~n19994 ;
  assign n24242 = n15486 ^ n5704 ^ 1'b0 ;
  assign n24243 = n24241 & ~n24242 ;
  assign n24244 = n8942 & n24243 ;
  assign n24245 = n24244 ^ n1865 ^ 1'b0 ;
  assign n24246 = n4085 | n8012 ;
  assign n24247 = n4471 ^ n1200 ^ 1'b0 ;
  assign n24248 = n9503 & ~n24247 ;
  assign n24249 = ~n10704 & n12936 ;
  assign n24250 = n24249 ^ n24188 ^ 1'b0 ;
  assign n24251 = n24250 ^ n12970 ^ n3479 ;
  assign n24252 = ( n16566 & n24248 ) | ( n16566 & ~n24251 ) | ( n24248 & ~n24251 ) ;
  assign n24253 = n18735 & n22500 ;
  assign n24259 = n16750 ^ n1655 ^ 1'b0 ;
  assign n24255 = n9338 ^ n7327 ^ 1'b0 ;
  assign n24256 = n20982 & ~n24255 ;
  assign n24254 = n13744 & ~n17118 ;
  assign n24257 = n24256 ^ n24254 ^ 1'b0 ;
  assign n24258 = n12688 | n24257 ;
  assign n24260 = n24259 ^ n24258 ^ n19516 ;
  assign n24261 = ~n13976 & n19313 ;
  assign n24262 = n24261 ^ n4090 ^ n3204 ;
  assign n24263 = ( n1605 & ~n20642 ) | ( n1605 & n20701 ) | ( ~n20642 & n20701 ) ;
  assign n24264 = n6597 | n15142 ;
  assign n24265 = n24264 ^ n4993 ^ 1'b0 ;
  assign n24266 = n24265 ^ n9827 ^ 1'b0 ;
  assign n24267 = n22606 ^ n5758 ^ 1'b0 ;
  assign n24268 = n20256 & ~n24267 ;
  assign n24269 = n12572 ^ n5832 ^ 1'b0 ;
  assign n24270 = n20067 ^ n19353 ^ 1'b0 ;
  assign n24271 = n8502 & ~n13917 ;
  assign n24272 = n6619 | n23968 ;
  assign n24273 = ( n2260 & ~n6502 ) | ( n2260 & n24272 ) | ( ~n6502 & n24272 ) ;
  assign n24274 = n3085 & ~n24273 ;
  assign n24275 = n24274 ^ n4631 ^ 1'b0 ;
  assign n24276 = n24275 ^ n1055 ^ 1'b0 ;
  assign n24277 = n24271 & ~n24276 ;
  assign n24278 = n3166 | n8050 ;
  assign n24279 = n6998 & n7386 ;
  assign n24280 = n6350 & n24279 ;
  assign n24281 = n24280 ^ n22386 ^ n15379 ;
  assign n24282 = ( n9018 & n9351 ) | ( n9018 & n22651 ) | ( n9351 & n22651 ) ;
  assign n24283 = n19294 ^ n5745 ^ 1'b0 ;
  assign n24284 = n15210 ^ n3630 ^ 1'b0 ;
  assign n24285 = n19346 & ~n24284 ;
  assign n24286 = n24285 ^ n18984 ^ 1'b0 ;
  assign n24287 = ( n6283 & n17326 ) | ( n6283 & n17519 ) | ( n17326 & n17519 ) ;
  assign n24288 = n24287 ^ n11758 ^ n1156 ;
  assign n24289 = n17073 ^ n8218 ^ 1'b0 ;
  assign n24290 = n12473 | n24289 ;
  assign n24292 = ~n3573 & n9886 ;
  assign n24293 = n24292 ^ n12294 ^ 1'b0 ;
  assign n24291 = n12752 & n16824 ;
  assign n24294 = n24293 ^ n24291 ^ n9952 ;
  assign n24295 = ( n5377 & ~n22822 ) | ( n5377 & n24038 ) | ( ~n22822 & n24038 ) ;
  assign n24296 = x162 | n21319 ;
  assign n24297 = n19114 ^ x182 ^ 1'b0 ;
  assign n24298 = n12672 | n24297 ;
  assign n24299 = n19230 ^ n16250 ^ 1'b0 ;
  assign n24300 = n3073 ^ x67 ^ 1'b0 ;
  assign n24301 = n9102 & n24300 ;
  assign n24302 = n24301 ^ n21420 ^ n1007 ;
  assign n24303 = n9553 ^ n5649 ^ 1'b0 ;
  assign n24304 = ~n8103 & n24303 ;
  assign n24305 = n5289 & n7513 ;
  assign n24306 = n7857 & ~n24305 ;
  assign n24307 = ~n14595 & n24306 ;
  assign n24308 = ( n8891 & n20097 ) | ( n8891 & n24307 ) | ( n20097 & n24307 ) ;
  assign n24309 = n19353 ^ n1504 ^ 1'b0 ;
  assign n24310 = ( ~n2314 & n17817 ) | ( ~n2314 & n24309 ) | ( n17817 & n24309 ) ;
  assign n24311 = n4198 & ~n24310 ;
  assign n24312 = n21228 ^ n11167 ^ 1'b0 ;
  assign n24313 = n10250 & ~n24312 ;
  assign n24314 = n22061 ^ n12684 ^ n4824 ;
  assign n24315 = n24314 ^ n5670 ^ 1'b0 ;
  assign n24316 = n9899 | n24315 ;
  assign n24317 = n7963 & n9983 ;
  assign n24318 = ~n838 & n24317 ;
  assign n24322 = n11148 ^ n10550 ^ 1'b0 ;
  assign n24323 = n9102 & ~n24322 ;
  assign n24324 = n11907 & n24323 ;
  assign n24321 = n6889 | n13857 ;
  assign n24319 = ( n4367 & ~n5485 ) | ( n4367 & n11028 ) | ( ~n5485 & n11028 ) ;
  assign n24320 = n9514 | n24319 ;
  assign n24325 = n24324 ^ n24321 ^ n24320 ;
  assign n24326 = n22451 & ~n24325 ;
  assign n24327 = n24326 ^ n8316 ^ 1'b0 ;
  assign n24328 = n16439 ^ n2401 ^ 1'b0 ;
  assign n24329 = x72 & n24328 ;
  assign n24330 = n16700 ^ n11434 ^ 1'b0 ;
  assign n24331 = n21944 & n22017 ;
  assign n24334 = n4407 ^ n1975 ^ n785 ;
  assign n24335 = ( ~n425 & n2262 ) | ( ~n425 & n24334 ) | ( n2262 & n24334 ) ;
  assign n24332 = n11302 | n21860 ;
  assign n24333 = n24332 ^ n4404 ^ 1'b0 ;
  assign n24336 = n24335 ^ n24333 ^ n12709 ;
  assign n24337 = n5795 ^ n3959 ^ 1'b0 ;
  assign n24338 = n11551 | n24337 ;
  assign n24339 = ( n482 & ~n13960 ) | ( n482 & n24338 ) | ( ~n13960 & n24338 ) ;
  assign n24340 = n8276 | n24339 ;
  assign n24341 = ~n13436 & n18768 ;
  assign n24342 = n24341 ^ n8144 ^ n7173 ;
  assign n24345 = ( n1470 & n3953 ) | ( n1470 & n23617 ) | ( n3953 & n23617 ) ;
  assign n24346 = n24345 ^ n1604 ^ 1'b0 ;
  assign n24347 = n5298 | n24346 ;
  assign n24343 = n4720 & n12733 ;
  assign n24344 = ( n8058 & n18718 ) | ( n8058 & n24343 ) | ( n18718 & n24343 ) ;
  assign n24348 = n24347 ^ n24344 ^ n20556 ;
  assign n24349 = n24230 ^ n19426 ^ 1'b0 ;
  assign n24350 = ~n16917 & n24349 ;
  assign n24351 = n4136 ^ n1557 ^ 1'b0 ;
  assign n24352 = n20772 ^ n1835 ^ 1'b0 ;
  assign n24353 = n24351 | n24352 ;
  assign n24354 = ~n3296 & n18936 ;
  assign n24355 = n3155 & ~n24354 ;
  assign n24356 = n24355 ^ n16919 ^ 1'b0 ;
  assign n24357 = n378 | n8158 ;
  assign n24358 = ( n8497 & n24356 ) | ( n8497 & ~n24357 ) | ( n24356 & ~n24357 ) ;
  assign n24359 = n13967 & n24358 ;
  assign n24360 = n24359 ^ n1538 ^ 1'b0 ;
  assign n24361 = n16847 | n24360 ;
  assign n24362 = n9152 ^ n4329 ^ 1'b0 ;
  assign n24363 = n24362 ^ n17450 ^ n15371 ;
  assign n24364 = n24363 ^ n18010 ^ 1'b0 ;
  assign n24365 = n24364 ^ n23614 ^ n23203 ;
  assign n24366 = n1891 ^ n1800 ^ 1'b0 ;
  assign n24367 = n6540 | n24366 ;
  assign n24368 = ( n8821 & n16969 ) | ( n8821 & n24367 ) | ( n16969 & n24367 ) ;
  assign n24369 = n8129 ^ n1895 ^ 1'b0 ;
  assign n24370 = n6246 | n24369 ;
  assign n24371 = n24370 ^ n4755 ^ n3794 ;
  assign n24372 = ( n7179 & n24368 ) | ( n7179 & ~n24371 ) | ( n24368 & ~n24371 ) ;
  assign n24374 = n15982 ^ n10162 ^ n2718 ;
  assign n24373 = ( n14600 & ~n19433 ) | ( n14600 & n19701 ) | ( ~n19433 & n19701 ) ;
  assign n24375 = n24374 ^ n24373 ^ n13947 ;
  assign n24376 = ( ~n11227 & n17795 ) | ( ~n11227 & n24375 ) | ( n17795 & n24375 ) ;
  assign n24377 = n4193 | n14487 ;
  assign n24378 = n3639 | n24377 ;
  assign n24379 = n7051 & ~n8480 ;
  assign n24380 = n14946 & ~n24379 ;
  assign n24381 = ~n17271 & n24380 ;
  assign n24382 = ( n1302 & ~n9194 ) | ( n1302 & n23206 ) | ( ~n9194 & n23206 ) ;
  assign n24383 = ( n9551 & ~n13783 ) | ( n9551 & n17146 ) | ( ~n13783 & n17146 ) ;
  assign n24384 = n20442 & n24383 ;
  assign n24385 = ~n14093 & n24384 ;
  assign n24386 = n20269 ^ n16946 ^ n3437 ;
  assign n24387 = ~n6246 & n8287 ;
  assign n24388 = n18785 ^ n10757 ^ 1'b0 ;
  assign n24389 = n19672 & ~n24388 ;
  assign n24390 = n24389 ^ n16139 ^ 1'b0 ;
  assign n24391 = ~n24387 & n24390 ;
  assign n24392 = ~n24386 & n24391 ;
  assign n24393 = n13424 ^ n6596 ^ n540 ;
  assign n24394 = n5424 | n9187 ;
  assign n24395 = n4239 | n24394 ;
  assign n24396 = n876 & n6439 ;
  assign n24397 = ~n11757 & n24396 ;
  assign n24398 = n9364 | n24397 ;
  assign n24399 = n10258 & ~n24398 ;
  assign n24400 = n24399 ^ n8734 ^ 1'b0 ;
  assign n24401 = n11163 ^ n6205 ^ 1'b0 ;
  assign n24402 = n12808 & n24401 ;
  assign n24403 = n24402 ^ n887 ^ 1'b0 ;
  assign n24404 = ( n24395 & n24400 ) | ( n24395 & n24403 ) | ( n24400 & n24403 ) ;
  assign n24405 = n6668 | n23159 ;
  assign n24406 = ~n4693 & n6351 ;
  assign n24407 = n10427 & n24406 ;
  assign n24408 = n11963 ^ n8843 ^ 1'b0 ;
  assign n24409 = n11484 & n24408 ;
  assign n24410 = n4395 & ~n7266 ;
  assign n24411 = n13877 & ~n24410 ;
  assign n24412 = ~n1227 & n6174 ;
  assign n24413 = n12133 & n24412 ;
  assign n24414 = n1486 & n24413 ;
  assign n24415 = n22355 & ~n24414 ;
  assign n24416 = n24415 ^ n352 ^ 1'b0 ;
  assign n24417 = ( n6436 & ~n21765 ) | ( n6436 & n24416 ) | ( ~n21765 & n24416 ) ;
  assign n24418 = n17999 ^ n10067 ^ n3083 ;
  assign n24419 = ( n5918 & ~n6149 ) | ( n5918 & n8075 ) | ( ~n6149 & n8075 ) ;
  assign n24420 = ( x108 & n9037 ) | ( x108 & n21456 ) | ( n9037 & n21456 ) ;
  assign n24421 = n24420 ^ n8378 ^ 1'b0 ;
  assign n24422 = n24419 & n24421 ;
  assign n24423 = ( n18127 & n24418 ) | ( n18127 & n24422 ) | ( n24418 & n24422 ) ;
  assign n24424 = n15941 ^ n9193 ^ n7919 ;
  assign n24425 = ( ~n7819 & n7840 ) | ( ~n7819 & n24424 ) | ( n7840 & n24424 ) ;
  assign n24426 = n20045 ^ n10165 ^ 1'b0 ;
  assign n24427 = n9283 & n9525 ;
  assign n24429 = n24129 ^ n17737 ^ 1'b0 ;
  assign n24428 = n4441 & n14889 ;
  assign n24430 = n24429 ^ n24428 ^ 1'b0 ;
  assign n24431 = n12438 & ~n24430 ;
  assign n24432 = n16652 ^ n5948 ^ 1'b0 ;
  assign n24433 = n24432 ^ n21133 ^ n13350 ;
  assign n24434 = n11733 & n22681 ;
  assign n24437 = ( n5384 & n6362 ) | ( n5384 & ~n19864 ) | ( n6362 & ~n19864 ) ;
  assign n24438 = n7899 & n24437 ;
  assign n24435 = x235 & ~n7073 ;
  assign n24436 = ~x235 & n24435 ;
  assign n24439 = n24438 ^ n24436 ^ n256 ;
  assign n24440 = n13271 ^ n731 ^ 1'b0 ;
  assign n24441 = n22959 & ~n24440 ;
  assign n24442 = ( ~n3996 & n6268 ) | ( ~n3996 & n19821 ) | ( n6268 & n19821 ) ;
  assign n24443 = ~n24441 & n24442 ;
  assign n24444 = n24443 ^ n5223 ^ 1'b0 ;
  assign n24449 = n4190 | n4909 ;
  assign n24450 = n22131 | n24449 ;
  assign n24445 = n5078 | n18990 ;
  assign n24446 = ~n4441 & n24445 ;
  assign n24447 = ~n4735 & n24446 ;
  assign n24448 = n24447 ^ n15198 ^ n8332 ;
  assign n24451 = n24450 ^ n24448 ^ 1'b0 ;
  assign n24452 = n22799 & ~n24451 ;
  assign n24453 = n4849 ^ n2007 ^ 1'b0 ;
  assign n24454 = n14005 | n24453 ;
  assign n24455 = n24454 ^ n14131 ^ n968 ;
  assign n24456 = ( n12396 & ~n22291 ) | ( n12396 & n24455 ) | ( ~n22291 & n24455 ) ;
  assign n24457 = n24456 ^ n12506 ^ n3426 ;
  assign n24458 = ( n11761 & n20739 ) | ( n11761 & n23665 ) | ( n20739 & n23665 ) ;
  assign n24459 = ( n7885 & n8407 ) | ( n7885 & ~n18980 ) | ( n8407 & ~n18980 ) ;
  assign n24460 = ( n8835 & n13885 ) | ( n8835 & ~n24459 ) | ( n13885 & ~n24459 ) ;
  assign n24461 = ( n11765 & ~n17823 ) | ( n11765 & n24460 ) | ( ~n17823 & n24460 ) ;
  assign n24462 = n18770 ^ n14562 ^ 1'b0 ;
  assign n24463 = ~n20066 & n24462 ;
  assign n24464 = n24463 ^ n15567 ^ 1'b0 ;
  assign n24465 = n24464 ^ n22520 ^ n21926 ;
  assign n24466 = n22571 ^ n11444 ^ n4487 ;
  assign n24467 = n24466 ^ n1441 ^ 1'b0 ;
  assign n24468 = n9323 | n12172 ;
  assign n24469 = n24468 ^ n22092 ^ n13268 ;
  assign n24470 = ( n2824 & ~n6960 ) | ( n2824 & n16396 ) | ( ~n6960 & n16396 ) ;
  assign n24471 = ~n964 & n24470 ;
  assign n24472 = ~n3794 & n24471 ;
  assign n24476 = n5157 & ~n5513 ;
  assign n24477 = n11846 & n24476 ;
  assign n24478 = ~n17061 & n24477 ;
  assign n24473 = n17930 ^ n11380 ^ 1'b0 ;
  assign n24474 = ( n16725 & n18569 ) | ( n16725 & ~n21179 ) | ( n18569 & ~n21179 ) ;
  assign n24475 = n24473 & ~n24474 ;
  assign n24479 = n24478 ^ n24475 ^ 1'b0 ;
  assign n24480 = n7767 & n17352 ;
  assign n24481 = n15030 ^ n9268 ^ 1'b0 ;
  assign n24482 = n6907 & ~n24481 ;
  assign n24483 = n9041 ^ n6611 ^ 1'b0 ;
  assign n24484 = n21748 | n24483 ;
  assign n24485 = n5526 ^ n1007 ^ 1'b0 ;
  assign n24486 = n3746 & n24485 ;
  assign n24487 = ( n2459 & n2720 ) | ( n2459 & n6808 ) | ( n2720 & n6808 ) ;
  assign n24488 = n22633 ^ n1966 ^ 1'b0 ;
  assign n24489 = ~n4195 & n12629 ;
  assign n24490 = n24489 ^ n9784 ^ 1'b0 ;
  assign n24491 = n10535 | n24490 ;
  assign n24492 = n24491 ^ n13555 ^ 1'b0 ;
  assign n24493 = x28 & ~n7088 ;
  assign n24494 = n9631 & n24493 ;
  assign n24495 = n15507 & ~n24494 ;
  assign n24496 = n24495 ^ n23602 ^ 1'b0 ;
  assign n24497 = n8225 ^ n7277 ^ 1'b0 ;
  assign n24498 = n19065 ^ n15121 ^ 1'b0 ;
  assign n24499 = n24497 & n24498 ;
  assign n24502 = ( n1486 & n8116 ) | ( n1486 & n8999 ) | ( n8116 & n8999 ) ;
  assign n24500 = n13855 ^ n6979 ^ n2392 ;
  assign n24501 = n15588 & ~n24500 ;
  assign n24503 = n24502 ^ n24501 ^ 1'b0 ;
  assign n24504 = x246 & ~n24503 ;
  assign n24505 = n716 & ~n826 ;
  assign n24506 = n24505 ^ n10559 ^ 1'b0 ;
  assign n24507 = n19089 | n24506 ;
  assign n24508 = n14430 ^ n13084 ^ 1'b0 ;
  assign n24509 = ~n820 & n8571 ;
  assign n24510 = n22879 & n24509 ;
  assign n24511 = n6094 & n12186 ;
  assign n24512 = ~n4854 & n10034 ;
  assign n24513 = ~n892 & n6647 ;
  assign n24514 = n18348 ^ n3959 ^ 1'b0 ;
  assign n24515 = ~n16627 & n20509 ;
  assign n24516 = ~n9421 & n12419 ;
  assign n24519 = n4844 ^ x146 ^ 1'b0 ;
  assign n24517 = n9232 ^ n1734 ^ 1'b0 ;
  assign n24518 = n18982 | n24517 ;
  assign n24520 = n24519 ^ n24518 ^ n8672 ;
  assign n24522 = n7277 & n10532 ;
  assign n24523 = ( n4528 & n6221 ) | ( n4528 & ~n24522 ) | ( n6221 & ~n24522 ) ;
  assign n24521 = n23852 ^ n932 ^ 1'b0 ;
  assign n24524 = n24523 ^ n24521 ^ n20224 ;
  assign n24525 = n10131 | n17629 ;
  assign n24526 = n24525 ^ n23019 ^ 1'b0 ;
  assign n24527 = n6063 | n15892 ;
  assign n24528 = n24527 ^ n10859 ^ 1'b0 ;
  assign n24529 = n24528 ^ n4776 ^ 1'b0 ;
  assign n24530 = n15012 ^ n13170 ^ 1'b0 ;
  assign n24531 = n24530 ^ n308 ^ 1'b0 ;
  assign n24532 = n13865 | n24531 ;
  assign n24533 = n20410 ^ n15634 ^ n3030 ;
  assign n24534 = n23089 & n24533 ;
  assign n24535 = ~n24532 & n24534 ;
  assign n24536 = n24535 ^ n2671 ^ 1'b0 ;
  assign n24537 = n7989 ^ n895 ^ 1'b0 ;
  assign n24538 = n24537 ^ n9583 ^ n2924 ;
  assign n24554 = n3998 & ~n11048 ;
  assign n24555 = n24554 ^ n3617 ^ 1'b0 ;
  assign n24539 = ~n8771 & n12566 ;
  assign n24540 = n24539 ^ n3093 ^ 1'b0 ;
  assign n24541 = n5565 & ~n24540 ;
  assign n24542 = n24541 ^ n19409 ^ 1'b0 ;
  assign n24550 = ( n2463 & n3464 ) | ( n2463 & ~n15817 ) | ( n3464 & ~n15817 ) ;
  assign n24549 = ~n10117 & n18992 ;
  assign n24551 = n24550 ^ n24549 ^ 1'b0 ;
  assign n24543 = n9345 ^ n8409 ^ n5515 ;
  assign n24546 = n8419 ^ n3932 ^ 1'b0 ;
  assign n24544 = n12917 ^ n1241 ^ 1'b0 ;
  assign n24545 = n1499 & ~n24544 ;
  assign n24547 = n24546 ^ n24545 ^ 1'b0 ;
  assign n24548 = n24543 | n24547 ;
  assign n24552 = n24551 ^ n24548 ^ 1'b0 ;
  assign n24553 = n24542 | n24552 ;
  assign n24556 = n24555 ^ n24553 ^ 1'b0 ;
  assign n24557 = n5795 ^ n4033 ^ n1301 ;
  assign n24558 = n24557 ^ n24418 ^ n21187 ;
  assign n24559 = n17514 & ~n24558 ;
  assign n24560 = n24559 ^ n15924 ^ 1'b0 ;
  assign n24561 = n8340 & ~n24560 ;
  assign n24562 = n13107 | n18191 ;
  assign n24563 = n21179 & ~n24562 ;
  assign n24564 = n17608 & ~n24563 ;
  assign n24565 = n8377 & n17311 ;
  assign n24566 = n6662 ^ n1013 ^ 1'b0 ;
  assign n24567 = n5541 & ~n24566 ;
  assign n24568 = n2705 ^ n1155 ^ 1'b0 ;
  assign n24569 = n6682 & n24568 ;
  assign n24570 = n8316 & n24569 ;
  assign n24571 = n24570 ^ n1037 ^ 1'b0 ;
  assign n24577 = n22927 ^ n2942 ^ 1'b0 ;
  assign n24572 = n3978 ^ n1206 ^ 1'b0 ;
  assign n24573 = n3967 | n24572 ;
  assign n24574 = n5405 ^ n2904 ^ 1'b0 ;
  assign n24575 = n18876 | n24574 ;
  assign n24576 = n24573 | n24575 ;
  assign n24578 = n24577 ^ n24576 ^ 1'b0 ;
  assign n24579 = n10303 | n24578 ;
  assign n24580 = n6027 & ~n24579 ;
  assign n24581 = n9864 & n10923 ;
  assign n24582 = n4720 & n24581 ;
  assign n24583 = n1206 & ~n11380 ;
  assign n24584 = n24582 & n24583 ;
  assign n24585 = n1312 & n19491 ;
  assign n24586 = n11630 & ~n24585 ;
  assign n24587 = n24584 & n24586 ;
  assign n24588 = ( ~n2993 & n3745 ) | ( ~n2993 & n24587 ) | ( n3745 & n24587 ) ;
  assign n24589 = n18045 | n24588 ;
  assign n24590 = n3231 & ~n24589 ;
  assign n24591 = n1166 & n15309 ;
  assign n24592 = ~n10562 & n24591 ;
  assign n24593 = n16157 ^ n13029 ^ 1'b0 ;
  assign n24594 = n18820 ^ n16817 ^ 1'b0 ;
  assign n24595 = n6972 ^ n4618 ^ 1'b0 ;
  assign n24596 = n15382 & ~n24595 ;
  assign n24597 = n15054 & n17787 ;
  assign n24598 = n5323 | n24597 ;
  assign n24599 = n12632 | n24598 ;
  assign n24600 = n24599 ^ n10053 ^ 1'b0 ;
  assign n24601 = n24232 | n24600 ;
  assign n24606 = n16365 ^ n12127 ^ n11587 ;
  assign n24607 = n24606 ^ n14847 ^ 1'b0 ;
  assign n24602 = n18208 ^ n2240 ^ 1'b0 ;
  assign n24603 = n2674 | n24602 ;
  assign n24604 = x50 & ~n24603 ;
  assign n24605 = ~n18176 & n24604 ;
  assign n24608 = n24607 ^ n24605 ^ n14433 ;
  assign n24609 = n21919 ^ n21433 ^ n12506 ;
  assign n24610 = n1597 ^ n702 ^ 1'b0 ;
  assign n24611 = ~n1222 & n24610 ;
  assign n24612 = ~n14374 & n24611 ;
  assign n24613 = n24612 ^ n8085 ^ 1'b0 ;
  assign n24614 = n9709 | n13303 ;
  assign n24615 = n24613 | n24614 ;
  assign n24616 = n24615 ^ n6664 ^ 1'b0 ;
  assign n24617 = ~n8188 & n17134 ;
  assign n24619 = n13407 ^ n9282 ^ n3305 ;
  assign n24618 = n1538 | n6434 ;
  assign n24620 = n24619 ^ n24618 ^ 1'b0 ;
  assign n24621 = n6896 & n8009 ;
  assign n24622 = n24621 ^ n18602 ^ 1'b0 ;
  assign n24623 = ~n9820 & n17535 ;
  assign n24624 = n24623 ^ n12099 ^ 1'b0 ;
  assign n24625 = n1300 & ~n24624 ;
  assign n24626 = n24622 & n24625 ;
  assign n24627 = n7554 & ~n18528 ;
  assign n24628 = ~n3322 & n4316 ;
  assign n24629 = n13792 & n14333 ;
  assign n24630 = n24629 ^ n17338 ^ n1497 ;
  assign n24631 = n24630 ^ n1217 ^ 1'b0 ;
  assign n24632 = n17517 ^ n535 ^ x75 ;
  assign n24633 = n17042 ^ n16878 ^ n16394 ;
  assign n24634 = ( ~n8488 & n9311 ) | ( ~n8488 & n15904 ) | ( n9311 & n15904 ) ;
  assign n24635 = ~n14327 & n24634 ;
  assign n24636 = ~n4356 & n24635 ;
  assign n24643 = ~n10453 & n13448 ;
  assign n24639 = ~n4045 & n8610 ;
  assign n24640 = n15068 | n24639 ;
  assign n24641 = n24420 | n24640 ;
  assign n24642 = n24641 ^ n15840 ^ 1'b0 ;
  assign n24637 = n18556 ^ n3694 ^ 1'b0 ;
  assign n24638 = n15157 & n24637 ;
  assign n24644 = n24643 ^ n24642 ^ n24638 ;
  assign n24645 = n5931 & n14543 ;
  assign n24646 = n24645 ^ n11011 ^ 1'b0 ;
  assign n24647 = ~x3 & n1680 ;
  assign n24648 = ( n1871 & ~n18528 ) | ( n1871 & n24647 ) | ( ~n18528 & n24647 ) ;
  assign n24649 = ~n5261 & n12296 ;
  assign n24650 = ( ~n1115 & n17371 ) | ( ~n1115 & n22004 ) | ( n17371 & n22004 ) ;
  assign n24651 = n4879 | n5230 ;
  assign n24652 = n7141 & ~n24651 ;
  assign n24653 = n3546 & n24652 ;
  assign n24654 = n15147 & n21385 ;
  assign n24655 = ~n21385 & n24654 ;
  assign n24656 = n21105 ^ n588 ^ 1'b0 ;
  assign n24657 = n18308 | n24656 ;
  assign n24658 = n11779 | n24657 ;
  assign n24659 = n16738 & ~n21780 ;
  assign n24660 = n24659 ^ n23021 ^ 1'b0 ;
  assign n24661 = n1412 & ~n3878 ;
  assign n24662 = ~n1040 & n24661 ;
  assign n24663 = ( ~n9117 & n10223 ) | ( ~n9117 & n24662 ) | ( n10223 & n24662 ) ;
  assign n24664 = ( n1687 & n16507 ) | ( n1687 & n24663 ) | ( n16507 & n24663 ) ;
  assign n24665 = n22619 ^ n3044 ^ 1'b0 ;
  assign n24666 = n2903 & n24665 ;
  assign n24667 = n16668 | n24666 ;
  assign n24668 = n15516 ^ n5797 ^ n3494 ;
  assign n24669 = n18134 ^ n14056 ^ 1'b0 ;
  assign n24670 = n4122 & ~n24669 ;
  assign n24671 = n24668 & n24670 ;
  assign n24672 = n21571 ^ n13895 ^ n10446 ;
  assign n24673 = n24672 ^ n15329 ^ n10056 ;
  assign n24674 = n7394 | n20221 ;
  assign n24675 = n12913 | n22728 ;
  assign n24676 = n24675 ^ n6847 ^ 1'b0 ;
  assign n24677 = n1217 ^ n1019 ^ 1'b0 ;
  assign n24678 = n12081 | n24677 ;
  assign n24679 = n22029 ^ n11273 ^ 1'b0 ;
  assign n24680 = ( n7035 & n24678 ) | ( n7035 & n24679 ) | ( n24678 & n24679 ) ;
  assign n24681 = n5923 & ~n16373 ;
  assign n24682 = n5185 & n24681 ;
  assign n24683 = n20674 & n24682 ;
  assign n24684 = ~n426 & n1928 ;
  assign n24685 = n15203 & n24684 ;
  assign n24686 = n21705 & n22361 ;
  assign n24687 = n24685 & n24686 ;
  assign n24688 = n18923 ^ n711 ^ 1'b0 ;
  assign n24689 = n9194 & ~n24688 ;
  assign n24690 = ~n694 & n16183 ;
  assign n24691 = n24690 ^ n2356 ^ 1'b0 ;
  assign n24692 = n24691 ^ n20693 ^ 1'b0 ;
  assign n24693 = n9924 & ~n24692 ;
  assign n24695 = n11289 | n18366 ;
  assign n24696 = n5961 | n24695 ;
  assign n24694 = n5389 | n21194 ;
  assign n24697 = n24696 ^ n24694 ^ n3170 ;
  assign n24698 = ~n922 & n8468 ;
  assign n24699 = n3375 & n24698 ;
  assign n24700 = n6814 & n24699 ;
  assign n24701 = n19065 ^ n7552 ^ 1'b0 ;
  assign n24702 = ~n24700 & n24701 ;
  assign n24703 = n24702 ^ n23405 ^ 1'b0 ;
  assign n24704 = ~n11211 & n16337 ;
  assign n24705 = n24704 ^ n5867 ^ 1'b0 ;
  assign n24711 = n11046 ^ n4199 ^ 1'b0 ;
  assign n24707 = ~n5052 & n19076 ;
  assign n24706 = n15361 ^ n11668 ^ n10760 ;
  assign n24708 = n24707 ^ n24706 ^ 1'b0 ;
  assign n24709 = n5425 & n24708 ;
  assign n24710 = ~n18639 & n24709 ;
  assign n24712 = n24711 ^ n24710 ^ 1'b0 ;
  assign n24713 = n12169 & ~n14446 ;
  assign n24714 = n11445 ^ n5878 ^ 1'b0 ;
  assign n24715 = n20893 ^ n13499 ^ 1'b0 ;
  assign n24716 = n5920 & n24715 ;
  assign n24717 = n15539 ^ n989 ^ 1'b0 ;
  assign n24718 = n6086 ^ x36 ^ 1'b0 ;
  assign n24719 = ~n6256 & n24718 ;
  assign n24720 = ~n14439 & n24719 ;
  assign n24721 = ( n10936 & n15557 ) | ( n10936 & ~n21689 ) | ( n15557 & ~n21689 ) ;
  assign n24722 = ~n4516 & n10814 ;
  assign n24723 = n24722 ^ n6422 ^ 1'b0 ;
  assign n24724 = n24723 ^ n19236 ^ n11762 ;
  assign n24725 = n23946 ^ n17168 ^ 1'b0 ;
  assign n24726 = n14216 & n24725 ;
  assign n24727 = n21010 ^ n16564 ^ n6410 ;
  assign n24728 = n7116 & ~n21122 ;
  assign n24729 = n16242 ^ n12015 ^ n1562 ;
  assign n24730 = n7200 ^ n4883 ^ 1'b0 ;
  assign n24731 = n8780 & n24730 ;
  assign n24732 = n21970 ^ n17169 ^ 1'b0 ;
  assign n24733 = ~n11782 & n24732 ;
  assign n24734 = n5920 ^ n2879 ^ 1'b0 ;
  assign n24735 = n14722 | n24734 ;
  assign n24736 = n3425 ^ n3296 ^ 1'b0 ;
  assign n24737 = n9336 & n20215 ;
  assign n24738 = n24736 & n24737 ;
  assign n24739 = n8654 ^ n1493 ^ 1'b0 ;
  assign n24740 = n24738 | n24739 ;
  assign n24742 = ( n1930 & ~n7881 ) | ( n1930 & n9134 ) | ( ~n7881 & n9134 ) ;
  assign n24741 = n3312 & ~n23054 ;
  assign n24743 = n24742 ^ n24741 ^ n21691 ;
  assign n24744 = n20601 ^ n7950 ^ 1'b0 ;
  assign n24745 = n13262 ^ n9184 ^ n599 ;
  assign n24746 = n24745 ^ n9068 ^ n8180 ;
  assign n24747 = n9772 & ~n9941 ;
  assign n24748 = n7124 | n24747 ;
  assign n24749 = n7669 & ~n24748 ;
  assign n24750 = ~n8277 & n24749 ;
  assign n24751 = n15291 ^ n7762 ^ 1'b0 ;
  assign n24752 = n24750 | n24751 ;
  assign n24753 = n13202 & n16695 ;
  assign n24754 = ( ~n6893 & n7522 ) | ( ~n6893 & n15191 ) | ( n7522 & n15191 ) ;
  assign n24755 = ~n3770 & n24754 ;
  assign n24756 = n24755 ^ n4114 ^ 1'b0 ;
  assign n24757 = ( n9493 & n24753 ) | ( n9493 & n24756 ) | ( n24753 & n24756 ) ;
  assign n24758 = n12592 ^ n8946 ^ 1'b0 ;
  assign n24759 = ~n13872 & n24758 ;
  assign n24760 = n24759 ^ n12771 ^ n3045 ;
  assign n24761 = n12042 ^ n9037 ^ 1'b0 ;
  assign n24762 = n17656 & n24761 ;
  assign n24763 = n24762 ^ n5572 ^ 1'b0 ;
  assign n24764 = ~n6516 & n14946 ;
  assign n24765 = n14754 | n24764 ;
  assign n24766 = ~n374 & n7859 ;
  assign n24769 = ~n5816 & n11163 ;
  assign n24767 = ( n14023 & ~n22946 ) | ( n14023 & n24070 ) | ( ~n22946 & n24070 ) ;
  assign n24768 = n8418 & n24767 ;
  assign n24770 = n24769 ^ n24768 ^ n15717 ;
  assign n24771 = n14215 | n24770 ;
  assign n24772 = n8665 & n10723 ;
  assign n24773 = n24772 ^ n4661 ^ 1'b0 ;
  assign n24774 = n7076 ^ n2534 ^ 1'b0 ;
  assign n24775 = n2837 & n19428 ;
  assign n24776 = n2523 & n24775 ;
  assign n24777 = ~n5927 & n15817 ;
  assign n24778 = n24777 ^ n19031 ^ 1'b0 ;
  assign n24779 = n24778 ^ n9857 ^ 1'b0 ;
  assign n24780 = n24779 ^ n18577 ^ n15136 ;
  assign n24781 = ~n15306 & n24780 ;
  assign n24782 = ( n2586 & ~n10153 ) | ( n2586 & n20448 ) | ( ~n10153 & n20448 ) ;
  assign n24783 = n24239 ^ n18915 ^ 1'b0 ;
  assign n24784 = n24782 & ~n24783 ;
  assign n24785 = ~n10095 & n24784 ;
  assign n24786 = n20786 & n24785 ;
  assign n24787 = n14157 ^ n10632 ^ n10005 ;
  assign n24788 = n22425 ^ n6398 ^ 1'b0 ;
  assign n24789 = n5475 & n24788 ;
  assign n24790 = n22542 ^ n18386 ^ n2140 ;
  assign n24791 = n19213 | n24790 ;
  assign n24792 = n24789 | n24791 ;
  assign n24793 = ( ~n15026 & n24787 ) | ( ~n15026 & n24792 ) | ( n24787 & n24792 ) ;
  assign n24794 = n9196 ^ n5242 ^ 1'b0 ;
  assign n24795 = n24793 & ~n24794 ;
  assign n24796 = n5873 ^ n485 ^ 1'b0 ;
  assign n24797 = n1197 | n24796 ;
  assign n24798 = n24797 ^ n16469 ^ 1'b0 ;
  assign n24799 = n24798 ^ n19049 ^ n11791 ;
  assign n24800 = n20688 ^ n949 ^ 1'b0 ;
  assign n24801 = ~n18305 & n24800 ;
  assign n24802 = n13913 ^ n8465 ^ 1'b0 ;
  assign n24803 = n4667 & ~n24802 ;
  assign n24804 = n23823 ^ n7400 ^ 1'b0 ;
  assign n24807 = n17250 ^ n11147 ^ 1'b0 ;
  assign n24808 = n4022 | n24807 ;
  assign n24805 = n24558 ^ n11137 ^ 1'b0 ;
  assign n24806 = ~n11194 & n24805 ;
  assign n24809 = n24808 ^ n24806 ^ n5190 ;
  assign n24810 = ( n10577 & n20708 ) | ( n10577 & ~n23449 ) | ( n20708 & ~n23449 ) ;
  assign n24811 = n7063 ^ n3633 ^ n661 ;
  assign n24812 = n3464 & n14819 ;
  assign n24813 = ~x166 & n24812 ;
  assign n24814 = n24813 ^ n7802 ^ 1'b0 ;
  assign n24815 = n5718 & ~n24814 ;
  assign n24816 = x20 & ~n9340 ;
  assign n24817 = ~n13040 & n24816 ;
  assign n24818 = n24817 ^ n20120 ^ 1'b0 ;
  assign n24819 = n8806 | n24818 ;
  assign n24820 = n24815 & n24819 ;
  assign n24821 = n4016 ^ n1353 ^ 1'b0 ;
  assign n24822 = n9908 ^ n2812 ^ 1'b0 ;
  assign n24823 = n23966 ^ n16617 ^ 1'b0 ;
  assign n24824 = n17881 | n24823 ;
  assign n24825 = ( n13640 & n24822 ) | ( n13640 & ~n24824 ) | ( n24822 & ~n24824 ) ;
  assign n24826 = n9351 ^ n8137 ^ 1'b0 ;
  assign n24827 = n1979 & ~n24826 ;
  assign n24828 = n17647 ^ n8760 ^ n8742 ;
  assign n24829 = ~n2179 & n24828 ;
  assign n24830 = n1228 & n24829 ;
  assign n24831 = n16846 ^ n15506 ^ 1'b0 ;
  assign n24832 = x158 & n24831 ;
  assign n24833 = ~n11288 & n21926 ;
  assign n24834 = n24833 ^ n5428 ^ 1'b0 ;
  assign n24835 = n24834 ^ n19879 ^ 1'b0 ;
  assign n24836 = n9521 | n24835 ;
  assign n24837 = ( n4868 & n6430 ) | ( n4868 & n9944 ) | ( n6430 & n9944 ) ;
  assign n24838 = n4585 | n8739 ;
  assign n24839 = n24838 ^ n4952 ^ 1'b0 ;
  assign n24840 = n24839 ^ n20870 ^ n11576 ;
  assign n24841 = n24837 | n24840 ;
  assign n24842 = n24841 ^ n7794 ^ 1'b0 ;
  assign n24843 = n20347 ^ n11714 ^ 1'b0 ;
  assign n24844 = n24843 ^ n2779 ^ 1'b0 ;
  assign n24845 = n19190 ^ n10982 ^ n4441 ;
  assign n24846 = ( n10236 & n17678 ) | ( n10236 & n24845 ) | ( n17678 & n24845 ) ;
  assign n24847 = n9832 & n24846 ;
  assign n24848 = ( ~n6351 & n18362 ) | ( ~n6351 & n21759 ) | ( n18362 & n21759 ) ;
  assign n24849 = ( n1237 & ~n11299 ) | ( n1237 & n24848 ) | ( ~n11299 & n24848 ) ;
  assign n24850 = n24849 ^ n18612 ^ 1'b0 ;
  assign n24851 = n3470 & ~n24850 ;
  assign n24852 = ~n5167 & n18818 ;
  assign n24853 = n22199 ^ n8357 ^ 1'b0 ;
  assign n24854 = n24746 & ~n24853 ;
  assign n24855 = n11447 ^ n6710 ^ n3967 ;
  assign n24856 = n24855 ^ n19315 ^ 1'b0 ;
  assign n24857 = n20115 ^ n10690 ^ 1'b0 ;
  assign n24858 = n7825 & n24857 ;
  assign n24859 = n24858 ^ n15731 ^ 1'b0 ;
  assign n24860 = n23699 ^ n22633 ^ n12933 ;
  assign n24861 = n7005 | n10346 ;
  assign n24862 = n24861 ^ n8143 ^ 1'b0 ;
  assign n24863 = ~n7769 & n24862 ;
  assign n24864 = ~n24860 & n24863 ;
  assign n24865 = n24864 ^ n17415 ^ 1'b0 ;
  assign n24866 = n4090 ^ n2729 ^ 1'b0 ;
  assign n24867 = ~n3054 & n24866 ;
  assign n24868 = n8794 ^ n7927 ^ 1'b0 ;
  assign n24869 = n24868 ^ n19063 ^ n1847 ;
  assign n24870 = ( ~n2194 & n9173 ) | ( ~n2194 & n10660 ) | ( n9173 & n10660 ) ;
  assign n24871 = n2307 & ~n18104 ;
  assign n24872 = ~n4992 & n9710 ;
  assign n24873 = n2937 & ~n4635 ;
  assign n24874 = n8598 & n9156 ;
  assign n24875 = n1561 ^ n1175 ^ 1'b0 ;
  assign n24876 = n1705 & n2688 ;
  assign n24877 = n24876 ^ n4029 ^ 1'b0 ;
  assign n24878 = ~n3607 & n12497 ;
  assign n24879 = n24878 ^ n3203 ^ 1'b0 ;
  assign n24880 = n24877 & n24879 ;
  assign n24881 = ~n6992 & n24880 ;
  assign n24882 = ( ~n24874 & n24875 ) | ( ~n24874 & n24881 ) | ( n24875 & n24881 ) ;
  assign n24883 = n1150 & n3469 ;
  assign n24884 = n24883 ^ n18967 ^ 1'b0 ;
  assign n24885 = ~n8660 & n24884 ;
  assign n24887 = x252 & ~n6650 ;
  assign n24888 = n24887 ^ n18074 ^ 1'b0 ;
  assign n24886 = ~n21466 & n24723 ;
  assign n24889 = n24888 ^ n24886 ^ 1'b0 ;
  assign n24890 = ( n829 & n9564 ) | ( n829 & n12814 ) | ( n9564 & n12814 ) ;
  assign n24891 = n24890 ^ n23703 ^ n7643 ;
  assign n24892 = n24891 ^ n3756 ^ 1'b0 ;
  assign n24893 = n22681 | n24892 ;
  assign n24894 = ( n9311 & ~n12351 ) | ( n9311 & n15981 ) | ( ~n12351 & n15981 ) ;
  assign n24895 = n13977 ^ n10923 ^ 1'b0 ;
  assign n24896 = ~n10016 & n24895 ;
  assign n24897 = n14980 & ~n24896 ;
  assign n24898 = n24897 ^ n5158 ^ 1'b0 ;
  assign n24899 = n18547 & ~n24898 ;
  assign n24900 = n9048 & ~n23136 ;
  assign n24901 = n4185 & n24900 ;
  assign n24902 = ( n1847 & n5768 ) | ( n1847 & ~n6654 ) | ( n5768 & ~n6654 ) ;
  assign n24903 = n24902 ^ n1690 ^ 1'b0 ;
  assign n24904 = n8116 & ~n24903 ;
  assign n24905 = n24904 ^ n12860 ^ 1'b0 ;
  assign n24906 = x129 | n5776 ;
  assign n24907 = n1032 | n6732 ;
  assign n24908 = n13873 ^ n3383 ^ 1'b0 ;
  assign n24909 = n4004 & n24908 ;
  assign n24912 = n973 | n7026 ;
  assign n24913 = n24912 ^ n18798 ^ 1'b0 ;
  assign n24910 = n4107 ^ n3677 ^ 1'b0 ;
  assign n24911 = n1083 & n24910 ;
  assign n24914 = n24913 ^ n24911 ^ n19191 ;
  assign n24915 = n15678 ^ n10942 ^ n1644 ;
  assign n24916 = n24915 ^ n7801 ^ 1'b0 ;
  assign n24917 = ( n21055 & n24914 ) | ( n21055 & ~n24916 ) | ( n24914 & ~n24916 ) ;
  assign n24918 = n11624 ^ n3731 ^ 1'b0 ;
  assign n24919 = n7395 ^ x103 ^ 1'b0 ;
  assign n24920 = n10096 ^ n5011 ^ 1'b0 ;
  assign n24921 = n24919 & n24920 ;
  assign n24923 = n1733 | n15073 ;
  assign n24924 = n1084 | n24923 ;
  assign n24922 = ~n17106 & n21800 ;
  assign n24925 = n24924 ^ n24922 ^ 1'b0 ;
  assign n24926 = n19446 ^ n13553 ^ 1'b0 ;
  assign n24927 = n24533 ^ n11765 ^ 1'b0 ;
  assign n24928 = ~n4963 & n7720 ;
  assign n24929 = n17053 & ~n24928 ;
  assign n24930 = n24929 ^ n10042 ^ 1'b0 ;
  assign n24931 = n22469 ^ n21477 ^ n10471 ;
  assign n24932 = n9941 ^ n1265 ^ 1'b0 ;
  assign n24933 = n6310 | n24932 ;
  assign n24934 = n24931 | n24933 ;
  assign n24935 = ~n5255 & n8339 ;
  assign n24936 = x90 & n24935 ;
  assign n24937 = ~n4280 & n10310 ;
  assign n24938 = n24937 ^ n9525 ^ 1'b0 ;
  assign n24939 = n24938 ^ n22836 ^ n14441 ;
  assign n24940 = n9972 & ~n22079 ;
  assign n24941 = n24393 & n24940 ;
  assign n24942 = n24941 ^ n3972 ^ 1'b0 ;
  assign n24943 = n12926 ^ n2411 ^ 1'b0 ;
  assign n24944 = ~n6280 & n12677 ;
  assign n24945 = n19762 & n24944 ;
  assign n24946 = ~n5177 & n11062 ;
  assign n24947 = n24946 ^ n8433 ^ 1'b0 ;
  assign n24948 = ( n17158 & ~n24860 ) | ( n17158 & n24947 ) | ( ~n24860 & n24947 ) ;
  assign n24949 = n20660 ^ n16148 ^ n9892 ;
  assign n24950 = n24949 ^ n7325 ^ n5376 ;
  assign n24951 = n24950 ^ n6063 ^ 1'b0 ;
  assign n24952 = n17188 ^ n13369 ^ 1'b0 ;
  assign n24953 = n3750 & ~n24952 ;
  assign n24954 = n24953 ^ n5047 ^ n3907 ;
  assign n24955 = n24954 ^ n9903 ^ 1'b0 ;
  assign n24956 = n10408 & n24955 ;
  assign n24957 = n24956 ^ n9933 ^ 1'b0 ;
  assign n24958 = n11875 | n18503 ;
  assign n24959 = n24958 ^ n15793 ^ 1'b0 ;
  assign n24960 = n3467 & ~n3645 ;
  assign n24961 = n13085 & n24960 ;
  assign n24962 = n24959 | n24961 ;
  assign n24963 = n22715 ^ n13968 ^ 1'b0 ;
  assign n24964 = ~n16402 & n24963 ;
  assign n24965 = n20731 ^ n7741 ^ n797 ;
  assign n24966 = n15035 ^ n5050 ^ 1'b0 ;
  assign n24967 = n9612 & ~n15101 ;
  assign n24968 = n24967 ^ n13675 ^ 1'b0 ;
  assign n24969 = n13643 | n24968 ;
  assign n24970 = n4097 | n24969 ;
  assign n24971 = n840 | n12080 ;
  assign n24972 = n24971 ^ n18204 ^ 1'b0 ;
  assign n24973 = n13046 | n21760 ;
  assign n24974 = n1178 & ~n2425 ;
  assign n24975 = n24974 ^ n1258 ^ 1'b0 ;
  assign n24976 = n16842 ^ n13172 ^ 1'b0 ;
  assign n24977 = n5855 & ~n24976 ;
  assign n24978 = n24977 ^ n8934 ^ 1'b0 ;
  assign n24979 = ( n19674 & n24975 ) | ( n19674 & ~n24978 ) | ( n24975 & ~n24978 ) ;
  assign n24980 = n6087 ^ n5437 ^ 1'b0 ;
  assign n24981 = n6364 | n24980 ;
  assign n24982 = n24981 ^ n17930 ^ 1'b0 ;
  assign n24983 = n3985 | n24982 ;
  assign n24984 = n11039 | n24983 ;
  assign n24985 = n11988 ^ n2386 ^ 1'b0 ;
  assign n24986 = n24984 & ~n24985 ;
  assign n24987 = n5334 & n24986 ;
  assign n24988 = n23884 ^ n9776 ^ n9714 ;
  assign n24989 = ~n18432 & n20438 ;
  assign n24990 = n19874 & n24989 ;
  assign n24991 = n9530 ^ n8204 ^ n4114 ;
  assign n24992 = ( n13785 & ~n17390 ) | ( n13785 & n24991 ) | ( ~n17390 & n24991 ) ;
  assign n24993 = n17375 ^ n14818 ^ n1651 ;
  assign n24994 = ~n3563 & n18525 ;
  assign n24995 = n7218 ^ n3107 ^ 1'b0 ;
  assign n24996 = n7835 & n24995 ;
  assign n24997 = x47 & n18182 ;
  assign n24998 = n24997 ^ n537 ^ 1'b0 ;
  assign n24999 = x197 & n3192 ;
  assign n25000 = n24998 & n24999 ;
  assign n25001 = ( ~n17094 & n24996 ) | ( ~n17094 & n25000 ) | ( n24996 & n25000 ) ;
  assign n25002 = n7145 ^ n2461 ^ 1'b0 ;
  assign n25003 = n25002 ^ n23690 ^ 1'b0 ;
  assign n25004 = n2473 | n12212 ;
  assign n25005 = n25004 ^ n2727 ^ 1'b0 ;
  assign n25006 = ~n1832 & n25005 ;
  assign n25007 = n25006 ^ n6484 ^ 1'b0 ;
  assign n25008 = ~n25003 & n25007 ;
  assign n25009 = n9309 & n13425 ;
  assign n25010 = n20135 ^ n7395 ^ n6656 ;
  assign n25011 = n1476 & ~n6802 ;
  assign n25012 = n25011 ^ n1842 ^ 1'b0 ;
  assign n25013 = n25010 & ~n25012 ;
  assign n25014 = n23383 ^ n663 ^ 1'b0 ;
  assign n25015 = n25014 ^ n17513 ^ n14971 ;
  assign n25016 = ~n3312 & n5436 ;
  assign n25017 = n25016 ^ n3056 ^ 1'b0 ;
  assign n25018 = ( n7652 & n11489 ) | ( n7652 & n25017 ) | ( n11489 & n25017 ) ;
  assign n25019 = ( n1931 & n5143 ) | ( n1931 & ~n17774 ) | ( n5143 & ~n17774 ) ;
  assign n25020 = n17159 ^ n12714 ^ 1'b0 ;
  assign n25021 = n25020 ^ n11557 ^ 1'b0 ;
  assign n25022 = n4260 | n25021 ;
  assign n25023 = n16921 & ~n25022 ;
  assign n25024 = ( ~n10361 & n10520 ) | ( ~n10361 & n19062 ) | ( n10520 & n19062 ) ;
  assign n25025 = n10016 ^ n2315 ^ 1'b0 ;
  assign n25026 = ( n2481 & n19975 ) | ( n2481 & ~n25025 ) | ( n19975 & ~n25025 ) ;
  assign n25027 = n13910 ^ n5580 ^ 1'b0 ;
  assign n25028 = n1150 & n13874 ;
  assign n25032 = n11462 | n20196 ;
  assign n25033 = n25032 ^ n5595 ^ 1'b0 ;
  assign n25034 = n25033 ^ n4489 ^ 1'b0 ;
  assign n25029 = ~n487 & n7223 ;
  assign n25030 = n16199 ^ n16154 ^ n3053 ;
  assign n25031 = n25029 | n25030 ;
  assign n25035 = n25034 ^ n25031 ^ 1'b0 ;
  assign n25036 = n25035 ^ n21319 ^ 1'b0 ;
  assign n25037 = x108 | n12198 ;
  assign n25038 = n25037 ^ n602 ^ 1'b0 ;
  assign n25039 = n5855 & n12153 ;
  assign n25040 = n25039 ^ n317 ^ 1'b0 ;
  assign n25041 = ( n18830 & n20297 ) | ( n18830 & ~n25040 ) | ( n20297 & ~n25040 ) ;
  assign n25042 = n12394 & ~n14476 ;
  assign n25043 = n25042 ^ n23541 ^ x115 ;
  assign n25044 = n2107 | n7287 ;
  assign n25045 = n7693 ^ n4915 ^ 1'b0 ;
  assign n25046 = ( n10218 & n25044 ) | ( n10218 & ~n25045 ) | ( n25044 & ~n25045 ) ;
  assign n25047 = n17305 & ~n25046 ;
  assign n25048 = n8356 & n13399 ;
  assign n25049 = n6239 | n8893 ;
  assign n25050 = n6068 & ~n25049 ;
  assign n25051 = n7754 ^ n6601 ^ 1'b0 ;
  assign n25052 = n16445 ^ n4805 ^ 1'b0 ;
  assign n25053 = n6988 | n25052 ;
  assign n25054 = n17517 ^ n11499 ^ 1'b0 ;
  assign n25055 = ~n15969 & n25054 ;
  assign n25056 = n813 | n4520 ;
  assign n25057 = n7568 ^ n2972 ^ n959 ;
  assign n25058 = n19126 & ~n25057 ;
  assign n25059 = n4611 | n5460 ;
  assign n25060 = ~n19849 & n25059 ;
  assign n25061 = n9552 & ~n22236 ;
  assign n25062 = n16382 & n25061 ;
  assign n25063 = n2808 ^ n378 ^ 1'b0 ;
  assign n25064 = n25063 ^ n2169 ^ 1'b0 ;
  assign n25065 = ~n18318 & n25064 ;
  assign n25066 = n25062 | n25065 ;
  assign n25067 = n1964 | n3037 ;
  assign n25068 = n9927 & ~n25067 ;
  assign n25069 = n25068 ^ n17649 ^ 1'b0 ;
  assign n25070 = n5328 & n25069 ;
  assign n25071 = x251 & n25070 ;
  assign n25072 = n7507 | n10820 ;
  assign n25073 = n15343 | n25072 ;
  assign n25074 = n21855 | n25073 ;
  assign n25075 = n25074 ^ n23512 ^ 1'b0 ;
  assign n25076 = n23148 ^ n3071 ^ 1'b0 ;
  assign n25077 = n20749 ^ n20168 ^ 1'b0 ;
  assign n25078 = n4311 & n15059 ;
  assign n25079 = n9082 ^ n3960 ^ n1519 ;
  assign n25080 = n1472 & n9132 ;
  assign n25081 = n25080 ^ n16551 ^ n4795 ;
  assign n25082 = n25079 | n25081 ;
  assign n25083 = n25082 ^ n15270 ^ 1'b0 ;
  assign n25084 = ( n22040 & ~n25078 ) | ( n22040 & n25083 ) | ( ~n25078 & n25083 ) ;
  assign n25085 = n21820 & ~n25084 ;
  assign n25088 = ( n16232 & ~n18321 ) | ( n16232 & n20168 ) | ( ~n18321 & n20168 ) ;
  assign n25086 = n20917 ^ n10971 ^ n6306 ;
  assign n25087 = n10816 | n25086 ;
  assign n25089 = n25088 ^ n25087 ^ 1'b0 ;
  assign n25090 = n8355 | n22107 ;
  assign n25091 = n7620 ^ n4601 ^ 1'b0 ;
  assign n25092 = n15954 & ~n25091 ;
  assign n25093 = n18147 & ~n25092 ;
  assign n25098 = n14672 ^ n3172 ^ 1'b0 ;
  assign n25096 = n305 & n3185 ;
  assign n25097 = n25096 ^ n7589 ^ 1'b0 ;
  assign n25094 = ~n9756 & n21478 ;
  assign n25095 = ~x194 & n25094 ;
  assign n25099 = n25098 ^ n25097 ^ n25095 ;
  assign n25100 = n11407 ^ n1387 ^ 1'b0 ;
  assign n25101 = n24908 | n25100 ;
  assign n25102 = n25101 ^ n10771 ^ n3080 ;
  assign n25103 = n6439 ^ n3429 ^ n741 ;
  assign n25104 = n10881 | n15195 ;
  assign n25105 = n25103 & ~n25104 ;
  assign n25108 = ~n1975 & n6875 ;
  assign n25109 = n25108 ^ n5991 ^ 1'b0 ;
  assign n25106 = n3267 & n17896 ;
  assign n25107 = ~n19449 & n25106 ;
  assign n25110 = n25109 ^ n25107 ^ 1'b0 ;
  assign n25111 = n8015 | n25110 ;
  assign n25112 = n25111 ^ n23423 ^ 1'b0 ;
  assign n25113 = n16342 ^ n2067 ^ 1'b0 ;
  assign n25114 = n461 & ~n25113 ;
  assign n25115 = n21194 & n25114 ;
  assign n25116 = ~n12839 & n25115 ;
  assign n25117 = n19968 ^ n16700 ^ 1'b0 ;
  assign n25118 = n10125 & ~n23703 ;
  assign n25119 = n25118 ^ n16923 ^ 1'b0 ;
  assign n25120 = n14415 ^ n6551 ^ 1'b0 ;
  assign n25121 = ( n25117 & n25119 ) | ( n25117 & ~n25120 ) | ( n25119 & ~n25120 ) ;
  assign n25122 = n10590 ^ n440 ^ 1'b0 ;
  assign n25123 = n1133 & n25122 ;
  assign n25124 = ( n1900 & n10106 ) | ( n1900 & n25123 ) | ( n10106 & n25123 ) ;
  assign n25125 = ( ~n5840 & n16673 ) | ( ~n5840 & n25124 ) | ( n16673 & n25124 ) ;
  assign n25126 = n9759 ^ n2094 ^ 1'b0 ;
  assign n25127 = x159 & n25126 ;
  assign n25128 = n25127 ^ n13420 ^ n5413 ;
  assign n25129 = n10507 & ~n25128 ;
  assign n25130 = n22089 ^ n6867 ^ 1'b0 ;
  assign n25131 = ( n596 & ~n1780 ) | ( n596 & n2233 ) | ( ~n1780 & n2233 ) ;
  assign n25132 = n25131 ^ n3370 ^ 1'b0 ;
  assign n25133 = n25130 | n25132 ;
  assign n25134 = n24037 ^ n7758 ^ 1'b0 ;
  assign n25135 = n13114 ^ n5285 ^ n4446 ;
  assign n25136 = n11327 & ~n22379 ;
  assign n25137 = ~n5396 & n25136 ;
  assign n25138 = n9448 ^ n8524 ^ 1'b0 ;
  assign n25139 = ~n1430 & n25138 ;
  assign n25140 = n25139 ^ n10449 ^ 1'b0 ;
  assign n25141 = n8572 & n9705 ;
  assign n25142 = n15313 | n25141 ;
  assign n25143 = ~n5406 & n10383 ;
  assign n25144 = n23550 ^ x95 ^ x80 ;
  assign n25145 = n25144 ^ n9637 ^ n2488 ;
  assign n25146 = n3707 & n11072 ;
  assign n25147 = n25145 & n25146 ;
  assign n25148 = n1536 | n25147 ;
  assign n25149 = n4589 ^ n4069 ^ 1'b0 ;
  assign n25150 = n9464 & n25149 ;
  assign n25151 = n4162 & n13877 ;
  assign n25152 = n22676 ^ n5840 ^ 1'b0 ;
  assign n25153 = ~x5 & n4107 ;
  assign n25154 = ( x146 & n2892 ) | ( x146 & ~n25153 ) | ( n2892 & ~n25153 ) ;
  assign n25155 = n3158 | n7942 ;
  assign n25156 = n14172 & ~n25155 ;
  assign n25157 = n7758 ^ n2598 ^ 1'b0 ;
  assign n25158 = ~n7425 & n25141 ;
  assign n25159 = ~n9902 & n25158 ;
  assign n25166 = ( n3376 & n6921 ) | ( n3376 & ~n23105 ) | ( n6921 & ~n23105 ) ;
  assign n25161 = n2645 & n5518 ;
  assign n25162 = n25161 ^ n11977 ^ 1'b0 ;
  assign n25163 = n10644 & n25162 ;
  assign n25164 = n25163 ^ n12222 ^ 1'b0 ;
  assign n25160 = n9746 & n17553 ;
  assign n25165 = n25164 ^ n25160 ^ 1'b0 ;
  assign n25167 = n25166 ^ n25165 ^ n13643 ;
  assign n25168 = n11324 ^ n4351 ^ 1'b0 ;
  assign n25169 = n2995 | n3887 ;
  assign n25170 = ( ~n2049 & n11229 ) | ( ~n2049 & n17042 ) | ( n11229 & n17042 ) ;
  assign n25171 = n12960 ^ n10122 ^ 1'b0 ;
  assign n25172 = n25170 & n25171 ;
  assign n25173 = ~n25169 & n25172 ;
  assign n25174 = ~n5588 & n5751 ;
  assign n25175 = n464 & n25174 ;
  assign n25176 = n16594 ^ n11068 ^ 1'b0 ;
  assign n25177 = ~n25175 & n25176 ;
  assign n25178 = ~n8537 & n16051 ;
  assign n25180 = n4115 ^ n3281 ^ 1'b0 ;
  assign n25181 = n25180 ^ n4081 ^ 1'b0 ;
  assign n25182 = n16152 & ~n25181 ;
  assign n25179 = n5191 ^ n3190 ^ 1'b0 ;
  assign n25183 = n25182 ^ n25179 ^ 1'b0 ;
  assign n25185 = ( n665 & n7556 ) | ( n665 & n16468 ) | ( n7556 & n16468 ) ;
  assign n25184 = n8683 | n24371 ;
  assign n25186 = n25185 ^ n25184 ^ n16841 ;
  assign n25187 = n3457 & n10775 ;
  assign n25188 = ~n21080 & n25187 ;
  assign n25191 = n9123 ^ n8659 ^ 1'b0 ;
  assign n25189 = n21851 ^ n3531 ^ 1'b0 ;
  assign n25190 = n12936 & ~n25189 ;
  assign n25192 = n25191 ^ n25190 ^ 1'b0 ;
  assign n25193 = n25188 | n25192 ;
  assign n25194 = n1678 | n6624 ;
  assign n25195 = n25194 ^ n3954 ^ 1'b0 ;
  assign n25196 = ~n290 & n22484 ;
  assign n25197 = n1038 | n13542 ;
  assign n25198 = n17091 & ~n25197 ;
  assign n25199 = ~n2648 & n11716 ;
  assign n25200 = n19581 ^ x57 ^ 1'b0 ;
  assign n25201 = n7051 & ~n25200 ;
  assign n25202 = n25201 ^ n4552 ^ 1'b0 ;
  assign n25203 = ~n8732 & n25202 ;
  assign n25204 = n22766 ^ n9512 ^ n5841 ;
  assign n25205 = n25203 & n25204 ;
  assign n25206 = ( n16417 & ~n16590 ) | ( n16417 & n16880 ) | ( ~n16590 & n16880 ) ;
  assign n25207 = n25206 ^ n18072 ^ n10706 ;
  assign n25208 = n11206 ^ n5081 ^ n1000 ;
  assign n25209 = n7782 & ~n17639 ;
  assign n25210 = x177 & n6308 ;
  assign n25211 = n25210 ^ x50 ^ 1'b0 ;
  assign n25212 = n23941 & ~n25211 ;
  assign n25213 = n18757 ^ n12963 ^ n9846 ;
  assign n25214 = n21793 & ~n25213 ;
  assign n25220 = ~n2471 & n6706 ;
  assign n25219 = n8719 | n9000 ;
  assign n25221 = n25220 ^ n25219 ^ 1'b0 ;
  assign n25222 = x0 & ~n5627 ;
  assign n25223 = n25222 ^ n2283 ^ 1'b0 ;
  assign n25224 = ( n887 & n12326 ) | ( n887 & ~n25223 ) | ( n12326 & ~n25223 ) ;
  assign n25225 = ( n4327 & ~n25221 ) | ( n4327 & n25224 ) | ( ~n25221 & n25224 ) ;
  assign n25215 = n8268 | n22444 ;
  assign n25216 = n24566 ^ n4461 ^ 1'b0 ;
  assign n25217 = ~n1425 & n25216 ;
  assign n25218 = ~n25215 & n25217 ;
  assign n25226 = n25225 ^ n25218 ^ 1'b0 ;
  assign n25230 = n1113 | n1322 ;
  assign n25231 = n25230 ^ n1450 ^ 1'b0 ;
  assign n25227 = n4298 & n13345 ;
  assign n25228 = ~n8895 & n25227 ;
  assign n25229 = n20923 & ~n25228 ;
  assign n25232 = n25231 ^ n25229 ^ 1'b0 ;
  assign n25233 = ( n6276 & n8954 ) | ( n6276 & ~n11236 ) | ( n8954 & ~n11236 ) ;
  assign n25234 = n21474 & n25233 ;
  assign n25235 = n7362 & n23608 ;
  assign n25236 = n18618 & ~n25070 ;
  assign n25237 = n14169 & ~n15451 ;
  assign n25238 = n9762 | n20798 ;
  assign n25239 = n19703 | n25238 ;
  assign n25240 = ~n12402 & n25239 ;
  assign n25241 = ~n2086 & n25240 ;
  assign n25242 = n4471 | n6983 ;
  assign n25243 = n4471 & ~n25242 ;
  assign n25244 = ( ~n2427 & n2452 ) | ( ~n2427 & n25243 ) | ( n2452 & n25243 ) ;
  assign n25245 = ( ~n3935 & n4013 ) | ( ~n3935 & n12390 ) | ( n4013 & n12390 ) ;
  assign n25246 = n9161 | n17607 ;
  assign n25247 = n25246 ^ n8569 ^ 1'b0 ;
  assign n25248 = n13537 | n20995 ;
  assign n25250 = n13562 ^ n11908 ^ 1'b0 ;
  assign n25252 = n8784 ^ n5692 ^ n1927 ;
  assign n25251 = n9067 ^ n8026 ^ n3585 ;
  assign n25253 = n25252 ^ n25251 ^ 1'b0 ;
  assign n25254 = n25250 & ~n25253 ;
  assign n25249 = n21213 ^ n9378 ^ 1'b0 ;
  assign n25255 = n25254 ^ n25249 ^ 1'b0 ;
  assign n25256 = n21827 & ~n25255 ;
  assign n25261 = n20861 ^ n8103 ^ n7212 ;
  assign n25257 = ~n7257 & n10340 ;
  assign n25258 = n25257 ^ n3874 ^ 1'b0 ;
  assign n25259 = n10303 & n17714 ;
  assign n25260 = n25258 | n25259 ;
  assign n25262 = n25261 ^ n25260 ^ 1'b0 ;
  assign n25263 = n385 & ~n20008 ;
  assign n25264 = n19495 & n25263 ;
  assign n25265 = n15032 ^ n9139 ^ 1'b0 ;
  assign n25266 = n5281 & ~n12365 ;
  assign n25267 = ( n3049 & ~n7354 ) | ( n3049 & n10806 ) | ( ~n7354 & n10806 ) ;
  assign n25268 = n20235 & ~n25267 ;
  assign n25274 = n19017 ^ n4699 ^ n2995 ;
  assign n25269 = n14905 ^ n3604 ^ n2052 ;
  assign n25270 = n25269 ^ n13015 ^ n10644 ;
  assign n25271 = n7601 & ~n25270 ;
  assign n25272 = n21792 | n25271 ;
  assign n25273 = n14730 & ~n25272 ;
  assign n25275 = n25274 ^ n25273 ^ 1'b0 ;
  assign n25276 = n958 | n25275 ;
  assign n25277 = n12522 ^ n7893 ^ n2465 ;
  assign n25278 = n25277 ^ n21340 ^ n5199 ;
  assign n25279 = n5609 & ~n10912 ;
  assign n25280 = n8300 | n25279 ;
  assign n25281 = n5351 & n25280 ;
  assign n25282 = n25281 ^ n4678 ^ 1'b0 ;
  assign n25283 = ~n17498 & n20433 ;
  assign n25284 = n17160 & n25283 ;
  assign n25285 = n20134 ^ n15520 ^ 1'b0 ;
  assign n25286 = n7029 & n12285 ;
  assign n25287 = n25286 ^ n23754 ^ n2824 ;
  assign n25288 = n4858 & ~n22108 ;
  assign n25289 = n25288 ^ n12285 ^ 1'b0 ;
  assign n25290 = ( n5398 & n20992 ) | ( n5398 & ~n24846 ) | ( n20992 & ~n24846 ) ;
  assign n25291 = n25290 ^ n20173 ^ 1'b0 ;
  assign n25292 = n5679 & n25291 ;
  assign n25293 = n23191 ^ n4179 ^ 1'b0 ;
  assign n25294 = ~n8325 & n25293 ;
  assign n25295 = n528 & n25294 ;
  assign n25296 = n25295 ^ n9941 ^ 1'b0 ;
  assign n25297 = ~n17916 & n25296 ;
  assign n25298 = ~n25292 & n25297 ;
  assign n25299 = n24210 ^ n16757 ^ n5827 ;
  assign n25300 = ~n5791 & n25299 ;
  assign n25301 = ~n5451 & n7859 ;
  assign n25302 = n25301 ^ n1156 ^ 1'b0 ;
  assign n25303 = ( ~n7037 & n12715 ) | ( ~n7037 & n25302 ) | ( n12715 & n25302 ) ;
  assign n25304 = n25303 ^ n11228 ^ 1'b0 ;
  assign n25305 = n24890 ^ n3714 ^ 1'b0 ;
  assign n25306 = n5269 & ~n25305 ;
  assign n25307 = ~n25304 & n25306 ;
  assign n25308 = ~n6649 & n17299 ;
  assign n25309 = ~n18525 & n25308 ;
  assign n25310 = n12550 ^ n8888 ^ 1'b0 ;
  assign n25311 = ~n25309 & n25310 ;
  assign n25312 = n1521 | n12164 ;
  assign n25313 = n25312 ^ n4069 ^ 1'b0 ;
  assign n25314 = ( n845 & n3855 ) | ( n845 & n24414 ) | ( n3855 & n24414 ) ;
  assign n25315 = n14881 ^ n3299 ^ 1'b0 ;
  assign n25316 = n854 & n25315 ;
  assign n25317 = ( n25313 & n25314 ) | ( n25313 & n25316 ) | ( n25314 & n25316 ) ;
  assign n25318 = n3152 & ~n18010 ;
  assign n25319 = n25318 ^ n14331 ^ 1'b0 ;
  assign n25320 = n25319 ^ n8816 ^ x135 ;
  assign n25321 = ( n11097 & n21221 ) | ( n11097 & n21261 ) | ( n21221 & n21261 ) ;
  assign n25322 = n3802 & ~n24852 ;
  assign n25323 = n12617 ^ n8787 ^ n3332 ;
  assign n25324 = n9086 ^ n2451 ^ 1'b0 ;
  assign n25325 = n1124 | n25324 ;
  assign n25326 = ~n6636 & n7871 ;
  assign n25327 = n25326 ^ n2650 ^ 1'b0 ;
  assign n25328 = n25327 ^ n14789 ^ 1'b0 ;
  assign n25329 = ( ~n25323 & n25325 ) | ( ~n25323 & n25328 ) | ( n25325 & n25328 ) ;
  assign n25330 = n12466 | n25329 ;
  assign n25331 = n25330 ^ n14311 ^ 1'b0 ;
  assign n25332 = n25068 ^ n22211 ^ n13251 ;
  assign n25333 = n12183 & n19908 ;
  assign n25334 = n25333 ^ n2229 ^ n1476 ;
  assign n25335 = n4395 & n4947 ;
  assign n25336 = n25334 | n25335 ;
  assign n25337 = n795 | n6506 ;
  assign n25338 = n797 | n25337 ;
  assign n25339 = n2844 | n11426 ;
  assign n25340 = n25338 | n25339 ;
  assign n25341 = ( n554 & n13314 ) | ( n554 & n25340 ) | ( n13314 & n25340 ) ;
  assign n25342 = n4827 | n13297 ;
  assign n25343 = n25341 & ~n25342 ;
  assign n25344 = n2192 & n16928 ;
  assign n25345 = n25344 ^ n3277 ^ 1'b0 ;
  assign n25346 = n25345 ^ n24673 ^ 1'b0 ;
  assign n25347 = n20384 | n25346 ;
  assign n25348 = n9687 ^ n8692 ^ 1'b0 ;
  assign n25349 = n4300 & n25348 ;
  assign n25350 = ~n16561 & n25349 ;
  assign n25351 = n25350 ^ n4495 ^ 1'b0 ;
  assign n25352 = n2243 & n25351 ;
  assign n25353 = n25352 ^ n20508 ^ 1'b0 ;
  assign n25354 = n16814 ^ n9226 ^ 1'b0 ;
  assign n25355 = n25354 ^ n1985 ^ 1'b0 ;
  assign n25356 = n25355 ^ n6689 ^ n1225 ;
  assign n25357 = n3349 | n25356 ;
  assign n25358 = n25353 | n25357 ;
  assign n25359 = n11670 & n12220 ;
  assign n25360 = n25359 ^ n6981 ^ n6046 ;
  assign n25361 = ~x198 & n3244 ;
  assign n25362 = n25361 ^ n5017 ^ 1'b0 ;
  assign n25363 = n5296 | n25362 ;
  assign n25364 = n25363 ^ n409 ^ 1'b0 ;
  assign n25365 = n5911 & ~n25364 ;
  assign n25366 = n25365 ^ n20334 ^ 1'b0 ;
  assign n25367 = n13950 ^ n13670 ^ 1'b0 ;
  assign n25368 = ~n5377 & n25367 ;
  assign n25369 = ~n8539 & n25368 ;
  assign n25370 = n14641 ^ n840 ^ 1'b0 ;
  assign n25371 = n25369 & ~n25370 ;
  assign n25372 = n2603 | n10541 ;
  assign n25373 = n17542 ^ n10739 ^ 1'b0 ;
  assign n25374 = n25372 | n25373 ;
  assign n25375 = n1023 & ~n5791 ;
  assign n25376 = ~n883 & n25375 ;
  assign n25377 = n23798 ^ n18436 ^ 1'b0 ;
  assign n25378 = ( ~n6157 & n25376 ) | ( ~n6157 & n25377 ) | ( n25376 & n25377 ) ;
  assign n25379 = n16001 ^ n12718 ^ n8597 ;
  assign n25380 = n15353 ^ n15256 ^ n2879 ;
  assign n25381 = ~n1350 & n25380 ;
  assign n25382 = ~n25379 & n25381 ;
  assign n25383 = n2173 & ~n12180 ;
  assign n25384 = ( x200 & ~n1543 ) | ( x200 & n25383 ) | ( ~n1543 & n25383 ) ;
  assign n25385 = n8001 & n25384 ;
  assign n25386 = ~n4411 & n25385 ;
  assign n25387 = n20009 ^ n11200 ^ 1'b0 ;
  assign n25388 = ~n14405 & n25387 ;
  assign n25389 = n3406 ^ n2649 ^ 1'b0 ;
  assign n25390 = n25389 ^ n20768 ^ 1'b0 ;
  assign n25391 = ~x85 & n24568 ;
  assign n25392 = ( n12273 & ~n13179 ) | ( n12273 & n18017 ) | ( ~n13179 & n18017 ) ;
  assign n25393 = n25392 ^ n621 ^ 1'b0 ;
  assign n25394 = n8149 ^ n2425 ^ 1'b0 ;
  assign n25395 = n8401 | n25394 ;
  assign n25396 = n4553 & ~n25395 ;
  assign n25397 = n22304 | n25396 ;
  assign n25398 = n16934 | n25397 ;
  assign n25399 = n15465 | n15715 ;
  assign n25400 = n6901 & ~n7787 ;
  assign n25403 = ( ~n15085 & n15493 ) | ( ~n15085 & n24321 ) | ( n15493 & n24321 ) ;
  assign n25401 = n4280 ^ n483 ^ 1'b0 ;
  assign n25402 = n3356 & ~n25401 ;
  assign n25404 = n25403 ^ n25402 ^ 1'b0 ;
  assign n25405 = ( n8767 & ~n25400 ) | ( n8767 & n25404 ) | ( ~n25400 & n25404 ) ;
  assign n25406 = n18217 ^ n15821 ^ n15273 ;
  assign n25407 = ~n501 & n3543 ;
  assign n25408 = ~n5840 & n25407 ;
  assign n25409 = n11450 | n25408 ;
  assign n25410 = n25409 ^ n10132 ^ 1'b0 ;
  assign n25411 = ( n13433 & n25406 ) | ( n13433 & n25410 ) | ( n25406 & n25410 ) ;
  assign n25412 = n18293 & ~n19894 ;
  assign n25413 = n15327 ^ n10835 ^ 1'b0 ;
  assign n25414 = n6894 | n25413 ;
  assign n25415 = n8603 | n14642 ;
  assign n25416 = ( n2416 & ~n14389 ) | ( n2416 & n25415 ) | ( ~n14389 & n25415 ) ;
  assign n25417 = ( n8984 & ~n16123 ) | ( n8984 & n25040 ) | ( ~n16123 & n25040 ) ;
  assign n25418 = n5437 ^ x224 ^ 1'b0 ;
  assign n25419 = n22553 & ~n25418 ;
  assign n25420 = n2875 & n4959 ;
  assign n25421 = n25420 ^ n17434 ^ 1'b0 ;
  assign n25422 = n5622 & n25421 ;
  assign n25423 = ~n25419 & n25422 ;
  assign n25424 = n12847 & ~n25423 ;
  assign n25425 = n3952 | n11425 ;
  assign n25426 = n11504 & ~n25425 ;
  assign n25427 = n5793 | n20650 ;
  assign n25428 = n25426 & ~n25427 ;
  assign n25429 = n5818 & n17375 ;
  assign n25430 = n25429 ^ n4170 ^ 1'b0 ;
  assign n25431 = n12123 ^ n9177 ^ 1'b0 ;
  assign n25432 = n25430 & n25431 ;
  assign n25437 = n1145 | n6986 ;
  assign n25438 = n17683 & ~n25437 ;
  assign n25435 = x120 & n1538 ;
  assign n25436 = ~n9690 & n25435 ;
  assign n25439 = n25438 ^ n25436 ^ n4088 ;
  assign n25433 = n3550 & n10285 ;
  assign n25434 = ( ~x215 & n5203 ) | ( ~x215 & n25433 ) | ( n5203 & n25433 ) ;
  assign n25440 = n25439 ^ n25434 ^ 1'b0 ;
  assign n25441 = n21647 ^ n16103 ^ 1'b0 ;
  assign n25442 = ~n663 & n25441 ;
  assign n25443 = n25442 ^ n15141 ^ 1'b0 ;
  assign n25444 = ~n25362 & n25443 ;
  assign n25445 = n25444 ^ n25404 ^ 1'b0 ;
  assign n25446 = n12505 | n15001 ;
  assign n25447 = n25446 ^ n15894 ^ 1'b0 ;
  assign n25448 = n4473 | n25447 ;
  assign n25449 = ( n11612 & n12721 ) | ( n11612 & n19615 ) | ( n12721 & n19615 ) ;
  assign n25450 = ~n1951 & n2019 ;
  assign n25451 = n7073 | n17295 ;
  assign n25452 = n25451 ^ n15039 ^ 1'b0 ;
  assign n25453 = n25450 | n25452 ;
  assign n25454 = n18007 ^ n4444 ^ 1'b0 ;
  assign n25455 = n11385 | n25454 ;
  assign n25456 = n2277 | n6130 ;
  assign n25457 = n25456 ^ n2085 ^ 1'b0 ;
  assign n25458 = ( x16 & n23448 ) | ( x16 & n25457 ) | ( n23448 & n25457 ) ;
  assign n25459 = n2221 & ~n6720 ;
  assign n25460 = ~n12828 & n25459 ;
  assign n25461 = n25460 ^ n9488 ^ n5053 ;
  assign n25462 = ~n11678 & n25461 ;
  assign n25463 = ~n1250 & n12003 ;
  assign n25464 = ( n1007 & n1205 ) | ( n1007 & ~n3368 ) | ( n1205 & ~n3368 ) ;
  assign n25465 = ( n4206 & n15572 ) | ( n4206 & ~n25464 ) | ( n15572 & ~n25464 ) ;
  assign n25466 = n24551 ^ n12836 ^ 1'b0 ;
  assign n25467 = n3094 & n25466 ;
  assign n25468 = ~n25465 & n25467 ;
  assign n25469 = n15415 & n25468 ;
  assign n25470 = n23884 & ~n25289 ;
  assign n25471 = n25470 ^ n11051 ^ 1'b0 ;
  assign n25472 = n440 | n7497 ;
  assign n25473 = n25472 ^ n1752 ^ 1'b0 ;
  assign n25474 = ~n10643 & n11956 ;
  assign n25475 = n25474 ^ n15336 ^ 1'b0 ;
  assign n25476 = x43 | n25475 ;
  assign n25477 = n16049 | n25476 ;
  assign n25478 = n25473 | n25477 ;
  assign n25479 = n8049 | n22207 ;
  assign n25480 = ( n6747 & n11338 ) | ( n6747 & n14721 ) | ( n11338 & n14721 ) ;
  assign n25481 = ~n2780 & n25366 ;
  assign n25482 = n25481 ^ n5764 ^ 1'b0 ;
  assign n25484 = n4550 & n9631 ;
  assign n25485 = n2264 & n3187 ;
  assign n25486 = ~n10285 & n25485 ;
  assign n25487 = n25484 | n25486 ;
  assign n25483 = n9958 & n24778 ;
  assign n25488 = n25487 ^ n25483 ^ 1'b0 ;
  assign n25489 = n5439 ^ n4823 ^ 1'b0 ;
  assign n25490 = n25489 ^ n6147 ^ 1'b0 ;
  assign n25491 = n6071 & ~n25490 ;
  assign n25492 = n25491 ^ n3758 ^ 1'b0 ;
  assign n25493 = n18395 ^ n18174 ^ n6432 ;
  assign n25494 = n24541 ^ n7701 ^ 1'b0 ;
  assign n25495 = n10068 ^ n4506 ^ 1'b0 ;
  assign n25496 = n18926 ^ n10986 ^ 1'b0 ;
  assign n25497 = n23351 | n25496 ;
  assign n25498 = ( n15159 & n24370 ) | ( n15159 & ~n25497 ) | ( n24370 & ~n25497 ) ;
  assign n25499 = n25498 ^ n10317 ^ n4059 ;
  assign n25500 = ( x118 & n7653 ) | ( x118 & n20577 ) | ( n7653 & n20577 ) ;
  assign n25501 = n10780 & n21987 ;
  assign n25502 = n9494 ^ n6196 ^ 1'b0 ;
  assign n25503 = n8572 & ~n25502 ;
  assign n25504 = n17627 ^ n7282 ^ 1'b0 ;
  assign n25505 = n5762 ^ x179 ^ 1'b0 ;
  assign n25506 = n2767 & n5850 ;
  assign n25507 = n25506 ^ n11381 ^ 1'b0 ;
  assign n25508 = n3905 & n8896 ;
  assign n25509 = n25508 ^ n16175 ^ 1'b0 ;
  assign n25510 = n24822 ^ n19696 ^ 1'b0 ;
  assign n25511 = n12877 ^ n1347 ^ 1'b0 ;
  assign n25512 = ~n14549 & n25511 ;
  assign n25513 = n25512 ^ n6105 ^ 1'b0 ;
  assign n25514 = n25510 & n25513 ;
  assign n25515 = n14859 ^ n8263 ^ 1'b0 ;
  assign n25516 = ( n15776 & n17880 ) | ( n15776 & ~n25515 ) | ( n17880 & ~n25515 ) ;
  assign n25517 = n1944 | n5516 ;
  assign n25518 = n25517 ^ n2073 ^ 1'b0 ;
  assign n25519 = ~n12261 & n25518 ;
  assign n25520 = n25519 ^ n11873 ^ 1'b0 ;
  assign n25521 = n17464 & n25520 ;
  assign n25522 = ( n4139 & ~n21593 ) | ( n4139 & n25521 ) | ( ~n21593 & n25521 ) ;
  assign n25523 = ~n3894 & n16569 ;
  assign n25524 = ~n6782 & n10738 ;
  assign n25525 = ~n3378 & n25524 ;
  assign n25526 = n14942 | n20627 ;
  assign n25527 = n7626 & ~n25526 ;
  assign n25530 = x7 & n2112 ;
  assign n25531 = n5929 ^ n5844 ^ 1'b0 ;
  assign n25532 = n15149 & ~n25531 ;
  assign n25533 = n25530 & n25532 ;
  assign n25528 = n19409 ^ n9257 ^ x57 ;
  assign n25529 = ~n16964 & n25528 ;
  assign n25534 = n25533 ^ n25529 ^ n2546 ;
  assign n25535 = n9413 | n25534 ;
  assign n25536 = n12317 & ~n25535 ;
  assign n25537 = n13312 ^ n3475 ^ 1'b0 ;
  assign n25538 = n6389 | n25537 ;
  assign n25539 = ( ~n10560 & n23049 ) | ( ~n10560 & n25538 ) | ( n23049 & n25538 ) ;
  assign n25540 = n23874 ^ n2680 ^ 1'b0 ;
  assign n25541 = n2964 ^ n1064 ^ 1'b0 ;
  assign n25542 = n18778 ^ n3454 ^ 1'b0 ;
  assign n25543 = n18617 ^ n13606 ^ 1'b0 ;
  assign n25544 = n885 | n25543 ;
  assign n25546 = n25442 ^ n3856 ^ n2038 ;
  assign n25545 = n6477 | n17579 ;
  assign n25547 = n25546 ^ n25545 ^ n22251 ;
  assign n25548 = ~n684 & n25547 ;
  assign n25549 = ( n385 & n3425 ) | ( n385 & ~n24422 ) | ( n3425 & ~n24422 ) ;
  assign n25550 = n25549 ^ n16253 ^ n6140 ;
  assign n25551 = n5869 ^ n1244 ^ 1'b0 ;
  assign n25552 = n2677 | n25551 ;
  assign n25553 = ~n2202 & n4614 ;
  assign n25554 = ~n12489 & n25553 ;
  assign n25555 = n766 & ~n25554 ;
  assign n25556 = n25555 ^ n4343 ^ 1'b0 ;
  assign n25557 = ~n25552 & n25556 ;
  assign n25558 = n2995 & ~n12589 ;
  assign n25559 = n3724 & n4744 ;
  assign n25560 = ~n25558 & n25559 ;
  assign n25561 = ( n3053 & n13333 ) | ( n3053 & ~n16419 ) | ( n13333 & ~n16419 ) ;
  assign n25562 = ( ~n2389 & n6644 ) | ( ~n2389 & n9889 ) | ( n6644 & n9889 ) ;
  assign n25563 = n6588 | n25562 ;
  assign n25564 = n25563 ^ n5301 ^ 1'b0 ;
  assign n25565 = n16829 & ~n25564 ;
  assign n25566 = n25565 ^ n12758 ^ 1'b0 ;
  assign n25567 = n16142 ^ x172 ^ 1'b0 ;
  assign n25568 = n3980 | n25567 ;
  assign n25569 = ( n8192 & n12099 ) | ( n8192 & n13604 ) | ( n12099 & n13604 ) ;
  assign n25570 = n25569 ^ n18162 ^ 1'b0 ;
  assign n25571 = n18641 | n25570 ;
  assign n25572 = n6056 ^ n5170 ^ 1'b0 ;
  assign n25573 = n25572 ^ n2832 ^ 1'b0 ;
  assign n25574 = n24305 & ~n25573 ;
  assign n25575 = n21691 ^ n10436 ^ n6514 ;
  assign n25576 = ( ~n6715 & n9274 ) | ( ~n6715 & n17161 ) | ( n9274 & n17161 ) ;
  assign n25577 = n24398 ^ n10950 ^ n5302 ;
  assign n25578 = ~n15885 & n25577 ;
  assign n25579 = n19100 ^ n12678 ^ 1'b0 ;
  assign n25580 = n25579 ^ n25498 ^ n19276 ;
  assign n25581 = n25580 ^ n21306 ^ 1'b0 ;
  assign n25582 = n8951 & ~n22958 ;
  assign n25583 = n21262 ^ n881 ^ 1'b0 ;
  assign n25584 = n9785 & n25583 ;
  assign n25585 = ~n5191 & n8632 ;
  assign n25586 = ( n25582 & n25584 ) | ( n25582 & n25585 ) | ( n25584 & n25585 ) ;
  assign n25587 = n25586 ^ n10631 ^ 1'b0 ;
  assign n25588 = n322 | n8924 ;
  assign n25589 = n25587 & ~n25588 ;
  assign n25590 = n20414 & ~n20836 ;
  assign n25591 = n14635 ^ n11714 ^ 1'b0 ;
  assign n25592 = n4827 & ~n14938 ;
  assign n25593 = ~n18908 & n25592 ;
  assign n25594 = n9206 & n25593 ;
  assign n25595 = n5778 | n25594 ;
  assign n25596 = n3156 & n10527 ;
  assign n25597 = n25596 ^ n7606 ^ 1'b0 ;
  assign n25598 = n25597 ^ n11889 ^ 1'b0 ;
  assign n25599 = n12772 | n25598 ;
  assign n25600 = ( ~n11157 & n25595 ) | ( ~n11157 & n25599 ) | ( n25595 & n25599 ) ;
  assign n25601 = n11448 & n11629 ;
  assign n25602 = n21434 ^ n1495 ^ 1'b0 ;
  assign n25603 = ~n23004 & n25602 ;
  assign n25604 = n2833 ^ n2216 ^ 1'b0 ;
  assign n25605 = n25604 ^ n4438 ^ n3054 ;
  assign n25606 = n25605 ^ n22941 ^ n870 ;
  assign n25607 = ( n5722 & n9795 ) | ( n5722 & ~n24402 ) | ( n9795 & ~n24402 ) ;
  assign n25608 = n1650 ^ n384 ^ x226 ;
  assign n25609 = ~n2223 & n6640 ;
  assign n25610 = n25608 & n25609 ;
  assign n25611 = n15049 & n25610 ;
  assign n25612 = n10686 & ~n19917 ;
  assign n25613 = ~n11541 & n25612 ;
  assign n25614 = ~n19192 & n25613 ;
  assign n25615 = n9588 ^ n519 ^ 1'b0 ;
  assign n25616 = ~n7197 & n25615 ;
  assign n25617 = n15046 ^ n8018 ^ 1'b0 ;
  assign n25618 = n1368 & ~n25617 ;
  assign n25619 = ( n684 & n3036 ) | ( n684 & n25618 ) | ( n3036 & n25618 ) ;
  assign n25620 = ( n11005 & n17290 ) | ( n11005 & n25619 ) | ( n17290 & n25619 ) ;
  assign n25621 = n25620 ^ n24446 ^ 1'b0 ;
  assign n25622 = n8363 & ~n25621 ;
  assign n25623 = n18077 ^ n7075 ^ 1'b0 ;
  assign n25624 = n994 & ~n6982 ;
  assign n25625 = n992 & n25624 ;
  assign n25626 = n7548 ^ n5754 ^ 1'b0 ;
  assign n25627 = ~n25625 & n25626 ;
  assign n25628 = n14889 & n25627 ;
  assign n25629 = n25628 ^ n24834 ^ 1'b0 ;
  assign n25630 = x73 & ~n9102 ;
  assign n25631 = n25630 ^ n651 ^ 1'b0 ;
  assign n25632 = ~n18825 & n25631 ;
  assign n25633 = n24786 & n25632 ;
  assign n25634 = n8590 & n19345 ;
  assign n25635 = n6612 & n25634 ;
  assign n25636 = n25635 ^ n7305 ^ 1'b0 ;
  assign n25637 = n12180 | n25636 ;
  assign n25638 = n25637 ^ n13582 ^ 1'b0 ;
  assign n25639 = n9295 ^ n8207 ^ 1'b0 ;
  assign n25640 = n7974 | n25639 ;
  assign n25641 = n9982 & ~n25640 ;
  assign n25642 = n25641 ^ n1727 ^ 1'b0 ;
  assign n25643 = n18390 ^ n5275 ^ n1425 ;
  assign n25650 = ( n1248 & ~n2016 ) | ( n1248 & n14753 ) | ( ~n2016 & n14753 ) ;
  assign n25651 = n906 & n25650 ;
  assign n25652 = n25651 ^ n5067 ^ 1'b0 ;
  assign n25653 = n3837 & n25652 ;
  assign n25654 = n25653 ^ n9378 ^ 1'b0 ;
  assign n25655 = n5741 & n25654 ;
  assign n25656 = n15366 & n25655 ;
  assign n25649 = n10339 | n10742 ;
  assign n25657 = n25656 ^ n25649 ^ 1'b0 ;
  assign n25646 = n4587 ^ n4311 ^ 1'b0 ;
  assign n25644 = n2488 | n10395 ;
  assign n25645 = n25644 ^ n14907 ^ 1'b0 ;
  assign n25647 = n25646 ^ n25645 ^ 1'b0 ;
  assign n25648 = ( ~n2259 & n19404 ) | ( ~n2259 & n25647 ) | ( n19404 & n25647 ) ;
  assign n25658 = n25657 ^ n25648 ^ n19112 ;
  assign n25659 = n24762 ^ n8867 ^ 1'b0 ;
  assign n25660 = n2137 | n25659 ;
  assign n25661 = n25660 ^ n18753 ^ 1'b0 ;
  assign n25664 = n1727 ^ n341 ^ 1'b0 ;
  assign n25665 = n25664 ^ n12061 ^ 1'b0 ;
  assign n25666 = n8588 | n25665 ;
  assign n25662 = ~n4068 & n7616 ;
  assign n25663 = n11242 & n25662 ;
  assign n25667 = n25666 ^ n25663 ^ 1'b0 ;
  assign n25668 = n17337 | n19916 ;
  assign n25669 = n9078 | n25668 ;
  assign n25671 = n7034 ^ n402 ^ 1'b0 ;
  assign n25672 = n5440 & n25671 ;
  assign n25673 = ~n24047 & n25672 ;
  assign n25674 = n25673 ^ n6005 ^ n580 ;
  assign n25670 = ~n4321 & n10412 ;
  assign n25675 = n25674 ^ n25670 ^ 1'b0 ;
  assign n25676 = n7521 ^ n3237 ^ 1'b0 ;
  assign n25677 = n1010 & ~n25676 ;
  assign n25678 = n14382 & n25677 ;
  assign n25679 = n21360 & ~n25678 ;
  assign n25684 = ~n6472 & n8683 ;
  assign n25685 = n25684 ^ n11192 ^ 1'b0 ;
  assign n25681 = x169 & n19100 ;
  assign n25680 = n22361 ^ n9645 ^ n8590 ;
  assign n25682 = n25681 ^ n25680 ^ 1'b0 ;
  assign n25683 = n462 & n25682 ;
  assign n25686 = n25685 ^ n25683 ^ 1'b0 ;
  assign n25687 = n22733 ^ n3952 ^ 1'b0 ;
  assign n25688 = ( ~n1267 & n7900 ) | ( ~n1267 & n25687 ) | ( n7900 & n25687 ) ;
  assign n25689 = n21794 ^ n2314 ^ 1'b0 ;
  assign n25690 = n25688 & n25689 ;
  assign n25691 = n25690 ^ n22430 ^ 1'b0 ;
  assign n25692 = n25691 ^ n3649 ^ n1002 ;
  assign n25693 = n20115 ^ n14856 ^ 1'b0 ;
  assign n25694 = n18509 | n25693 ;
  assign n25695 = n20021 & ~n25694 ;
  assign n25703 = n10239 | n13563 ;
  assign n25704 = n10239 & ~n25703 ;
  assign n25696 = ~n550 & n7983 ;
  assign n25697 = ~n7983 & n25696 ;
  assign n25698 = n7901 & n25697 ;
  assign n25699 = n7839 ^ n6437 ^ 1'b0 ;
  assign n25700 = n4097 & ~n25699 ;
  assign n25701 = n7315 & n25700 ;
  assign n25702 = n25698 & n25701 ;
  assign n25705 = n25704 ^ n25702 ^ 1'b0 ;
  assign n25706 = ~n8693 & n25705 ;
  assign n25707 = ~n4924 & n6524 ;
  assign n25708 = ( n14966 & ~n22788 ) | ( n14966 & n25707 ) | ( ~n22788 & n25707 ) ;
  assign n25709 = n1196 & n8831 ;
  assign n25710 = n24171 ^ n14235 ^ 1'b0 ;
  assign n25711 = n4695 | n12476 ;
  assign n25712 = n25710 & ~n25711 ;
  assign n25713 = n18797 ^ n978 ^ 1'b0 ;
  assign n25714 = n17525 ^ n1586 ^ 1'b0 ;
  assign n25715 = ~n19279 & n24077 ;
  assign n25716 = n1979 & n25715 ;
  assign n25717 = ~n850 & n24103 ;
  assign n25718 = n25717 ^ n971 ^ 1'b0 ;
  assign n25719 = n21669 ^ n6239 ^ 1'b0 ;
  assign n25720 = ~n25718 & n25719 ;
  assign n25721 = n7747 & n11108 ;
  assign n25722 = n25721 ^ n15240 ^ n1482 ;
  assign n25723 = n7044 & ~n16786 ;
  assign n25724 = n21385 ^ n15572 ^ n10248 ;
  assign n25725 = ( ~n2900 & n4965 ) | ( ~n2900 & n5027 ) | ( n4965 & n5027 ) ;
  assign n25726 = ~n4462 & n25725 ;
  assign n25727 = ( n10243 & ~n25654 ) | ( n10243 & n25726 ) | ( ~n25654 & n25726 ) ;
  assign n25728 = n7037 ^ n3817 ^ 1'b0 ;
  assign n25729 = n6077 | n25728 ;
  assign n25730 = n25729 ^ n14469 ^ n3158 ;
  assign n25731 = n25730 ^ n6322 ^ 1'b0 ;
  assign n25732 = ( n6332 & n11418 ) | ( n6332 & n25731 ) | ( n11418 & n25731 ) ;
  assign n25733 = n25732 ^ n11043 ^ 1'b0 ;
  assign n25734 = ( n1100 & ~n9410 ) | ( n1100 & n15917 ) | ( ~n9410 & n15917 ) ;
  assign n25738 = ( n9861 & n16218 ) | ( n9861 & n17051 ) | ( n16218 & n17051 ) ;
  assign n25735 = ~n2680 & n5506 ;
  assign n25736 = n25735 ^ n9370 ^ 1'b0 ;
  assign n25737 = n13818 & ~n25736 ;
  assign n25739 = n25738 ^ n25737 ^ 1'b0 ;
  assign n25740 = n15766 & n25739 ;
  assign n25741 = ~n14085 & n25740 ;
  assign n25742 = ~n588 & n8507 ;
  assign n25743 = ( n11349 & n21763 ) | ( n11349 & ~n25742 ) | ( n21763 & ~n25742 ) ;
  assign n25744 = n10162 ^ n7468 ^ n5740 ;
  assign n25745 = n23513 ^ n21465 ^ 1'b0 ;
  assign n25746 = n21888 | n25745 ;
  assign n25747 = n13114 | n25746 ;
  assign n25748 = n25747 ^ n347 ^ 1'b0 ;
  assign n25749 = ~n3081 & n25748 ;
  assign n25750 = n21222 ^ n6377 ^ n3016 ;
  assign n25751 = ~n12529 & n14765 ;
  assign n25752 = ~n13438 & n25751 ;
  assign n25753 = n9547 | n23366 ;
  assign n25754 = n25752 & ~n25753 ;
  assign n25755 = n24356 ^ n19479 ^ n13617 ;
  assign n25756 = n7810 ^ n4336 ^ 1'b0 ;
  assign n25757 = n25755 | n25756 ;
  assign n25762 = n3406 ^ n1285 ^ 1'b0 ;
  assign n25763 = n1174 & ~n5546 ;
  assign n25764 = n25762 & n25763 ;
  assign n25758 = ( x91 & ~n1467 ) | ( x91 & n17635 ) | ( ~n1467 & n17635 ) ;
  assign n25759 = ~n1350 & n25758 ;
  assign n25760 = n25759 ^ n21177 ^ 1'b0 ;
  assign n25761 = n18374 & ~n25760 ;
  assign n25765 = n25764 ^ n25761 ^ 1'b0 ;
  assign n25766 = n24062 ^ n11039 ^ 1'b0 ;
  assign n25767 = n25765 & ~n25766 ;
  assign n25768 = n9100 ^ n1140 ^ 1'b0 ;
  assign n25769 = n403 | n25768 ;
  assign n25770 = n25769 ^ n17735 ^ 1'b0 ;
  assign n25771 = n18114 ^ n13545 ^ 1'b0 ;
  assign n25772 = n2800 & n25771 ;
  assign n25773 = n21190 & n25772 ;
  assign n25774 = n18972 & n25773 ;
  assign n25775 = n15230 ^ n4432 ^ 1'b0 ;
  assign n25776 = n2314 ^ n509 ^ 1'b0 ;
  assign n25777 = ~n20422 & n25776 ;
  assign n25778 = n25777 ^ n19261 ^ 1'b0 ;
  assign n25779 = n10632 | n10863 ;
  assign n25780 = n951 & ~n25779 ;
  assign n25781 = n6652 & ~n13008 ;
  assign n25782 = ( n10326 & n12726 ) | ( n10326 & n25781 ) | ( n12726 & n25781 ) ;
  assign n25783 = ( ~n14587 & n25191 ) | ( ~n14587 & n25782 ) | ( n25191 & n25782 ) ;
  assign n25784 = n23351 ^ n12502 ^ 1'b0 ;
  assign n25785 = ( n15719 & ~n25783 ) | ( n15719 & n25784 ) | ( ~n25783 & n25784 ) ;
  assign n25787 = n6473 ^ n6368 ^ 1'b0 ;
  assign n25788 = n9587 | n25787 ;
  assign n25789 = n12595 | n23096 ;
  assign n25790 = n25788 & ~n25789 ;
  assign n25786 = ~n3320 & n16992 ;
  assign n25791 = n25790 ^ n25786 ^ n18534 ;
  assign n25792 = n10986 & n25791 ;
  assign n25793 = n6665 & n15398 ;
  assign n25794 = n5592 ^ n5109 ^ 1'b0 ;
  assign n25795 = n25793 | n25794 ;
  assign n25796 = n20768 ^ n7589 ^ 1'b0 ;
  assign n25797 = n17931 | n25796 ;
  assign n25798 = n11199 ^ n1002 ^ 1'b0 ;
  assign n25799 = n25798 ^ n637 ^ 1'b0 ;
  assign n25800 = n25799 ^ n9069 ^ 1'b0 ;
  assign n25801 = n8432 & ~n17237 ;
  assign n25805 = n1304 | n14889 ;
  assign n25802 = ~x218 & n12084 ;
  assign n25803 = ~n8675 & n25802 ;
  assign n25804 = n25803 ^ n23837 ^ n14140 ;
  assign n25806 = n25805 ^ n25804 ^ 1'b0 ;
  assign n25807 = ~n6750 & n25806 ;
  assign n25809 = ~n11663 & n19754 ;
  assign n25810 = n25809 ^ n11568 ^ 1'b0 ;
  assign n25808 = n4579 | n24618 ;
  assign n25811 = n25810 ^ n25808 ^ 1'b0 ;
  assign n25812 = n9569 ^ n3475 ^ 1'b0 ;
  assign n25813 = ~n2754 & n25812 ;
  assign n25814 = n25813 ^ n21898 ^ n6881 ;
  assign n25815 = n21674 ^ n14870 ^ 1'b0 ;
  assign n25816 = n25814 & ~n25815 ;
  assign n25817 = n20470 ^ n10416 ^ n4139 ;
  assign n25818 = n2089 | n25817 ;
  assign n25819 = n8089 | n25818 ;
  assign n25820 = n21840 & n25819 ;
  assign n25823 = n11443 & n21319 ;
  assign n25824 = ( ~n8466 & n16972 ) | ( ~n8466 & n25823 ) | ( n16972 & n25823 ) ;
  assign n25825 = ( n9897 & ~n23355 ) | ( n9897 & n25824 ) | ( ~n23355 & n25824 ) ;
  assign n25821 = n15054 ^ n3588 ^ 1'b0 ;
  assign n25822 = n12438 & ~n25821 ;
  assign n25826 = n25825 ^ n25822 ^ 1'b0 ;
  assign n25827 = n25528 ^ n24897 ^ n11156 ;
  assign n25834 = n6177 ^ n5988 ^ 1'b0 ;
  assign n25828 = ~n4489 & n15094 ;
  assign n25829 = n25828 ^ n2551 ^ 1'b0 ;
  assign n25830 = n25829 ^ n3899 ^ n3847 ;
  assign n25831 = ~n21898 & n25830 ;
  assign n25832 = n25831 ^ n9864 ^ 1'b0 ;
  assign n25833 = n13345 & ~n25832 ;
  assign n25835 = n25834 ^ n25833 ^ n3049 ;
  assign n25836 = n4788 & n15404 ;
  assign n25837 = n3608 & ~n6989 ;
  assign n25838 = n2665 & n25837 ;
  assign n25839 = ( n16078 & ~n20157 ) | ( n16078 & n25838 ) | ( ~n20157 & n25838 ) ;
  assign n25840 = n25839 ^ n4553 ^ 1'b0 ;
  assign n25841 = ( n5353 & n15744 ) | ( n5353 & n20631 ) | ( n15744 & n20631 ) ;
  assign n25842 = ~n2794 & n19488 ;
  assign n25843 = n25841 & n25842 ;
  assign n25844 = n8926 ^ n1487 ^ 1'b0 ;
  assign n25845 = n3728 & ~n25844 ;
  assign n25846 = n1725 & n25845 ;
  assign n25847 = n23114 & n25846 ;
  assign n25848 = n7932 ^ n3364 ^ 1'b0 ;
  assign n25849 = n25848 ^ n19437 ^ n6669 ;
  assign n25852 = n11177 ^ n3009 ^ 1'b0 ;
  assign n25853 = ~n16122 & n25852 ;
  assign n25850 = n7285 | n17345 ;
  assign n25851 = n5191 | n25850 ;
  assign n25854 = n25853 ^ n25851 ^ 1'b0 ;
  assign n25855 = n6130 | n25854 ;
  assign n25856 = n25849 & ~n25855 ;
  assign n25857 = n25856 ^ n4154 ^ 1'b0 ;
  assign n25858 = ( ~n3063 & n3314 ) | ( ~n3063 & n25857 ) | ( n3314 & n25857 ) ;
  assign n25859 = n1202 & n7030 ;
  assign n25860 = n25859 ^ n12259 ^ 1'b0 ;
  assign n25861 = n13189 ^ n1923 ^ 1'b0 ;
  assign n25862 = ~x226 & n19595 ;
  assign n25863 = n8525 | n13736 ;
  assign n25864 = n25863 ^ n6002 ^ 1'b0 ;
  assign n25865 = n25864 ^ n15892 ^ n1647 ;
  assign n25866 = ( n2818 & n6649 ) | ( n2818 & ~n18888 ) | ( n6649 & ~n18888 ) ;
  assign n25867 = ~n2798 & n7212 ;
  assign n25868 = n7699 | n25867 ;
  assign n25869 = n25866 | n25868 ;
  assign n25875 = ( n12723 & n16867 ) | ( n12723 & ~n22412 ) | ( n16867 & ~n22412 ) ;
  assign n25870 = ~n7562 & n8197 ;
  assign n25871 = n9987 | n17886 ;
  assign n25872 = n25871 ^ n2611 ^ 1'b0 ;
  assign n25873 = n25870 & ~n25872 ;
  assign n25874 = ~n3683 & n25873 ;
  assign n25876 = n25875 ^ n25874 ^ 1'b0 ;
  assign n25877 = x218 & n1013 ;
  assign n25878 = ( n11883 & ~n22775 ) | ( n11883 & n25877 ) | ( ~n22775 & n25877 ) ;
  assign n25881 = n10318 ^ n7842 ^ n263 ;
  assign n25879 = ( ~x82 & n11898 ) | ( ~x82 & n16113 ) | ( n11898 & n16113 ) ;
  assign n25880 = n3315 & ~n25879 ;
  assign n25882 = n25881 ^ n25880 ^ 1'b0 ;
  assign n25883 = n13369 ^ n5363 ^ n5128 ;
  assign n25884 = n20096 & n25883 ;
  assign n25885 = n25884 ^ n23293 ^ 1'b0 ;
  assign n25886 = n9084 | n10218 ;
  assign n25887 = n25886 ^ n2818 ^ 1'b0 ;
  assign n25888 = n9985 ^ n8424 ^ 1'b0 ;
  assign n25889 = n10089 ^ n9952 ^ 1'b0 ;
  assign n25892 = n23258 ^ n8368 ^ n1202 ;
  assign n25893 = n25892 ^ n22784 ^ n21452 ;
  assign n25894 = n25893 ^ n5771 ^ 1'b0 ;
  assign n25890 = n21285 | n25147 ;
  assign n25891 = n25890 ^ n3994 ^ 1'b0 ;
  assign n25895 = n25894 ^ n25891 ^ 1'b0 ;
  assign n25896 = n25889 | n25895 ;
  assign n25897 = n722 | n7068 ;
  assign n25898 = n1079 & ~n25897 ;
  assign n25899 = ~n24511 & n25898 ;
  assign n25900 = n25899 ^ n25213 ^ n22678 ;
  assign n25901 = n16444 ^ n3992 ^ 1'b0 ;
  assign n25902 = n25901 ^ n23180 ^ 1'b0 ;
  assign n25903 = n1739 & n3984 ;
  assign n25904 = ~n5193 & n25903 ;
  assign n25905 = ( n1105 & ~n21540 ) | ( n1105 & n25904 ) | ( ~n21540 & n25904 ) ;
  assign n25907 = x239 & ~n1981 ;
  assign n25908 = n25907 ^ n8565 ^ 1'b0 ;
  assign n25906 = n20747 ^ n8317 ^ n7260 ;
  assign n25909 = n25908 ^ n25906 ^ 1'b0 ;
  assign n25910 = n862 & n11347 ;
  assign n25911 = n25910 ^ n3523 ^ 1'b0 ;
  assign n25912 = ( ~n1055 & n25909 ) | ( ~n1055 & n25911 ) | ( n25909 & n25911 ) ;
  assign n25913 = ( ~n1037 & n11435 ) | ( ~n1037 & n16269 ) | ( n11435 & n16269 ) ;
  assign n25914 = n25913 ^ n3770 ^ n2619 ;
  assign n25915 = n25914 ^ n18977 ^ n12731 ;
  assign n25916 = n3674 & ~n25915 ;
  assign n25917 = ~n25912 & n25916 ;
  assign n25918 = n10527 | n25917 ;
  assign n25919 = n25918 ^ n22065 ^ 1'b0 ;
  assign n25920 = n12836 & ~n16939 ;
  assign n25921 = n8818 & n25920 ;
  assign n25922 = n13341 ^ n7958 ^ 1'b0 ;
  assign n25923 = ( n15703 & ~n16199 ) | ( n15703 & n25057 ) | ( ~n16199 & n25057 ) ;
  assign n25924 = n13545 ^ n1120 ^ 1'b0 ;
  assign n25925 = n22961 ^ n9519 ^ 1'b0 ;
  assign n25926 = ( n24555 & ~n25924 ) | ( n24555 & n25925 ) | ( ~n25924 & n25925 ) ;
  assign n25927 = ~n6330 & n8021 ;
  assign n25928 = n18643 ^ n3447 ^ 1'b0 ;
  assign n25929 = ~n25927 & n25928 ;
  assign n25932 = ( n4925 & n6093 ) | ( n4925 & ~n17397 ) | ( n6093 & ~n17397 ) ;
  assign n25933 = ~n4332 & n25932 ;
  assign n25934 = n25933 ^ n7948 ^ 1'b0 ;
  assign n25930 = n13050 ^ n5986 ^ 1'b0 ;
  assign n25931 = ( ~n816 & n22431 ) | ( ~n816 & n25930 ) | ( n22431 & n25930 ) ;
  assign n25935 = n25934 ^ n25931 ^ 1'b0 ;
  assign n25936 = n25929 & ~n25935 ;
  assign n25937 = n8360 ^ n2334 ^ 1'b0 ;
  assign n25938 = ~n21479 & n23631 ;
  assign n25939 = ~n25937 & n25938 ;
  assign n25943 = n2422 & n11699 ;
  assign n25941 = ~n800 & n4071 ;
  assign n25942 = n8129 & n25941 ;
  assign n25940 = ( n3100 & n4237 ) | ( n3100 & n14772 ) | ( n4237 & n14772 ) ;
  assign n25944 = n25943 ^ n25942 ^ n25940 ;
  assign n25945 = n7665 | n15177 ;
  assign n25946 = n16872 & ~n25945 ;
  assign n25947 = n23696 ^ n18723 ^ 1'b0 ;
  assign n25948 = n2235 | n25947 ;
  assign n25949 = n21160 ^ n10372 ^ 1'b0 ;
  assign n25950 = n14567 ^ x184 ^ 1'b0 ;
  assign n25951 = n20216 | n25950 ;
  assign n25952 = x104 & n1074 ;
  assign n25953 = n7543 & n25952 ;
  assign n25954 = n25953 ^ n4557 ^ 1'b0 ;
  assign n25955 = n25954 ^ n21023 ^ n403 ;
  assign n25956 = n17860 ^ n10928 ^ 1'b0 ;
  assign n25957 = n24358 ^ n718 ^ 1'b0 ;
  assign n25958 = n1675 & ~n1736 ;
  assign n25959 = ~n17934 & n25958 ;
  assign n25960 = ~n19571 & n25959 ;
  assign n25961 = n10076 | n25960 ;
  assign n25962 = n25961 ^ n18635 ^ 1'b0 ;
  assign n25963 = n15692 ^ n4958 ^ 1'b0 ;
  assign n25964 = n19449 ^ n10145 ^ 1'b0 ;
  assign n25965 = ~n25879 & n25964 ;
  assign n25966 = n19723 ^ n6218 ^ 1'b0 ;
  assign n25967 = n4296 | n25966 ;
  assign n25968 = n24928 ^ n7369 ^ n6509 ;
  assign n25969 = n25968 ^ n21060 ^ n3607 ;
  assign n25970 = n1586 | n20323 ;
  assign n25971 = n25970 ^ n20023 ^ 1'b0 ;
  assign n25972 = n25969 | n25971 ;
  assign n25973 = n14112 ^ n10892 ^ 1'b0 ;
  assign n25974 = ( n10922 & ~n10982 ) | ( n10922 & n25973 ) | ( ~n10982 & n25973 ) ;
  assign n25975 = n25972 | n25974 ;
  assign n25976 = ( ~n8690 & n15311 ) | ( ~n8690 & n23968 ) | ( n15311 & n23968 ) ;
  assign n25978 = n10727 & n11317 ;
  assign n25977 = ( n13862 & ~n22733 ) | ( n13862 & n23082 ) | ( ~n22733 & n23082 ) ;
  assign n25979 = n25978 ^ n25977 ^ n13279 ;
  assign n25980 = n16416 & n19816 ;
  assign n25981 = n25980 ^ n6502 ^ 1'b0 ;
  assign n25982 = n3875 | n20031 ;
  assign n25983 = n25982 ^ n4581 ^ 1'b0 ;
  assign n25984 = ( n1634 & n3389 ) | ( n1634 & ~n4814 ) | ( n3389 & ~n4814 ) ;
  assign n25985 = n10637 ^ n360 ^ 1'b0 ;
  assign n25986 = n4156 & ~n25985 ;
  assign n25987 = ~n3345 & n8679 ;
  assign n25988 = n25987 ^ n4434 ^ 1'b0 ;
  assign n25989 = ( n6075 & n25986 ) | ( n6075 & n25988 ) | ( n25986 & n25988 ) ;
  assign n25990 = n25988 ^ n22406 ^ n3329 ;
  assign n25992 = n16737 ^ n5850 ^ 1'b0 ;
  assign n25993 = ~n1951 & n25992 ;
  assign n25991 = ~n6934 & n20771 ;
  assign n25994 = n25993 ^ n25991 ^ 1'b0 ;
  assign n25995 = n2407 & n7063 ;
  assign n25996 = ~n19814 & n25995 ;
  assign n25997 = n3766 & n25996 ;
  assign n25998 = n9173 ^ n6888 ^ 1'b0 ;
  assign n25999 = n25998 ^ n7342 ^ n1286 ;
  assign n26000 = n25997 & ~n25999 ;
  assign n26003 = n7732 | n10361 ;
  assign n26001 = n16779 | n19580 ;
  assign n26002 = n10471 & ~n26001 ;
  assign n26004 = n26003 ^ n26002 ^ 1'b0 ;
  assign n26005 = ~n25141 & n26004 ;
  assign n26006 = n7736 | n12839 ;
  assign n26007 = ( ~n15157 & n22590 ) | ( ~n15157 & n26006 ) | ( n22590 & n26006 ) ;
  assign n26008 = n1290 & n21486 ;
  assign n26009 = n26008 ^ n19556 ^ n18235 ;
  assign n26010 = n26009 ^ n19876 ^ 1'b0 ;
  assign n26011 = n8208 | n9551 ;
  assign n26012 = n26011 ^ n6186 ^ n3851 ;
  assign n26013 = n6403 & n9592 ;
  assign n26014 = ~n26012 & n26013 ;
  assign n26015 = ( n8914 & ~n23086 ) | ( n8914 & n25042 ) | ( ~n23086 & n25042 ) ;
  assign n26016 = n6826 ^ n2219 ^ 1'b0 ;
  assign n26017 = n13278 ^ n8161 ^ 1'b0 ;
  assign n26018 = n26017 ^ n22913 ^ 1'b0 ;
  assign n26019 = n10081 | n26018 ;
  assign n26020 = n8755 ^ n4107 ^ 1'b0 ;
  assign n26021 = n4487 & n26020 ;
  assign n26022 = n8309 & n11401 ;
  assign n26023 = ~n26021 & n26022 ;
  assign n26025 = n1260 & ~n12447 ;
  assign n26024 = ~n21647 & n22407 ;
  assign n26026 = n26025 ^ n26024 ^ 1'b0 ;
  assign n26027 = n15971 ^ n4904 ^ 1'b0 ;
  assign n26028 = ( n2326 & ~n10138 ) | ( n2326 & n14689 ) | ( ~n10138 & n14689 ) ;
  assign n26029 = n25415 ^ n16301 ^ 1'b0 ;
  assign n26030 = ~n807 & n8616 ;
  assign n26031 = n12874 | n17415 ;
  assign n26032 = n26031 ^ n6784 ^ 1'b0 ;
  assign n26033 = n26030 | n26032 ;
  assign n26034 = n1069 | n15917 ;
  assign n26035 = n23427 & ~n26034 ;
  assign n26036 = n26035 ^ n4224 ^ 1'b0 ;
  assign n26037 = n6710 ^ n5768 ^ n1284 ;
  assign n26038 = n7804 ^ n7550 ^ 1'b0 ;
  assign n26039 = n9644 | n17294 ;
  assign n26040 = n4561 | n26039 ;
  assign n26041 = n13184 ^ n10117 ^ n5368 ;
  assign n26042 = n6889 ^ n4673 ^ 1'b0 ;
  assign n26043 = n23868 ^ n7466 ^ 1'b0 ;
  assign n26044 = ~n26042 & n26043 ;
  assign n26045 = n9337 & ~n20813 ;
  assign n26046 = n2886 & n26045 ;
  assign n26047 = n24815 ^ n15754 ^ n10311 ;
  assign n26048 = n6039 | n24573 ;
  assign n26049 = n26048 ^ n8662 ^ 1'b0 ;
  assign n26050 = n26049 ^ n19249 ^ n1465 ;
  assign n26051 = ( n15864 & ~n26047 ) | ( n15864 & n26050 ) | ( ~n26047 & n26050 ) ;
  assign n26052 = n24166 ^ n18713 ^ 1'b0 ;
  assign n26053 = n23343 ^ n7958 ^ n2233 ;
  assign n26054 = ( n4835 & n9948 ) | ( n4835 & ~n10211 ) | ( n9948 & ~n10211 ) ;
  assign n26055 = n6795 ^ n1077 ^ 1'b0 ;
  assign n26056 = ~n26054 & n26055 ;
  assign n26057 = n26056 ^ n3376 ^ 1'b0 ;
  assign n26058 = ( n1827 & n21726 ) | ( n1827 & ~n24629 ) | ( n21726 & ~n24629 ) ;
  assign n26059 = ( n2236 & ~n23110 ) | ( n2236 & n23841 ) | ( ~n23110 & n23841 ) ;
  assign n26060 = n7223 & n10053 ;
  assign n26061 = n20936 & n26060 ;
  assign n26062 = n20353 & n23207 ;
  assign n26063 = n13756 & n14360 ;
  assign n26064 = n15410 & n26063 ;
  assign n26065 = n2974 & n13171 ;
  assign n26066 = ~n12435 & n26065 ;
  assign n26067 = n22469 ^ n11967 ^ n1728 ;
  assign n26068 = ( n5810 & ~n26066 ) | ( n5810 & n26067 ) | ( ~n26066 & n26067 ) ;
  assign n26069 = n8186 ^ n4723 ^ 1'b0 ;
  assign n26070 = n11154 & n14947 ;
  assign n26071 = n26070 ^ n4495 ^ 1'b0 ;
  assign n26072 = ~n6764 & n26071 ;
  assign n26073 = ~n8343 & n26072 ;
  assign n26074 = n26073 ^ n8872 ^ 1'b0 ;
  assign n26075 = n15954 ^ n7145 ^ 1'b0 ;
  assign n26076 = ( n6812 & ~n7557 ) | ( n6812 & n26075 ) | ( ~n7557 & n26075 ) ;
  assign n26078 = ( n2204 & ~n5622 ) | ( n2204 & n10189 ) | ( ~n5622 & n10189 ) ;
  assign n26079 = n6267 & n26078 ;
  assign n26080 = n10888 & n26079 ;
  assign n26077 = x88 & n19828 ;
  assign n26081 = n26080 ^ n26077 ^ 1'b0 ;
  assign n26082 = n12768 ^ n1998 ^ 1'b0 ;
  assign n26083 = n23397 & ~n26082 ;
  assign n26084 = ~n1691 & n26083 ;
  assign n26085 = n8685 & n26084 ;
  assign n26086 = n26085 ^ n8390 ^ 1'b0 ;
  assign n26087 = n24046 & ~n26086 ;
  assign n26088 = n26087 ^ n21326 ^ 1'b0 ;
  assign n26090 = x57 | n1948 ;
  assign n26089 = ~n3080 & n22799 ;
  assign n26091 = n26090 ^ n26089 ^ 1'b0 ;
  assign n26096 = n4298 & ~n17433 ;
  assign n26097 = n26096 ^ n8060 ^ 1'b0 ;
  assign n26092 = n1217 & n8780 ;
  assign n26093 = ~n2705 & n26092 ;
  assign n26094 = n4327 & n26093 ;
  assign n26095 = ( n4869 & n6711 ) | ( n4869 & ~n26094 ) | ( n6711 & ~n26094 ) ;
  assign n26098 = n26097 ^ n26095 ^ 1'b0 ;
  assign n26099 = n23455 ^ n1492 ^ 1'b0 ;
  assign n26100 = n26099 ^ n16254 ^ n4105 ;
  assign n26101 = n2164 | n24310 ;
  assign n26102 = n26101 ^ n24211 ^ 1'b0 ;
  assign n26103 = n26102 ^ n22633 ^ n3761 ;
  assign n26104 = n26103 ^ n17326 ^ 1'b0 ;
  assign n26105 = n6831 & n26104 ;
  assign n26106 = n26105 ^ n7627 ^ 1'b0 ;
  assign n26107 = n691 & n2699 ;
  assign n26108 = n17015 & n26107 ;
  assign n26109 = n26108 ^ n22029 ^ 1'b0 ;
  assign n26110 = n17997 ^ n7686 ^ 1'b0 ;
  assign n26111 = ~n8962 & n11620 ;
  assign n26112 = n26111 ^ n11601 ^ 1'b0 ;
  assign n26113 = n24150 ^ n15644 ^ 1'b0 ;
  assign n26116 = ~n3279 & n5506 ;
  assign n26117 = ~n14372 & n26116 ;
  assign n26114 = ~n5554 & n7189 ;
  assign n26115 = n26114 ^ n1907 ^ 1'b0 ;
  assign n26118 = n26117 ^ n26115 ^ n2067 ;
  assign n26119 = n10851 ^ n3106 ^ 1'b0 ;
  assign n26120 = ~n740 & n26119 ;
  assign n26121 = ( n287 & n1170 ) | ( n287 & n26120 ) | ( n1170 & n26120 ) ;
  assign n26122 = n20104 & n20916 ;
  assign n26123 = n6221 ^ n4653 ^ 1'b0 ;
  assign n26124 = ~n19984 & n26123 ;
  assign n26125 = n17353 ^ n1178 ^ 1'b0 ;
  assign n26126 = n26125 ^ n18575 ^ 1'b0 ;
  assign n26129 = n8111 & ~n8112 ;
  assign n26127 = n15448 ^ n7141 ^ 1'b0 ;
  assign n26128 = n26127 ^ n10909 ^ 1'b0 ;
  assign n26130 = n26129 ^ n26128 ^ n9475 ;
  assign n26131 = n19101 ^ n8732 ^ 1'b0 ;
  assign n26132 = n16927 ^ n10445 ^ n6110 ;
  assign n26133 = n26132 ^ n7071 ^ n4763 ;
  assign n26134 = n26133 ^ n26132 ^ n14670 ;
  assign n26135 = n9437 & n11013 ;
  assign n26136 = ~n16449 & n26135 ;
  assign n26137 = ~n26134 & n26136 ;
  assign n26138 = n26137 ^ n8810 ^ 1'b0 ;
  assign n26139 = n26131 & ~n26138 ;
  assign n26140 = n1386 & ~n6881 ;
  assign n26141 = n18273 ^ n3088 ^ 1'b0 ;
  assign n26142 = x159 & n4654 ;
  assign n26143 = n7552 & n26142 ;
  assign n26144 = ~n26141 & n26143 ;
  assign n26145 = ~n17826 & n26144 ;
  assign n26146 = n12912 ^ n10969 ^ 1'b0 ;
  assign n26147 = ~n8505 & n26146 ;
  assign n26148 = n26147 ^ n9030 ^ x246 ;
  assign n26150 = n15058 & ~n16755 ;
  assign n26151 = n26150 ^ n7496 ^ 1'b0 ;
  assign n26152 = ~n814 & n26151 ;
  assign n26149 = ~n10672 & n25321 ;
  assign n26153 = n26152 ^ n26149 ^ 1'b0 ;
  assign n26154 = n11854 ^ n11176 ^ 1'b0 ;
  assign n26155 = n26153 & ~n26154 ;
  assign n26161 = ( n1203 & n2809 ) | ( n1203 & n7379 ) | ( n2809 & n7379 ) ;
  assign n26156 = n16205 ^ n310 ^ 1'b0 ;
  assign n26157 = n343 | n5557 ;
  assign n26158 = n26157 ^ n7231 ^ 1'b0 ;
  assign n26159 = n23443 & n26158 ;
  assign n26160 = ~n26156 & n26159 ;
  assign n26162 = n26161 ^ n26160 ^ n262 ;
  assign n26163 = n4768 & n26162 ;
  assign n26164 = n8049 & n15526 ;
  assign n26165 = n26164 ^ n12617 ^ 1'b0 ;
  assign n26166 = ~n2026 & n26165 ;
  assign n26167 = ~n5379 & n5982 ;
  assign n26168 = n26167 ^ n25201 ^ 1'b0 ;
  assign n26169 = ~n5981 & n19171 ;
  assign n26170 = ( ~n6711 & n15157 ) | ( ~n6711 & n24267 ) | ( n15157 & n24267 ) ;
  assign n26171 = n10593 ^ n2865 ^ 1'b0 ;
  assign n26172 = ~n4495 & n26171 ;
  assign n26173 = n26172 ^ n11367 ^ 1'b0 ;
  assign n26174 = n26173 ^ n19101 ^ n14270 ;
  assign n26175 = n11377 ^ n567 ^ x57 ;
  assign n26176 = n1104 ^ x212 ^ 1'b0 ;
  assign n26177 = x200 & n26176 ;
  assign n26178 = ~n6908 & n26177 ;
  assign n26179 = n26175 & n26178 ;
  assign n26180 = n1413 & n9024 ;
  assign n26181 = ~n9370 & n20584 ;
  assign n26182 = n26181 ^ n4705 ^ 1'b0 ;
  assign n26183 = n6636 | n26182 ;
  assign n26184 = n5963 & ~n26183 ;
  assign n26185 = n13738 ^ n2064 ^ 1'b0 ;
  assign n26186 = n679 & ~n26185 ;
  assign n26187 = n3153 & ~n26186 ;
  assign n26188 = n8490 | n23860 ;
  assign n26189 = n6597 & ~n18617 ;
  assign n26190 = n7135 ^ n6816 ^ 1'b0 ;
  assign n26191 = n2643 & n26190 ;
  assign n26192 = n26191 ^ n19742 ^ 1'b0 ;
  assign n26193 = ~n3794 & n26192 ;
  assign n26194 = n26193 ^ n14363 ^ 1'b0 ;
  assign n26195 = n26189 | n26194 ;
  assign n26196 = n279 & ~n4696 ;
  assign n26197 = ~n11928 & n26196 ;
  assign n26198 = ~n16066 & n19739 ;
  assign n26199 = n26198 ^ n20475 ^ 1'b0 ;
  assign n26201 = n6886 & ~n6897 ;
  assign n26200 = n9834 ^ n1663 ^ 1'b0 ;
  assign n26202 = n26201 ^ n26200 ^ n21835 ;
  assign n26203 = n11722 ^ n11415 ^ 1'b0 ;
  assign n26204 = n18518 ^ n1636 ^ 1'b0 ;
  assign n26205 = n4471 | n10928 ;
  assign n26206 = n26205 ^ n15224 ^ 1'b0 ;
  assign n26207 = n20323 ^ n8732 ^ 1'b0 ;
  assign n26208 = ( n14186 & n19692 ) | ( n14186 & ~n26207 ) | ( n19692 & ~n26207 ) ;
  assign n26209 = n26206 & n26208 ;
  assign n26210 = n26209 ^ n11027 ^ 1'b0 ;
  assign n26211 = n26210 ^ n14901 ^ 1'b0 ;
  assign n26212 = ~n8465 & n26211 ;
  assign n26213 = n26099 ^ n20473 ^ 1'b0 ;
  assign n26214 = n13134 & ~n26213 ;
  assign n26215 = ~n9244 & n13766 ;
  assign n26216 = n26215 ^ n17252 ^ 1'b0 ;
  assign n26217 = n26216 ^ n14529 ^ n12700 ;
  assign n26219 = ~n13873 & n17716 ;
  assign n26218 = n7012 & ~n7915 ;
  assign n26220 = n26219 ^ n26218 ^ n3335 ;
  assign n26221 = n26220 ^ n23019 ^ n5740 ;
  assign n26222 = n13735 & n22172 ;
  assign n26223 = ~n4153 & n26222 ;
  assign n26224 = n7764 & n20927 ;
  assign n26225 = n10774 & n12836 ;
  assign n26226 = n18608 & n26225 ;
  assign n26227 = n3259 & n21485 ;
  assign n26228 = n26227 ^ n24914 ^ n413 ;
  assign n26229 = ~n7497 & n26228 ;
  assign n26230 = n16551 | n21037 ;
  assign n26231 = n1074 & ~n1759 ;
  assign n26232 = n26231 ^ n7657 ^ 1'b0 ;
  assign n26233 = n25489 ^ n1444 ^ 1'b0 ;
  assign n26234 = n14553 | n26233 ;
  assign n26235 = n26234 ^ n8067 ^ 1'b0 ;
  assign n26236 = n8149 ^ n5215 ^ 1'b0 ;
  assign n26237 = ( ~n26232 & n26235 ) | ( ~n26232 & n26236 ) | ( n26235 & n26236 ) ;
  assign n26238 = n5771 & n8227 ;
  assign n26239 = ( n8158 & n23994 ) | ( n8158 & n26238 ) | ( n23994 & n26238 ) ;
  assign n26241 = n15854 ^ n10989 ^ 1'b0 ;
  assign n26240 = n10310 & ~n14965 ;
  assign n26242 = n26241 ^ n26240 ^ 1'b0 ;
  assign n26243 = n18861 & n24919 ;
  assign n26244 = n17033 & ~n19721 ;
  assign n26245 = n14382 | n26244 ;
  assign n26246 = n1639 | n26245 ;
  assign n26247 = n24383 ^ n15747 ^ 1'b0 ;
  assign n26251 = n8365 ^ n1590 ^ 1'b0 ;
  assign n26252 = n4134 | n26251 ;
  assign n26253 = n8302 ^ n1407 ^ 1'b0 ;
  assign n26254 = ~n26252 & n26253 ;
  assign n26255 = n26254 ^ n8772 ^ 1'b0 ;
  assign n26256 = x225 & n26255 ;
  assign n26248 = n3029 & n22766 ;
  assign n26249 = n21413 ^ n15703 ^ n3887 ;
  assign n26250 = n26248 & n26249 ;
  assign n26257 = n26256 ^ n26250 ^ n16806 ;
  assign n26258 = n2489 ^ n1166 ^ 1'b0 ;
  assign n26259 = n3568 | n20389 ;
  assign n26260 = n12815 | n26259 ;
  assign n26261 = ( n1040 & n1950 ) | ( n1040 & ~n5914 ) | ( n1950 & ~n5914 ) ;
  assign n26262 = ( n6352 & ~n21765 ) | ( n6352 & n26261 ) | ( ~n21765 & n26261 ) ;
  assign n26263 = ( ~n525 & n5042 ) | ( ~n525 & n10685 ) | ( n5042 & n10685 ) ;
  assign n26264 = ( ~n19680 & n26262 ) | ( ~n19680 & n26263 ) | ( n26262 & n26263 ) ;
  assign n26265 = n5432 & ~n14955 ;
  assign n26266 = ~n4490 & n11926 ;
  assign n26267 = n8453 & n26266 ;
  assign n26269 = n9478 ^ n7460 ^ n6944 ;
  assign n26270 = ~n9054 & n26269 ;
  assign n26271 = ~n22854 & n26270 ;
  assign n26268 = n23057 ^ n21396 ^ 1'b0 ;
  assign n26272 = n26271 ^ n26268 ^ n4997 ;
  assign n26273 = n9005 ^ n7801 ^ 1'b0 ;
  assign n26274 = n9484 | n26273 ;
  assign n26275 = n5078 | n26274 ;
  assign n26276 = n10185 ^ n888 ^ 1'b0 ;
  assign n26277 = ( ~n22483 & n24083 ) | ( ~n22483 & n26276 ) | ( n24083 & n26276 ) ;
  assign n26278 = n10296 ^ n3304 ^ 1'b0 ;
  assign n26279 = ~n22284 & n26278 ;
  assign n26280 = n9038 & ~n11390 ;
  assign n26281 = n18008 ^ n10358 ^ n4398 ;
  assign n26282 = n26281 ^ n20094 ^ 1'b0 ;
  assign n26283 = n26280 | n26282 ;
  assign n26284 = n25710 ^ n17346 ^ n3259 ;
  assign n26285 = n7775 | n12303 ;
  assign n26286 = n26284 | n26285 ;
  assign n26287 = n17300 ^ n8302 ^ n2818 ;
  assign n26288 = n19278 ^ n15876 ^ 1'b0 ;
  assign n26289 = n8539 | n26288 ;
  assign n26290 = ( ~n6450 & n26287 ) | ( ~n6450 & n26289 ) | ( n26287 & n26289 ) ;
  assign n26291 = n11612 ^ n3466 ^ 1'b0 ;
  assign n26292 = n5326 ^ n2572 ^ 1'b0 ;
  assign n26293 = n14386 | n26292 ;
  assign n26294 = n19916 | n26293 ;
  assign n26295 = n26294 ^ n22287 ^ 1'b0 ;
  assign n26296 = n15074 ^ n3996 ^ n1150 ;
  assign n26297 = n19726 | n26296 ;
  assign n26298 = n26297 ^ n7044 ^ 1'b0 ;
  assign n26299 = ~n21029 & n26298 ;
  assign n26300 = n26295 & n26299 ;
  assign n26301 = n21027 ^ n16113 ^ 1'b0 ;
  assign n26302 = n26301 ^ n1222 ^ 1'b0 ;
  assign n26306 = n13423 & ~n18560 ;
  assign n26305 = ~n17888 & n20797 ;
  assign n26307 = n26306 ^ n26305 ^ 1'b0 ;
  assign n26303 = n366 & ~n15677 ;
  assign n26304 = ~n7959 & n26303 ;
  assign n26308 = n26307 ^ n26304 ^ 1'b0 ;
  assign n26309 = ~n1082 & n17167 ;
  assign n26310 = n5525 & n8608 ;
  assign n26311 = ~n13273 & n26310 ;
  assign n26312 = n26311 ^ n9562 ^ n6710 ;
  assign n26313 = n1675 & ~n26312 ;
  assign n26314 = ~n26309 & n26313 ;
  assign n26315 = n5358 & n16811 ;
  assign n26316 = n26315 ^ n8563 ^ 1'b0 ;
  assign n26317 = n14171 ^ n807 ^ 1'b0 ;
  assign n26318 = n6052 | n16653 ;
  assign n26319 = n26318 ^ n1603 ^ 1'b0 ;
  assign n26320 = ( n26316 & ~n26317 ) | ( n26316 & n26319 ) | ( ~n26317 & n26319 ) ;
  assign n26321 = ~n4158 & n8969 ;
  assign n26322 = n26321 ^ n6048 ^ 1'b0 ;
  assign n26323 = ( n2799 & ~n11933 ) | ( n2799 & n26322 ) | ( ~n11933 & n26322 ) ;
  assign n26324 = n12102 & ~n14304 ;
  assign n26325 = n307 | n11985 ;
  assign n26326 = ~n4419 & n14941 ;
  assign n26327 = n26325 & n26326 ;
  assign n26329 = ~n2838 & n10067 ;
  assign n26328 = ~n3756 & n4977 ;
  assign n26330 = n26329 ^ n26328 ^ 1'b0 ;
  assign n26331 = n18190 & n19525 ;
  assign n26332 = ~n26330 & n26331 ;
  assign n26333 = ~n17029 & n25758 ;
  assign n26334 = n20067 & n26333 ;
  assign n26335 = n26334 ^ n20626 ^ 1'b0 ;
  assign n26336 = n25647 ^ n20679 ^ n6051 ;
  assign n26337 = ~n16806 & n26336 ;
  assign n26338 = n22214 ^ n4078 ^ 1'b0 ;
  assign n26339 = ~n3165 & n7824 ;
  assign n26340 = n10918 ^ n2024 ^ 1'b0 ;
  assign n26341 = n26340 ^ n9764 ^ 1'b0 ;
  assign n26342 = n6111 & ~n25080 ;
  assign n26343 = n1107 | n5214 ;
  assign n26344 = n7084 | n26343 ;
  assign n26345 = n26344 ^ n13156 ^ 1'b0 ;
  assign n26347 = n7329 & ~n12666 ;
  assign n26348 = n6638 & n26347 ;
  assign n26349 = n26348 ^ n1274 ^ 1'b0 ;
  assign n26346 = n24875 ^ n2746 ^ 1'b0 ;
  assign n26350 = n26349 ^ n26346 ^ 1'b0 ;
  assign n26353 = n13003 ^ n10348 ^ 1'b0 ;
  assign n26354 = n26353 ^ n8722 ^ x25 ;
  assign n26351 = n3160 & n25338 ;
  assign n26352 = n9165 & ~n26351 ;
  assign n26355 = n26354 ^ n26352 ^ n6449 ;
  assign n26356 = n13111 ^ n11402 ^ 1'b0 ;
  assign n26357 = ~n10606 & n26356 ;
  assign n26358 = ~n9757 & n26357 ;
  assign n26359 = n22728 & n26358 ;
  assign n26360 = ~n21306 & n26359 ;
  assign n26361 = ~n14855 & n18420 ;
  assign n26362 = n21356 ^ n15484 ^ 1'b0 ;
  assign n26363 = n8764 & n26362 ;
  assign n26364 = n22291 ^ n881 ^ 1'b0 ;
  assign n26365 = ~n3990 & n26364 ;
  assign n26366 = n26365 ^ n2367 ^ 1'b0 ;
  assign n26367 = ~n19698 & n26366 ;
  assign n26368 = ( x93 & x202 ) | ( x93 & n329 ) | ( x202 & n329 ) ;
  assign n26369 = n6686 & n26368 ;
  assign n26370 = n25203 ^ n9714 ^ n4215 ;
  assign n26371 = n26370 ^ n20815 ^ 1'b0 ;
  assign n26372 = n26369 & ~n26371 ;
  assign n26373 = n23874 & ~n24808 ;
  assign n26374 = ~n6786 & n26373 ;
  assign n26375 = n26372 | n26374 ;
  assign n26376 = n3716 ^ x26 ^ 1'b0 ;
  assign n26377 = ( n1152 & n17971 ) | ( n1152 & ~n26376 ) | ( n17971 & ~n26376 ) ;
  assign n26378 = n10891 & ~n24041 ;
  assign n26379 = n4995 ^ n922 ^ 1'b0 ;
  assign n26380 = n26379 ^ n7923 ^ 1'b0 ;
  assign n26382 = n10708 & n14753 ;
  assign n26383 = n26382 ^ n9990 ^ 1'b0 ;
  assign n26381 = ( n7151 & ~n10909 ) | ( n7151 & n15707 ) | ( ~n10909 & n15707 ) ;
  assign n26384 = n26383 ^ n26381 ^ n3581 ;
  assign n26385 = n26384 ^ n22990 ^ n18409 ;
  assign n26386 = n19757 ^ n8130 ^ n1858 ;
  assign n26387 = ~n20158 & n26386 ;
  assign n26388 = x164 & ~n22056 ;
  assign n26389 = ~n22898 & n26388 ;
  assign n26390 = n26389 ^ n1228 ^ 1'b0 ;
  assign n26391 = n20950 ^ n5448 ^ 1'b0 ;
  assign n26392 = n13263 | n26391 ;
  assign n26393 = n5751 & n12131 ;
  assign n26394 = n26393 ^ n15350 ^ 1'b0 ;
  assign n26395 = n15575 ^ n11401 ^ 1'b0 ;
  assign n26396 = n12872 & ~n26395 ;
  assign n26397 = n24605 ^ n11527 ^ 1'b0 ;
  assign n26399 = n12550 | n14294 ;
  assign n26398 = n13460 & ~n14943 ;
  assign n26400 = n26399 ^ n26398 ^ 1'b0 ;
  assign n26401 = n26400 ^ n22482 ^ n15557 ;
  assign n26402 = n19188 ^ n6543 ^ n635 ;
  assign n26403 = n4041 ^ n2660 ^ 1'b0 ;
  assign n26404 = n10564 & ~n26403 ;
  assign n26405 = n26404 ^ n16638 ^ n14770 ;
  assign n26406 = n3439 & ~n20840 ;
  assign n26408 = n13625 ^ n1985 ^ n1465 ;
  assign n26407 = n5138 & n14128 ;
  assign n26409 = n26408 ^ n26407 ^ n6018 ;
  assign n26410 = n21035 ^ n3331 ^ 1'b0 ;
  assign n26411 = ( n13527 & n18337 ) | ( n13527 & n26410 ) | ( n18337 & n26410 ) ;
  assign n26412 = n2691 & n15320 ;
  assign n26413 = n10778 ^ n6011 ^ 1'b0 ;
  assign n26414 = n11750 & n23030 ;
  assign n26415 = n26413 & n26414 ;
  assign n26416 = n4996 | n26415 ;
  assign n26417 = n26412 & ~n26416 ;
  assign n26418 = n3881 & ~n23686 ;
  assign n26419 = ~n23678 & n26418 ;
  assign n26420 = n22680 ^ n18359 ^ 1'b0 ;
  assign n26421 = n3119 | n26420 ;
  assign n26422 = ~n5916 & n9438 ;
  assign n26423 = ~n797 & n26422 ;
  assign n26424 = n18091 & ~n18997 ;
  assign n26425 = n26424 ^ n4569 ^ 1'b0 ;
  assign n26426 = n2939 & ~n6395 ;
  assign n26427 = ~x69 & n26426 ;
  assign n26428 = n2510 ^ x120 ^ 1'b0 ;
  assign n26429 = n21493 ^ n18822 ^ n496 ;
  assign n26430 = ~n8181 & n19136 ;
  assign n26431 = ( n1729 & ~n11486 ) | ( n1729 & n15361 ) | ( ~n11486 & n15361 ) ;
  assign n26432 = n26431 ^ n25864 ^ 1'b0 ;
  assign n26433 = ( n6063 & ~n17405 ) | ( n6063 & n19234 ) | ( ~n17405 & n19234 ) ;
  assign n26434 = n489 | n6727 ;
  assign n26437 = n22257 ^ n7602 ^ 1'b0 ;
  assign n26435 = ( x211 & n14892 ) | ( x211 & n16341 ) | ( n14892 & n16341 ) ;
  assign n26436 = n4498 & ~n26435 ;
  assign n26438 = n26437 ^ n26436 ^ 1'b0 ;
  assign n26439 = ~n4234 & n26438 ;
  assign n26440 = n18573 & n26439 ;
  assign n26441 = n16328 | n20819 ;
  assign n26442 = n26441 ^ n2688 ^ 1'b0 ;
  assign n26443 = ~n18106 & n26442 ;
  assign n26444 = n933 | n8941 ;
  assign n26445 = n26444 ^ n1939 ^ 1'b0 ;
  assign n26446 = n11668 & n26445 ;
  assign n26447 = ~n4067 & n26446 ;
  assign n26448 = n26447 ^ n25063 ^ 1'b0 ;
  assign n26449 = ~x234 & n1175 ;
  assign n26450 = n26449 ^ n3259 ^ 1'b0 ;
  assign n26451 = n1666 & n26450 ;
  assign n26452 = n21264 ^ n18483 ^ 1'b0 ;
  assign n26453 = n26452 ^ n21573 ^ n4588 ;
  assign n26454 = n11251 & n24378 ;
  assign n26455 = ~n10064 & n26454 ;
  assign n26456 = n12291 & n12896 ;
  assign n26457 = n26456 ^ n11441 ^ 1'b0 ;
  assign n26458 = ( ~n6534 & n12525 ) | ( ~n6534 & n26457 ) | ( n12525 & n26457 ) ;
  assign n26459 = n26458 ^ n16371 ^ 1'b0 ;
  assign n26460 = n8189 | n26459 ;
  assign n26461 = n5229 ^ x43 ^ 1'b0 ;
  assign n26462 = n6853 & n26461 ;
  assign n26463 = n12498 ^ n9201 ^ n7362 ;
  assign n26464 = n15815 & ~n26463 ;
  assign n26465 = ~n12968 & n26464 ;
  assign n26466 = n10980 & ~n14318 ;
  assign n26467 = n12392 ^ n9532 ^ 1'b0 ;
  assign n26468 = n26286 & n26467 ;
  assign n26469 = n22783 ^ n7131 ^ 1'b0 ;
  assign n26470 = n8357 ^ n1236 ^ 1'b0 ;
  assign n26471 = ~n4378 & n26470 ;
  assign n26472 = n7976 ^ n3865 ^ 1'b0 ;
  assign n26473 = n8930 | n26472 ;
  assign n26474 = n2661 | n26473 ;
  assign n26475 = n26474 ^ n8542 ^ 1'b0 ;
  assign n26476 = n24150 ^ n14930 ^ n1937 ;
  assign n26477 = n20466 ^ n19672 ^ 1'b0 ;
  assign n26478 = n2938 & ~n26477 ;
  assign n26479 = n17654 ^ n17052 ^ n5467 ;
  assign n26480 = ( n843 & n8045 ) | ( n843 & ~n20785 ) | ( n8045 & ~n20785 ) ;
  assign n26481 = n3578 & n26480 ;
  assign n26482 = ~n26479 & n26481 ;
  assign n26483 = n9186 & n10770 ;
  assign n26484 = n26483 ^ n856 ^ 1'b0 ;
  assign n26485 = n16099 | n26484 ;
  assign n26486 = n6410 & n11232 ;
  assign n26487 = n26486 ^ n20610 ^ 1'b0 ;
  assign n26488 = ~n8345 & n13717 ;
  assign n26489 = n12190 & n26488 ;
  assign n26490 = x119 & n3155 ;
  assign n26491 = n13450 & n26490 ;
  assign n26492 = n2744 & ~n24298 ;
  assign n26493 = ~n14495 & n26492 ;
  assign n26494 = n15557 & n22167 ;
  assign n26495 = n1185 | n2491 ;
  assign n26496 = n26495 ^ n5710 ^ n3191 ;
  assign n26497 = n26496 ^ n19242 ^ n12408 ;
  assign n26498 = n26497 ^ n24643 ^ 1'b0 ;
  assign n26499 = n10621 & n26498 ;
  assign n26500 = ~n10416 & n26499 ;
  assign n26501 = n26500 ^ n15431 ^ 1'b0 ;
  assign n26502 = ( n3244 & n12911 ) | ( n3244 & n13226 ) | ( n12911 & n13226 ) ;
  assign n26503 = ~n1935 & n26502 ;
  assign n26504 = n26503 ^ n24582 ^ 1'b0 ;
  assign n26505 = ~n2454 & n26504 ;
  assign n26506 = ~n1465 & n10900 ;
  assign n26507 = n26506 ^ n10088 ^ 1'b0 ;
  assign n26509 = n6283 ^ n4572 ^ n4101 ;
  assign n26508 = n2762 | n6791 ;
  assign n26510 = n26509 ^ n26508 ^ 1'b0 ;
  assign n26511 = n6098 ^ n2504 ^ 1'b0 ;
  assign n26512 = n538 | n26511 ;
  assign n26513 = ( n17596 & n26510 ) | ( n17596 & n26512 ) | ( n26510 & n26512 ) ;
  assign n26514 = n6995 ^ n3576 ^ 1'b0 ;
  assign n26515 = ~n3939 & n16605 ;
  assign n26516 = n1705 & n13172 ;
  assign n26517 = ~n9276 & n26516 ;
  assign n26518 = n26517 ^ n3547 ^ 1'b0 ;
  assign n26519 = ~n5666 & n7346 ;
  assign n26520 = n1257 & n26519 ;
  assign n26521 = n20632 | n26520 ;
  assign n26522 = n26521 ^ n25447 ^ 1'b0 ;
  assign n26523 = ( n26515 & n26518 ) | ( n26515 & ~n26522 ) | ( n26518 & ~n26522 ) ;
  assign n26524 = ~n5297 & n24088 ;
  assign n26525 = n15033 | n22236 ;
  assign n26526 = n9439 & ~n26525 ;
  assign n26527 = ( n1142 & n8192 ) | ( n1142 & n8900 ) | ( n8192 & n8900 ) ;
  assign n26528 = ( n639 & ~n9083 ) | ( n639 & n26527 ) | ( ~n9083 & n26527 ) ;
  assign n26529 = n23781 ^ n8193 ^ n6857 ;
  assign n26530 = n2781 | n5377 ;
  assign n26531 = n3262 & ~n26530 ;
  assign n26532 = n20252 ^ n9443 ^ 1'b0 ;
  assign n26533 = ~n26531 & n26532 ;
  assign n26534 = n4705 & n26533 ;
  assign n26535 = ~n13389 & n26534 ;
  assign n26536 = n18156 ^ n13189 ^ n2793 ;
  assign n26537 = n26536 ^ n4675 ^ n4153 ;
  assign n26538 = n14542 ^ n1534 ^ 1'b0 ;
  assign n26540 = n15972 ^ n8882 ^ n5366 ;
  assign n26541 = n26540 ^ n16017 ^ 1'b0 ;
  assign n26539 = n2050 | n16653 ;
  assign n26542 = n26541 ^ n26539 ^ 1'b0 ;
  assign n26543 = n2996 & ~n3080 ;
  assign n26544 = n24039 & n26543 ;
  assign n26551 = n15542 ^ n2616 ^ n2106 ;
  assign n26547 = ~x90 & n25109 ;
  assign n26548 = n26547 ^ n668 ^ 1'b0 ;
  assign n26549 = ~n4854 & n26548 ;
  assign n26550 = ~n14758 & n26549 ;
  assign n26545 = n2836 & n13701 ;
  assign n26546 = n9041 | n26545 ;
  assign n26552 = n26551 ^ n26550 ^ n26546 ;
  assign n26553 = n17889 ^ n11532 ^ 1'b0 ;
  assign n26554 = ~n3112 & n26553 ;
  assign n26555 = n7462 ^ n4920 ^ 1'b0 ;
  assign n26556 = n10543 ^ x172 ^ 1'b0 ;
  assign n26557 = n26403 & n26556 ;
  assign n26558 = ( n3322 & ~n26555 ) | ( n3322 & n26557 ) | ( ~n26555 & n26557 ) ;
  assign n26559 = ~n26554 & n26558 ;
  assign n26560 = n3447 ^ n2844 ^ 1'b0 ;
  assign n26561 = n5752 | n26560 ;
  assign n26562 = n26561 ^ n22165 ^ n7427 ;
  assign n26563 = n10889 & n12370 ;
  assign n26564 = ~n3952 & n26563 ;
  assign n26565 = n1403 & ~n22219 ;
  assign n26572 = n3097 ^ n1650 ^ 1'b0 ;
  assign n26568 = n7494 | n9688 ;
  assign n26569 = n16656 | n26568 ;
  assign n26566 = n1658 | n3471 ;
  assign n26567 = n2764 | n26566 ;
  assign n26570 = n26569 ^ n26567 ^ 1'b0 ;
  assign n26571 = n6917 & n26570 ;
  assign n26573 = n26572 ^ n26571 ^ 1'b0 ;
  assign n26574 = n14327 | n15109 ;
  assign n26575 = n440 & ~n26574 ;
  assign n26578 = ~n10949 & n22073 ;
  assign n26576 = n13511 | n16643 ;
  assign n26577 = n26576 ^ n24035 ^ 1'b0 ;
  assign n26579 = n26578 ^ n26577 ^ 1'b0 ;
  assign n26580 = n20780 | n26579 ;
  assign n26582 = n4301 & ~n14786 ;
  assign n26583 = n5188 & n26582 ;
  assign n26584 = ~n19692 & n26583 ;
  assign n26581 = n11842 & ~n13725 ;
  assign n26585 = n26584 ^ n26581 ^ 1'b0 ;
  assign n26594 = n2275 | n22544 ;
  assign n26595 = n26594 ^ n4703 ^ 1'b0 ;
  assign n26586 = n11032 ^ n5417 ^ 1'b0 ;
  assign n26587 = n6251 & n26586 ;
  assign n26588 = n26587 ^ n2800 ^ 1'b0 ;
  assign n26590 = n7180 ^ n3518 ^ 1'b0 ;
  assign n26589 = n18176 & n19112 ;
  assign n26591 = n26590 ^ n26589 ^ 1'b0 ;
  assign n26592 = n26591 ^ n17472 ^ 1'b0 ;
  assign n26593 = n26588 & ~n26592 ;
  assign n26596 = n26595 ^ n26593 ^ 1'b0 ;
  assign n26597 = n12361 & n14137 ;
  assign n26598 = n23300 & n26597 ;
  assign n26599 = n10221 & n15128 ;
  assign n26600 = ~n25090 & n26599 ;
  assign n26601 = ( n5179 & ~n15881 ) | ( n5179 & n16759 ) | ( ~n15881 & n16759 ) ;
  assign n26602 = ( n1757 & ~n7618 ) | ( n1757 & n18728 ) | ( ~n7618 & n18728 ) ;
  assign n26603 = n3138 | n26602 ;
  assign n26604 = n26603 ^ n12508 ^ 1'b0 ;
  assign n26605 = ( n1804 & ~n8321 ) | ( n1804 & n26604 ) | ( ~n8321 & n26604 ) ;
  assign n26611 = n9008 ^ n4456 ^ n3133 ;
  assign n26612 = n8681 & ~n26611 ;
  assign n26613 = ( x202 & n6706 ) | ( x202 & ~n26612 ) | ( n6706 & ~n26612 ) ;
  assign n26608 = n10134 ^ n7696 ^ 1'b0 ;
  assign n26609 = n13996 & ~n26608 ;
  assign n26610 = n26609 ^ n13789 ^ 1'b0 ;
  assign n26614 = n26613 ^ n26610 ^ 1'b0 ;
  assign n26606 = n7307 | n17422 ;
  assign n26607 = n1598 & n26606 ;
  assign n26615 = n26614 ^ n26607 ^ 1'b0 ;
  assign n26616 = n13833 ^ n8865 ^ 1'b0 ;
  assign n26617 = ~n19425 & n26616 ;
  assign n26618 = ( n4187 & n11105 ) | ( n4187 & n13135 ) | ( n11105 & n13135 ) ;
  assign n26619 = ( x47 & n7265 ) | ( x47 & n13000 ) | ( n7265 & n13000 ) ;
  assign n26620 = ( n15929 & ~n26618 ) | ( n15929 & n26619 ) | ( ~n26618 & n26619 ) ;
  assign n26621 = ( n405 & ~n4484 ) | ( n405 & n5233 ) | ( ~n4484 & n5233 ) ;
  assign n26622 = n26621 ^ n18945 ^ 1'b0 ;
  assign n26623 = ( n4097 & ~n7051 ) | ( n4097 & n14448 ) | ( ~n7051 & n14448 ) ;
  assign n26624 = n18516 & n22335 ;
  assign n26625 = n3014 & n26624 ;
  assign n26626 = n7395 ^ n5591 ^ n4437 ;
  assign n26627 = n2811 & n6611 ;
  assign n26628 = n26626 & n26627 ;
  assign n26629 = ( ~n23024 & n26625 ) | ( ~n23024 & n26628 ) | ( n26625 & n26628 ) ;
  assign n26630 = n5810 ^ n891 ^ 1'b0 ;
  assign n26631 = n21782 | n26630 ;
  assign n26632 = n26631 ^ n9004 ^ 1'b0 ;
  assign n26633 = n22174 ^ n2277 ^ 1'b0 ;
  assign n26634 = n24781 ^ n16241 ^ n9198 ;
  assign n26635 = n1322 & ~n26495 ;
  assign n26636 = n13086 & ~n26635 ;
  assign n26637 = ( n8357 & n8551 ) | ( n8357 & n15076 ) | ( n8551 & n15076 ) ;
  assign n26638 = n26637 ^ n2341 ^ 1'b0 ;
  assign n26639 = n11664 & n20426 ;
  assign n26640 = ~n22696 & n26639 ;
  assign n26641 = n18726 & n26640 ;
  assign n26642 = n26638 | n26641 ;
  assign n26643 = n11546 | n26642 ;
  assign n26644 = ~n26636 & n26643 ;
  assign n26645 = n26644 ^ x163 ^ 1'b0 ;
  assign n26646 = n4777 ^ n3786 ^ 1'b0 ;
  assign n26647 = n26646 ^ n7624 ^ n3755 ;
  assign n26648 = n11567 ^ n7326 ^ 1'b0 ;
  assign n26649 = n26648 ^ n25400 ^ n20895 ;
  assign n26650 = n16911 | n18321 ;
  assign n26653 = n4672 | n7132 ;
  assign n26654 = n26653 ^ n4214 ^ 1'b0 ;
  assign n26655 = ~n3848 & n4707 ;
  assign n26656 = n26654 & ~n26655 ;
  assign n26657 = n576 & n26656 ;
  assign n26651 = n9846 ^ n9180 ^ 1'b0 ;
  assign n26652 = n22309 & n26651 ;
  assign n26658 = n26657 ^ n26652 ^ n1465 ;
  assign n26659 = n26658 ^ n16290 ^ 1'b0 ;
  assign n26662 = n11296 ^ n410 ^ 1'b0 ;
  assign n26660 = n16643 & ~n17894 ;
  assign n26661 = ~n19287 & n26660 ;
  assign n26663 = n26662 ^ n26661 ^ n16060 ;
  assign n26664 = n9141 & ~n9783 ;
  assign n26665 = n26664 ^ n11521 ^ 1'b0 ;
  assign n26666 = n26665 ^ n17387 ^ 1'b0 ;
  assign n26667 = ( n21404 & n24143 ) | ( n21404 & n26666 ) | ( n24143 & n26666 ) ;
  assign n26668 = ( n13791 & n15546 ) | ( n13791 & n22888 ) | ( n15546 & n22888 ) ;
  assign n26669 = n26668 ^ n23037 ^ n20067 ;
  assign n26670 = n14121 | n19640 ;
  assign n26671 = n14438 ^ n5186 ^ 1'b0 ;
  assign n26672 = n6410 & ~n17556 ;
  assign n26673 = n2487 | n26672 ;
  assign n26675 = ( n9235 & n11997 ) | ( n9235 & ~n16714 ) | ( n11997 & ~n16714 ) ;
  assign n26674 = ( n5712 & n19540 ) | ( n5712 & n24798 ) | ( n19540 & n24798 ) ;
  assign n26676 = n26675 ^ n26674 ^ n16743 ;
  assign n26677 = ( ~n442 & n7049 ) | ( ~n442 & n13712 ) | ( n7049 & n13712 ) ;
  assign n26678 = n26677 ^ n11447 ^ 1'b0 ;
  assign n26679 = n18807 & n22916 ;
  assign n26680 = n14107 ^ n8001 ^ 1'b0 ;
  assign n26681 = ~n26164 & n26680 ;
  assign n26682 = n5833 & n19068 ;
  assign n26683 = n1129 & ~n4578 ;
  assign n26684 = n15524 | n26683 ;
  assign n26685 = n10026 ^ n4570 ^ n610 ;
  assign n26686 = ( n574 & n8071 ) | ( n574 & n15954 ) | ( n8071 & n15954 ) ;
  assign n26687 = n26686 ^ n20572 ^ 1'b0 ;
  assign n26688 = n15746 | n26687 ;
  assign n26689 = ~n1896 & n21664 ;
  assign n26690 = n26689 ^ n3972 ^ 1'b0 ;
  assign n26691 = n2816 & n12136 ;
  assign n26692 = n26691 ^ n2532 ^ 1'b0 ;
  assign n26693 = n26692 ^ x199 ^ 1'b0 ;
  assign n26694 = n974 & ~n4726 ;
  assign n26695 = n5443 & n26694 ;
  assign n26696 = n8502 & ~n26695 ;
  assign n26697 = ( n5023 & n25978 ) | ( n5023 & ~n26696 ) | ( n25978 & ~n26696 ) ;
  assign n26698 = n26693 & ~n26697 ;
  assign n26699 = n7447 & n26698 ;
  assign n26700 = n11636 & ~n13211 ;
  assign n26701 = n26700 ^ n3342 ^ 1'b0 ;
  assign n26702 = n4381 & n14407 ;
  assign n26703 = n8490 ^ n1454 ^ 1'b0 ;
  assign n26704 = ~n6283 & n26703 ;
  assign n26707 = n14936 ^ n6103 ^ 1'b0 ;
  assign n26708 = x27 & ~n26707 ;
  assign n26705 = n15326 & ~n18522 ;
  assign n26706 = ~n19238 & n26705 ;
  assign n26709 = n26708 ^ n26706 ^ n5275 ;
  assign n26712 = n4963 & n11665 ;
  assign n26713 = n26712 ^ n22861 ^ n7812 ;
  assign n26710 = n4323 | n25334 ;
  assign n26711 = n26710 ^ n4760 ^ 1'b0 ;
  assign n26714 = n26713 ^ n26711 ^ 1'b0 ;
  assign n26715 = n24404 | n26714 ;
  assign n26716 = n19594 ^ n741 ^ 1'b0 ;
  assign n26724 = n22554 ^ n775 ^ 1'b0 ;
  assign n26717 = n5333 ^ n1187 ^ 1'b0 ;
  assign n26718 = n8163 & n26717 ;
  assign n26719 = n2443 | n5349 ;
  assign n26720 = n1927 & ~n26719 ;
  assign n26721 = ( n12933 & n26718 ) | ( n12933 & n26720 ) | ( n26718 & n26720 ) ;
  assign n26722 = n11151 & n26721 ;
  assign n26723 = n4783 & n26722 ;
  assign n26725 = n26724 ^ n26723 ^ 1'b0 ;
  assign n26726 = n24862 & n26725 ;
  assign n26727 = n25819 ^ n21135 ^ 1'b0 ;
  assign n26728 = ( ~n5855 & n26726 ) | ( ~n5855 & n26727 ) | ( n26726 & n26727 ) ;
  assign n26729 = n9538 ^ x54 ^ 1'b0 ;
  assign n26730 = n12888 & ~n26729 ;
  assign n26731 = n1899 | n26730 ;
  assign n26732 = ~n16555 & n17379 ;
  assign n26733 = ~n26731 & n26732 ;
  assign n26734 = n26733 ^ n26041 ^ n10697 ;
  assign n26735 = n13816 ^ n13368 ^ 1'b0 ;
  assign n26736 = n12363 & n26735 ;
  assign n26737 = n7333 & ~n26736 ;
  assign n26738 = ( ~n7872 & n10491 ) | ( ~n7872 & n19333 ) | ( n10491 & n19333 ) ;
  assign n26739 = n15185 ^ n13734 ^ n12061 ;
  assign n26740 = n1983 & ~n5337 ;
  assign n26741 = n7923 | n26740 ;
  assign n26742 = n26741 ^ n11997 ^ 1'b0 ;
  assign n26743 = n2358 & ~n22440 ;
  assign n26744 = n26743 ^ n15772 ^ 1'b0 ;
  assign n26745 = n13538 & ~n19254 ;
  assign n26746 = n26745 ^ n14810 ^ 1'b0 ;
  assign n26747 = ( ~n4080 & n19789 ) | ( ~n4080 & n21991 ) | ( n19789 & n21991 ) ;
  assign n26748 = n1821 & n11317 ;
  assign n26749 = ( x221 & n4432 ) | ( x221 & n15397 ) | ( n4432 & n15397 ) ;
  assign n26750 = n13961 & ~n26749 ;
  assign n26751 = n26750 ^ n18590 ^ 1'b0 ;
  assign n26752 = n4291 ^ n1979 ^ n1320 ;
  assign n26753 = n17199 | n26752 ;
  assign n26754 = ~n7169 & n17083 ;
  assign n26755 = n900 & n2562 ;
  assign n26756 = n16792 | n26755 ;
  assign n26757 = n26756 ^ n23443 ^ n6097 ;
  assign n26758 = n310 | n3744 ;
  assign n26759 = n26758 ^ n2529 ^ 1'b0 ;
  assign n26760 = n26759 ^ n15693 ^ n6857 ;
  assign n26761 = n19974 | n26760 ;
  assign n26762 = n26761 ^ n8032 ^ 1'b0 ;
  assign n26763 = ~n857 & n26762 ;
  assign n26764 = n16714 ^ n15906 ^ n9337 ;
  assign n26765 = n26389 ^ n7917 ^ n4915 ;
  assign n26766 = n14433 & n26765 ;
  assign n26767 = ~n26764 & n26766 ;
  assign n26768 = n12676 & ~n13816 ;
  assign n26772 = n10618 & ~n15023 ;
  assign n26773 = n26772 ^ n25490 ^ 1'b0 ;
  assign n26769 = ( n5174 & ~n11011 ) | ( n5174 & n17307 ) | ( ~n11011 & n17307 ) ;
  assign n26770 = ~n7867 & n26769 ;
  assign n26771 = n6302 & n26770 ;
  assign n26774 = n26773 ^ n26771 ^ 1'b0 ;
  assign n26775 = n10261 | n12757 ;
  assign n26776 = n26775 ^ n15524 ^ 1'b0 ;
  assign n26777 = ~n16230 & n26776 ;
  assign n26778 = n26777 ^ n21261 ^ 1'b0 ;
  assign n26779 = ~x63 & n20531 ;
  assign n26780 = ( n341 & n6184 ) | ( n341 & ~n26779 ) | ( n6184 & ~n26779 ) ;
  assign n26781 = n24051 | n26780 ;
  assign n26782 = n17581 ^ n16586 ^ 1'b0 ;
  assign n26783 = n8343 & n26782 ;
  assign n26784 = n12169 ^ n740 ^ 1'b0 ;
  assign n26785 = n26783 & ~n26784 ;
  assign n26786 = x119 & ~n7055 ;
  assign n26787 = n5363 & n26786 ;
  assign n26788 = n16202 ^ n8387 ^ 1'b0 ;
  assign n26789 = n15462 ^ n3331 ^ 1'b0 ;
  assign n26792 = n5128 | n9910 ;
  assign n26793 = n26792 ^ n20727 ^ 1'b0 ;
  assign n26790 = n3649 & n21354 ;
  assign n26791 = ( ~n5825 & n24172 ) | ( ~n5825 & n26790 ) | ( n24172 & n26790 ) ;
  assign n26794 = n26793 ^ n26791 ^ 1'b0 ;
  assign n26795 = n684 & ~n5198 ;
  assign n26796 = n26795 ^ n3974 ^ 1'b0 ;
  assign n26797 = ( n2693 & n17738 ) | ( n2693 & ~n20446 ) | ( n17738 & ~n20446 ) ;
  assign n26798 = n6534 | n26797 ;
  assign n26799 = n6523 & ~n26798 ;
  assign n26800 = ( n19037 & n20513 ) | ( n19037 & n26799 ) | ( n20513 & n26799 ) ;
  assign n26801 = n13012 | n26800 ;
  assign n26802 = n26801 ^ n16548 ^ 1'b0 ;
  assign n26803 = n20193 ^ n10152 ^ 1'b0 ;
  assign n26804 = n23047 ^ n5014 ^ 1'b0 ;
  assign n26805 = n3042 & ~n6904 ;
  assign n26806 = n26805 ^ n640 ^ 1'b0 ;
  assign n26807 = n1999 & n26806 ;
  assign n26808 = n26807 ^ n387 ^ 1'b0 ;
  assign n26810 = n5462 ^ n733 ^ 1'b0 ;
  assign n26811 = n4902 & ~n26810 ;
  assign n26812 = ~n21799 & n26811 ;
  assign n26809 = ( n1981 & n13375 ) | ( n1981 & n20055 ) | ( n13375 & n20055 ) ;
  assign n26813 = n26812 ^ n26809 ^ 1'b0 ;
  assign n26814 = n26808 | n26813 ;
  assign n26815 = ~n6699 & n9444 ;
  assign n26816 = n22580 & n26815 ;
  assign n26817 = ( ~n6733 & n7376 ) | ( ~n6733 & n25153 ) | ( n7376 & n25153 ) ;
  assign n26818 = n26817 ^ n20240 ^ n7213 ;
  assign n26819 = n24981 ^ n4528 ^ 1'b0 ;
  assign n26820 = x63 & n26819 ;
  assign n26821 = ~n5762 & n19910 ;
  assign n26822 = ~n8742 & n26821 ;
  assign n26823 = ( n10050 & n12962 ) | ( n10050 & n22050 ) | ( n12962 & n22050 ) ;
  assign n26824 = n1174 & ~n10817 ;
  assign n26825 = n26824 ^ n7921 ^ 1'b0 ;
  assign n26826 = ~n18306 & n26825 ;
  assign n26827 = n2196 & n26826 ;
  assign n26828 = n26827 ^ n25078 ^ n10805 ;
  assign n26829 = n26823 & n26828 ;
  assign n26830 = ~n2977 & n26829 ;
  assign n26831 = n26830 ^ n2489 ^ 1'b0 ;
  assign n26832 = n11771 ^ n10402 ^ n7554 ;
  assign n26833 = ( x248 & n9600 ) | ( x248 & ~n26832 ) | ( n9600 & ~n26832 ) ;
  assign n26834 = n26833 ^ n5649 ^ 1'b0 ;
  assign n26835 = n26831 & n26834 ;
  assign n26841 = n981 & n6695 ;
  assign n26839 = n8709 ^ n1298 ^ 1'b0 ;
  assign n26840 = n2846 | n26839 ;
  assign n26842 = n26841 ^ n26840 ^ n6854 ;
  assign n26843 = ~n13314 & n26842 ;
  assign n26844 = n26843 ^ n19610 ^ 1'b0 ;
  assign n26836 = n12853 ^ n10922 ^ 1'b0 ;
  assign n26837 = n6420 & ~n26836 ;
  assign n26838 = ~n14424 & n26837 ;
  assign n26845 = n26844 ^ n26838 ^ 1'b0 ;
  assign n26848 = n21699 ^ n7994 ^ 1'b0 ;
  assign n26849 = n25943 & n26848 ;
  assign n26846 = n2645 | n10917 ;
  assign n26847 = ( ~n4938 & n9552 ) | ( ~n4938 & n26846 ) | ( n9552 & n26846 ) ;
  assign n26850 = n26849 ^ n26847 ^ 1'b0 ;
  assign n26851 = n727 & ~n13843 ;
  assign n26852 = n26851 ^ n7317 ^ 1'b0 ;
  assign n26853 = n8524 ^ n1886 ^ 1'b0 ;
  assign n26854 = ( n9937 & n18145 ) | ( n9937 & ~n26853 ) | ( n18145 & ~n26853 ) ;
  assign n26855 = ~n16722 & n24487 ;
  assign n26856 = n1761 & n16175 ;
  assign n26857 = ~n2484 & n26856 ;
  assign n26858 = n6411 & n26857 ;
  assign n26859 = n10826 ^ n1115 ^ 1'b0 ;
  assign n26860 = ~n26858 & n26859 ;
  assign n26861 = n15621 ^ n6065 ^ 1'b0 ;
  assign n26862 = ( n19121 & ~n26256 ) | ( n19121 & n26861 ) | ( ~n26256 & n26861 ) ;
  assign n26863 = n20723 ^ n17095 ^ 1'b0 ;
  assign n26864 = ( n457 & n26862 ) | ( n457 & ~n26863 ) | ( n26862 & ~n26863 ) ;
  assign n26865 = n6505 & n14224 ;
  assign n26866 = n23084 & ~n26865 ;
  assign n26867 = n26866 ^ n1434 ^ 1'b0 ;
  assign n26868 = n11114 & n26867 ;
  assign n26869 = ( n2439 & ~n5583 ) | ( n2439 & n9173 ) | ( ~n5583 & n9173 ) ;
  assign n26870 = n19311 ^ n3840 ^ 1'b0 ;
  assign n26871 = n23967 ^ n3578 ^ 1'b0 ;
  assign n26872 = n16693 ^ n3042 ^ 1'b0 ;
  assign n26873 = n26872 ^ n12811 ^ 1'b0 ;
  assign n26874 = n26871 | n26873 ;
  assign n26875 = n17526 ^ n13875 ^ 1'b0 ;
  assign n26876 = n5149 & n26875 ;
  assign n26877 = n1976 & n26876 ;
  assign n26878 = n21868 ^ n12268 ^ 1'b0 ;
  assign n26879 = ( n1770 & ~n26877 ) | ( n1770 & n26878 ) | ( ~n26877 & n26878 ) ;
  assign n26880 = n6086 ^ n4159 ^ n1674 ;
  assign n26881 = n949 & n23132 ;
  assign n26882 = n1310 & ~n26881 ;
  assign n26883 = ~n18386 & n26882 ;
  assign n26884 = ~n10067 & n18612 ;
  assign n26885 = n3688 & n4276 ;
  assign n26886 = n26885 ^ n14348 ^ 1'b0 ;
  assign n26887 = n14786 | n26886 ;
  assign n26888 = n6402 & ~n13446 ;
  assign n26889 = n8945 & n26888 ;
  assign n26890 = n21416 | n26889 ;
  assign n26891 = n26887 & ~n26890 ;
  assign n26892 = n12233 & n15424 ;
  assign n26893 = n26892 ^ n19123 ^ 1'b0 ;
  assign n26894 = n3403 & n26893 ;
  assign n26895 = ( n4237 & n9226 ) | ( n4237 & ~n26779 ) | ( n9226 & ~n26779 ) ;
  assign n26896 = n26895 ^ n7854 ^ 1'b0 ;
  assign n26897 = n8606 | n13150 ;
  assign n26898 = ~n4234 & n26507 ;
  assign n26899 = n1755 & ~n7209 ;
  assign n26900 = n26899 ^ n3705 ^ 1'b0 ;
  assign n26901 = ( n14734 & n23503 ) | ( n14734 & ~n26900 ) | ( n23503 & ~n26900 ) ;
  assign n26902 = x237 & ~n782 ;
  assign n26903 = n26902 ^ n1110 ^ 1'b0 ;
  assign n26904 = n26903 ^ n3583 ^ 1'b0 ;
  assign n26905 = n26901 & ~n26904 ;
  assign n26906 = n2118 ^ x137 ^ 1'b0 ;
  assign n26907 = n18416 ^ n15440 ^ n8343 ;
  assign n26908 = n26906 | n26907 ;
  assign n26909 = n17810 ^ n13257 ^ 1'b0 ;
  assign n26910 = n5049 ^ n4909 ^ 1'b0 ;
  assign n26911 = ~n1327 & n26910 ;
  assign n26912 = n26911 ^ x24 ^ 1'b0 ;
  assign n26913 = n18156 & n26912 ;
  assign n26914 = n26909 & ~n26913 ;
  assign n26915 = ( n676 & n2893 ) | ( n676 & ~n4341 ) | ( n2893 & ~n4341 ) ;
  assign n26916 = n26915 ^ n12682 ^ n5918 ;
  assign n26917 = n26916 ^ n18626 ^ 1'b0 ;
  assign n26918 = n1026 | n17562 ;
  assign n26919 = n26918 ^ n5972 ^ 1'b0 ;
  assign n26920 = n23182 ^ n20017 ^ 1'b0 ;
  assign n26921 = n26920 ^ n7426 ^ 1'b0 ;
  assign n26922 = ~n6480 & n26921 ;
  assign n26923 = ~n5267 & n12874 ;
  assign n26924 = n7741 & ~n12800 ;
  assign n26925 = n3351 | n13820 ;
  assign n26926 = n26925 ^ n18049 ^ n15098 ;
  assign n26927 = n4317 & n20979 ;
  assign n26928 = n6716 ^ n1196 ^ 1'b0 ;
  assign n26929 = n11140 & ~n12966 ;
  assign n26930 = n16767 & n26929 ;
  assign n26931 = n2560 | n3328 ;
  assign n26932 = n26930 & ~n26931 ;
  assign n26933 = n7489 ^ n7017 ^ 1'b0 ;
  assign n26934 = n1453 & n26933 ;
  assign n26935 = n26934 ^ n21715 ^ 1'b0 ;
  assign n26936 = n11853 & n12416 ;
  assign n26937 = n19868 ^ n16817 ^ 1'b0 ;
  assign n26938 = n26936 | n26937 ;
  assign n26939 = n9266 & ~n24085 ;
  assign n26940 = ~n24787 & n26939 ;
  assign n26941 = n5550 & ~n9158 ;
  assign n26942 = n26941 ^ n14924 ^ 1'b0 ;
  assign n26943 = n23874 ^ n5471 ^ 1'b0 ;
  assign n26944 = n26942 & ~n26943 ;
  assign n26945 = n26944 ^ n13735 ^ 1'b0 ;
  assign n26947 = n4954 ^ n3396 ^ 1'b0 ;
  assign n26948 = n23631 & ~n26947 ;
  assign n26949 = n26948 ^ n13057 ^ 1'b0 ;
  assign n26946 = n656 & n9215 ;
  assign n26950 = n26949 ^ n26946 ^ n18545 ;
  assign n26952 = n3050 ^ n2057 ^ 1'b0 ;
  assign n26953 = ~n3494 & n26952 ;
  assign n26954 = n14170 | n26953 ;
  assign n26955 = x200 & n26954 ;
  assign n26951 = n7950 & n16290 ;
  assign n26956 = n26955 ^ n26951 ^ 1'b0 ;
  assign n26957 = n13051 ^ n3667 ^ n3634 ;
  assign n26958 = n6669 ^ n3758 ^ 1'b0 ;
  assign n26959 = n26957 & ~n26958 ;
  assign n26960 = n1586 & n9318 ;
  assign n26961 = n1852 | n22717 ;
  assign n26962 = n26960 | n26961 ;
  assign n26963 = n21318 | n21522 ;
  assign n26964 = n6910 & ~n26963 ;
  assign n26965 = ~n3404 & n17335 ;
  assign n26966 = n4867 & n26965 ;
  assign n26967 = n26966 ^ n9025 ^ 1'b0 ;
  assign n26968 = n2662 & n26967 ;
  assign n26969 = n18944 ^ n17209 ^ 1'b0 ;
  assign n26970 = n26969 ^ n25522 ^ n6563 ;
  assign n26971 = n3343 | n6133 ;
  assign n26972 = n4083 | n15517 ;
  assign n26973 = ~n4752 & n26972 ;
  assign n26974 = n26973 ^ n10435 ^ n438 ;
  assign n26975 = n26974 ^ n23417 ^ n612 ;
  assign n26976 = n17063 | n25825 ;
  assign n26977 = n26976 ^ n12358 ^ 1'b0 ;
  assign n26978 = n2394 & n12036 ;
  assign n26979 = ( n5075 & n6351 ) | ( n5075 & ~n14567 ) | ( n6351 & ~n14567 ) ;
  assign n26980 = n24613 ^ n3432 ^ 1'b0 ;
  assign n26981 = n26979 & n26980 ;
  assign n26982 = n5114 ^ n3024 ^ 1'b0 ;
  assign n26983 = ~n5746 & n19677 ;
  assign n26984 = n26982 & n26983 ;
  assign n26985 = n26984 ^ n26966 ^ n16536 ;
  assign n26986 = n13748 ^ n1463 ^ 1'b0 ;
  assign n26987 = n10056 & n26747 ;
  assign n26988 = ~n26986 & n26987 ;
  assign n26989 = n14251 & n16938 ;
  assign n26990 = n11048 | n14082 ;
  assign n26991 = n2502 | n10877 ;
  assign n26992 = n11873 | n26991 ;
  assign n26993 = ( n7444 & n9960 ) | ( n7444 & n26992 ) | ( n9960 & n26992 ) ;
  assign n26994 = n14926 ^ n853 ^ 1'b0 ;
  assign n26995 = ( n14248 & n26993 ) | ( n14248 & n26994 ) | ( n26993 & n26994 ) ;
  assign n26996 = n2500 & ~n20091 ;
  assign n26997 = n26996 ^ n3062 ^ 1'b0 ;
  assign n26998 = ( n1813 & ~n26995 ) | ( n1813 & n26997 ) | ( ~n26995 & n26997 ) ;
  assign n26999 = n15766 ^ n5499 ^ 1'b0 ;
  assign n27000 = n17042 | n26999 ;
  assign n27001 = n3378 & ~n19598 ;
  assign n27002 = n27001 ^ n16619 ^ 1'b0 ;
  assign n27005 = n1486 & ~n4525 ;
  assign n27004 = ( n4940 & ~n7925 ) | ( n4940 & n15139 ) | ( ~n7925 & n15139 ) ;
  assign n27003 = n7389 | n11680 ;
  assign n27006 = n27005 ^ n27004 ^ n27003 ;
  assign n27007 = n307 & ~n12458 ;
  assign n27008 = n13786 & ~n14279 ;
  assign n27009 = n27007 & n27008 ;
  assign n27010 = ~n12062 & n13556 ;
  assign n27011 = ~n10636 & n27010 ;
  assign n27012 = n27011 ^ n8306 ^ 1'b0 ;
  assign n27016 = n991 & ~n9295 ;
  assign n27017 = n27016 ^ n7762 ^ 1'b0 ;
  assign n27018 = n27017 ^ n6164 ^ n1862 ;
  assign n27013 = ( n1105 & n1853 ) | ( n1105 & ~n2133 ) | ( n1853 & ~n2133 ) ;
  assign n27014 = n15660 ^ n2026 ^ 1'b0 ;
  assign n27015 = n27013 | n27014 ;
  assign n27019 = n27018 ^ n27015 ^ n10695 ;
  assign n27020 = n3853 & ~n16060 ;
  assign n27021 = n1597 & n27020 ;
  assign n27022 = ( n22135 & n23138 ) | ( n22135 & ~n27021 ) | ( n23138 & ~n27021 ) ;
  assign n27023 = ( n3768 & n21875 ) | ( n3768 & ~n23635 ) | ( n21875 & ~n23635 ) ;
  assign n27024 = n8552 | n11686 ;
  assign n27025 = n4059 | n27024 ;
  assign n27026 = n27025 ^ n2992 ^ 1'b0 ;
  assign n27027 = n6839 & ~n27026 ;
  assign n27028 = n15423 & n27027 ;
  assign n27029 = n13884 ^ n11291 ^ 1'b0 ;
  assign n27030 = n27029 ^ n19386 ^ n10212 ;
  assign n27031 = n27030 ^ n10123 ^ n906 ;
  assign n27032 = n7486 ^ n5749 ^ 1'b0 ;
  assign n27033 = n3096 & n6750 ;
  assign n27034 = ~n27032 & n27033 ;
  assign n27035 = n8193 & n27034 ;
  assign n27036 = n27035 ^ n19333 ^ n6546 ;
  assign n27037 = ( ~n559 & n10292 ) | ( ~n559 & n19700 ) | ( n10292 & n19700 ) ;
  assign n27038 = n6280 | n24550 ;
  assign n27039 = n12450 | n27038 ;
  assign n27041 = n13102 | n20271 ;
  assign n27040 = n11909 | n12664 ;
  assign n27042 = n27041 ^ n27040 ^ 1'b0 ;
  assign n27043 = n17896 ^ n7296 ^ n1862 ;
  assign n27044 = n27043 ^ n1616 ^ 1'b0 ;
  assign n27045 = n27044 ^ n6473 ^ 1'b0 ;
  assign n27046 = n11173 & ~n11365 ;
  assign n27047 = ~n10925 & n27046 ;
  assign n27048 = n27047 ^ n11045 ^ 1'b0 ;
  assign n27049 = n11588 & ~n11880 ;
  assign n27050 = n27049 ^ n19669 ^ x24 ;
  assign n27051 = n27050 ^ n14427 ^ 1'b0 ;
  assign n27052 = n5269 & n8416 ;
  assign n27053 = n23468 & n27052 ;
  assign n27054 = n15972 ^ n4115 ^ 1'b0 ;
  assign n27055 = n3227 | n27054 ;
  assign n27056 = n26054 ^ n18985 ^ n15572 ;
  assign n27058 = n10271 & n10866 ;
  assign n27059 = n20980 ^ n951 ^ 1'b0 ;
  assign n27060 = n27058 & ~n27059 ;
  assign n27057 = n21869 ^ n5726 ^ n518 ;
  assign n27061 = n27060 ^ n27057 ^ n3002 ;
  assign n27062 = n4664 & ~n12866 ;
  assign n27063 = n18992 & ~n27062 ;
  assign n27064 = ~n10437 & n27063 ;
  assign n27065 = n27064 ^ n3954 ^ 1'b0 ;
  assign n27066 = n10947 | n27065 ;
  assign n27067 = ~n1406 & n22967 ;
  assign n27068 = n7881 & n27067 ;
  assign n27069 = n9838 | n27068 ;
  assign n27070 = n13317 | n23052 ;
  assign n27071 = n27070 ^ n9732 ^ 1'b0 ;
  assign n27073 = n19078 ^ n907 ^ 1'b0 ;
  assign n27074 = ( n7568 & n12360 ) | ( n7568 & n27073 ) | ( n12360 & n27073 ) ;
  assign n27072 = n8264 ^ n3732 ^ 1'b0 ;
  assign n27075 = n27074 ^ n27072 ^ 1'b0 ;
  assign n27076 = ( n5107 & ~n6326 ) | ( n5107 & n8589 ) | ( ~n6326 & n8589 ) ;
  assign n27077 = n5288 & ~n27076 ;
  assign n27078 = n8787 ^ n3121 ^ 1'b0 ;
  assign n27079 = n10850 & n27078 ;
  assign n27080 = n27079 ^ n4441 ^ 1'b0 ;
  assign n27081 = ( n15654 & n23355 ) | ( n15654 & ~n26374 ) | ( n23355 & ~n26374 ) ;
  assign n27083 = n2523 | n20248 ;
  assign n27084 = n1831 & ~n27083 ;
  assign n27082 = n14596 & ~n22617 ;
  assign n27085 = n27084 ^ n27082 ^ 1'b0 ;
  assign n27086 = n27085 ^ n13630 ^ 1'b0 ;
  assign n27087 = ~n565 & n10518 ;
  assign n27088 = n27087 ^ n15221 ^ 1'b0 ;
  assign n27089 = n19911 ^ n15590 ^ 1'b0 ;
  assign n27090 = ( n11048 & n27088 ) | ( n11048 & ~n27089 ) | ( n27088 & ~n27089 ) ;
  assign n27091 = ~n9829 & n19897 ;
  assign n27092 = n5012 ^ x126 ^ 1'b0 ;
  assign n27093 = n27092 ^ n21473 ^ n16761 ;
  assign n27098 = n7775 | n20654 ;
  assign n27099 = n27098 ^ n15436 ^ 1'b0 ;
  assign n27096 = n4449 | n15114 ;
  assign n27097 = n15299 | n27096 ;
  assign n27100 = n27099 ^ n27097 ^ 1'b0 ;
  assign n27101 = n27100 ^ n6619 ^ 1'b0 ;
  assign n27102 = n27101 ^ n427 ^ 1'b0 ;
  assign n27103 = n10323 & ~n27102 ;
  assign n27094 = n4342 & ~n18557 ;
  assign n27095 = n6060 & ~n27094 ;
  assign n27104 = n27103 ^ n27095 ^ 1'b0 ;
  assign n27105 = n22306 ^ n8406 ^ 1'b0 ;
  assign n27106 = n27105 ^ n21119 ^ 1'b0 ;
  assign n27107 = n10296 | n11590 ;
  assign n27108 = n6434 & ~n27107 ;
  assign n27109 = n27108 ^ n7647 ^ 1'b0 ;
  assign n27110 = n6636 | n12194 ;
  assign n27111 = n5065 & n27110 ;
  assign n27112 = n8716 & n27111 ;
  assign n27113 = n9314 | n27112 ;
  assign n27114 = n4817 ^ n1472 ^ 1'b0 ;
  assign n27115 = n21311 | n27114 ;
  assign n27116 = n27115 ^ n6910 ^ 1'b0 ;
  assign n27117 = n1452 & ~n3793 ;
  assign n27118 = ~n27116 & n27117 ;
  assign n27122 = n6853 ^ n6093 ^ 1'b0 ;
  assign n27123 = n27122 ^ n1624 ^ 1'b0 ;
  assign n27119 = n1689 | n4591 ;
  assign n27120 = n27119 ^ n9497 ^ 1'b0 ;
  assign n27121 = n12664 & ~n27120 ;
  assign n27124 = n27123 ^ n27121 ^ 1'b0 ;
  assign n27125 = n18916 & n21121 ;
  assign n27126 = ~n18590 & n27125 ;
  assign n27127 = n12721 ^ n5956 ^ 1'b0 ;
  assign n27128 = n9280 & n26752 ;
  assign n27129 = ~n4776 & n27128 ;
  assign n27130 = n9845 | n27129 ;
  assign n27131 = ~n7958 & n27130 ;
  assign n27132 = n27131 ^ n21651 ^ 1'b0 ;
  assign n27133 = ( ~n12828 & n18576 ) | ( ~n12828 & n24537 ) | ( n18576 & n24537 ) ;
  assign n27134 = ~n7665 & n24446 ;
  assign n27135 = n7035 | n13508 ;
  assign n27136 = n1386 & ~n27135 ;
  assign n27137 = n4714 & ~n24691 ;
  assign n27138 = n14711 ^ n5368 ^ n4400 ;
  assign n27139 = n18482 & ~n27138 ;
  assign n27140 = n10712 & n27139 ;
  assign n27141 = ( n3368 & n7335 ) | ( n3368 & n8948 ) | ( n7335 & n8948 ) ;
  assign n27142 = n27141 ^ n26808 ^ n11187 ;
  assign n27143 = n24707 ^ n8975 ^ 1'b0 ;
  assign n27144 = n24858 ^ n21715 ^ 1'b0 ;
  assign n27145 = ~n8657 & n27144 ;
  assign n27146 = n3436 | n26006 ;
  assign n27147 = n27146 ^ n16840 ^ 1'b0 ;
  assign n27148 = n23306 | n27147 ;
  assign n27149 = n9615 ^ n1134 ^ 1'b0 ;
  assign n27150 = n27149 ^ n13810 ^ n5895 ;
  assign n27153 = ( n704 & ~n5291 ) | ( n704 & n10317 ) | ( ~n5291 & n10317 ) ;
  assign n27151 = n17396 ^ n16643 ^ n12035 ;
  assign n27152 = ~n22120 & n27151 ;
  assign n27154 = n27153 ^ n27152 ^ 1'b0 ;
  assign n27155 = n14606 ^ n2578 ^ n1378 ;
  assign n27156 = n13041 ^ n8887 ^ 1'b0 ;
  assign n27157 = n13107 | n27156 ;
  assign n27158 = n9467 | n27157 ;
  assign n27159 = n17808 & ~n27158 ;
  assign n27160 = ~n16292 & n21205 ;
  assign n27161 = n1304 | n12826 ;
  assign n27162 = n27160 | n27161 ;
  assign n27163 = n3962 & n8150 ;
  assign n27164 = n3338 & n8711 ;
  assign n27165 = n1628 & n6105 ;
  assign n27166 = n27165 ^ n6034 ^ 1'b0 ;
  assign n27167 = n27166 ^ n17615 ^ n6446 ;
  assign n27168 = n9486 ^ n7580 ^ 1'b0 ;
  assign n27169 = n26657 | n27168 ;
  assign n27170 = ~n12270 & n19919 ;
  assign n27171 = ~n27169 & n27170 ;
  assign n27172 = ( n5767 & n15707 ) | ( n5767 & n22679 ) | ( n15707 & n22679 ) ;
  assign n27173 = n4265 & ~n15029 ;
  assign n27174 = n1746 & n27173 ;
  assign n27175 = n27174 ^ n5191 ^ 1'b0 ;
  assign n27176 = ( ~n6534 & n9206 ) | ( ~n6534 & n9645 ) | ( n9206 & n9645 ) ;
  assign n27177 = n11635 ^ n5002 ^ 1'b0 ;
  assign n27178 = n27176 & n27177 ;
  assign n27179 = n26353 ^ n18165 ^ 1'b0 ;
  assign n27180 = n27178 & n27179 ;
  assign n27181 = n27180 ^ n8588 ^ 1'b0 ;
  assign n27182 = n3073 & ~n16022 ;
  assign n27183 = ( n7266 & ~n12956 ) | ( n7266 & n27182 ) | ( ~n12956 & n27182 ) ;
  assign n27184 = n27183 ^ n15599 ^ 1'b0 ;
  assign n27185 = n24968 | n27184 ;
  assign n27186 = ( n15240 & ~n16948 ) | ( n15240 & n27185 ) | ( ~n16948 & n27185 ) ;
  assign n27192 = n9936 & ~n13215 ;
  assign n27193 = ~n1174 & n27192 ;
  assign n27194 = n27193 ^ n10824 ^ n9422 ;
  assign n27187 = n11969 & n24164 ;
  assign n27188 = n13062 & n27187 ;
  assign n27189 = n19947 ^ n962 ^ 1'b0 ;
  assign n27190 = ~n27188 & n27189 ;
  assign n27191 = ~n17916 & n27190 ;
  assign n27195 = n27194 ^ n27191 ^ 1'b0 ;
  assign n27196 = n3300 ^ n1374 ^ 1'b0 ;
  assign n27197 = n20065 & ~n27196 ;
  assign n27198 = n10303 ^ n5444 ^ 1'b0 ;
  assign n27199 = n11481 ^ n9366 ^ 1'b0 ;
  assign n27200 = ( n15461 & n16703 ) | ( n15461 & ~n27199 ) | ( n16703 & ~n27199 ) ;
  assign n27201 = n27200 ^ n22977 ^ 1'b0 ;
  assign n27202 = n27198 | n27201 ;
  assign n27203 = n15039 ^ n11591 ^ n10646 ;
  assign n27204 = n2466 | n12341 ;
  assign n27205 = n9059 & n17203 ;
  assign n27206 = n424 & n27205 ;
  assign n27207 = ( n4264 & ~n18534 ) | ( n4264 & n27206 ) | ( ~n18534 & n27206 ) ;
  assign n27208 = ( x0 & ~n23198 ) | ( x0 & n27207 ) | ( ~n23198 & n27207 ) ;
  assign n27209 = ( n421 & ~n10585 ) | ( n421 & n13972 ) | ( ~n10585 & n13972 ) ;
  assign n27210 = n3366 & ~n27209 ;
  assign n27211 = n27210 ^ n9985 ^ 1'b0 ;
  assign n27212 = n4190 & n27211 ;
  assign n27213 = n18875 ^ n7503 ^ 1'b0 ;
  assign n27214 = n8760 ^ n3417 ^ n1058 ;
  assign n27215 = ~n13437 & n27214 ;
  assign n27216 = n6476 & n27215 ;
  assign n27217 = n27216 ^ n2838 ^ 1'b0 ;
  assign n27218 = n1821 & ~n27217 ;
  assign n27219 = n27218 ^ n3712 ^ 1'b0 ;
  assign n27220 = n27219 ^ n2230 ^ 1'b0 ;
  assign n27221 = n3722 & n12156 ;
  assign n27222 = n13797 ^ n1175 ^ 1'b0 ;
  assign n27223 = ( ~n1776 & n7542 ) | ( ~n1776 & n27222 ) | ( n7542 & n27222 ) ;
  assign n27224 = ~n12354 & n27223 ;
  assign n27225 = n27224 ^ n13344 ^ 1'b0 ;
  assign n27226 = ~n4176 & n27225 ;
  assign n27227 = ~n27221 & n27226 ;
  assign n27228 = n27227 ^ x172 ^ 1'b0 ;
  assign n27229 = x64 & n2468 ;
  assign n27230 = n3156 & n27229 ;
  assign n27231 = n24907 & ~n27230 ;
  assign n27232 = ~n17039 & n27231 ;
  assign n27233 = n262 & n5793 ;
  assign n27234 = n4544 & n7950 ;
  assign n27235 = n27233 & n27234 ;
  assign n27236 = ~n10906 & n20965 ;
  assign n27237 = n5773 ^ n4173 ^ 1'b0 ;
  assign n27238 = n21004 ^ n8781 ^ n7716 ;
  assign n27239 = n18453 & n19058 ;
  assign n27240 = n27239 ^ n20453 ^ 1'b0 ;
  assign n27241 = n27240 ^ n20772 ^ n8985 ;
  assign n27242 = n19604 ^ n2406 ^ 1'b0 ;
  assign n27243 = n19555 & n27242 ;
  assign n27244 = n1219 | n25002 ;
  assign n27245 = n24220 | n27244 ;
  assign n27246 = n6812 ^ n2551 ^ n814 ;
  assign n27247 = n9075 | n27246 ;
  assign n27248 = n19353 ^ n7823 ^ n2729 ;
  assign n27249 = ( n4553 & n6462 ) | ( n4553 & ~n11007 ) | ( n6462 & ~n11007 ) ;
  assign n27250 = ( n27247 & n27248 ) | ( n27247 & n27249 ) | ( n27248 & n27249 ) ;
  assign n27251 = ( ~n12650 & n16366 ) | ( ~n12650 & n18915 ) | ( n16366 & n18915 ) ;
  assign n27252 = ( n6894 & n14905 ) | ( n6894 & ~n27251 ) | ( n14905 & ~n27251 ) ;
  assign n27253 = n3999 ^ n3770 ^ 1'b0 ;
  assign n27254 = n18372 ^ n10245 ^ 1'b0 ;
  assign n27256 = n8381 ^ n3591 ^ n330 ;
  assign n27255 = n10226 | n10345 ;
  assign n27257 = n27256 ^ n27255 ^ n6626 ;
  assign n27258 = n12515 & n15451 ;
  assign n27259 = n20781 & n27258 ;
  assign n27260 = n21487 ^ n7275 ^ 1'b0 ;
  assign n27261 = n25448 & n27260 ;
  assign n27262 = n27261 ^ n2859 ^ 1'b0 ;
  assign n27263 = ( ~n3986 & n9643 ) | ( ~n3986 & n20568 ) | ( n9643 & n20568 ) ;
  assign n27264 = ( n7359 & ~n15981 ) | ( n7359 & n27263 ) | ( ~n15981 & n27263 ) ;
  assign n27265 = n27264 ^ n7265 ^ n4308 ;
  assign n27266 = n4223 & n25261 ;
  assign n27267 = n13127 & n27266 ;
  assign n27268 = ( n7305 & ~n10798 ) | ( n7305 & n11202 ) | ( ~n10798 & n11202 ) ;
  assign n27269 = n16737 & ~n21003 ;
  assign n27270 = n27269 ^ n10231 ^ 1'b0 ;
  assign n27271 = ( n9163 & n14304 ) | ( n9163 & ~n27270 ) | ( n14304 & ~n27270 ) ;
  assign n27272 = ~n5973 & n21987 ;
  assign n27273 = n27272 ^ n12231 ^ 1'b0 ;
  assign n27274 = n24796 ^ n19947 ^ 1'b0 ;
  assign n27275 = n8572 & n27274 ;
  assign n27276 = n1956 | n8978 ;
  assign n27283 = n2045 ^ n286 ^ 1'b0 ;
  assign n27284 = n3905 & n27283 ;
  assign n27279 = n3510 | n17649 ;
  assign n27280 = n9857 & ~n27279 ;
  assign n27277 = n7064 | n10520 ;
  assign n27278 = n27277 ^ n3693 ^ 1'b0 ;
  assign n27281 = n27280 ^ n27278 ^ 1'b0 ;
  assign n27282 = n7485 & ~n27281 ;
  assign n27285 = n27284 ^ n27282 ^ 1'b0 ;
  assign n27286 = n5077 & ~n18529 ;
  assign n27287 = n27286 ^ n13753 ^ 1'b0 ;
  assign n27288 = n2504 ^ x150 ^ 1'b0 ;
  assign n27289 = ~n18610 & n19810 ;
  assign n27290 = n27289 ^ n9800 ^ 1'b0 ;
  assign n27291 = n27290 ^ n20310 ^ 1'b0 ;
  assign n27292 = n2023 | n8076 ;
  assign n27293 = n27291 | n27292 ;
  assign n27299 = n11154 & ~n20291 ;
  assign n27300 = n27299 ^ n7745 ^ 1'b0 ;
  assign n27294 = n18836 ^ n7607 ^ 1'b0 ;
  assign n27295 = n13703 ^ n2877 ^ 1'b0 ;
  assign n27296 = n4191 & n27295 ;
  assign n27297 = n27294 & n27296 ;
  assign n27298 = n8116 & n27297 ;
  assign n27301 = n27300 ^ n27298 ^ n25093 ;
  assign n27305 = n15870 ^ n15287 ^ n4083 ;
  assign n27302 = n12828 ^ n961 ^ 1'b0 ;
  assign n27303 = ~n16542 & n27302 ;
  assign n27304 = ~n9711 & n27303 ;
  assign n27306 = n27305 ^ n27304 ^ n25235 ;
  assign n27307 = n945 & ~n3071 ;
  assign n27308 = n27307 ^ n14407 ^ 1'b0 ;
  assign n27309 = n27308 ^ n19438 ^ n14225 ;
  assign n27310 = n6512 | n13643 ;
  assign n27311 = n9592 & n13962 ;
  assign n27312 = ~n27310 & n27311 ;
  assign n27313 = n27312 ^ n1657 ^ 1'b0 ;
  assign n27315 = x252 & ~n10732 ;
  assign n27314 = n11589 & ~n21153 ;
  assign n27316 = n27315 ^ n27314 ^ 1'b0 ;
  assign n27317 = n14348 & n27316 ;
  assign n27318 = ~n1962 & n6050 ;
  assign n27319 = n19490 ^ n7410 ^ n2090 ;
  assign n27320 = ( n4489 & n8675 ) | ( n4489 & ~n24723 ) | ( n8675 & ~n24723 ) ;
  assign n27321 = ( n18713 & n27319 ) | ( n18713 & ~n27320 ) | ( n27319 & ~n27320 ) ;
  assign n27322 = ~n27318 & n27321 ;
  assign n27323 = n1435 & n27322 ;
  assign n27324 = n13996 ^ n2086 ^ 1'b0 ;
  assign n27325 = ( n1249 & ~n2657 ) | ( n1249 & n10171 ) | ( ~n2657 & n10171 ) ;
  assign n27326 = ~n13951 & n27325 ;
  assign n27327 = n23024 & n27326 ;
  assign n27328 = n11515 | n27327 ;
  assign n27329 = n27328 ^ n24736 ^ n6532 ;
  assign n27332 = n24817 ^ n23073 ^ 1'b0 ;
  assign n27333 = n6688 & ~n27332 ;
  assign n27330 = ( n717 & ~n2199 ) | ( n717 & n2287 ) | ( ~n2199 & n2287 ) ;
  assign n27331 = ~n1882 & n27330 ;
  assign n27334 = n27333 ^ n27331 ^ 1'b0 ;
  assign n27335 = n436 & ~n8837 ;
  assign n27336 = ~n7382 & n27335 ;
  assign n27337 = n27336 ^ n4343 ^ 1'b0 ;
  assign n27338 = n14498 ^ n1455 ^ 1'b0 ;
  assign n27339 = ( ~n18255 & n18950 ) | ( ~n18255 & n27338 ) | ( n18950 & n27338 ) ;
  assign n27340 = n10675 ^ n7749 ^ 1'b0 ;
  assign n27341 = n7339 ^ n1438 ^ 1'b0 ;
  assign n27342 = n27341 ^ n9176 ^ 1'b0 ;
  assign n27343 = ~n27340 & n27342 ;
  assign n27344 = n2701 & ~n4916 ;
  assign n27345 = n17625 & n27344 ;
  assign n27347 = n15035 ^ n6103 ^ n5911 ;
  assign n27346 = n6592 & n16890 ;
  assign n27348 = n27347 ^ n27346 ^ 1'b0 ;
  assign n27349 = n13168 ^ n8524 ^ 1'b0 ;
  assign n27350 = n27349 ^ n24494 ^ n14510 ;
  assign n27352 = n4088 & n4199 ;
  assign n27351 = n5236 | n15744 ;
  assign n27353 = n27352 ^ n27351 ^ 1'b0 ;
  assign n27354 = ( ~n2449 & n5658 ) | ( ~n2449 & n13535 ) | ( n5658 & n13535 ) ;
  assign n27355 = n1585 | n1846 ;
  assign n27356 = n5377 & ~n27355 ;
  assign n27357 = n10283 | n27356 ;
  assign n27358 = n12145 | n25026 ;
  assign n27359 = n15577 ^ n10688 ^ n6382 ;
  assign n27360 = n17161 ^ n1260 ^ 1'b0 ;
  assign n27361 = n6730 & n27360 ;
  assign n27362 = n27359 & n27361 ;
  assign n27363 = n8416 & n27362 ;
  assign n27364 = n27363 ^ n19114 ^ 1'b0 ;
  assign n27365 = n27364 ^ n17874 ^ 1'b0 ;
  assign n27366 = n19305 ^ n6179 ^ 1'b0 ;
  assign n27367 = n11777 ^ n2333 ^ 1'b0 ;
  assign n27368 = n3146 ^ n476 ^ 1'b0 ;
  assign n27369 = n4373 & n27368 ;
  assign n27370 = n4954 ^ x75 ^ 1'b0 ;
  assign n27371 = n1178 & n27370 ;
  assign n27372 = ( n7322 & ~n9417 ) | ( n7322 & n27371 ) | ( ~n9417 & n27371 ) ;
  assign n27373 = ~n4070 & n7327 ;
  assign n27374 = n3263 | n27373 ;
  assign n27375 = n27374 ^ n16569 ^ 1'b0 ;
  assign n27376 = n27375 ^ n8343 ^ 1'b0 ;
  assign n27377 = n27372 & ~n27376 ;
  assign n27378 = n8964 & n27377 ;
  assign n27379 = n27378 ^ n22681 ^ 1'b0 ;
  assign n27380 = n27110 & n27379 ;
  assign n27381 = n5778 ^ n1863 ^ x210 ;
  assign n27382 = ~n27380 & n27381 ;
  assign n27383 = n12778 ^ n5436 ^ 1'b0 ;
  assign n27384 = n26675 ^ n10339 ^ n2391 ;
  assign n27385 = n6152 & ~n9160 ;
  assign n27386 = n27385 ^ n5606 ^ 1'b0 ;
  assign n27387 = n27384 | n27386 ;
  assign n27388 = n27387 ^ n6154 ^ 1'b0 ;
  assign n27389 = ~n27383 & n27388 ;
  assign n27390 = n9154 ^ n6915 ^ 1'b0 ;
  assign n27391 = n1306 | n27390 ;
  assign n27392 = ~n2062 & n27391 ;
  assign n27393 = ~n6260 & n21259 ;
  assign n27394 = n5387 & ~n27393 ;
  assign n27395 = n11546 & ~n27394 ;
  assign n27396 = n5475 ^ n892 ^ x68 ;
  assign n27397 = n27396 ^ n7019 ^ 1'b0 ;
  assign n27398 = n7726 & n27397 ;
  assign n27399 = ~n7568 & n9957 ;
  assign n27400 = n4361 & n27399 ;
  assign n27401 = n8585 & n27400 ;
  assign n27405 = n11114 & n11990 ;
  assign n27406 = ~n11227 & n27405 ;
  assign n27402 = n7248 & ~n8072 ;
  assign n27403 = n26066 & n27402 ;
  assign n27404 = n2650 | n27403 ;
  assign n27407 = n27406 ^ n27404 ^ 1'b0 ;
  assign n27408 = n10030 | n17191 ;
  assign n27409 = n19874 | n27408 ;
  assign n27410 = n19363 & n20722 ;
  assign n27411 = n3978 & n27410 ;
  assign n27412 = n22155 ^ n8420 ^ 1'b0 ;
  assign n27413 = n27411 | n27412 ;
  assign n27418 = n3093 & ~n7179 ;
  assign n27419 = ~n279 & n27418 ;
  assign n27420 = ( n5803 & n12391 ) | ( n5803 & n27419 ) | ( n12391 & n27419 ) ;
  assign n27414 = n8871 ^ n7892 ^ 1'b0 ;
  assign n27415 = ~n9903 & n27414 ;
  assign n27416 = n1116 & n27415 ;
  assign n27417 = ~n12155 & n27416 ;
  assign n27421 = n27420 ^ n27417 ^ n9836 ;
  assign n27422 = ( n13130 & n16876 ) | ( n13130 & n18825 ) | ( n16876 & n18825 ) ;
  assign n27423 = n8612 & n27243 ;
  assign n27424 = n27422 & n27423 ;
  assign n27425 = n13542 ^ n7320 ^ n5225 ;
  assign n27426 = n27425 ^ n3187 ^ n2199 ;
  assign n27427 = n8799 & ~n27426 ;
  assign n27428 = n1927 & ~n18654 ;
  assign n27429 = n27428 ^ n9277 ^ 1'b0 ;
  assign n27430 = n27427 & n27429 ;
  assign n27431 = n10439 & ~n11995 ;
  assign n27432 = n27431 ^ n11059 ^ 1'b0 ;
  assign n27434 = n6711 | n11365 ;
  assign n27435 = n27434 ^ n692 ^ 1'b0 ;
  assign n27433 = n11059 | n27362 ;
  assign n27436 = n27435 ^ n27433 ^ 1'b0 ;
  assign n27437 = n8721 | n22012 ;
  assign n27438 = n18848 & ~n27437 ;
  assign n27439 = ( n3539 & ~n6931 ) | ( n3539 & n13341 ) | ( ~n6931 & n13341 ) ;
  assign n27440 = ( n2418 & n17608 ) | ( n2418 & n27439 ) | ( n17608 & n27439 ) ;
  assign n27441 = n2630 ^ n2344 ^ n1274 ;
  assign n27442 = n27441 ^ n9632 ^ 1'b0 ;
  assign n27443 = n23988 ^ n10489 ^ n1349 ;
  assign n27444 = ~n2205 & n10288 ;
  assign n27445 = n15073 ^ n2942 ^ 1'b0 ;
  assign n27447 = n2172 ^ n981 ^ 1'b0 ;
  assign n27448 = ~n2511 & n27447 ;
  assign n27449 = n27448 ^ n3518 ^ 1'b0 ;
  assign n27446 = n2731 & ~n9944 ;
  assign n27450 = n27449 ^ n27446 ^ 1'b0 ;
  assign n27451 = n1162 & n27450 ;
  assign n27453 = n18984 ^ n15109 ^ 1'b0 ;
  assign n27452 = n3247 & ~n17278 ;
  assign n27454 = n27453 ^ n27452 ^ n15893 ;
  assign n27455 = n16125 | n22294 ;
  assign n27456 = n2966 | n27455 ;
  assign n27457 = n25688 ^ n12957 ^ 1'b0 ;
  assign n27458 = n13407 ^ n13340 ^ 1'b0 ;
  assign n27459 = n4577 & n27458 ;
  assign n27460 = n398 & n27459 ;
  assign n27461 = x74 & ~n7355 ;
  assign n27462 = n27461 ^ n945 ^ 1'b0 ;
  assign n27463 = n9309 | n27462 ;
  assign n27464 = n14560 | n27463 ;
  assign n27465 = ( n4329 & n10134 ) | ( n4329 & ~n21851 ) | ( n10134 & ~n21851 ) ;
  assign n27466 = ( n8690 & n16487 ) | ( n8690 & ~n27465 ) | ( n16487 & ~n27465 ) ;
  assign n27467 = n27466 ^ n9957 ^ 1'b0 ;
  assign n27468 = n27464 & ~n27467 ;
  assign n27469 = n27468 ^ n25190 ^ 1'b0 ;
  assign n27470 = n6775 & ~n12539 ;
  assign n27471 = n27470 ^ n10281 ^ 1'b0 ;
  assign n27472 = ~n10963 & n27471 ;
  assign n27473 = n8122 & ~n8382 ;
  assign n27474 = n557 & n8219 ;
  assign n27475 = n27474 ^ n9388 ^ 1'b0 ;
  assign n27476 = n27473 & n27475 ;
  assign n27477 = n27476 ^ n11775 ^ n7092 ;
  assign n27478 = ~n12183 & n22469 ;
  assign n27479 = ( n1374 & n3232 ) | ( n1374 & n10010 ) | ( n3232 & n10010 ) ;
  assign n27480 = n2722 & ~n27479 ;
  assign n27481 = n1541 & n27480 ;
  assign n27482 = n15532 ^ n5241 ^ 1'b0 ;
  assign n27484 = n2914 | n3139 ;
  assign n27485 = n27484 ^ n16213 ^ 1'b0 ;
  assign n27483 = n7128 | n15661 ;
  assign n27486 = n27485 ^ n27483 ^ n16565 ;
  assign n27487 = n8008 ^ n4286 ^ 1'b0 ;
  assign n27490 = n7835 & n17185 ;
  assign n27488 = n6053 ^ n5411 ^ 1'b0 ;
  assign n27489 = n4153 & ~n27488 ;
  assign n27491 = n27490 ^ n27489 ^ 1'b0 ;
  assign n27492 = ~n17836 & n27491 ;
  assign n27493 = n14757 ^ n12500 ^ 1'b0 ;
  assign n27494 = n19159 & ~n27493 ;
  assign n27495 = ( n552 & n5199 ) | ( n552 & ~n8261 ) | ( n5199 & ~n8261 ) ;
  assign n27496 = n15489 & n27495 ;
  assign n27497 = n2645 | n8142 ;
  assign n27498 = n16470 & n26008 ;
  assign n27499 = n21941 ^ n8545 ^ 1'b0 ;
  assign n27500 = n1613 & n27499 ;
  assign n27501 = n17778 | n23192 ;
  assign n27502 = n27501 ^ n20213 ^ 1'b0 ;
  assign n27503 = ( ~n4271 & n7812 ) | ( ~n4271 & n27502 ) | ( n7812 & n27502 ) ;
  assign n27504 = n4550 | n4645 ;
  assign n27505 = n27504 ^ n4785 ^ 1'b0 ;
  assign n27506 = ( ~n5712 & n13550 ) | ( ~n5712 & n27505 ) | ( n13550 & n27505 ) ;
  assign n27507 = n14116 ^ n8626 ^ 1'b0 ;
  assign n27508 = n1574 | n16066 ;
  assign n27509 = x38 | n27508 ;
  assign n27510 = ( n5518 & ~n27507 ) | ( n5518 & n27509 ) | ( ~n27507 & n27509 ) ;
  assign n27511 = x146 & ~n9176 ;
  assign n27512 = ~n3604 & n27511 ;
  assign n27513 = x141 & ~n1497 ;
  assign n27514 = n27513 ^ n3543 ^ 1'b0 ;
  assign n27515 = n27514 ^ n13062 ^ n7380 ;
  assign n27516 = n23526 | n27515 ;
  assign n27517 = n24356 ^ n14984 ^ 1'b0 ;
  assign n27518 = n27517 ^ n7361 ^ 1'b0 ;
  assign n27519 = ~n15704 & n27518 ;
  assign n27520 = ( n354 & n14045 ) | ( n354 & ~n16668 ) | ( n14045 & ~n16668 ) ;
  assign n27521 = n23947 & ~n27520 ;
  assign n27524 = ~n6789 & n9640 ;
  assign n27525 = ~n4467 & n17273 ;
  assign n27526 = n27524 & n27525 ;
  assign n27527 = n27130 & n27526 ;
  assign n27522 = n1216 | n1576 ;
  assign n27523 = n27522 ^ n12300 ^ 1'b0 ;
  assign n27528 = n27527 ^ n27523 ^ 1'b0 ;
  assign n27529 = ~n6272 & n8900 ;
  assign n27530 = n27529 ^ n13619 ^ 1'b0 ;
  assign n27531 = n1133 | n27530 ;
  assign n27532 = ~n11187 & n27531 ;
  assign n27533 = n27532 ^ n19104 ^ 1'b0 ;
  assign n27534 = n27533 ^ n1046 ^ 1'b0 ;
  assign n27536 = n22291 ^ n12034 ^ 1'b0 ;
  assign n27537 = n4269 & n27536 ;
  assign n27538 = n25002 | n27537 ;
  assign n27535 = n4639 | n13887 ;
  assign n27539 = n27538 ^ n27535 ^ 1'b0 ;
  assign n27540 = n20572 ^ n1951 ^ 1'b0 ;
  assign n27541 = n23570 & ~n27540 ;
  assign n27542 = n13249 & n27541 ;
  assign n27543 = n1442 ^ x39 ^ 1'b0 ;
  assign n27544 = n9637 | n27543 ;
  assign n27545 = n27544 ^ n15161 ^ 1'b0 ;
  assign n27546 = n16652 & n27545 ;
  assign n27547 = n9148 ^ n2722 ^ 1'b0 ;
  assign n27548 = n27547 ^ n12610 ^ 1'b0 ;
  assign n27549 = n7915 ^ n2762 ^ 1'b0 ;
  assign n27550 = n20694 | n27549 ;
  assign n27551 = ~n5580 & n17531 ;
  assign n27552 = n1407 & ~n3899 ;
  assign n27553 = n27551 & n27552 ;
  assign n27554 = n10535 & n27553 ;
  assign n27555 = n10859 | n27554 ;
  assign n27556 = n21020 & ~n27555 ;
  assign n27557 = n18832 ^ n17764 ^ 1'b0 ;
  assign n27558 = n6565 & ~n14877 ;
  assign n27559 = n27557 & n27558 ;
  assign n27563 = ~n519 & n13368 ;
  assign n27560 = n22154 ^ n14948 ^ 1'b0 ;
  assign n27561 = n19701 & ~n27560 ;
  assign n27562 = n8494 & n27561 ;
  assign n27564 = n27563 ^ n27562 ^ 1'b0 ;
  assign n27565 = n17507 ^ n6538 ^ n507 ;
  assign n27566 = ( n7674 & n11457 ) | ( n7674 & ~n27565 ) | ( n11457 & ~n27565 ) ;
  assign n27567 = n5308 & ~n7661 ;
  assign n27568 = ~n2638 & n27567 ;
  assign n27569 = ( n9373 & n27566 ) | ( n9373 & n27568 ) | ( n27566 & n27568 ) ;
  assign n27570 = n11796 ^ n4668 ^ 1'b0 ;
  assign n27571 = n27570 ^ n24224 ^ n5072 ;
  assign n27572 = n5112 | n12899 ;
  assign n27573 = n6913 & ~n27572 ;
  assign n27574 = n13094 | n27573 ;
  assign n27575 = n14781 & ~n27574 ;
  assign n27576 = n20518 ^ n12646 ^ 1'b0 ;
  assign n27577 = n9576 | n10821 ;
  assign n27578 = n18347 | n27577 ;
  assign n27579 = n9498 ^ x141 ^ 1'b0 ;
  assign n27580 = ( n10086 & ~n17041 ) | ( n10086 & n27579 ) | ( ~n17041 & n27579 ) ;
  assign n27581 = ( ~n3900 & n13340 ) | ( ~n3900 & n17357 ) | ( n13340 & n17357 ) ;
  assign n27582 = n18225 & ~n27581 ;
  assign n27583 = n27582 ^ n25256 ^ n5780 ;
  assign n27584 = n12421 & ~n17735 ;
  assign n27585 = n2541 & n19710 ;
  assign n27586 = n27585 ^ n1002 ^ 1'b0 ;
  assign n27587 = n13129 & n27586 ;
  assign n27588 = n1800 | n15940 ;
  assign n27589 = n27587 | n27588 ;
  assign n27590 = n13017 ^ n10220 ^ n8608 ;
  assign n27591 = ( n7554 & n16346 ) | ( n7554 & ~n20933 ) | ( n16346 & ~n20933 ) ;
  assign n27592 = n10998 ^ n10422 ^ 1'b0 ;
  assign n27594 = n1880 & n10056 ;
  assign n27595 = n12193 ^ n3609 ^ 1'b0 ;
  assign n27596 = ( n22679 & n27594 ) | ( n22679 & ~n27595 ) | ( n27594 & ~n27595 ) ;
  assign n27597 = ~n3288 & n6926 ;
  assign n27598 = n27596 & n27597 ;
  assign n27593 = n1124 | n14978 ;
  assign n27599 = n27598 ^ n27593 ^ 1'b0 ;
  assign n27600 = ~n1225 & n26841 ;
  assign n27601 = n21349 & ~n27600 ;
  assign n27604 = n2312 ^ x118 ^ 1'b0 ;
  assign n27605 = ~n4193 & n27604 ;
  assign n27602 = n4890 & n7197 ;
  assign n27603 = n22110 | n27602 ;
  assign n27606 = n27605 ^ n27603 ^ 1'b0 ;
  assign n27607 = n1991 ^ n1228 ^ 1'b0 ;
  assign n27608 = n25221 & ~n27607 ;
  assign n27609 = n1789 | n3869 ;
  assign n27610 = n27609 ^ n7269 ^ n3197 ;
  assign n27611 = n904 | n19430 ;
  assign n27612 = n27611 ^ n9149 ^ 1'b0 ;
  assign n27613 = n3088 & ~n27612 ;
  assign n27614 = n27610 & n27613 ;
  assign n27615 = ( n7382 & n26120 ) | ( n7382 & ~n27614 ) | ( n26120 & ~n27614 ) ;
  assign n27616 = n27615 ^ n4365 ^ 1'b0 ;
  assign n27617 = n13701 ^ n5815 ^ 1'b0 ;
  assign n27618 = n9312 & n27617 ;
  assign n27619 = n24301 ^ n17001 ^ 1'b0 ;
  assign n27620 = n2240 & ~n27619 ;
  assign n27621 = n27620 ^ n22337 ^ n14951 ;
  assign n27622 = n6528 ^ n3590 ^ n3512 ;
  assign n27623 = n8833 ^ n7978 ^ 1'b0 ;
  assign n27624 = n8044 & n21530 ;
  assign n27625 = ~n27623 & n27624 ;
  assign n27628 = ~n6260 & n7787 ;
  assign n27629 = n27628 ^ n4690 ^ 1'b0 ;
  assign n27626 = n7566 ^ n3452 ^ 1'b0 ;
  assign n27627 = ~n1323 & n27626 ;
  assign n27630 = n27629 ^ n27627 ^ 1'b0 ;
  assign n27631 = n559 | n2590 ;
  assign n27632 = n2038 & ~n27631 ;
  assign n27633 = n27632 ^ n14773 ^ n7573 ;
  assign n27634 = n27633 ^ n24504 ^ n22358 ;
  assign n27635 = x169 & n3755 ;
  assign n27636 = n27635 ^ n2416 ^ 1'b0 ;
  assign n27637 = n16788 & ~n27636 ;
  assign n27638 = n15617 | n27637 ;
  assign n27639 = n7604 ^ n1155 ^ 1'b0 ;
  assign n27640 = ( n752 & ~n1754 ) | ( n752 & n27639 ) | ( ~n1754 & n27639 ) ;
  assign n27641 = ~n1197 & n10403 ;
  assign n27642 = n20585 ^ n5440 ^ n3190 ;
  assign n27643 = n6291 & n26057 ;
  assign n27644 = n13138 ^ n9498 ^ 1'b0 ;
  assign n27645 = n6703 & n20899 ;
  assign n27646 = ~n27644 & n27645 ;
  assign n27647 = ( n4278 & ~n9675 ) | ( n4278 & n27646 ) | ( ~n9675 & n27646 ) ;
  assign n27648 = n27647 ^ n19247 ^ 1'b0 ;
  assign n27649 = n9736 & ~n22234 ;
  assign n27650 = n8430 & n27649 ;
  assign n27651 = n5801 & n11489 ;
  assign n27652 = n27651 ^ n16817 ^ 1'b0 ;
  assign n27653 = n7380 & ~n14013 ;
  assign n27654 = n27652 & n27653 ;
  assign n27655 = n27654 ^ n2333 ^ 1'b0 ;
  assign n27656 = ~n1321 & n14018 ;
  assign n27657 = n22009 ^ n19711 ^ 1'b0 ;
  assign n27658 = n27656 & n27657 ;
  assign n27659 = n18954 ^ n3125 ^ 1'b0 ;
  assign n27660 = n27659 ^ n10234 ^ 1'b0 ;
  assign n27661 = n27615 & n27660 ;
  assign n27662 = n19869 ^ n5593 ^ 1'b0 ;
  assign n27663 = n21022 | n26241 ;
  assign n27664 = n2771 & ~n27663 ;
  assign n27665 = n27664 ^ n24931 ^ 1'b0 ;
  assign n27666 = n15469 & ~n27665 ;
  assign n27667 = n15031 & ~n27666 ;
  assign n27668 = ~n1842 & n24890 ;
  assign n27669 = ( n4675 & n10984 ) | ( n4675 & ~n25327 ) | ( n10984 & ~n25327 ) ;
  assign n27670 = n10611 & ~n27669 ;
  assign n27671 = n27668 & n27670 ;
  assign n27672 = n27667 & n27671 ;
  assign n27673 = n27672 ^ n27149 ^ n15625 ;
  assign n27674 = ( n4371 & ~n12558 ) | ( n4371 & n15924 ) | ( ~n12558 & n15924 ) ;
  assign n27675 = n6669 | n27674 ;
  assign n27676 = n7159 | n12422 ;
  assign n27677 = ~n3172 & n17663 ;
  assign n27678 = n18962 & n27677 ;
  assign n27679 = n5261 & ~n16497 ;
  assign n27680 = n27679 ^ n18192 ^ 1'b0 ;
  assign n27681 = n10764 ^ n1936 ^ 1'b0 ;
  assign n27682 = n16255 & n27681 ;
  assign n27683 = n13896 & ~n27682 ;
  assign n27684 = n6485 ^ n6444 ^ 1'b0 ;
  assign n27685 = ~n2875 & n27684 ;
  assign n27686 = n13853 ^ n12885 ^ 1'b0 ;
  assign n27687 = n14489 & n27686 ;
  assign n27688 = ( n26386 & n27685 ) | ( n26386 & n27687 ) | ( n27685 & n27687 ) ;
  assign n27691 = n13135 ^ n6056 ^ n2940 ;
  assign n27689 = n1671 ^ n914 ^ x124 ;
  assign n27690 = n23483 | n27689 ;
  assign n27692 = n27691 ^ n27690 ^ 1'b0 ;
  assign n27693 = n8129 ^ n4455 ^ 1'b0 ;
  assign n27694 = n4072 & ~n27693 ;
  assign n27695 = n5690 & n27694 ;
  assign n27696 = n8045 | n27695 ;
  assign n27697 = ( n11076 & n14246 ) | ( n11076 & ~n16581 ) | ( n14246 & ~n16581 ) ;
  assign n27698 = n27697 ^ n20678 ^ 1'b0 ;
  assign n27699 = n6511 | n27698 ;
  assign n27700 = n4670 & ~n17906 ;
  assign n27701 = ~n5936 & n27700 ;
  assign n27702 = n11331 ^ n7747 ^ n3045 ;
  assign n27703 = n27702 ^ n8683 ^ 1'b0 ;
  assign n27704 = n22124 ^ n7626 ^ n344 ;
  assign n27705 = n1763 | n13559 ;
  assign n27706 = n7293 & ~n18306 ;
  assign n27707 = n27706 ^ n7440 ^ 1'b0 ;
  assign n27708 = n20707 & ~n27707 ;
  assign n27709 = n27708 ^ n15183 ^ 1'b0 ;
  assign n27710 = ( ~n7715 & n27705 ) | ( ~n7715 & n27709 ) | ( n27705 & n27709 ) ;
  assign n27711 = n14796 ^ n9411 ^ 1'b0 ;
  assign n27712 = n26697 ^ n3496 ^ 1'b0 ;
  assign n27713 = n23898 & ~n26755 ;
  assign n27714 = ( n3568 & ~n12511 ) | ( n3568 & n27713 ) | ( ~n12511 & n27713 ) ;
  assign n27715 = n25730 ^ n13174 ^ n8799 ;
  assign n27716 = n12543 & ~n21892 ;
  assign n27717 = n18053 & n27716 ;
  assign n27718 = n3455 & n26303 ;
  assign n27719 = n27718 ^ n23013 ^ 1'b0 ;
  assign n27720 = n11321 & n26230 ;
  assign n27721 = n4882 & n27720 ;
  assign n27722 = n9823 ^ n1367 ^ 1'b0 ;
  assign n27723 = n9944 | n27722 ;
  assign n27724 = n27723 ^ n2722 ^ 1'b0 ;
  assign n27725 = n8764 & n27724 ;
  assign n27726 = n21259 & n27725 ;
  assign n27727 = ~n12191 & n27726 ;
  assign n27728 = n8533 | n27727 ;
  assign n27729 = n6195 | n9732 ;
  assign n27730 = n27729 ^ n649 ^ 1'b0 ;
  assign n27731 = ( n1432 & ~n5862 ) | ( n1432 & n27730 ) | ( ~n5862 & n27730 ) ;
  assign n27733 = n17108 ^ n13309 ^ n1035 ;
  assign n27734 = ~n10945 & n27733 ;
  assign n27732 = n15010 ^ n4034 ^ 1'b0 ;
  assign n27735 = n27734 ^ n27732 ^ 1'b0 ;
  assign n27736 = ~n23387 & n27735 ;
  assign n27737 = ~n2133 & n23468 ;
  assign n27738 = n27736 & n27737 ;
  assign n27739 = n7308 ^ n4480 ^ 1'b0 ;
  assign n27740 = n16452 & ~n27739 ;
  assign n27741 = n27740 ^ n21830 ^ 1'b0 ;
  assign n27742 = n16385 ^ n5066 ^ 1'b0 ;
  assign n27743 = n14217 ^ n3567 ^ n1626 ;
  assign n27744 = n16809 ^ n16032 ^ 1'b0 ;
  assign n27745 = ~n13935 & n27744 ;
  assign n27746 = ~n994 & n27745 ;
  assign n27747 = n27746 ^ n14302 ^ 1'b0 ;
  assign n27748 = n27747 ^ n14971 ^ n4282 ;
  assign n27749 = n16624 ^ n1357 ^ 1'b0 ;
  assign n27750 = n5335 | n27749 ;
  assign n27751 = n5506 | n27750 ;
  assign n27752 = n22080 & ~n27751 ;
  assign n27753 = n18552 ^ n18383 ^ 1'b0 ;
  assign n27754 = ( n1468 & n5303 ) | ( n1468 & n27753 ) | ( n5303 & n27753 ) ;
  assign n27755 = n15500 ^ n1037 ^ 1'b0 ;
  assign n27756 = n1237 & n27755 ;
  assign n27757 = n13399 & n23504 ;
  assign n27758 = n5459 & ~n27757 ;
  assign n27759 = n12938 & n27758 ;
  assign n27760 = n27073 ^ n14135 ^ n1996 ;
  assign n27761 = n2961 & ~n27760 ;
  assign n27762 = n8613 & ~n27761 ;
  assign n27763 = n27762 ^ n8327 ^ 1'b0 ;
  assign n27764 = n8829 ^ n2897 ^ 1'b0 ;
  assign n27765 = n27764 ^ n5624 ^ n1000 ;
  assign n27766 = n13346 ^ n1005 ^ 1'b0 ;
  assign n27767 = ~n15109 & n27766 ;
  assign n27768 = n27767 ^ n8509 ^ n7850 ;
  assign n27769 = n7226 ^ n5069 ^ n1635 ;
  assign n27770 = n3052 & n7182 ;
  assign n27771 = n27769 & n27770 ;
  assign n27772 = n13761 ^ n12935 ^ 1'b0 ;
  assign n27773 = ( ~n17271 & n27771 ) | ( ~n17271 & n27772 ) | ( n27771 & n27772 ) ;
  assign n27774 = n6528 ^ n3452 ^ 1'b0 ;
  assign n27775 = ~n5377 & n27774 ;
  assign n27776 = ( n19987 & n26558 ) | ( n19987 & ~n27775 ) | ( n26558 & ~n27775 ) ;
  assign n27777 = ~n2709 & n14685 ;
  assign n27778 = n4724 & n9676 ;
  assign n27779 = n27778 ^ n10667 ^ 1'b0 ;
  assign n27780 = n27223 ^ n4345 ^ 1'b0 ;
  assign n27781 = n15732 | n27780 ;
  assign n27782 = n26295 ^ n17963 ^ n3312 ;
  assign n27784 = n3262 & ~n14726 ;
  assign n27783 = ~n1487 & n25145 ;
  assign n27785 = n27784 ^ n27783 ^ 1'b0 ;
  assign n27786 = x28 & n14661 ;
  assign n27787 = n27786 ^ n16641 ^ 1'b0 ;
  assign n27788 = ~n20107 & n27787 ;
  assign n27789 = n14870 ^ n11623 ^ n7564 ;
  assign n27790 = n14781 ^ n5926 ^ 1'b0 ;
  assign n27791 = ~n27789 & n27790 ;
  assign n27792 = n9352 ^ n5761 ^ 1'b0 ;
  assign n27793 = n21594 ^ n7368 ^ 1'b0 ;
  assign n27794 = ~n27792 & n27793 ;
  assign n27796 = n10449 ^ n3742 ^ n1928 ;
  assign n27797 = ~n9811 & n27796 ;
  assign n27798 = n27797 ^ n21664 ^ n591 ;
  assign n27799 = n27798 ^ n22797 ^ 1'b0 ;
  assign n27800 = n13677 | n27799 ;
  assign n27795 = n18049 & n18917 ;
  assign n27801 = n27800 ^ n27795 ^ 1'b0 ;
  assign n27802 = ~n20333 & n27801 ;
  assign n27803 = n27802 ^ n12760 ^ n6817 ;
  assign n27805 = n1202 & ~n3093 ;
  assign n27804 = n3425 ^ n1082 ^ 1'b0 ;
  assign n27806 = n27805 ^ n27804 ^ n18270 ;
  assign n27807 = ( x215 & ~n15123 ) | ( x215 & n27806 ) | ( ~n15123 & n27806 ) ;
  assign n27809 = n1717 & ~n6578 ;
  assign n27810 = n2680 & n27809 ;
  assign n27808 = n556 & n25476 ;
  assign n27811 = n27810 ^ n27808 ^ 1'b0 ;
  assign n27812 = n22325 ^ n1964 ^ 1'b0 ;
  assign n27813 = n14575 | n27812 ;
  assign n27816 = n10859 | n25572 ;
  assign n27814 = n8598 ^ n1605 ^ 1'b0 ;
  assign n27815 = n15274 & ~n27814 ;
  assign n27817 = n27816 ^ n27815 ^ 1'b0 ;
  assign n27818 = n12457 ^ n11631 ^ 1'b0 ;
  assign n27819 = n27817 & ~n27818 ;
  assign n27820 = n18443 ^ x104 ^ 1'b0 ;
  assign n27821 = n10904 & n15606 ;
  assign n27822 = n15327 ^ n13915 ^ 1'b0 ;
  assign n27823 = n23265 & ~n27822 ;
  assign n27824 = ( n27820 & ~n27821 ) | ( n27820 & n27823 ) | ( ~n27821 & n27823 ) ;
  assign n27825 = n21755 & ~n27674 ;
  assign n27826 = ~n895 & n27825 ;
  assign n27827 = n4202 & ~n5263 ;
  assign n27828 = n27827 ^ n1672 ^ 1'b0 ;
  assign n27829 = ~n9762 & n27828 ;
  assign n27830 = ~n12804 & n27829 ;
  assign n27831 = n3500 & n8900 ;
  assign n27832 = n15110 & n27831 ;
  assign n27833 = ( n21164 & n27654 ) | ( n21164 & ~n27832 ) | ( n27654 & ~n27832 ) ;
  assign n27834 = n787 | n12843 ;
  assign n27835 = n27834 ^ n19926 ^ 1'b0 ;
  assign n27836 = n8999 | n27835 ;
  assign n27837 = n21387 | n27836 ;
  assign n27838 = ~n1961 & n2822 ;
  assign n27839 = n27838 ^ n844 ^ 1'b0 ;
  assign n27840 = n12479 & n27839 ;
  assign n27842 = ~n1397 & n3237 ;
  assign n27841 = ~n13244 & n20548 ;
  assign n27843 = n27842 ^ n27841 ^ n14870 ;
  assign n27844 = n23072 ^ n6240 ^ 1'b0 ;
  assign n27845 = n21557 ^ n3640 ^ 1'b0 ;
  assign n27846 = n17558 ^ n6300 ^ 1'b0 ;
  assign n27847 = n1398 & n27846 ;
  assign n27848 = n18293 & n27847 ;
  assign n27849 = n27848 ^ n23096 ^ 1'b0 ;
  assign n27850 = ( n9743 & n15527 ) | ( n9743 & ~n16819 ) | ( n15527 & ~n16819 ) ;
  assign n27852 = n13988 ^ n12848 ^ n2904 ;
  assign n27851 = ~n5073 & n6335 ;
  assign n27853 = n27852 ^ n27851 ^ 1'b0 ;
  assign n27854 = n14002 | n27853 ;
  assign n27855 = n1847 & n5199 ;
  assign n27856 = ~n18092 & n27855 ;
  assign n27857 = n26323 ^ n13974 ^ 1'b0 ;
  assign n27858 = n16669 | n27857 ;
  assign n27859 = n1979 ^ n390 ^ 1'b0 ;
  assign n27860 = n27859 ^ n12691 ^ n10531 ;
  assign n27861 = ( ~n13895 & n17447 ) | ( ~n13895 & n27860 ) | ( n17447 & n27860 ) ;
  assign n27862 = n27861 ^ n10226 ^ 1'b0 ;
  assign n27863 = n15991 ^ n13390 ^ n10448 ;
  assign n27864 = n6225 | n26407 ;
  assign n27865 = n11435 ^ n4332 ^ 1'b0 ;
  assign n27866 = ( n966 & ~n12504 ) | ( n966 & n27865 ) | ( ~n12504 & n27865 ) ;
  assign n27867 = n27866 ^ n7210 ^ 1'b0 ;
  assign n27868 = n26319 | n27867 ;
  assign n27869 = n27868 ^ n20634 ^ 1'b0 ;
  assign n27870 = n7732 ^ n4519 ^ n3267 ;
  assign n27871 = n17617 ^ n15542 ^ n1729 ;
  assign n27872 = n15018 | n27871 ;
  assign n27873 = n27872 ^ n6674 ^ 1'b0 ;
  assign n27874 = n19580 ^ n7503 ^ 1'b0 ;
  assign n27875 = n539 & ~n7746 ;
  assign n27876 = n18256 | n27875 ;
  assign n27877 = n12930 & n20164 ;
  assign n27878 = n8457 ^ n3188 ^ 1'b0 ;
  assign n27879 = n3919 | n27878 ;
  assign n27880 = ( n945 & n9271 ) | ( n945 & n27879 ) | ( n9271 & n27879 ) ;
  assign n27881 = n27880 ^ n3312 ^ 1'b0 ;
  assign n27882 = ~x167 & n1563 ;
  assign n27883 = n14878 & n27435 ;
  assign n27884 = ( n14011 & n21671 ) | ( n14011 & n27883 ) | ( n21671 & n27883 ) ;
  assign n27886 = n14188 & n17023 ;
  assign n27885 = n602 & ~n9659 ;
  assign n27887 = n27886 ^ n27885 ^ 1'b0 ;
  assign n27888 = n21603 ^ n15662 ^ n459 ;
  assign n27889 = n27887 & ~n27888 ;
  assign n27890 = n25497 ^ n10323 ^ 1'b0 ;
  assign n27891 = n22154 ^ n9331 ^ 1'b0 ;
  assign n27892 = n7468 & ~n12895 ;
  assign n27893 = n27892 ^ n6399 ^ 1'b0 ;
  assign n27894 = n27893 ^ n8922 ^ 1'b0 ;
  assign n27895 = ( n827 & n4694 ) | ( n827 & ~n27894 ) | ( n4694 & ~n27894 ) ;
  assign n27896 = ( n27890 & ~n27891 ) | ( n27890 & n27895 ) | ( ~n27891 & n27895 ) ;
  assign n27897 = n11063 ^ n6827 ^ n4080 ;
  assign n27898 = ~n5858 & n17531 ;
  assign n27899 = n12503 & ~n27898 ;
  assign n27900 = n2359 & n7001 ;
  assign n27901 = n18303 ^ n17963 ^ n16627 ;
  assign n27902 = n21190 ^ n8051 ^ n7904 ;
  assign n27903 = n27902 ^ n382 ^ 1'b0 ;
  assign n27904 = n11172 & ~n27903 ;
  assign n27905 = n9604 ^ n3648 ^ 1'b0 ;
  assign n27906 = n7697 & n27905 ;
  assign n27907 = ( n10191 & n21027 ) | ( n10191 & ~n23427 ) | ( n21027 & ~n23427 ) ;
  assign n27908 = n27906 & ~n27907 ;
  assign n27909 = n5938 & n27908 ;
  assign n27910 = n2860 | n14382 ;
  assign n27911 = n27910 ^ n2267 ^ 1'b0 ;
  assign n27912 = n13012 | n27911 ;
  assign n27913 = n9797 ^ n1975 ^ 1'b0 ;
  assign n27914 = n27912 | n27913 ;
  assign n27915 = n25671 ^ n12491 ^ 1'b0 ;
  assign n27916 = ~n956 & n3081 ;
  assign n27917 = n13066 | n27916 ;
  assign n27918 = n27917 ^ n2596 ^ 1'b0 ;
  assign n27919 = n8908 & ~n26657 ;
  assign n27920 = ( ~n8348 & n19409 ) | ( ~n8348 & n27919 ) | ( n19409 & n27919 ) ;
  assign n27922 = ~n17303 & n21351 ;
  assign n27923 = n1284 & n27922 ;
  assign n27921 = ( n3414 & n5637 ) | ( n3414 & ~n20275 ) | ( n5637 & ~n20275 ) ;
  assign n27924 = n27923 ^ n27921 ^ 1'b0 ;
  assign n27925 = n6082 | n9118 ;
  assign n27926 = n21762 ^ n12685 ^ n5189 ;
  assign n27927 = n12451 & n27926 ;
  assign n27928 = n4477 & n27927 ;
  assign n27929 = n27928 ^ n671 ^ 1'b0 ;
  assign n27930 = n17033 ^ n10230 ^ 1'b0 ;
  assign n27931 = n6193 & n27930 ;
  assign n27932 = n4630 & ~n5524 ;
  assign n27933 = n18416 & ~n27932 ;
  assign n27934 = n12478 & ~n27933 ;
  assign n27935 = n4388 | n7929 ;
  assign n27936 = ( ~n2560 & n4744 ) | ( ~n2560 & n27935 ) | ( n4744 & n27935 ) ;
  assign n27937 = n27936 ^ n3792 ^ 1'b0 ;
  assign n27938 = n2215 & ~n27937 ;
  assign n27939 = n27938 ^ n12744 ^ 1'b0 ;
  assign n27940 = ~n4189 & n7002 ;
  assign n27941 = n10713 & n27940 ;
  assign n27942 = n27941 ^ n22912 ^ n8755 ;
  assign n27943 = n3731 & n27942 ;
  assign n27944 = ~n27939 & n27943 ;
  assign n27945 = n18240 ^ n7570 ^ 1'b0 ;
  assign n27946 = n17257 ^ n11679 ^ 1'b0 ;
  assign n27947 = ~n4114 & n27946 ;
  assign n27948 = ~n3414 & n5351 ;
  assign n27949 = n3320 & ~n27948 ;
  assign n27950 = n5573 & ~n5699 ;
  assign n27951 = ~n3792 & n27950 ;
  assign n27952 = n27951 ^ n14781 ^ n4290 ;
  assign n27953 = n19709 ^ n15865 ^ 1'b0 ;
  assign n27954 = ~n3526 & n27953 ;
  assign n27955 = n27954 ^ n10021 ^ 1'b0 ;
  assign n27956 = n23862 ^ n8000 ^ 1'b0 ;
  assign n27957 = n1727 & n23885 ;
  assign n27958 = ~n20501 & n27957 ;
  assign n27959 = n898 & ~n3042 ;
  assign n27962 = n12587 ^ n11211 ^ 1'b0 ;
  assign n27963 = n18862 & ~n27962 ;
  assign n27964 = ~n22923 & n27963 ;
  assign n27965 = ~n1452 & n27964 ;
  assign n27960 = ~n297 & n11276 ;
  assign n27961 = n12362 & ~n27960 ;
  assign n27966 = n27965 ^ n27961 ^ 1'b0 ;
  assign n27967 = x189 & ~n10092 ;
  assign n27968 = n27967 ^ n15638 ^ 1'b0 ;
  assign n27969 = n6175 | n27968 ;
  assign n27970 = n27969 ^ n15590 ^ 1'b0 ;
  assign n27971 = n9868 ^ n5926 ^ 1'b0 ;
  assign n27972 = ( n16293 & n22701 ) | ( n16293 & ~n27971 ) | ( n22701 & ~n27971 ) ;
  assign n27973 = n27921 & ~n27972 ;
  assign n27974 = n27973 ^ n22680 ^ 1'b0 ;
  assign n27975 = ( ~n256 & n6846 ) | ( ~n256 & n17542 ) | ( n6846 & n17542 ) ;
  assign n27976 = n13147 ^ n3338 ^ 1'b0 ;
  assign n27977 = ~n27975 & n27976 ;
  assign n27978 = ( x189 & n27974 ) | ( x189 & n27977 ) | ( n27974 & n27977 ) ;
  assign n27979 = ~n20332 & n27978 ;
  assign n27980 = ( n5850 & n9840 ) | ( n5850 & ~n12837 ) | ( n9840 & ~n12837 ) ;
  assign n27981 = n27980 ^ n16103 ^ x23 ;
  assign n27982 = n6213 | n21108 ;
  assign n27983 = n2118 ^ n1543 ^ 1'b0 ;
  assign n27984 = n2083 & ~n27983 ;
  assign n27985 = ( ~n17375 & n20680 ) | ( ~n17375 & n27984 ) | ( n20680 & n27984 ) ;
  assign n27986 = n12147 ^ n8936 ^ 1'b0 ;
  assign n27987 = n27986 ^ n1650 ^ x207 ;
  assign n27988 = ~n26833 & n27987 ;
  assign n27989 = n19565 | n24927 ;
  assign n27999 = n26903 ^ n24541 ^ n7855 ;
  assign n28000 = n27999 ^ n18057 ^ 1'b0 ;
  assign n27990 = n5387 | n7762 ;
  assign n27991 = ( n6006 & n19174 ) | ( n6006 & n27990 ) | ( n19174 & n27990 ) ;
  assign n27992 = n15257 & ~n27991 ;
  assign n27993 = ~n8740 & n27992 ;
  assign n27994 = n16397 & ~n27993 ;
  assign n27995 = ~n3140 & n27994 ;
  assign n27996 = n8813 ^ n424 ^ 1'b0 ;
  assign n27997 = n27996 ^ n23154 ^ n2005 ;
  assign n27998 = n27995 | n27997 ;
  assign n28001 = n28000 ^ n27998 ^ 1'b0 ;
  assign n28002 = n17848 & ~n18852 ;
  assign n28003 = n8903 & n28002 ;
  assign n28004 = n2191 & ~n26908 ;
  assign n28005 = ~n6448 & n20252 ;
  assign n28006 = n21343 & n27415 ;
  assign n28007 = n18366 & n28006 ;
  assign n28008 = ~n15167 & n28007 ;
  assign n28009 = ~n5178 & n5809 ;
  assign n28010 = n12281 & n28009 ;
  assign n28011 = ( n7471 & n21985 ) | ( n7471 & n28010 ) | ( n21985 & n28010 ) ;
  assign n28012 = ~n2887 & n19124 ;
  assign n28013 = n28012 ^ n27185 ^ 1'b0 ;
  assign n28014 = ~n11701 & n23822 ;
  assign n28015 = n20603 ^ n10680 ^ n7282 ;
  assign n28016 = ( n1487 & n8907 ) | ( n1487 & ~n18628 ) | ( n8907 & ~n18628 ) ;
  assign n28019 = n7990 ^ n3261 ^ 1'b0 ;
  assign n28017 = n1350 | n5679 ;
  assign n28018 = n22948 | n28017 ;
  assign n28020 = n28019 ^ n28018 ^ n8754 ;
  assign n28026 = n15971 ^ n2705 ^ 1'b0 ;
  assign n28027 = n17825 & n28026 ;
  assign n28021 = n10629 ^ n7827 ^ n391 ;
  assign n28022 = n7883 & ~n28021 ;
  assign n28023 = ~n17493 & n28022 ;
  assign n28024 = n10010 & n28023 ;
  assign n28025 = n7024 | n28024 ;
  assign n28028 = n28027 ^ n28025 ^ 1'b0 ;
  assign n28029 = ( ~n5891 & n28020 ) | ( ~n5891 & n28028 ) | ( n28020 & n28028 ) ;
  assign n28030 = n2661 & ~n28029 ;
  assign n28031 = n3848 & n15707 ;
  assign n28032 = n1807 & n28031 ;
  assign n28033 = n17763 ^ n6065 ^ 1'b0 ;
  assign n28034 = n28033 ^ n18715 ^ n18139 ;
  assign n28035 = n2764 & n10606 ;
  assign n28036 = n28035 ^ n26588 ^ n21955 ;
  assign n28038 = n20665 ^ n2536 ^ 1'b0 ;
  assign n28039 = n7795 & n28038 ;
  assign n28037 = n2359 | n20544 ;
  assign n28040 = n28039 ^ n28037 ^ 1'b0 ;
  assign n28041 = n1761 & n21339 ;
  assign n28042 = ~n12939 & n28041 ;
  assign n28043 = n3335 | n11852 ;
  assign n28044 = n28043 ^ n645 ^ 1'b0 ;
  assign n28045 = n8099 ^ n7670 ^ 1'b0 ;
  assign n28046 = n28045 ^ n14322 ^ n13793 ;
  assign n28047 = ( ~n26856 & n28044 ) | ( ~n26856 & n28046 ) | ( n28044 & n28046 ) ;
  assign n28048 = n25726 ^ n18961 ^ 1'b0 ;
  assign n28049 = ~n3211 & n20023 ;
  assign n28050 = n18091 & ~n28049 ;
  assign n28051 = ~n4454 & n28050 ;
  assign n28052 = ( n1838 & n27341 ) | ( n1838 & n28051 ) | ( n27341 & n28051 ) ;
  assign n28053 = n13622 ^ n12029 ^ n10351 ;
  assign n28054 = n13046 | n28053 ;
  assign n28055 = n28054 ^ n11750 ^ 1'b0 ;
  assign n28056 = ~n3610 & n18189 ;
  assign n28057 = ~n21283 & n28056 ;
  assign n28058 = ~n1729 & n3541 ;
  assign n28059 = ( ~n17769 & n19167 ) | ( ~n17769 & n28058 ) | ( n19167 & n28058 ) ;
  assign n28060 = n11342 & n11366 ;
  assign n28061 = n16044 ^ n10396 ^ 1'b0 ;
  assign n28062 = n22131 & ~n28061 ;
  assign n28063 = ( n2950 & ~n21474 ) | ( n2950 & n28062 ) | ( ~n21474 & n28062 ) ;
  assign n28064 = ~n6816 & n28063 ;
  assign n28065 = n28064 ^ n8165 ^ 1'b0 ;
  assign n28066 = n16731 ^ n9048 ^ n3269 ;
  assign n28067 = n26033 & ~n28066 ;
  assign n28068 = n24726 & n24899 ;
  assign n28069 = n1356 | n9302 ;
  assign n28070 = n12084 | n28069 ;
  assign n28071 = n4600 | n13892 ;
  assign n28072 = n28070 | n28071 ;
  assign n28073 = n18725 ^ n14654 ^ 1'b0 ;
  assign n28074 = n17894 | n28073 ;
  assign n28075 = n2985 ^ n503 ^ 1'b0 ;
  assign n28076 = n11397 ^ n2050 ^ 1'b0 ;
  assign n28077 = n5975 & ~n28076 ;
  assign n28078 = n28077 ^ n11437 ^ 1'b0 ;
  assign n28079 = n28075 & n28078 ;
  assign n28080 = n28079 ^ n1048 ^ 1'b0 ;
  assign n28081 = n21015 & n25358 ;
  assign n28082 = n20166 ^ n4464 ^ 1'b0 ;
  assign n28083 = n28082 ^ n10171 ^ 1'b0 ;
  assign n28084 = n27335 & n28083 ;
  assign n28085 = ~n25613 & n28084 ;
  assign n28086 = n8682 & n28085 ;
  assign n28087 = n28086 ^ n10708 ^ n7345 ;
  assign n28088 = n17874 ^ n5681 ^ 1'b0 ;
  assign n28089 = n3069 | n18519 ;
  assign n28090 = n10899 | n28089 ;
  assign n28091 = n28090 ^ n7619 ^ n1550 ;
  assign n28092 = n20486 ^ n16409 ^ 1'b0 ;
  assign n28093 = ~n5998 & n28092 ;
  assign n28094 = n5193 ^ n2136 ^ 1'b0 ;
  assign n28095 = n9498 ^ n2784 ^ 1'b0 ;
  assign n28098 = ~n17301 & n19388 ;
  assign n28099 = n28098 ^ n8111 ^ 1'b0 ;
  assign n28096 = n21792 ^ n14903 ^ n8657 ;
  assign n28097 = n1702 & n28096 ;
  assign n28100 = n28099 ^ n28097 ^ 1'b0 ;
  assign n28101 = ~n28095 & n28100 ;
  assign n28102 = n8578 ^ n801 ^ 1'b0 ;
  assign n28103 = n17275 & n28102 ;
  assign n28104 = n10189 ^ n10145 ^ 1'b0 ;
  assign n28105 = n14436 | n28104 ;
  assign n28106 = n28105 ^ n2644 ^ 1'b0 ;
  assign n28107 = ~n9506 & n11554 ;
  assign n28108 = n28107 ^ n18251 ^ n8114 ;
  assign n28109 = ~n4861 & n21319 ;
  assign n28110 = n24344 ^ n5003 ^ 1'b0 ;
  assign n28111 = n1578 & ~n28110 ;
  assign n28112 = n16085 ^ n427 ^ 1'b0 ;
  assign n28113 = n16508 ^ n15988 ^ 1'b0 ;
  assign n28114 = ( ~n1593 & n6315 ) | ( ~n1593 & n28113 ) | ( n6315 & n28113 ) ;
  assign n28115 = n12032 ^ n3632 ^ 1'b0 ;
  assign n28117 = n8745 & ~n17042 ;
  assign n28118 = n12561 & n28117 ;
  assign n28116 = ~n15407 & n19066 ;
  assign n28119 = n28118 ^ n28116 ^ 1'b0 ;
  assign n28121 = n1863 | n10598 ;
  assign n28122 = n28121 ^ n14798 ^ 1'b0 ;
  assign n28120 = n8386 | n11028 ;
  assign n28123 = n28122 ^ n28120 ^ 1'b0 ;
  assign n28124 = n2494 | n10134 ;
  assign n28125 = n28124 ^ n7812 ^ 1'b0 ;
  assign n28126 = n18092 & ~n28125 ;
  assign n28127 = n8693 ^ n3447 ^ n3375 ;
  assign n28128 = n8774 & ~n20399 ;
  assign n28129 = ~n28127 & n28128 ;
  assign n28130 = n12104 | n28129 ;
  assign n28131 = n28130 ^ n6677 ^ 1'b0 ;
  assign n28132 = ( n3472 & n10659 ) | ( n3472 & ~n28131 ) | ( n10659 & ~n28131 ) ;
  assign n28133 = n2502 ^ n604 ^ 1'b0 ;
  assign n28134 = n28132 | n28133 ;
  assign n28135 = n18635 ^ n7974 ^ 1'b0 ;
  assign n28136 = n702 & n28135 ;
  assign n28137 = n22770 & ~n26008 ;
  assign n28138 = ~n28136 & n28137 ;
  assign n28139 = n1067 & n10694 ;
  assign n28140 = n6734 & n28139 ;
  assign n28141 = n28140 ^ n15750 ^ 1'b0 ;
  assign n28142 = n10135 & n23738 ;
  assign n28145 = n14334 & n16898 ;
  assign n28146 = ~n11545 & n28145 ;
  assign n28147 = n28146 ^ n11920 ^ 1'b0 ;
  assign n28148 = n9778 | n28147 ;
  assign n28143 = n14762 ^ n7298 ^ 1'b0 ;
  assign n28144 = n2883 | n28143 ;
  assign n28149 = n28148 ^ n28144 ^ 1'b0 ;
  assign n28150 = n3847 & n7869 ;
  assign n28151 = n9868 & n27919 ;
  assign n28152 = n20143 & n28151 ;
  assign n28156 = n8473 | n11767 ;
  assign n28157 = n28156 ^ n8897 ^ 1'b0 ;
  assign n28153 = n358 | n7483 ;
  assign n28154 = n28153 ^ n1742 ^ 1'b0 ;
  assign n28155 = n23360 & ~n28154 ;
  assign n28158 = n28157 ^ n28155 ^ 1'b0 ;
  assign n28159 = n706 & n1634 ;
  assign n28160 = n10178 & n28159 ;
  assign n28161 = ( n4686 & n22693 ) | ( n4686 & n23335 ) | ( n22693 & n23335 ) ;
  assign n28162 = ( n2468 & ~n4931 ) | ( n2468 & n25045 ) | ( ~n4931 & n25045 ) ;
  assign n28163 = n14878 & ~n25220 ;
  assign n28164 = n7772 ^ n409 ^ 1'b0 ;
  assign n28165 = n14907 & ~n28164 ;
  assign n28166 = n20979 ^ n7794 ^ 1'b0 ;
  assign n28167 = n16627 & n28166 ;
  assign n28168 = n26789 | n28167 ;
  assign n28169 = n13050 & ~n28168 ;
  assign n28170 = n750 | n1489 ;
  assign n28171 = n22626 & ~n28170 ;
  assign n28172 = ~n1521 & n24270 ;
  assign n28173 = ( n5781 & n12129 ) | ( n5781 & ~n28172 ) | ( n12129 & ~n28172 ) ;
  assign n28174 = n9809 | n15722 ;
  assign n28175 = n28174 ^ n21154 ^ 1'b0 ;
  assign n28176 = n7897 ^ n4039 ^ x11 ;
  assign n28177 = n22852 ^ n323 ^ 1'b0 ;
  assign n28178 = n3923 | n13967 ;
  assign n28179 = ( n16197 & ~n20519 ) | ( n16197 & n28178 ) | ( ~n20519 & n28178 ) ;
  assign n28180 = n28179 ^ n21154 ^ 1'b0 ;
  assign n28181 = ~n14497 & n28180 ;
  assign n28182 = n28181 ^ x230 ^ 1'b0 ;
  assign n28183 = ~n19397 & n28182 ;
  assign n28184 = n12582 & n22743 ;
  assign n28185 = n8398 & n28184 ;
  assign n28189 = n12776 ^ n1129 ^ n286 ;
  assign n28190 = n3070 & ~n28189 ;
  assign n28186 = n21372 ^ n9431 ^ 1'b0 ;
  assign n28187 = n1024 | n28186 ;
  assign n28188 = ( n11161 & ~n17124 ) | ( n11161 & n28187 ) | ( ~n17124 & n28187 ) ;
  assign n28191 = n28190 ^ n28188 ^ n3057 ;
  assign n28192 = n7366 & ~n28191 ;
  assign n28193 = n28185 & n28192 ;
  assign n28196 = n1045 & n3693 ;
  assign n28194 = n9153 ^ n2513 ^ 1'b0 ;
  assign n28195 = n3102 & n28194 ;
  assign n28197 = n28196 ^ n28195 ^ 1'b0 ;
  assign n28198 = n16128 ^ n11054 ^ n2788 ;
  assign n28199 = ( n11767 & ~n27385 ) | ( n11767 & n28198 ) | ( ~n27385 & n28198 ) ;
  assign n28200 = n8004 ^ n1791 ^ 1'b0 ;
  assign n28201 = n300 & n28200 ;
  assign n28202 = n2427 & n7208 ;
  assign n28203 = n19940 & n28202 ;
  assign n28204 = ( n6689 & n28201 ) | ( n6689 & n28203 ) | ( n28201 & n28203 ) ;
  assign n28205 = x121 | n4612 ;
  assign n28206 = n2551 ^ n1452 ^ 1'b0 ;
  assign n28207 = n27537 & n28206 ;
  assign n28208 = ~n3746 & n8132 ;
  assign n28209 = n9241 | n28208 ;
  assign n28210 = n28209 ^ n7395 ^ 1'b0 ;
  assign n28211 = ( n2240 & ~n26652 ) | ( n2240 & n28210 ) | ( ~n26652 & n28210 ) ;
  assign n28212 = ( n10573 & ~n17129 ) | ( n10573 & n28211 ) | ( ~n17129 & n28211 ) ;
  assign n28213 = n3810 | n19440 ;
  assign n28214 = n27151 | n28213 ;
  assign n28215 = n28214 ^ n5368 ^ n4182 ;
  assign n28216 = ~n326 & n14506 ;
  assign n28217 = ~n2236 & n28216 ;
  assign n28218 = n28217 ^ n4583 ^ 1'b0 ;
  assign n28219 = n28218 ^ n22701 ^ n19269 ;
  assign n28220 = n27542 ^ n12577 ^ 1'b0 ;
  assign n28221 = ~n28219 & n28220 ;
  assign n28222 = n1120 | n4032 ;
  assign n28223 = ( n2594 & n2693 ) | ( n2594 & n28222 ) | ( n2693 & n28222 ) ;
  assign n28224 = n16066 ^ n11311 ^ 1'b0 ;
  assign n28225 = n28224 ^ n5729 ^ n4473 ;
  assign n28226 = n28223 & n28225 ;
  assign n28227 = n19553 ^ n17843 ^ n13538 ;
  assign n28228 = n28227 ^ n8924 ^ n1534 ;
  assign n28229 = n14216 ^ n14021 ^ n3024 ;
  assign n28230 = n1150 & n28229 ;
  assign n28231 = n21994 & n28230 ;
  assign n28232 = n13460 ^ n10292 ^ 1'b0 ;
  assign n28233 = ~n5965 & n26192 ;
  assign n28234 = n28233 ^ n8393 ^ 1'b0 ;
  assign n28236 = n9866 ^ n629 ^ 1'b0 ;
  assign n28235 = n20883 ^ n5539 ^ 1'b0 ;
  assign n28237 = n28236 ^ n28235 ^ n2440 ;
  assign n28238 = n10239 | n28237 ;
  assign n28239 = n7410 & ~n10028 ;
  assign n28240 = ( n6839 & n8672 ) | ( n6839 & ~n11045 ) | ( n8672 & ~n11045 ) ;
  assign n28241 = ( n5801 & ~n9647 ) | ( n5801 & n28240 ) | ( ~n9647 & n28240 ) ;
  assign n28242 = ~n28239 & n28241 ;
  assign n28244 = n3768 & ~n4465 ;
  assign n28245 = n28244 ^ n2494 ^ 1'b0 ;
  assign n28246 = n28245 ^ n13494 ^ 1'b0 ;
  assign n28247 = n3065 & ~n28246 ;
  assign n28243 = n6051 & ~n9461 ;
  assign n28248 = n28247 ^ n28243 ^ n14659 ;
  assign n28249 = n5102 & ~n28248 ;
  assign n28250 = ~n15211 & n28249 ;
  assign n28251 = n28250 ^ n26103 ^ 1'b0 ;
  assign n28252 = n16897 ^ n16123 ^ n1517 ;
  assign n28254 = n8286 & ~n9453 ;
  assign n28255 = n28159 & n28254 ;
  assign n28253 = n12595 | n15186 ;
  assign n28256 = n28255 ^ n28253 ^ 1'b0 ;
  assign n28257 = ( n5444 & n15338 ) | ( n5444 & ~n28256 ) | ( n15338 & ~n28256 ) ;
  assign n28258 = n4227 | n8275 ;
  assign n28259 = n28258 ^ n7723 ^ 1'b0 ;
  assign n28260 = n3423 | n28259 ;
  assign n28261 = n2662 & n27932 ;
  assign n28262 = ~n11525 & n28261 ;
  assign n28263 = n10231 & ~n28262 ;
  assign n28264 = n28263 ^ n20801 ^ 1'b0 ;
  assign n28265 = ( x59 & ~n6565 ) | ( x59 & n28264 ) | ( ~n6565 & n28264 ) ;
  assign n28266 = n28265 ^ n23973 ^ n20216 ;
  assign n28267 = x82 & n1111 ;
  assign n28268 = n25170 ^ n13937 ^ 1'b0 ;
  assign n28269 = n3431 & ~n17886 ;
  assign n28270 = ( ~x6 & n12168 ) | ( ~x6 & n28269 ) | ( n12168 & n28269 ) ;
  assign n28271 = n28270 ^ n23840 ^ 1'b0 ;
  assign n28272 = n16012 ^ n15275 ^ 1'b0 ;
  assign n28274 = ( n782 & ~n4623 ) | ( n782 & n7044 ) | ( ~n4623 & n7044 ) ;
  assign n28273 = n8088 & ~n8370 ;
  assign n28275 = n28274 ^ n28273 ^ 1'b0 ;
  assign n28276 = n1558 ^ x52 ^ 1'b0 ;
  assign n28277 = n6802 | n28276 ;
  assign n28278 = n28277 ^ n11606 ^ 1'b0 ;
  assign n28279 = n656 & n1655 ;
  assign n28280 = n28279 ^ n5270 ^ 1'b0 ;
  assign n28281 = ( n1586 & n9545 ) | ( n1586 & n28280 ) | ( n9545 & n28280 ) ;
  assign n28282 = n28281 ^ n19929 ^ 1'b0 ;
  assign n28283 = n24210 & n28282 ;
  assign n28284 = ( n5535 & n28278 ) | ( n5535 & ~n28283 ) | ( n28278 & ~n28283 ) ;
  assign n28285 = n13064 | n15282 ;
  assign n28286 = ~n3211 & n6228 ;
  assign n28287 = n28286 ^ n11022 ^ 1'b0 ;
  assign n28288 = n2141 & ~n5925 ;
  assign n28289 = n28287 & n28288 ;
  assign n28290 = n12801 ^ n5502 ^ 1'b0 ;
  assign n28291 = n28290 ^ n22602 ^ n9852 ;
  assign n28292 = n18413 | n21362 ;
  assign n28293 = n5111 & ~n28292 ;
  assign n28294 = ( n7311 & ~n10839 ) | ( n7311 & n19324 ) | ( ~n10839 & n19324 ) ;
  assign n28295 = n28294 ^ n8038 ^ 1'b0 ;
  assign n28296 = n28293 | n28295 ;
  assign n28297 = n28296 ^ n17749 ^ n17452 ;
  assign n28298 = n14045 & n15130 ;
  assign n28299 = ~n13198 & n28298 ;
  assign n28300 = n5974 ^ n1910 ^ 1'b0 ;
  assign n28301 = n9416 | n28300 ;
  assign n28302 = n14253 & n21151 ;
  assign n28303 = n3217 | n4645 ;
  assign n28304 = n6240 & ~n28303 ;
  assign n28305 = n28304 ^ x108 ^ 1'b0 ;
  assign n28306 = n3219 & n28305 ;
  assign n28307 = ~n6723 & n16525 ;
  assign n28308 = ~n3687 & n10113 ;
  assign n28309 = ( n16897 & ~n28307 ) | ( n16897 & n28308 ) | ( ~n28307 & n28308 ) ;
  assign n28310 = n7973 & n28309 ;
  assign n28311 = n6870 & n8290 ;
  assign n28312 = n28311 ^ n18874 ^ 1'b0 ;
  assign n28313 = n18238 ^ n8411 ^ 1'b0 ;
  assign n28314 = x143 | n28313 ;
  assign n28315 = n23518 | n28314 ;
  assign n28316 = n12546 ^ n6005 ^ 1'b0 ;
  assign n28317 = n13967 ^ n7342 ^ n5503 ;
  assign n28318 = ( n4115 & ~n18800 ) | ( n4115 & n28317 ) | ( ~n18800 & n28317 ) ;
  assign n28319 = n25700 ^ n5520 ^ n4638 ;
  assign n28320 = n6113 | n8690 ;
  assign n28321 = n10628 | n28320 ;
  assign n28322 = n19138 ^ x57 ^ 1'b0 ;
  assign n28323 = ( n15206 & ~n28321 ) | ( n15206 & n28322 ) | ( ~n28321 & n28322 ) ;
  assign n28324 = n11963 ^ n9515 ^ 1'b0 ;
  assign n28325 = n13905 | n28324 ;
  assign n28326 = n28325 ^ n12314 ^ 1'b0 ;
  assign n28327 = n7810 & ~n10535 ;
  assign n28328 = n14113 ^ n11627 ^ 1'b0 ;
  assign n28329 = ( n2489 & ~n26208 ) | ( n2489 & n28328 ) | ( ~n26208 & n28328 ) ;
  assign n28330 = n24949 ^ n4173 ^ 1'b0 ;
  assign n28331 = n8945 | n28330 ;
  assign n28332 = n28331 ^ n14415 ^ 1'b0 ;
  assign n28333 = ~n6477 & n28332 ;
  assign n28334 = n17223 & n28333 ;
  assign n28335 = n5588 ^ n1120 ^ 1'b0 ;
  assign n28336 = n2174 & n5344 ;
  assign n28337 = n10140 & n13762 ;
  assign n28338 = n21784 & n28337 ;
  assign n28339 = n22467 ^ n14848 ^ 1'b0 ;
  assign n28340 = n19182 ^ n14093 ^ 1'b0 ;
  assign n28341 = n5620 & n27615 ;
  assign n28342 = n14969 ^ n769 ^ 1'b0 ;
  assign n28343 = n9235 | n28342 ;
  assign n28344 = n512 & n28343 ;
  assign n28345 = n18772 & n28344 ;
  assign n28346 = n28345 ^ n18456 ^ 1'b0 ;
  assign n28347 = ~n4852 & n10498 ;
  assign n28348 = n19157 & n26901 ;
  assign n28349 = n26641 & n28348 ;
  assign n28350 = ( n14116 & ~n25228 ) | ( n14116 & n28339 ) | ( ~n25228 & n28339 ) ;
  assign n28351 = ~n654 & n3662 ;
  assign n28352 = n24559 ^ n15087 ^ 1'b0 ;
  assign n28353 = n28352 ^ n13144 ^ 1'b0 ;
  assign n28354 = ~n28351 & n28353 ;
  assign n28355 = ~n13548 & n18342 ;
  assign n28356 = n28355 ^ n13968 ^ 1'b0 ;
  assign n28357 = ( x159 & n2185 ) | ( x159 & n28356 ) | ( n2185 & n28356 ) ;
  assign n28358 = n3421 ^ n1091 ^ 1'b0 ;
  assign n28359 = n28357 & n28358 ;
  assign n28360 = ( n1397 & n6488 ) | ( n1397 & n28359 ) | ( n6488 & n28359 ) ;
  assign n28361 = n5789 | n22183 ;
  assign n28362 = n28361 ^ n16886 ^ 1'b0 ;
  assign n28363 = n28362 ^ n16390 ^ 1'b0 ;
  assign n28364 = n5903 & n7812 ;
  assign n28365 = n17045 & n28364 ;
  assign n28366 = n28363 & n28365 ;
  assign n28367 = n1336 ^ x254 ^ 1'b0 ;
  assign n28368 = n10304 & n17275 ;
  assign n28369 = ~n28367 & n28368 ;
  assign n28370 = n27551 ^ n7573 ^ 1'b0 ;
  assign n28371 = n14791 ^ n10928 ^ 1'b0 ;
  assign n28372 = ~n6266 & n28371 ;
  assign n28373 = n28370 & n28372 ;
  assign n28374 = n12899 ^ n9795 ^ n747 ;
  assign n28375 = n28374 ^ n8415 ^ 1'b0 ;
  assign n28376 = n10697 | n28375 ;
  assign n28377 = ~n14173 & n23437 ;
  assign n28378 = ~n26669 & n28377 ;
  assign n28379 = n5415 & ~n6306 ;
  assign n28380 = n18934 & ~n28379 ;
  assign n28381 = ~n9067 & n18764 ;
  assign n28382 = n28381 ^ n21795 ^ 1'b0 ;
  assign n28383 = ( n679 & n3791 ) | ( n679 & ~n10378 ) | ( n3791 & ~n10378 ) ;
  assign n28384 = n28383 ^ n19674 ^ n11837 ;
  assign n28385 = n28384 ^ n27820 ^ 1'b0 ;
  assign n28386 = n18106 | n28385 ;
  assign n28387 = n28386 ^ n16758 ^ 1'b0 ;
  assign n28388 = n15590 ^ n12245 ^ n2197 ;
  assign n28389 = n11920 ^ n7182 ^ 1'b0 ;
  assign n28390 = ~n10116 & n28389 ;
  assign n28391 = n350 & ~n28390 ;
  assign n28392 = ~n16630 & n18453 ;
  assign n28394 = n14555 | n21311 ;
  assign n28395 = n28394 ^ n12249 ^ 1'b0 ;
  assign n28396 = n28395 ^ n21656 ^ n14358 ;
  assign n28393 = n19186 ^ n3572 ^ 1'b0 ;
  assign n28397 = n28396 ^ n28393 ^ 1'b0 ;
  assign n28398 = n28397 ^ n23301 ^ n20213 ;
  assign n28399 = n10744 ^ n3859 ^ 1'b0 ;
  assign n28400 = n10073 | n28399 ;
  assign n28401 = n23562 ^ n4602 ^ 1'b0 ;
  assign n28402 = n9402 & ~n28401 ;
  assign n28403 = ~n4242 & n28402 ;
  assign n28404 = n28403 ^ n22483 ^ n18187 ;
  assign n28405 = n22905 | n28404 ;
  assign n28406 = n9575 | n22135 ;
  assign n28407 = n25320 & ~n28406 ;
  assign n28408 = n19858 ^ n5669 ^ 1'b0 ;
  assign n28409 = n10621 ^ n4847 ^ 1'b0 ;
  assign n28410 = n14130 & ~n28409 ;
  assign n28411 = n4294 & n14051 ;
  assign n28412 = n11054 & ~n14091 ;
  assign n28413 = ~n9472 & n28412 ;
  assign n28414 = ~n27618 & n28413 ;
  assign n28415 = ( n20789 & n22608 ) | ( n20789 & n27247 ) | ( n22608 & n27247 ) ;
  assign n28416 = x63 & ~n20180 ;
  assign n28417 = ( n10331 & n19104 ) | ( n10331 & ~n28416 ) | ( n19104 & ~n28416 ) ;
  assign n28418 = n1217 & n2709 ;
  assign n28419 = n2441 & ~n25458 ;
  assign n28420 = n5424 ^ n2994 ^ n1816 ;
  assign n28421 = ( ~n13589 & n19068 ) | ( ~n13589 & n28420 ) | ( n19068 & n28420 ) ;
  assign n28422 = n1909 & n1962 ;
  assign n28423 = n28422 ^ n567 ^ 1'b0 ;
  assign n28424 = n28423 ^ n22606 ^ 1'b0 ;
  assign n28425 = n16723 | n28424 ;
  assign n28427 = n4921 | n10982 ;
  assign n28426 = n5443 | n15885 ;
  assign n28428 = n28427 ^ n28426 ^ 1'b0 ;
  assign n28429 = n7801 ^ n5603 ^ 1'b0 ;
  assign n28430 = ~n16927 & n28429 ;
  assign n28431 = n27127 ^ n17865 ^ n15290 ;
  assign n28432 = n1061 & ~n22004 ;
  assign n28433 = n25332 & ~n28432 ;
  assign n28434 = n12649 & n28433 ;
  assign n28435 = n1998 & n25987 ;
  assign n28436 = n7794 | n13099 ;
  assign n28437 = n5878 & ~n28436 ;
  assign n28438 = ( n8862 & n16858 ) | ( n8862 & n28437 ) | ( n16858 & n28437 ) ;
  assign n28439 = n28438 ^ n3142 ^ 1'b0 ;
  assign n28440 = n3042 & ~n10405 ;
  assign n28441 = n13905 & n28440 ;
  assign n28442 = n292 & n7758 ;
  assign n28443 = n11232 & n26995 ;
  assign n28444 = ~n2871 & n28443 ;
  assign n28445 = ( n17896 & ~n19876 ) | ( n17896 & n27313 ) | ( ~n19876 & n27313 ) ;
  assign n28446 = n1271 & n27899 ;
  assign n28447 = n28446 ^ n22481 ^ 1'b0 ;
  assign n28448 = n1102 & n5424 ;
  assign n28449 = ~n13659 & n28448 ;
  assign n28450 = n14510 | n16238 ;
  assign n28451 = n28450 ^ n15414 ^ 1'b0 ;
  assign n28453 = n17607 ^ n4876 ^ 1'b0 ;
  assign n28452 = n16128 | n21622 ;
  assign n28454 = n28453 ^ n28452 ^ 1'b0 ;
  assign n28455 = n6345 ^ n6186 ^ 1'b0 ;
  assign n28458 = n3965 & ~n4979 ;
  assign n28459 = n2722 & n28458 ;
  assign n28456 = ~n9494 & n11873 ;
  assign n28457 = ~n14316 & n28456 ;
  assign n28460 = n28459 ^ n28457 ^ 1'b0 ;
  assign n28461 = n13822 | n14762 ;
  assign n28462 = n28461 ^ n14297 ^ 1'b0 ;
  assign n28463 = n28462 ^ n12321 ^ 1'b0 ;
  assign n28464 = x122 & ~n9783 ;
  assign n28465 = n4237 & n28464 ;
  assign n28466 = n6062 | n8973 ;
  assign n28467 = n12416 ^ n6408 ^ n5950 ;
  assign n28468 = ~n20721 & n21277 ;
  assign n28469 = n21782 ^ n11723 ^ 1'b0 ;
  assign n28470 = ~n6980 & n28469 ;
  assign n28471 = n18181 ^ n15539 ^ n14621 ;
  assign n28472 = n28470 & n28471 ;
  assign n28473 = n1269 & ~n18109 ;
  assign n28474 = n28473 ^ n4202 ^ 1'b0 ;
  assign n28475 = ( n5810 & n7708 ) | ( n5810 & ~n24067 ) | ( n7708 & ~n24067 ) ;
  assign n28476 = n4987 & n7223 ;
  assign n28477 = n28476 ^ n18752 ^ 1'b0 ;
  assign n28478 = n28477 ^ n18011 ^ 1'b0 ;
  assign n28479 = n9492 ^ n3502 ^ 1'b0 ;
  assign n28480 = n9063 & n25258 ;
  assign n28481 = n15665 & n20262 ;
  assign n28482 = n28481 ^ n18106 ^ n15001 ;
  assign n28483 = n22092 ^ n20835 ^ n18459 ;
  assign n28484 = n26567 | n28483 ;
  assign n28485 = ~n3007 & n28484 ;
  assign n28486 = ( ~x90 & n2822 ) | ( ~x90 & n6050 ) | ( n2822 & n6050 ) ;
  assign n28487 = n28486 ^ n4787 ^ n2244 ;
  assign n28488 = n1848 & ~n17770 ;
  assign n28489 = n28487 & n28488 ;
  assign n28490 = n2998 ^ n2915 ^ 1'b0 ;
  assign n28491 = n19323 & ~n28490 ;
  assign n28492 = n10753 & ~n11916 ;
  assign n28493 = ~n8598 & n14714 ;
  assign n28494 = n1316 & n28493 ;
  assign n28495 = n21823 & ~n28494 ;
  assign n28499 = ~n1258 & n3723 ;
  assign n28500 = n28499 ^ n22050 ^ 1'b0 ;
  assign n28501 = n13503 ^ n2105 ^ 1'b0 ;
  assign n28502 = n28500 | n28501 ;
  assign n28498 = n11682 | n17825 ;
  assign n28496 = n12098 & n12962 ;
  assign n28497 = ~n8036 & n28496 ;
  assign n28503 = n28502 ^ n28498 ^ n28497 ;
  assign n28504 = n15423 | n20735 ;
  assign n28505 = n5434 | n9468 ;
  assign n28506 = n28504 & ~n28505 ;
  assign n28508 = n27221 ^ n18350 ^ n1701 ;
  assign n28507 = x144 | n1269 ;
  assign n28509 = n28508 ^ n28507 ^ n26833 ;
  assign n28510 = n15536 ^ n3146 ^ 1'b0 ;
  assign n28511 = n8641 & ~n28510 ;
  assign n28512 = n6232 & n13500 ;
  assign n28513 = ~n28511 & n28512 ;
  assign n28514 = n10583 & ~n15615 ;
  assign n28515 = x137 & n13168 ;
  assign n28516 = ~n28514 & n28515 ;
  assign n28520 = n5408 | n6065 ;
  assign n28521 = n28520 ^ n10577 ^ 1'b0 ;
  assign n28517 = n864 | n9840 ;
  assign n28518 = n28517 ^ n25597 ^ 1'b0 ;
  assign n28519 = n4471 | n28518 ;
  assign n28522 = n28521 ^ n28519 ^ n10364 ;
  assign n28523 = n28522 ^ n22030 ^ 1'b0 ;
  assign n28524 = ( n15831 & n23437 ) | ( n15831 & n26585 ) | ( n23437 & n26585 ) ;
  assign n28526 = n9890 | n12826 ;
  assign n28527 = n28526 ^ n2680 ^ 1'b0 ;
  assign n28525 = n7740 & ~n18007 ;
  assign n28528 = n28527 ^ n28525 ^ 1'b0 ;
  assign n28529 = ~n26210 & n28528 ;
  assign n28530 = ~n2772 & n9156 ;
  assign n28531 = ~n5934 & n28530 ;
  assign n28532 = n8318 & ~n28531 ;
  assign n28533 = n28532 ^ n20549 ^ 1'b0 ;
  assign n28534 = n10372 & n28533 ;
  assign n28535 = ( n13046 & n13685 ) | ( n13046 & n14553 ) | ( n13685 & n14553 ) ;
  assign n28536 = n14279 ^ n6417 ^ 1'b0 ;
  assign n28537 = n28535 | n28536 ;
  assign n28538 = n10334 ^ n5098 ^ 1'b0 ;
  assign n28539 = n12072 & n28538 ;
  assign n28540 = n28539 ^ n13064 ^ 1'b0 ;
  assign n28541 = n12784 ^ n10921 ^ 1'b0 ;
  assign n28542 = ~n4398 & n28541 ;
  assign n28543 = n28542 ^ n8773 ^ 1'b0 ;
  assign n28544 = x106 & n28543 ;
  assign n28545 = n15343 | n28544 ;
  assign n28546 = n16508 ^ n3257 ^ 1'b0 ;
  assign n28547 = n441 | n28546 ;
  assign n28548 = n11010 | n26345 ;
  assign n28549 = n5622 & ~n5766 ;
  assign n28550 = n28549 ^ n11455 ^ 1'b0 ;
  assign n28551 = n19394 ^ n7856 ^ 1'b0 ;
  assign n28552 = n28551 ^ n5662 ^ 1'b0 ;
  assign n28553 = n28550 & ~n28552 ;
  assign n28554 = ( n2964 & n5119 ) | ( n2964 & n7517 ) | ( n5119 & n7517 ) ;
  assign n28555 = ~n379 & n17987 ;
  assign n28556 = n28555 ^ n5934 ^ 1'b0 ;
  assign n28557 = n9385 | n28556 ;
  assign n28558 = n15347 | n28557 ;
  assign n28559 = n28558 ^ n5485 ^ 1'b0 ;
  assign n28560 = ( n7568 & n13246 ) | ( n7568 & ~n28559 ) | ( n13246 & ~n28559 ) ;
  assign n28565 = ~n9453 & n13006 ;
  assign n28563 = n764 & ~n18061 ;
  assign n28564 = ~n9206 & n28563 ;
  assign n28561 = n19621 | n27373 ;
  assign n28562 = n13189 | n28561 ;
  assign n28566 = n28565 ^ n28564 ^ n28562 ;
  assign n28567 = n5496 | n7016 ;
  assign n28568 = n28567 ^ n4050 ^ 1'b0 ;
  assign n28569 = n11370 ^ n2197 ^ n823 ;
  assign n28570 = n28569 ^ n4203 ^ n2830 ;
  assign n28571 = n6897 ^ n577 ^ 1'b0 ;
  assign n28572 = n28570 & n28571 ;
  assign n28573 = n825 | n4305 ;
  assign n28574 = n28573 ^ n2123 ^ 1'b0 ;
  assign n28576 = n16596 ^ n7729 ^ 1'b0 ;
  assign n28575 = ( n8175 & ~n10333 ) | ( n8175 & n10419 ) | ( ~n10333 & n10419 ) ;
  assign n28577 = n28576 ^ n28575 ^ 1'b0 ;
  assign n28578 = n28574 & ~n28577 ;
  assign n28579 = n24867 ^ n10237 ^ 1'b0 ;
  assign n28580 = ( n1750 & n4948 ) | ( n1750 & ~n23798 ) | ( n4948 & ~n23798 ) ;
  assign n28581 = ~n16140 & n22361 ;
  assign n28582 = ~n28580 & n28581 ;
  assign n28583 = ~n6043 & n25484 ;
  assign n28584 = ( n28256 & ~n28582 ) | ( n28256 & n28583 ) | ( ~n28582 & n28583 ) ;
  assign n28585 = n28584 ^ n5768 ^ n3749 ;
  assign n28586 = n9165 | n27911 ;
  assign n28587 = n28586 ^ n5307 ^ 1'b0 ;
  assign n28588 = n23439 & n28547 ;
  assign n28589 = n24345 ^ n23284 ^ 1'b0 ;
  assign n28590 = n17075 ^ n17002 ^ n5011 ;
  assign n28594 = x29 & n6634 ;
  assign n28595 = ~n3021 & n28594 ;
  assign n28591 = n6727 & ~n7833 ;
  assign n28592 = n28591 ^ n5682 ^ 1'b0 ;
  assign n28593 = n434 & ~n28592 ;
  assign n28596 = n28595 ^ n28593 ^ n10680 ;
  assign n28597 = n28596 ^ n27313 ^ 1'b0 ;
  assign n28598 = n26485 ^ n13437 ^ n7629 ;
  assign n28599 = n14336 & n18250 ;
  assign n28600 = ~n11441 & n28599 ;
  assign n28601 = n28600 ^ n6170 ^ 1'b0 ;
  assign n28602 = n14186 ^ n3877 ^ 1'b0 ;
  assign n28603 = n1791 & ~n28602 ;
  assign n28604 = n24454 & ~n28603 ;
  assign n28605 = ~n13214 & n28604 ;
  assign n28610 = ~n5090 & n5488 ;
  assign n28611 = n28610 ^ n1709 ^ 1'b0 ;
  assign n28612 = n1394 & ~n4612 ;
  assign n28613 = ~n7620 & n28612 ;
  assign n28614 = ( n25911 & n28611 ) | ( n25911 & n28613 ) | ( n28611 & n28613 ) ;
  assign n28606 = n15839 ^ n8073 ^ 1'b0 ;
  assign n28607 = n12291 & ~n28606 ;
  assign n28608 = n28607 ^ n3069 ^ 1'b0 ;
  assign n28609 = n17452 & n28608 ;
  assign n28615 = n28614 ^ n28609 ^ 1'b0 ;
  assign n28616 = n12010 & ~n18865 ;
  assign n28617 = n28616 ^ x24 ^ 1'b0 ;
  assign n28618 = n15430 & ~n28617 ;
  assign n28619 = ( ~n1010 & n9921 ) | ( ~n1010 & n11576 ) | ( n9921 & n11576 ) ;
  assign n28620 = n28619 ^ n10705 ^ n5931 ;
  assign n28621 = n23200 ^ n20135 ^ n5257 ;
  assign n28622 = n944 | n8961 ;
  assign n28623 = n8851 & ~n28622 ;
  assign n28624 = ~n21715 & n28623 ;
  assign n28625 = ( n290 & n7199 ) | ( n290 & ~n16547 ) | ( n7199 & ~n16547 ) ;
  assign n28626 = n28625 ^ n21637 ^ n16550 ;
  assign n28628 = n9188 & ~n11332 ;
  assign n28629 = n28628 ^ n6065 ^ 1'b0 ;
  assign n28627 = n16707 ^ n8947 ^ n4845 ;
  assign n28630 = n28629 ^ n28627 ^ n18509 ;
  assign n28631 = n684 | n14300 ;
  assign n28632 = n1176 & ~n28631 ;
  assign n28633 = n28632 ^ n7192 ^ n4520 ;
  assign n28634 = n16633 | n28633 ;
  assign n28635 = n28481 ^ n9398 ^ 1'b0 ;
  assign n28636 = ( ~n7754 & n21750 ) | ( ~n7754 & n28635 ) | ( n21750 & n28635 ) ;
  assign n28639 = ( x72 & n2319 ) | ( x72 & n8130 ) | ( n2319 & n8130 ) ;
  assign n28637 = n10959 ^ n4454 ^ 1'b0 ;
  assign n28638 = n2945 & n28637 ;
  assign n28640 = n28639 ^ n28638 ^ 1'b0 ;
  assign n28641 = n4498 & n26407 ;
  assign n28642 = ~n3938 & n23900 ;
  assign n28643 = n28642 ^ n5133 ^ 1'b0 ;
  assign n28644 = n22216 | n28643 ;
  assign n28645 = n27538 | n28644 ;
  assign n28647 = ( n6050 & n23312 ) | ( n6050 & n24500 ) | ( n23312 & n24500 ) ;
  assign n28646 = n17346 & ~n17810 ;
  assign n28648 = n28647 ^ n28646 ^ n20378 ;
  assign n28651 = n12438 ^ n647 ^ 1'b0 ;
  assign n28650 = ~n6927 & n8257 ;
  assign n28649 = n4041 | n9507 ;
  assign n28652 = n28651 ^ n28650 ^ n28649 ;
  assign n28653 = ~n19630 & n25646 ;
  assign n28654 = n28653 ^ n4824 ^ 1'b0 ;
  assign n28655 = n18982 ^ n18871 ^ 1'b0 ;
  assign n28656 = ( n4041 & n18029 ) | ( n4041 & n28655 ) | ( n18029 & n28655 ) ;
  assign n28657 = n4528 | n10072 ;
  assign n28658 = n21084 | n28657 ;
  assign n28659 = n28658 ^ n4940 ^ 1'b0 ;
  assign n28660 = n26936 | n28659 ;
  assign n28661 = n22701 & ~n28660 ;
  assign n28662 = ( n14946 & ~n26551 ) | ( n14946 & n28661 ) | ( ~n26551 & n28661 ) ;
  assign n28663 = n9690 ^ n3479 ^ 1'b0 ;
  assign n28664 = ~n19294 & n28663 ;
  assign n28665 = n3998 & n28664 ;
  assign n28666 = n2399 & n28665 ;
  assign n28667 = ( n780 & n6846 ) | ( n780 & ~n14863 ) | ( n6846 & ~n14863 ) ;
  assign n28668 = n8440 | n28667 ;
  assign n28669 = n28668 ^ n9459 ^ 1'b0 ;
  assign n28670 = ( n4553 & n23926 ) | ( n4553 & n24494 ) | ( n23926 & n24494 ) ;
  assign n28671 = n25175 ^ n2423 ^ 1'b0 ;
  assign n28672 = ~n2051 & n28671 ;
  assign n28676 = n2227 | n19371 ;
  assign n28677 = ~n7973 & n28676 ;
  assign n28673 = ~n944 & n3216 ;
  assign n28674 = n28673 ^ n4789 ^ 1'b0 ;
  assign n28675 = n4614 & ~n28674 ;
  assign n28678 = n28677 ^ n28675 ^ n1534 ;
  assign n28679 = n27902 | n28678 ;
  assign n28680 = n8539 ^ n4940 ^ 1'b0 ;
  assign n28681 = ~n12066 & n28680 ;
  assign n28682 = n4209 ^ n3010 ^ n2645 ;
  assign n28683 = n28681 & n28682 ;
  assign n28684 = n14744 & n28683 ;
  assign n28692 = n4756 & n24314 ;
  assign n28686 = n13359 ^ n13308 ^ 1'b0 ;
  assign n28687 = n20603 & ~n28686 ;
  assign n28685 = n13916 & ~n24915 ;
  assign n28688 = n28687 ^ n28685 ^ 1'b0 ;
  assign n28689 = ~n9422 & n28688 ;
  assign n28690 = n28689 ^ n3985 ^ 1'b0 ;
  assign n28691 = ~n22434 & n28690 ;
  assign n28693 = n28692 ^ n28691 ^ 1'b0 ;
  assign n28694 = ~n27030 & n28693 ;
  assign n28701 = n4048 & ~n10375 ;
  assign n28702 = n28701 ^ n16663 ^ 1'b0 ;
  assign n28699 = n13607 | n18224 ;
  assign n28698 = ~n6118 & n13147 ;
  assign n28700 = n28699 ^ n28698 ^ 1'b0 ;
  assign n28695 = n14217 ^ n3675 ^ 1'b0 ;
  assign n28696 = n12087 | n28695 ;
  assign n28697 = n18186 & ~n28696 ;
  assign n28703 = n28702 ^ n28700 ^ n28697 ;
  assign n28704 = n12709 ^ n2278 ^ 1'b0 ;
  assign n28705 = ~n11256 & n16682 ;
  assign n28706 = n28704 & n28705 ;
  assign n28707 = n23142 ^ n263 ^ 1'b0 ;
  assign n28708 = n22114 ^ n2238 ^ 1'b0 ;
  assign n28709 = n9511 & ~n28708 ;
  assign n28710 = n271 & n2656 ;
  assign n28711 = ~n2885 & n28710 ;
  assign n28712 = n14887 ^ n1266 ^ 1'b0 ;
  assign n28713 = ~n28711 & n28712 ;
  assign n28714 = ~n1684 & n28713 ;
  assign n28715 = ~n28709 & n28714 ;
  assign n28716 = n7961 & n12483 ;
  assign n28720 = n11905 ^ n4592 ^ x240 ;
  assign n28717 = n10067 ^ n6978 ^ 1'b0 ;
  assign n28718 = n28717 ^ n13954 ^ 1'b0 ;
  assign n28719 = n3810 & n28718 ;
  assign n28721 = n28720 ^ n28719 ^ n16812 ;
  assign n28722 = n12874 & ~n15237 ;
  assign n28723 = n821 & ~n28722 ;
  assign n28724 = n13448 ^ n4717 ^ 1'b0 ;
  assign n28725 = ~n19907 & n28724 ;
  assign n28726 = n4374 | n4817 ;
  assign n28727 = n2178 | n28726 ;
  assign n28728 = n10005 ^ n2334 ^ 1'b0 ;
  assign n28729 = n28728 ^ n14846 ^ 1'b0 ;
  assign n28730 = n28727 & n28729 ;
  assign n28731 = n17116 ^ n16181 ^ 1'b0 ;
  assign n28732 = x252 & n28731 ;
  assign n28733 = n22430 ^ n16739 ^ n14029 ;
  assign n28734 = n28733 ^ n3023 ^ 1'b0 ;
  assign n28735 = ~n7385 & n28734 ;
  assign n28736 = n2962 & ~n4752 ;
  assign n28737 = ~n4714 & n28736 ;
  assign n28738 = n28737 ^ n7761 ^ 1'b0 ;
  assign n28739 = n28735 & n28738 ;
  assign n28740 = n10322 ^ n8056 ^ 1'b0 ;
  assign n28741 = n28740 ^ n27338 ^ 1'b0 ;
  assign n28742 = n27131 ^ n25931 ^ n4989 ;
  assign n28743 = ( n5203 & ~n11972 ) | ( n5203 & n18781 ) | ( ~n11972 & n18781 ) ;
  assign n28744 = n1818 & n18666 ;
  assign n28745 = n28744 ^ n25313 ^ 1'b0 ;
  assign n28746 = n1789 & ~n17727 ;
  assign n28747 = n14185 | n28746 ;
  assign n28748 = n3693 | n28747 ;
  assign n28749 = n18846 ^ n15108 ^ 1'b0 ;
  assign n28750 = n3749 ^ n2774 ^ 1'b0 ;
  assign n28751 = n22687 & n28750 ;
  assign n28752 = n3235 ^ n1424 ^ 1'b0 ;
  assign n28753 = n4145 & n28752 ;
  assign n28754 = n28753 ^ n18703 ^ 1'b0 ;
  assign n28755 = ( n1629 & n3239 ) | ( n1629 & n28754 ) | ( n3239 & n28754 ) ;
  assign n28756 = ~x226 & n14774 ;
  assign n28757 = n28756 ^ n9852 ^ 1'b0 ;
  assign n28758 = ( n22557 & n24824 ) | ( n22557 & n26780 ) | ( n24824 & n26780 ) ;
  assign n28759 = n20446 & ~n21872 ;
  assign n28760 = n2562 & n20357 ;
  assign n28761 = n11495 | n24166 ;
  assign n28762 = n6053 | n28761 ;
  assign n28763 = n264 | n7394 ;
  assign n28764 = n28763 ^ n1919 ^ 1'b0 ;
  assign n28765 = n1688 & ~n28764 ;
  assign n28766 = n28765 ^ n6479 ^ 1'b0 ;
  assign n28767 = n28766 ^ n5903 ^ n1582 ;
  assign n28768 = ( n1425 & n18410 ) | ( n1425 & n28767 ) | ( n18410 & n28767 ) ;
  assign n28769 = ( n8175 & n14811 ) | ( n8175 & ~n28768 ) | ( n14811 & ~n28768 ) ;
  assign n28770 = ( n10617 & ~n28762 ) | ( n10617 & n28769 ) | ( ~n28762 & n28769 ) ;
  assign n28771 = n14593 & n19557 ;
  assign n28772 = n9096 & n11163 ;
  assign n28773 = ~n17631 & n28772 ;
  assign n28774 = n9052 & ~n20706 ;
  assign n28775 = n20591 ^ n4547 ^ n3434 ;
  assign n28776 = n4311 | n23798 ;
  assign n28777 = ~n410 & n28776 ;
  assign n28778 = n28777 ^ n9383 ^ 1'b0 ;
  assign n28779 = ( n1617 & n3379 ) | ( n1617 & ~n12906 ) | ( n3379 & ~n12906 ) ;
  assign n28780 = ( ~n4314 & n22783 ) | ( ~n4314 & n28779 ) | ( n22783 & n28779 ) ;
  assign n28781 = n20649 & n25360 ;
  assign n28782 = n28780 & n28781 ;
  assign n28783 = n7647 & n17880 ;
  assign n28784 = n2506 & ~n28351 ;
  assign n28785 = n28784 ^ n21270 ^ 1'b0 ;
  assign n28786 = ~n745 & n10287 ;
  assign n28787 = ( n9378 & ~n10264 ) | ( n9378 & n28786 ) | ( ~n10264 & n28786 ) ;
  assign n28788 = n7189 & ~n18476 ;
  assign n28789 = ( n10416 & n24762 ) | ( n10416 & n28788 ) | ( n24762 & n28788 ) ;
  assign n28790 = n7416 & ~n28789 ;
  assign n28795 = n16852 ^ n11357 ^ n1776 ;
  assign n28791 = n10711 ^ n4007 ^ 1'b0 ;
  assign n28792 = n15475 ^ n13267 ^ 1'b0 ;
  assign n28793 = ~n27951 & n28792 ;
  assign n28794 = n28791 & n28793 ;
  assign n28796 = n28795 ^ n28794 ^ 1'b0 ;
  assign n28797 = n6308 & n17690 ;
  assign n28798 = n28797 ^ n9542 ^ 1'b0 ;
  assign n28799 = n8375 ^ n4285 ^ n2867 ;
  assign n28800 = n4498 ^ n1727 ^ 1'b0 ;
  assign n28801 = ( n1035 & n10801 ) | ( n1035 & n13979 ) | ( n10801 & n13979 ) ;
  assign n28802 = n28801 ^ n13591 ^ 1'b0 ;
  assign n28803 = n18222 & ~n28802 ;
  assign n28804 = n28800 & n28803 ;
  assign n28805 = n2630 | n28804 ;
  assign n28806 = n12970 ^ n11937 ^ n11874 ;
  assign n28807 = n9234 & n28806 ;
  assign n28808 = ( n5914 & n7379 ) | ( n5914 & n23082 ) | ( n7379 & n23082 ) ;
  assign n28809 = n8553 & n19077 ;
  assign n28810 = n7425 & n28809 ;
  assign n28811 = x100 & ~n28810 ;
  assign n28812 = n28811 ^ n21886 ^ 1'b0 ;
  assign n28813 = n28812 ^ n19762 ^ 1'b0 ;
  assign n28814 = n20043 & n28813 ;
  assign n28815 = n28814 ^ n14709 ^ 1'b0 ;
  assign n28816 = ( n12114 & n14760 ) | ( n12114 & n28167 ) | ( n14760 & n28167 ) ;
  assign n28817 = n28816 ^ n25128 ^ n5622 ;
  assign n28818 = n10212 & n14201 ;
  assign n28819 = n3433 ^ n1337 ^ 1'b0 ;
  assign n28820 = n21557 & ~n28819 ;
  assign n28821 = n4112 & n28820 ;
  assign n28822 = ~n8762 & n28821 ;
  assign n28823 = ~n4226 & n16640 ;
  assign n28824 = n22715 | n28823 ;
  assign n28825 = n28824 ^ n13316 ^ 1'b0 ;
  assign n28826 = ~n28504 & n28825 ;
  assign n28827 = n7148 ^ n4347 ^ 1'b0 ;
  assign n28828 = n4740 & n28827 ;
  assign n28829 = ( n7617 & n14314 ) | ( n7617 & ~n28828 ) | ( n14314 & ~n28828 ) ;
  assign n28830 = ~n3019 & n23904 ;
  assign n28831 = n21373 | n26954 ;
  assign n28832 = n27723 & ~n28831 ;
  assign n28833 = ~n8088 & n18123 ;
  assign n28834 = n15081 & n24033 ;
  assign n28835 = n28834 ^ n20544 ^ 1'b0 ;
  assign n28836 = n18121 ^ n10405 ^ n7702 ;
  assign n28837 = n2976 & ~n28836 ;
  assign n28838 = ~n24160 & n28837 ;
  assign n28839 = ( n1213 & n13189 ) | ( n1213 & ~n15054 ) | ( n13189 & ~n15054 ) ;
  assign n28840 = n22236 ^ n19408 ^ 1'b0 ;
  assign n28841 = n27935 ^ n22816 ^ n14317 ;
  assign n28842 = n28840 | n28841 ;
  assign n28843 = n7273 & ~n27202 ;
  assign n28844 = n28843 ^ n18270 ^ 1'b0 ;
  assign n28845 = n9583 | n12721 ;
  assign n28846 = n12010 | n28845 ;
  assign n28847 = n25605 ^ n23290 ^ 1'b0 ;
  assign n28848 = n28846 | n28847 ;
  assign n28849 = n23586 ^ n11365 ^ n7561 ;
  assign n28850 = n22443 ^ n9770 ^ n7473 ;
  assign n28851 = ( ~n4952 & n5158 ) | ( ~n4952 & n22653 ) | ( n5158 & n22653 ) ;
  assign n28852 = ( n4273 & n16328 ) | ( n4273 & ~n28851 ) | ( n16328 & ~n28851 ) ;
  assign n28853 = n14321 ^ n8335 ^ n3825 ;
  assign n28854 = ( ~n19268 & n26472 ) | ( ~n19268 & n28853 ) | ( n26472 & n28853 ) ;
  assign n28855 = n3259 & ~n4973 ;
  assign n28856 = n28855 ^ n3297 ^ 1'b0 ;
  assign n28857 = n28856 ^ n19241 ^ n7801 ;
  assign n28858 = ~n26522 & n28857 ;
  assign n28859 = n17466 & n28858 ;
  assign n28860 = n26247 ^ n13835 ^ n9163 ;
  assign n28861 = n5190 & n9779 ;
  assign n28862 = n12158 ^ n2403 ^ 1'b0 ;
  assign n28863 = n28861 & n28862 ;
  assign n28864 = n21982 ^ n9932 ^ 1'b0 ;
  assign n28865 = n2036 | n28864 ;
  assign n28866 = n12978 ^ n3833 ^ 1'b0 ;
  assign n28867 = ( n27215 & n28865 ) | ( n27215 & n28866 ) | ( n28865 & n28866 ) ;
  assign n28868 = n1576 | n22736 ;
  assign n28869 = n1635 & ~n17496 ;
  assign n28870 = n9917 & ~n22258 ;
  assign n28871 = n28870 ^ n22389 ^ n21790 ;
  assign n28872 = ( n2348 & n5456 ) | ( n2348 & ~n5483 ) | ( n5456 & ~n5483 ) ;
  assign n28875 = n18884 ^ n6540 ^ n2387 ;
  assign n28873 = n10093 ^ n7029 ^ 1'b0 ;
  assign n28874 = n28873 ^ n3817 ^ 1'b0 ;
  assign n28876 = n28875 ^ n28874 ^ n10899 ;
  assign n28877 = ( n10873 & n28872 ) | ( n10873 & ~n28876 ) | ( n28872 & ~n28876 ) ;
  assign n28880 = n7902 & n9176 ;
  assign n28878 = n12110 ^ n8962 ^ n5153 ;
  assign n28879 = n26818 | n28878 ;
  assign n28881 = n28880 ^ n28879 ^ 1'b0 ;
  assign n28882 = n28881 ^ n21785 ^ 1'b0 ;
  assign n28883 = n10857 & ~n28882 ;
  assign n28884 = ~n25124 & n27443 ;
  assign n28885 = n28884 ^ n18676 ^ 1'b0 ;
  assign n28889 = n663 & ~n5848 ;
  assign n28886 = n8363 & n17206 ;
  assign n28887 = n1933 & n28886 ;
  assign n28888 = ( n10086 & n22648 ) | ( n10086 & n28887 ) | ( n22648 & n28887 ) ;
  assign n28890 = n28889 ^ n28888 ^ 1'b0 ;
  assign n28891 = ( n14688 & n23724 ) | ( n14688 & n26935 ) | ( n23724 & n26935 ) ;
  assign n28892 = n3995 & n24657 ;
  assign n28893 = n28892 ^ n14761 ^ 1'b0 ;
  assign n28894 = n14057 ^ n11366 ^ 1'b0 ;
  assign n28895 = n28551 | n28894 ;
  assign n28896 = ( n1051 & n5953 ) | ( n1051 & ~n7336 ) | ( n5953 & ~n7336 ) ;
  assign n28897 = n20559 | n28896 ;
  assign n28898 = n23811 ^ n13236 ^ 1'b0 ;
  assign n28899 = ( ~n798 & n27812 ) | ( ~n798 & n28898 ) | ( n27812 & n28898 ) ;
  assign n28900 = ( n6699 & n28897 ) | ( n6699 & ~n28899 ) | ( n28897 & ~n28899 ) ;
  assign n28908 = n24019 ^ n6965 ^ 1'b0 ;
  assign n28904 = n1736 | n14921 ;
  assign n28905 = n28904 ^ n3248 ^ 1'b0 ;
  assign n28901 = n20459 ^ n5012 ^ n3260 ;
  assign n28902 = n28901 ^ n2146 ^ 1'b0 ;
  assign n28903 = n21481 & ~n28902 ;
  assign n28906 = n28905 ^ n28903 ^ 1'b0 ;
  assign n28907 = n17338 & n28906 ;
  assign n28909 = n28908 ^ n28907 ^ 1'b0 ;
  assign n28915 = n7850 | n14805 ;
  assign n28911 = n18378 ^ n6776 ^ 1'b0 ;
  assign n28912 = ~n11210 & n28911 ;
  assign n28910 = n7089 | n9451 ;
  assign n28913 = n28912 ^ n28910 ^ 1'b0 ;
  assign n28914 = n350 & ~n28913 ;
  assign n28916 = n28915 ^ n28914 ^ 1'b0 ;
  assign n28917 = n17995 ^ x90 ^ 1'b0 ;
  assign n28918 = n7720 ^ n5969 ^ 1'b0 ;
  assign n28919 = n10628 & ~n28918 ;
  assign n28920 = ( n1067 & ~n28917 ) | ( n1067 & n28919 ) | ( ~n28917 & n28919 ) ;
  assign n28921 = n12412 & ~n19954 ;
  assign n28922 = x20 & ~n3288 ;
  assign n28923 = ~n1928 & n28922 ;
  assign n28924 = n24870 & ~n28923 ;
  assign n28925 = x148 & ~x251 ;
  assign n28926 = n12138 & ~n28925 ;
  assign n28927 = n26885 ^ n16842 ^ n7540 ;
  assign n28928 = ( n2130 & ~n8492 ) | ( n2130 & n28927 ) | ( ~n8492 & n28927 ) ;
  assign n28929 = n12234 | n28928 ;
  assign n28930 = n28929 ^ n27987 ^ 1'b0 ;
  assign n28931 = ~n13954 & n28930 ;
  assign n28932 = ~n28926 & n28931 ;
  assign n28933 = ( n6086 & n21456 ) | ( n6086 & n26995 ) | ( n21456 & n26995 ) ;
  assign n28934 = n16478 ^ n4049 ^ 1'b0 ;
  assign n28935 = ~n409 & n25320 ;
  assign n28936 = ~n27464 & n28935 ;
  assign n28937 = ( n1182 & n1321 ) | ( n1182 & ~n17921 ) | ( n1321 & ~n17921 ) ;
  assign n28938 = n28937 ^ n8066 ^ 1'b0 ;
  assign n28939 = n1884 & n4291 ;
  assign n28940 = ~n1409 & n11334 ;
  assign n28941 = n28940 ^ n11849 ^ 1'b0 ;
  assign n28942 = ~n24234 & n28941 ;
  assign n28943 = n28939 & n28942 ;
  assign n28944 = n24146 ^ n6003 ^ n3475 ;
  assign n28945 = n28944 ^ n10909 ^ 1'b0 ;
  assign n28946 = ( n6813 & ~n8012 ) | ( n6813 & n19433 ) | ( ~n8012 & n19433 ) ;
  assign n28947 = ~n2488 & n14867 ;
  assign n28948 = n28947 ^ n6157 ^ 1'b0 ;
  assign n28949 = ( n3782 & ~n9247 ) | ( n3782 & n28948 ) | ( ~n9247 & n28948 ) ;
  assign n28950 = ~n8106 & n24500 ;
  assign n28951 = n12429 ^ n8533 ^ 1'b0 ;
  assign n28952 = n3965 & n28951 ;
  assign n28953 = n13138 ^ n595 ^ 1'b0 ;
  assign n28954 = n6312 | n20424 ;
  assign n28955 = n9257 & ~n28954 ;
  assign n28956 = n28955 ^ n15051 ^ n8818 ;
  assign n28957 = ~n832 & n10253 ;
  assign n28958 = ~n28956 & n28957 ;
  assign n28959 = n5437 | n26415 ;
  assign n28960 = n28635 & ~n28959 ;
  assign n28961 = n17486 ^ n1397 ^ 1'b0 ;
  assign n28962 = n5593 | n18617 ;
  assign n28963 = ~n813 & n16038 ;
  assign n28964 = n7331 & n28963 ;
  assign n28966 = n1196 & ~n6683 ;
  assign n28967 = ~n12859 & n28966 ;
  assign n28968 = n5751 & n14158 ;
  assign n28969 = n28967 & n28968 ;
  assign n28970 = ( n18379 & n27971 ) | ( n18379 & n28969 ) | ( n27971 & n28969 ) ;
  assign n28965 = n10105 | n19584 ;
  assign n28971 = n28970 ^ n28965 ^ 1'b0 ;
  assign n28972 = x197 & n19233 ;
  assign n28973 = ~n7830 & n28972 ;
  assign n28974 = n16078 ^ n5492 ^ 1'b0 ;
  assign n28975 = n27736 | n28974 ;
  assign n28976 = ( ~n500 & n7764 ) | ( ~n500 & n26552 ) | ( n7764 & n26552 ) ;
  assign n28977 = n7512 | n14589 ;
  assign n28978 = n28977 ^ n10052 ^ 1'b0 ;
  assign n28979 = n3708 & ~n5884 ;
  assign n28980 = n5709 & n28979 ;
  assign n28981 = n22053 ^ n5863 ^ 1'b0 ;
  assign n28982 = ( n4641 & ~n4645 ) | ( n4641 & n12539 ) | ( ~n4645 & n12539 ) ;
  assign n28983 = ( n20846 & ~n25460 ) | ( n20846 & n28982 ) | ( ~n25460 & n28982 ) ;
  assign n28984 = n28983 ^ n10346 ^ 1'b0 ;
  assign n28985 = n28437 ^ n16903 ^ 1'b0 ;
  assign n28986 = ~n8321 & n28985 ;
  assign n28987 = n13120 | n22294 ;
  assign n28988 = n24173 & ~n28987 ;
  assign n28989 = ( n928 & n19041 ) | ( n928 & ~n28988 ) | ( n19041 & ~n28988 ) ;
  assign n28990 = n9709 | n28989 ;
  assign n28991 = n16060 & ~n24570 ;
  assign n28992 = ~n7148 & n28044 ;
  assign n28993 = n8658 & n18356 ;
  assign n28994 = n28993 ^ n19842 ^ 1'b0 ;
  assign n28996 = n1550 & n3158 ;
  assign n28997 = n28996 ^ n5134 ^ 1'b0 ;
  assign n28998 = n28997 ^ n2683 ^ 1'b0 ;
  assign n28999 = n12026 & n28998 ;
  assign n29000 = n1950 & n28999 ;
  assign n29001 = n29000 ^ n3786 ^ 1'b0 ;
  assign n29002 = n29001 ^ n18229 ^ n6749 ;
  assign n28995 = n10484 | n23371 ;
  assign n29003 = n29002 ^ n28995 ^ n13730 ;
  assign n29004 = n29003 ^ n17960 ^ 1'b0 ;
  assign n29005 = n9454 ^ n329 ^ 1'b0 ;
  assign n29006 = n8079 ^ n1393 ^ 1'b0 ;
  assign n29007 = n9943 | n17833 ;
  assign n29008 = ~n20980 & n29007 ;
  assign n29009 = n29008 ^ n28423 ^ n1495 ;
  assign n29010 = ( n2993 & ~n21369 ) | ( n2993 & n22737 ) | ( ~n21369 & n22737 ) ;
  assign n29011 = n27531 ^ n10341 ^ 1'b0 ;
  assign n29012 = n2243 & n29011 ;
  assign n29013 = n29012 ^ n12277 ^ 1'b0 ;
  assign n29019 = n1987 & n4975 ;
  assign n29017 = n26177 ^ n6808 ^ 1'b0 ;
  assign n29018 = n20193 & n29017 ;
  assign n29020 = n29019 ^ n29018 ^ 1'b0 ;
  assign n29014 = n16956 ^ n11277 ^ n8049 ;
  assign n29015 = n29014 ^ n19217 ^ 1'b0 ;
  assign n29016 = n18410 & ~n29015 ;
  assign n29021 = n29020 ^ n29016 ^ n4654 ;
  assign n29022 = n2836 | n13303 ;
  assign n29023 = n29022 ^ n2049 ^ 1'b0 ;
  assign n29024 = ( ~n12241 & n18624 ) | ( ~n12241 & n29023 ) | ( n18624 & n29023 ) ;
  assign n29025 = n1680 | n10473 ;
  assign n29026 = n5208 | n12232 ;
  assign n29027 = n29026 ^ n7535 ^ 1'b0 ;
  assign n29028 = ( n20412 & ~n29025 ) | ( n20412 & n29027 ) | ( ~n29025 & n29027 ) ;
  assign n29029 = n10662 ^ n861 ^ 1'b0 ;
  assign n29030 = n29029 ^ n9308 ^ 1'b0 ;
  assign n29031 = ( ~x220 & n24248 ) | ( ~x220 & n26762 ) | ( n24248 & n26762 ) ;
  assign n29032 = ( n1359 & n1890 ) | ( n1359 & n11813 ) | ( n1890 & n11813 ) ;
  assign n29034 = ( n4317 & ~n15529 ) | ( n4317 & n26811 ) | ( ~n15529 & n26811 ) ;
  assign n29033 = n337 & ~n2077 ;
  assign n29035 = n29034 ^ n29033 ^ 1'b0 ;
  assign n29037 = n8351 ^ n6468 ^ 1'b0 ;
  assign n29038 = ( ~x29 & n14779 ) | ( ~x29 & n29037 ) | ( n14779 & n29037 ) ;
  assign n29036 = ( n10919 & n21759 ) | ( n10919 & n27333 ) | ( n21759 & n27333 ) ;
  assign n29039 = n29038 ^ n29036 ^ 1'b0 ;
  assign n29040 = n9320 & ~n14696 ;
  assign n29041 = n29040 ^ n13139 ^ x229 ;
  assign n29042 = ( n12235 & n14606 ) | ( n12235 & ~n15760 ) | ( n14606 & ~n15760 ) ;
  assign n29043 = n24760 | n29042 ;
  assign n29044 = n29043 ^ n7921 ^ 1'b0 ;
  assign n29046 = n4469 & n13346 ;
  assign n29047 = n29046 ^ n1519 ^ 1'b0 ;
  assign n29045 = n5405 ^ n530 ^ 1'b0 ;
  assign n29048 = n29047 ^ n29045 ^ x196 ;
  assign n29049 = n12469 | n29048 ;
  assign n29050 = n7088 & ~n29049 ;
  assign n29051 = n17387 ^ n6555 ^ 1'b0 ;
  assign n29052 = n11627 & n29051 ;
  assign n29053 = n29052 ^ n8526 ^ n6854 ;
  assign n29054 = ( ~n13250 & n14013 ) | ( ~n13250 & n29053 ) | ( n14013 & n29053 ) ;
  assign n29056 = n19608 ^ n17129 ^ 1'b0 ;
  assign n29057 = n2885 & ~n29056 ;
  assign n29055 = n28058 ^ n12875 ^ n4280 ;
  assign n29058 = n29057 ^ n29055 ^ n27605 ;
  assign n29059 = ( n1912 & ~n7113 ) | ( n1912 & n10808 ) | ( ~n7113 & n10808 ) ;
  assign n29060 = n3410 & n29059 ;
  assign n29061 = ( ~n6670 & n19646 ) | ( ~n6670 & n29060 ) | ( n19646 & n29060 ) ;
  assign n29062 = ( n5439 & n11430 ) | ( n5439 & ~n29061 ) | ( n11430 & ~n29061 ) ;
  assign n29063 = n29062 ^ n5162 ^ 1'b0 ;
  assign n29064 = ( n2680 & n18449 ) | ( n2680 & n29063 ) | ( n18449 & n29063 ) ;
  assign n29065 = n25849 ^ n23494 ^ 1'b0 ;
  assign n29066 = ~n2766 & n29065 ;
  assign n29067 = n8683 ^ n2972 ^ 1'b0 ;
  assign n29068 = n5070 | n29067 ;
  assign n29069 = ~x70 & n1261 ;
  assign n29070 = n5302 | n17230 ;
  assign n29071 = n29070 ^ n19992 ^ 1'b0 ;
  assign n29072 = ~n29069 & n29071 ;
  assign n29073 = n29068 & n29072 ;
  assign n29074 = n27928 ^ n20470 ^ n10365 ;
  assign n29075 = n11655 | n12341 ;
  assign n29076 = n13583 ^ n1677 ^ 1'b0 ;
  assign n29077 = n19265 & n29076 ;
  assign n29078 = n20034 ^ n8052 ^ 1'b0 ;
  assign n29079 = n325 & n29078 ;
  assign n29080 = n29079 ^ n3965 ^ 1'b0 ;
  assign n29081 = n29077 & n29080 ;
  assign n29082 = n18247 ^ n7460 ^ 1'b0 ;
  assign n29083 = ~n27383 & n29082 ;
  assign n29084 = n3633 ^ n2149 ^ 1'b0 ;
  assign n29085 = n29084 ^ n23697 ^ 1'b0 ;
  assign n29086 = n13498 ^ n6468 ^ 1'b0 ;
  assign n29087 = n10709 | n14705 ;
  assign n29088 = n8769 & ~n29087 ;
  assign n29089 = n29088 ^ n24152 ^ 1'b0 ;
  assign n29090 = n29086 & ~n29089 ;
  assign n29091 = n8651 ^ n3402 ^ n2654 ;
  assign n29092 = n15557 ^ n8191 ^ 1'b0 ;
  assign n29093 = ~n21132 & n29092 ;
  assign n29094 = ( n8760 & n29091 ) | ( n8760 & n29093 ) | ( n29091 & n29093 ) ;
  assign n29095 = n12860 ^ n12051 ^ 1'b0 ;
  assign n29096 = ( n3437 & ~n27615 ) | ( n3437 & n29095 ) | ( ~n27615 & n29095 ) ;
  assign n29097 = n2227 | n5697 ;
  assign n29098 = n29097 ^ n8418 ^ 1'b0 ;
  assign n29099 = ( n13204 & n20358 ) | ( n13204 & n29098 ) | ( n20358 & n29098 ) ;
  assign n29100 = n14026 ^ n2574 ^ 1'b0 ;
  assign n29101 = n29099 | n29100 ;
  assign n29102 = n15704 | n29101 ;
  assign n29103 = n21057 | n29102 ;
  assign n29104 = ( n7637 & ~n27018 ) | ( n7637 & n29103 ) | ( ~n27018 & n29103 ) ;
  assign n29105 = ~n7394 & n7948 ;
  assign n29106 = n29105 ^ n5532 ^ 1'b0 ;
  assign n29107 = n29106 ^ n11857 ^ 1'b0 ;
  assign n29108 = n20025 ^ n14845 ^ n7218 ;
  assign n29109 = n29108 ^ n27476 ^ 1'b0 ;
  assign n29110 = n12991 & n29109 ;
  assign n29111 = n29107 & n29110 ;
  assign n29112 = n13678 & ~n29111 ;
  assign n29113 = n26516 & ~n29112 ;
  assign n29114 = n29113 ^ n25367 ^ 1'b0 ;
  assign n29115 = n8548 ^ n4965 ^ 1'b0 ;
  assign n29116 = ~n17015 & n29115 ;
  assign n29117 = ( n3941 & ~n8048 ) | ( n3941 & n24097 ) | ( ~n8048 & n24097 ) ;
  assign n29121 = n10445 & ~n21884 ;
  assign n29120 = ( x47 & x59 ) | ( x47 & ~n6446 ) | ( x59 & ~n6446 ) ;
  assign n29118 = n23418 ^ n16668 ^ n15239 ;
  assign n29119 = n18622 & ~n29118 ;
  assign n29122 = n29121 ^ n29120 ^ n29119 ;
  assign n29123 = n821 & ~n857 ;
  assign n29124 = ( n9627 & n17268 ) | ( n9627 & ~n29123 ) | ( n17268 & ~n29123 ) ;
  assign n29125 = x219 & ~n1995 ;
  assign n29126 = n29125 ^ n14261 ^ 1'b0 ;
  assign n29127 = n29126 ^ n20386 ^ 1'b0 ;
  assign n29128 = ( n11046 & ~n29124 ) | ( n11046 & n29127 ) | ( ~n29124 & n29127 ) ;
  assign n29130 = n21888 ^ n10169 ^ n9529 ;
  assign n29129 = ~n7559 & n27300 ;
  assign n29131 = n29130 ^ n29129 ^ n9898 ;
  assign n29132 = ( n4924 & n5024 ) | ( n4924 & ~n7212 ) | ( n5024 & ~n7212 ) ;
  assign n29133 = n4351 | n5926 ;
  assign n29134 = n12162 & ~n29133 ;
  assign n29135 = n3421 & ~n29134 ;
  assign n29136 = ~n9814 & n29135 ;
  assign n29137 = ~n9273 & n29136 ;
  assign n29138 = n29132 & n29137 ;
  assign n29139 = n16761 ^ n11942 ^ 1'b0 ;
  assign n29140 = n7294 | n14236 ;
  assign n29141 = n29140 ^ n8629 ^ 1'b0 ;
  assign n29142 = n4701 & n29141 ;
  assign n29143 = n29142 ^ n8128 ^ 1'b0 ;
  assign n29144 = ~n3119 & n5459 ;
  assign n29145 = n29144 ^ n3507 ^ 1'b0 ;
  assign n29146 = n16008 | n29145 ;
  assign n29147 = n26572 | n29146 ;
  assign n29148 = x131 & ~n10260 ;
  assign n29149 = n29148 ^ n26989 ^ 1'b0 ;
  assign n29150 = n7881 | n23239 ;
  assign n29151 = n28825 ^ n25738 ^ 1'b0 ;
  assign n29152 = n29150 | n29151 ;
  assign n29153 = n15449 & n16222 ;
  assign n29154 = n5837 & n29153 ;
  assign n29155 = n29154 ^ n26749 ^ 1'b0 ;
  assign n29156 = n27279 ^ n10748 ^ 1'b0 ;
  assign n29157 = n22098 | n29156 ;
  assign n29158 = ( n6904 & n29077 ) | ( n6904 & n29157 ) | ( n29077 & n29157 ) ;
  assign n29159 = ( n2094 & ~n3108 ) | ( n2094 & n3715 ) | ( ~n3108 & n3715 ) ;
  assign n29160 = n29159 ^ n28172 ^ 1'b0 ;
  assign n29161 = n3464 | n29160 ;
  assign n29162 = n29158 & ~n29161 ;
  assign n29163 = n9836 ^ n2408 ^ n1420 ;
  assign n29164 = n29163 ^ n2722 ^ n861 ;
  assign n29165 = ( ~n1377 & n10614 ) | ( ~n1377 & n11313 ) | ( n10614 & n11313 ) ;
  assign n29167 = n2621 ^ n1083 ^ 1'b0 ;
  assign n29168 = n2680 | n29167 ;
  assign n29166 = ~n7324 & n17428 ;
  assign n29169 = n29168 ^ n29166 ^ n1204 ;
  assign n29170 = ~n10199 & n29169 ;
  assign n29171 = n2141 & ~n26849 ;
  assign n29172 = n22430 ^ n10501 ^ 1'b0 ;
  assign n29173 = ~n29171 & n29172 ;
  assign n29174 = n26483 ^ n10844 ^ 1'b0 ;
  assign n29175 = n2142 & ~n29174 ;
  assign n29176 = n2321 & n10641 ;
  assign n29177 = n29175 & n29176 ;
  assign n29178 = n9261 & n29177 ;
  assign n29179 = n25302 ^ n5739 ^ 1'b0 ;
  assign n29180 = n26847 ^ n26046 ^ n3268 ;
  assign n29181 = n19068 ^ n17718 ^ 1'b0 ;
  assign n29182 = n20592 | n29181 ;
  assign n29183 = n17102 ^ n1533 ^ 1'b0 ;
  assign n29184 = n29183 ^ n5567 ^ 1'b0 ;
  assign n29185 = n5843 | n29184 ;
  assign n29186 = ~n5384 & n28189 ;
  assign n29187 = n13405 | n29186 ;
  assign n29189 = n12857 & n13184 ;
  assign n29190 = n29189 ^ n6403 ^ 1'b0 ;
  assign n29188 = n3494 | n27185 ;
  assign n29191 = n29190 ^ n29188 ^ 1'b0 ;
  assign n29192 = n11522 ^ n2344 ^ 1'b0 ;
  assign n29193 = n18614 ^ n12297 ^ 1'b0 ;
  assign n29194 = n21588 & n29193 ;
  assign n29195 = n29194 ^ n16702 ^ 1'b0 ;
  assign n29196 = n29192 & n29195 ;
  assign n29197 = n17007 & ~n29196 ;
  assign n29198 = n29197 ^ n15563 ^ 1'b0 ;
  assign n29199 = n24815 ^ n22948 ^ 1'b0 ;
  assign n29200 = n29199 ^ n430 ^ 1'b0 ;
  assign n29201 = ~n631 & n29200 ;
  assign n29202 = n19382 ^ n5347 ^ 1'b0 ;
  assign n29203 = n5628 & n15149 ;
  assign n29204 = ( n12287 & ~n22175 ) | ( n12287 & n24172 ) | ( ~n22175 & n24172 ) ;
  assign n29205 = n9600 & ~n12300 ;
  assign n29206 = n10695 & n29205 ;
  assign n29207 = n29204 & n29206 ;
  assign n29208 = n11173 ^ n10909 ^ 1'b0 ;
  assign n29209 = ~n4855 & n29208 ;
  assign n29210 = n29209 ^ n7250 ^ 1'b0 ;
  assign n29211 = ~n22583 & n29210 ;
  assign n29212 = ~n7989 & n29211 ;
  assign n29213 = n29212 ^ n5613 ^ 1'b0 ;
  assign n29214 = n29213 ^ n20031 ^ 1'b0 ;
  assign n29215 = n22190 & n26762 ;
  assign n29216 = n29215 ^ n28757 ^ n13566 ;
  assign n29217 = n1548 ^ n1082 ^ 1'b0 ;
  assign n29218 = ~n6723 & n29217 ;
  assign n29219 = n12026 & ~n15573 ;
  assign n29220 = n8850 & n29219 ;
  assign n29221 = x184 & n5358 ;
  assign n29222 = n29221 ^ n2816 ^ 1'b0 ;
  assign n29223 = n14648 ^ n2680 ^ 1'b0 ;
  assign n29224 = n4982 & ~n18598 ;
  assign n29225 = n14841 ^ n1888 ^ 1'b0 ;
  assign n29226 = n29224 | n29225 ;
  assign n29227 = n9986 ^ n7966 ^ n5021 ;
  assign n29228 = n17562 ^ x107 ^ 1'b0 ;
  assign n29229 = n21314 & ~n29228 ;
  assign n29230 = n29229 ^ n4948 ^ 1'b0 ;
  assign n29231 = ( n16040 & n29227 ) | ( n16040 & ~n29230 ) | ( n29227 & ~n29230 ) ;
  assign n29232 = ( ~n5986 & n9005 ) | ( ~n5986 & n29231 ) | ( n9005 & n29231 ) ;
  assign n29233 = n11791 & ~n15224 ;
  assign n29234 = n29233 ^ n14148 ^ 1'b0 ;
  assign n29235 = n9641 ^ n3975 ^ n3640 ;
  assign n29236 = n8966 | n19640 ;
  assign n29237 = n15240 & ~n15872 ;
  assign n29238 = ~n22163 & n29237 ;
  assign n29241 = n27217 ^ n13795 ^ 1'b0 ;
  assign n29239 = n11936 ^ n950 ^ n402 ;
  assign n29240 = n6507 & n29239 ;
  assign n29242 = n29241 ^ n29240 ^ 1'b0 ;
  assign n29243 = n10822 & n20668 ;
  assign n29244 = n23116 ^ n20968 ^ 1'b0 ;
  assign n29245 = ~n29243 & n29244 ;
  assign n29246 = ~n1361 & n23663 ;
  assign n29247 = n3487 & n29246 ;
  assign n29248 = ( n13959 & n17496 ) | ( n13959 & n29247 ) | ( n17496 & n29247 ) ;
  assign n29249 = n24476 & n29248 ;
  assign n29250 = ( n3207 & n18606 ) | ( n3207 & n25960 ) | ( n18606 & n25960 ) ;
  assign n29251 = n14069 ^ n3777 ^ 1'b0 ;
  assign n29252 = n12498 ^ n8449 ^ 1'b0 ;
  assign n29253 = n8519 & ~n9974 ;
  assign n29254 = n29253 ^ n6403 ^ 1'b0 ;
  assign n29256 = n7165 & n7649 ;
  assign n29257 = n29256 ^ n8114 ^ 1'b0 ;
  assign n29255 = n12910 ^ n4326 ^ 1'b0 ;
  assign n29258 = n29257 ^ n29255 ^ 1'b0 ;
  assign n29261 = n4592 | n13498 ;
  assign n29262 = n3640 & ~n29261 ;
  assign n29259 = n3097 | n13097 ;
  assign n29260 = n1816 & ~n29259 ;
  assign n29263 = n29262 ^ n29260 ^ n27757 ;
  assign n29275 = n2012 | n19076 ;
  assign n29269 = n3564 & ~n8823 ;
  assign n29270 = n29269 ^ n1337 ^ 1'b0 ;
  assign n29271 = ( ~n7243 & n12126 ) | ( ~n7243 & n29270 ) | ( n12126 & n29270 ) ;
  assign n29272 = n8855 & ~n29271 ;
  assign n29273 = n29272 ^ n23116 ^ 1'b0 ;
  assign n29274 = n29273 ^ n28820 ^ 1'b0 ;
  assign n29264 = n2897 | n20104 ;
  assign n29265 = ~n9948 & n29264 ;
  assign n29266 = ~n26021 & n29265 ;
  assign n29267 = n11804 & ~n29266 ;
  assign n29268 = n29267 ^ n23358 ^ 1'b0 ;
  assign n29276 = n29275 ^ n29274 ^ n29268 ;
  assign n29277 = n13452 ^ n11232 ^ n7242 ;
  assign n29278 = n29277 ^ n23967 ^ n16487 ;
  assign n29279 = n12059 & ~n29278 ;
  assign n29280 = n29279 ^ n10367 ^ 1'b0 ;
  assign n29281 = n22771 | n29280 ;
  assign n29282 = x160 & n20313 ;
  assign n29283 = n27466 ^ n25083 ^ n14618 ;
  assign n29284 = ~n15379 & n20233 ;
  assign n29285 = n5433 ^ n3439 ^ 1'b0 ;
  assign n29286 = n10360 ^ n10230 ^ 1'b0 ;
  assign n29287 = n14366 | n29286 ;
  assign n29288 = n659 & n26868 ;
  assign n29289 = ~n25707 & n29288 ;
  assign n29290 = n3347 | n23897 ;
  assign n29291 = n13642 | n26233 ;
  assign n29292 = n18818 | n29291 ;
  assign n29293 = n10555 & n29292 ;
  assign n29294 = n14658 ^ n729 ^ 1'b0 ;
  assign n29295 = n19673 & n29294 ;
  assign n29296 = n29293 & n29295 ;
  assign n29297 = n18934 ^ n12627 ^ 1'b0 ;
  assign n29301 = n7218 & ~n8217 ;
  assign n29302 = n2112 & n29301 ;
  assign n29303 = n29302 ^ n9929 ^ 1'b0 ;
  assign n29300 = n2644 & n11211 ;
  assign n29298 = n9226 | n14597 ;
  assign n29299 = ( ~n18518 & n28828 ) | ( ~n18518 & n29298 ) | ( n28828 & n29298 ) ;
  assign n29304 = n29303 ^ n29300 ^ n29299 ;
  assign n29305 = n10483 & n15294 ;
  assign n29306 = ( n798 & n10361 ) | ( n798 & ~n11880 ) | ( n10361 & ~n11880 ) ;
  assign n29307 = x159 & n5628 ;
  assign n29308 = ~n27119 & n29307 ;
  assign n29309 = n29308 ^ n11765 ^ 1'b0 ;
  assign n29310 = n11285 & n12296 ;
  assign n29311 = n9300 & n29310 ;
  assign n29313 = n9100 & ~n11908 ;
  assign n29314 = n29313 ^ n7102 ^ 1'b0 ;
  assign n29315 = n22656 | n29314 ;
  assign n29316 = n29315 ^ n21679 ^ 1'b0 ;
  assign n29312 = n895 | n17227 ;
  assign n29317 = n29316 ^ n29312 ^ 1'b0 ;
  assign n29322 = n3649 & ~n15306 ;
  assign n29318 = n4072 & n4261 ;
  assign n29319 = n16094 & n29318 ;
  assign n29320 = n12783 | n29319 ;
  assign n29321 = n29320 ^ n4520 ^ 1'b0 ;
  assign n29323 = n29322 ^ n29321 ^ 1'b0 ;
  assign n29324 = n3543 | n29323 ;
  assign n29325 = n12363 ^ n9054 ^ 1'b0 ;
  assign n29326 = n29325 ^ n22697 ^ 1'b0 ;
  assign n29327 = n3097 ^ n2998 ^ 1'b0 ;
  assign n29328 = n23587 ^ n312 ^ 1'b0 ;
  assign n29329 = n29327 & n29328 ;
  assign n29330 = n29329 ^ n27517 ^ 1'b0 ;
  assign n29331 = n4411 & ~n10780 ;
  assign n29332 = n11655 & n29331 ;
  assign n29333 = n21201 | n29332 ;
  assign n29335 = n11844 ^ n11152 ^ 1'b0 ;
  assign n29334 = ~n11329 & n26349 ;
  assign n29336 = n29335 ^ n29334 ^ 1'b0 ;
  assign n29337 = ~n4298 & n22609 ;
  assign n29338 = ~x107 & n29337 ;
  assign n29339 = n12636 & n17104 ;
  assign n29340 = ~n1933 & n29339 ;
  assign n29341 = n29338 & n29340 ;
  assign n29342 = n3912 ^ n2463 ^ 1'b0 ;
  assign n29343 = n22259 | n26271 ;
  assign n29344 = n20335 ^ n15951 ^ 1'b0 ;
  assign n29345 = ~n18872 & n29344 ;
  assign n29346 = n4277 | n11168 ;
  assign n29347 = ~n12198 & n29346 ;
  assign n29348 = n29347 ^ n411 ^ 1'b0 ;
  assign n29349 = n29348 ^ n21271 ^ n5181 ;
  assign n29350 = n4421 & n29349 ;
  assign n29351 = n22810 ^ n8858 ^ 1'b0 ;
  assign n29352 = n14663 & n23874 ;
  assign n29353 = n29352 ^ n4019 ^ 1'b0 ;
  assign n29354 = n29353 ^ n17902 ^ 1'b0 ;
  assign n29355 = ~n29351 & n29354 ;
  assign n29356 = n3683 & n4707 ;
  assign n29357 = n17806 & n29356 ;
  assign n29358 = n14514 ^ n8144 ^ 1'b0 ;
  assign n29359 = n13894 ^ n6461 ^ 1'b0 ;
  assign n29360 = n15854 & n29359 ;
  assign n29361 = n7806 ^ n4216 ^ 1'b0 ;
  assign n29362 = n26164 ^ n12127 ^ n9780 ;
  assign n29363 = ( ~n1666 & n17285 ) | ( ~n1666 & n29362 ) | ( n17285 & n29362 ) ;
  assign n29364 = n16993 ^ n9591 ^ 1'b0 ;
  assign n29365 = n14017 & n24047 ;
  assign n29366 = n11252 & ~n13677 ;
  assign n29367 = x183 | n21522 ;
  assign n29368 = ( n1181 & ~n11793 ) | ( n1181 & n18350 ) | ( ~n11793 & n18350 ) ;
  assign n29369 = n28943 & n29368 ;
  assign n29370 = n11105 & ~n29000 ;
  assign n29371 = n29370 ^ n27787 ^ 1'b0 ;
  assign n29372 = n10274 ^ n2341 ^ 1'b0 ;
  assign n29373 = n16185 | n29372 ;
  assign n29374 = n4367 & ~n24367 ;
  assign n29375 = ~n29373 & n29374 ;
  assign n29376 = n18448 ^ n11441 ^ n7708 ;
  assign n29377 = n23140 ^ n20708 ^ n9666 ;
  assign n29378 = ~n13074 & n29377 ;
  assign n29379 = n5535 & n18980 ;
  assign n29380 = ~n5030 & n29379 ;
  assign n29381 = n28863 & ~n29380 ;
  assign n29382 = n4933 ^ n4898 ^ 1'b0 ;
  assign n29383 = n9802 | n29382 ;
  assign n29384 = n2616 | n29383 ;
  assign n29385 = n12078 ^ n10634 ^ 1'b0 ;
  assign n29386 = n14906 & n20654 ;
  assign n29387 = ( n1058 & n2645 ) | ( n1058 & n29386 ) | ( n2645 & n29386 ) ;
  assign n29388 = n15818 & ~n22400 ;
  assign n29389 = ~n12098 & n29388 ;
  assign n29390 = ( ~n14400 & n17826 ) | ( ~n14400 & n29389 ) | ( n17826 & n29389 ) ;
  assign n29391 = n2419 | n12256 ;
  assign n29392 = n20606 & ~n29391 ;
  assign n29393 = n1607 | n29392 ;
  assign n29394 = ( ~n11961 & n13280 ) | ( ~n11961 & n27926 ) | ( n13280 & n27926 ) ;
  assign n29395 = n29394 ^ n27026 ^ n5731 ;
  assign n29396 = ~n5065 & n11072 ;
  assign n29397 = x125 & ~n8664 ;
  assign n29398 = ~n12582 & n29397 ;
  assign n29399 = ( n15161 & n18963 ) | ( n15161 & ~n29398 ) | ( n18963 & ~n29398 ) ;
  assign n29400 = n29399 ^ n11043 ^ 1'b0 ;
  assign n29401 = n2748 & ~n4548 ;
  assign n29402 = n26726 ^ n22991 ^ 1'b0 ;
  assign n29403 = n13209 | n29402 ;
  assign n29404 = n29403 ^ n9353 ^ 1'b0 ;
  assign n29405 = ( n9156 & n29401 ) | ( n9156 & n29404 ) | ( n29401 & n29404 ) ;
  assign n29406 = n4749 ^ n4654 ^ 1'b0 ;
  assign n29408 = n17051 ^ n1258 ^ 1'b0 ;
  assign n29407 = n2551 & ~n15392 ;
  assign n29409 = n29408 ^ n29407 ^ 1'b0 ;
  assign n29410 = n29409 ^ n21332 ^ 1'b0 ;
  assign n29411 = x224 & n29410 ;
  assign n29412 = n19757 ^ n7277 ^ 1'b0 ;
  assign n29413 = n29412 ^ n16391 ^ n9217 ;
  assign n29414 = n29413 ^ n12809 ^ 1'b0 ;
  assign n29415 = n9219 | n18029 ;
  assign n29416 = ~n15033 & n17609 ;
  assign n29417 = n20494 ^ n5832 ^ 1'b0 ;
  assign n29418 = n11243 & n11795 ;
  assign n29419 = n14869 ^ x129 ^ 1'b0 ;
  assign n29422 = ~n6723 & n7447 ;
  assign n29420 = ~n12621 & n14439 ;
  assign n29421 = ~n14439 & n29420 ;
  assign n29423 = n29422 ^ n29421 ^ n4657 ;
  assign n29424 = n4115 & n14502 ;
  assign n29425 = n909 | n4666 ;
  assign n29426 = n29424 & n29425 ;
  assign n29427 = n29426 ^ n21249 ^ 1'b0 ;
  assign n29428 = n7444 | n29427 ;
  assign n29429 = ( n14044 & n24013 ) | ( n14044 & ~n29428 ) | ( n24013 & ~n29428 ) ;
  assign n29430 = n28269 ^ n600 ^ 1'b0 ;
  assign n29431 = ~n3305 & n29430 ;
  assign n29432 = n20958 ^ n14753 ^ n8466 ;
  assign n29433 = n8194 | n29432 ;
  assign n29434 = n29431 | n29433 ;
  assign n29435 = n4592 | n20293 ;
  assign n29436 = n29435 ^ n9030 ^ 1'b0 ;
  assign n29437 = ~n9414 & n24216 ;
  assign n29438 = n29437 ^ n9538 ^ 1'b0 ;
  assign n29443 = n1224 & ~n12478 ;
  assign n29444 = ( n631 & n2717 ) | ( n631 & n29443 ) | ( n2717 & n29443 ) ;
  assign n29440 = ( n6758 & n6990 ) | ( n6758 & n7161 ) | ( n6990 & n7161 ) ;
  assign n29439 = n5862 ^ n3433 ^ 1'b0 ;
  assign n29441 = n29440 ^ n29439 ^ 1'b0 ;
  assign n29442 = n26595 | n29441 ;
  assign n29445 = n29444 ^ n29442 ^ 1'b0 ;
  assign n29446 = n21970 ^ n1374 ^ n1079 ;
  assign n29447 = ( ~n7403 & n14909 ) | ( ~n7403 & n25664 ) | ( n14909 & n25664 ) ;
  assign n29448 = ~n16066 & n28983 ;
  assign n29449 = ~n1136 & n22227 ;
  assign n29450 = ~n26946 & n29449 ;
  assign n29451 = x224 & n28593 ;
  assign n29454 = n16862 ^ n12091 ^ 1'b0 ;
  assign n29452 = n300 & n4814 ;
  assign n29453 = n6376 & n29452 ;
  assign n29455 = n29454 ^ n29453 ^ n17635 ;
  assign n29456 = ( n7322 & n9642 ) | ( n7322 & ~n18798 ) | ( n9642 & ~n18798 ) ;
  assign n29457 = ~n29166 & n29456 ;
  assign n29458 = ~n5619 & n29457 ;
  assign n29459 = ( ~n1944 & n6678 ) | ( ~n1944 & n20982 ) | ( n6678 & n20982 ) ;
  assign n29460 = n29459 ^ n23592 ^ n2111 ;
  assign n29463 = n16115 ^ n8810 ^ 1'b0 ;
  assign n29464 = n11806 | n29463 ;
  assign n29465 = ( ~x177 & n10052 ) | ( ~x177 & n29464 ) | ( n10052 & n29464 ) ;
  assign n29461 = n1251 | n6300 ;
  assign n29462 = n29461 ^ n5458 ^ 1'b0 ;
  assign n29466 = n29465 ^ n29462 ^ 1'b0 ;
  assign n29467 = ~n8721 & n29466 ;
  assign n29468 = n20613 ^ n13686 ^ n6968 ;
  assign n29469 = n18791 ^ n13670 ^ n3390 ;
  assign n29470 = n29469 ^ n3255 ^ 1'b0 ;
  assign n29471 = ~n29468 & n29470 ;
  assign n29472 = n11454 & n29471 ;
  assign n29473 = ~n6247 & n6865 ;
  assign n29474 = n12394 & ~n29473 ;
  assign n29475 = n29474 ^ n7113 ^ 1'b0 ;
  assign n29476 = n279 & n7647 ;
  assign n29477 = n29476 ^ n24740 ^ n5269 ;
  assign n29478 = n2630 & n22398 ;
  assign n29479 = n29478 ^ n12124 ^ 1'b0 ;
  assign n29480 = n12483 & n29479 ;
  assign n29481 = ~n15179 & n29480 ;
  assign n29482 = n29481 ^ n25878 ^ 1'b0 ;
  assign n29483 = ( n3529 & n3657 ) | ( n3529 & n4350 ) | ( n3657 & n4350 ) ;
  assign n29484 = ( n10116 & n13198 ) | ( n10116 & ~n29483 ) | ( n13198 & ~n29483 ) ;
  assign n29485 = n29484 ^ n13957 ^ n8614 ;
  assign n29486 = n3320 & n10754 ;
  assign n29487 = n29486 ^ n21473 ^ n337 ;
  assign n29488 = n29487 ^ n13688 ^ n3207 ;
  assign n29489 = ( n2695 & ~n29485 ) | ( n2695 & n29488 ) | ( ~n29485 & n29488 ) ;
  assign n29491 = ~n12305 & n21508 ;
  assign n29490 = n2601 ^ n1576 ^ 1'b0 ;
  assign n29492 = n29491 ^ n29490 ^ 1'b0 ;
  assign n29493 = n29489 & n29492 ;
  assign n29494 = n18729 ^ n7235 ^ 1'b0 ;
  assign n29495 = n18830 ^ n11680 ^ n10208 ;
  assign n29496 = n13933 ^ n3956 ^ 1'b0 ;
  assign n29497 = n7747 & ~n9837 ;
  assign n29498 = n13129 ^ n11223 ^ 1'b0 ;
  assign n29499 = ( n15445 & ~n27972 ) | ( n15445 & n29498 ) | ( ~n27972 & n29498 ) ;
  assign n29500 = n11401 & n13260 ;
  assign n29501 = n28767 ^ n5485 ^ 1'b0 ;
  assign n29502 = n14859 | n29501 ;
  assign n29503 = n12400 | n29502 ;
  assign n29504 = n20512 ^ n18610 ^ n2608 ;
  assign n29505 = n24844 | n25831 ;
  assign n29507 = n18015 ^ n1296 ^ n507 ;
  assign n29506 = n3637 & n5476 ;
  assign n29508 = n29507 ^ n29506 ^ n16550 ;
  assign n29509 = ~n4383 & n14998 ;
  assign n29510 = ~n464 & n9780 ;
  assign n29511 = n29510 ^ n13453 ^ 1'b0 ;
  assign n29512 = n27340 ^ n7380 ^ 1'b0 ;
  assign n29513 = n4778 & n29512 ;
  assign n29514 = ( n19364 & n20465 ) | ( n19364 & n29513 ) | ( n20465 & n29513 ) ;
  assign n29515 = n26441 ^ n4500 ^ 1'b0 ;
  assign n29516 = n13270 & n29515 ;
  assign n29520 = n9292 ^ n6728 ^ 1'b0 ;
  assign n29521 = ( n6361 & ~n14796 ) | ( n6361 & n29520 ) | ( ~n14796 & n29520 ) ;
  assign n29518 = ~n1372 & n12094 ;
  assign n29519 = n18968 & n29518 ;
  assign n29522 = n29521 ^ n29519 ^ 1'b0 ;
  assign n29517 = x176 & ~n28219 ;
  assign n29523 = n29522 ^ n29517 ^ 1'b0 ;
  assign n29524 = ( ~n4720 & n6888 ) | ( ~n4720 & n8473 ) | ( n6888 & n8473 ) ;
  assign n29525 = ( n2216 & n4022 ) | ( n2216 & ~n16829 ) | ( n4022 & ~n16829 ) ;
  assign n29526 = ~n29524 & n29525 ;
  assign n29527 = n9737 & ~n14655 ;
  assign n29528 = n8158 & ~n19304 ;
  assign n29529 = n29528 ^ n16940 ^ 1'b0 ;
  assign n29530 = n15730 ^ n4553 ^ 1'b0 ;
  assign n29531 = n10884 ^ n8573 ^ 1'b0 ;
  assign n29532 = n17197 & ~n18004 ;
  assign n29533 = n29532 ^ n19795 ^ 1'b0 ;
  assign n29536 = n5287 ^ n5028 ^ 1'b0 ;
  assign n29537 = n29536 ^ n8209 ^ n1452 ;
  assign n29534 = n7837 ^ n5736 ^ 1'b0 ;
  assign n29535 = n1717 & ~n29534 ;
  assign n29538 = n29537 ^ n29535 ^ 1'b0 ;
  assign n29542 = ~n4641 & n5358 ;
  assign n29543 = n4447 & n29542 ;
  assign n29544 = n29543 ^ n10581 ^ n3274 ;
  assign n29539 = n7758 ^ n6912 ^ 1'b0 ;
  assign n29540 = ~n18732 & n29539 ;
  assign n29541 = n23337 & n29540 ;
  assign n29545 = n29544 ^ n29541 ^ 1'b0 ;
  assign n29549 = n528 & n1936 ;
  assign n29550 = n4966 & n29549 ;
  assign n29546 = n2961 | n8101 ;
  assign n29547 = n8201 | n29546 ;
  assign n29548 = n8091 & n29547 ;
  assign n29551 = n29550 ^ n29548 ^ 1'b0 ;
  assign n29552 = n18956 & n29551 ;
  assign n29553 = n13682 & ~n23609 ;
  assign n29554 = n29553 ^ n6738 ^ n2077 ;
  assign n29555 = n11135 & ~n15208 ;
  assign n29556 = n29555 ^ n2419 ^ 1'b0 ;
  assign n29557 = n9533 | n16709 ;
  assign n29558 = n29556 | n29557 ;
  assign n29559 = n23123 ^ n12667 ^ 1'b0 ;
  assign n29560 = ( n19907 & n29558 ) | ( n19907 & ~n29559 ) | ( n29558 & ~n29559 ) ;
  assign n29561 = ~n7799 & n23391 ;
  assign n29562 = ( ~n12616 & n20031 ) | ( ~n12616 & n22381 ) | ( n20031 & n22381 ) ;
  assign n29563 = ~n7385 & n27238 ;
  assign n29564 = n29562 & n29563 ;
  assign n29565 = n9184 ^ n1082 ^ 1'b0 ;
  assign n29566 = n10922 & ~n29565 ;
  assign n29567 = n13212 & n13506 ;
  assign n29568 = ~n4150 & n29567 ;
  assign n29569 = ( ~n6357 & n29566 ) | ( ~n6357 & n29568 ) | ( n29566 & n29568 ) ;
  assign n29570 = n1420 | n9452 ;
  assign n29571 = n29570 ^ n26590 ^ n4542 ;
  assign n29572 = n10264 | n27609 ;
  assign n29573 = n7078 & ~n29572 ;
  assign n29574 = n18635 ^ n876 ^ 1'b0 ;
  assign n29575 = n16011 | n29574 ;
  assign n29576 = n6255 & ~n29575 ;
  assign n29577 = n29573 & n29576 ;
  assign n29578 = n2959 & ~n6581 ;
  assign n29579 = n7792 | n29578 ;
  assign n29580 = n29579 ^ n26668 ^ 1'b0 ;
  assign n29581 = n18849 ^ n1132 ^ 1'b0 ;
  assign n29582 = n10129 ^ n5206 ^ 1'b0 ;
  assign n29583 = n15435 | n29582 ;
  assign n29584 = ( n4709 & n5535 ) | ( n4709 & ~n7948 ) | ( n5535 & ~n7948 ) ;
  assign n29585 = n29584 ^ n11076 ^ 1'b0 ;
  assign n29586 = n8611 | n22655 ;
  assign n29587 = n2142 | n29586 ;
  assign n29588 = n4700 & ~n28066 ;
  assign n29589 = ~n29587 & n29588 ;
  assign n29590 = n3745 & ~n29589 ;
  assign n29591 = n8435 & ~n29590 ;
  assign n29592 = n29585 & n29591 ;
  assign n29593 = n5800 ^ n1922 ^ 1'b0 ;
  assign n29594 = ~n13010 & n29593 ;
  assign n29595 = n23109 ^ n14618 ^ 1'b0 ;
  assign n29596 = n29594 & ~n29595 ;
  assign n29597 = n1031 ^ n973 ^ 1'b0 ;
  assign n29598 = n2608 & ~n29597 ;
  assign n29599 = n7769 & n29598 ;
  assign n29600 = ~n4020 & n22155 ;
  assign n29601 = n29600 ^ n6127 ^ n300 ;
  assign n29602 = n7470 & n18350 ;
  assign n29603 = n16964 | n29602 ;
  assign n29604 = ( ~n7433 & n24976 ) | ( ~n7433 & n29603 ) | ( n24976 & n29603 ) ;
  assign n29605 = n14790 | n21762 ;
  assign n29606 = n25525 ^ x235 ^ 1'b0 ;
  assign n29607 = n29605 & ~n29606 ;
  assign n29608 = n23396 & ~n25831 ;
  assign n29609 = n13321 ^ n5981 ^ n1148 ;
  assign n29610 = n11201 & n21035 ;
  assign n29614 = ~n3947 & n8218 ;
  assign n29615 = n29614 ^ n1595 ^ 1'b0 ;
  assign n29611 = n18945 ^ n6910 ^ 1'b0 ;
  assign n29612 = n2372 & n29611 ;
  assign n29613 = n11471 & ~n29612 ;
  assign n29616 = n29615 ^ n29613 ^ 1'b0 ;
  assign n29617 = n339 & n2680 ;
  assign n29618 = n2827 | n9547 ;
  assign n29619 = n2740 & ~n10443 ;
  assign n29620 = n29619 ^ n11617 ^ 1'b0 ;
  assign n29621 = n13317 | n29620 ;
  assign n29622 = n13255 ^ n13177 ^ 1'b0 ;
  assign n29623 = n9139 & ~n29622 ;
  assign n29624 = n7983 ^ x41 ^ 1'b0 ;
  assign n29625 = ( n7197 & n7887 ) | ( n7197 & ~n17514 ) | ( n7887 & ~n17514 ) ;
  assign n29626 = n29624 & ~n29625 ;
  assign n29627 = ~n29624 & n29626 ;
  assign n29628 = n2133 ^ n1486 ^ 1'b0 ;
  assign n29629 = n17414 | n29628 ;
  assign n29630 = n5462 | n29629 ;
  assign n29631 = n29630 ^ n6528 ^ 1'b0 ;
  assign n29632 = n29627 | n29631 ;
  assign n29633 = n3259 & n17396 ;
  assign n29634 = ~n7063 & n29633 ;
  assign n29635 = ~n13526 & n26731 ;
  assign n29636 = n29635 ^ n3059 ^ 1'b0 ;
  assign n29637 = n29636 ^ n6914 ^ 1'b0 ;
  assign n29638 = n469 | n6024 ;
  assign n29639 = n19060 & ~n29638 ;
  assign n29641 = ~n3452 & n5873 ;
  assign n29640 = n10806 ^ n2573 ^ 1'b0 ;
  assign n29642 = n29641 ^ n29640 ^ n8965 ;
  assign n29643 = n18606 | n29642 ;
  assign n29644 = n10087 ^ n7475 ^ 1'b0 ;
  assign n29652 = n15180 & ~n25270 ;
  assign n29653 = n5215 ^ n5198 ^ 1'b0 ;
  assign n29654 = ( n14637 & ~n24086 ) | ( n14637 & n29653 ) | ( ~n24086 & n29653 ) ;
  assign n29655 = n29652 & ~n29654 ;
  assign n29656 = n29655 ^ n7560 ^ 1'b0 ;
  assign n29645 = n11349 ^ n2052 ^ 1'b0 ;
  assign n29646 = n7513 & n29645 ;
  assign n29648 = n5705 ^ n2013 ^ 1'b0 ;
  assign n29649 = n1387 & n29648 ;
  assign n29647 = n20905 ^ n18419 ^ 1'b0 ;
  assign n29650 = n29649 ^ n29647 ^ 1'b0 ;
  assign n29651 = ( n1037 & n29646 ) | ( n1037 & ~n29650 ) | ( n29646 & ~n29650 ) ;
  assign n29657 = n29656 ^ n29651 ^ n27302 ;
  assign n29658 = n29657 ^ n24101 ^ n3590 ;
  assign n29659 = n19075 ^ n3045 ^ 1'b0 ;
  assign n29660 = ~n11034 & n29659 ;
  assign n29661 = n10918 ^ n10439 ^ n2758 ;
  assign n29662 = n29661 ^ n14163 ^ 1'b0 ;
  assign n29663 = ~n12480 & n29662 ;
  assign n29664 = ( n18138 & n24169 ) | ( n18138 & n29663 ) | ( n24169 & n29663 ) ;
  assign n29665 = n16067 ^ n9858 ^ 1'b0 ;
  assign n29666 = n29664 & ~n29665 ;
  assign n29667 = ( n1111 & ~n29660 ) | ( n1111 & n29666 ) | ( ~n29660 & n29666 ) ;
  assign n29668 = n19425 ^ n9065 ^ 1'b0 ;
  assign n29669 = n20367 & ~n29668 ;
  assign n29670 = n8284 ^ n2315 ^ 1'b0 ;
  assign n29671 = n24243 & ~n29670 ;
  assign n29672 = n7800 & n11084 ;
  assign n29673 = n6854 & n10667 ;
  assign n29674 = n2506 ^ n1688 ^ 1'b0 ;
  assign n29675 = n29673 & ~n29674 ;
  assign n29676 = n15721 ^ n1217 ^ n759 ;
  assign n29677 = n29676 ^ n19092 ^ n9207 ;
  assign n29678 = n14102 ^ n12863 ^ 1'b0 ;
  assign n29679 = ~n5067 & n29678 ;
  assign n29680 = n29679 ^ n19519 ^ 1'b0 ;
  assign n29681 = n4766 | n29680 ;
  assign n29682 = ( n7670 & n11708 ) | ( n7670 & n29681 ) | ( n11708 & n29681 ) ;
  assign n29683 = n5022 & n11416 ;
  assign n29684 = n29683 ^ n27393 ^ 1'b0 ;
  assign n29685 = ( n6324 & n8362 ) | ( n6324 & n12127 ) | ( n8362 & n12127 ) ;
  assign n29686 = n29685 ^ n24985 ^ 1'b0 ;
  assign n29687 = n29684 & ~n29686 ;
  assign n29688 = n29687 ^ n19840 ^ n9776 ;
  assign n29689 = n394 & n17870 ;
  assign n29690 = n2504 & n29689 ;
  assign n29691 = n29690 ^ n6950 ^ n349 ;
  assign n29692 = n2764 & ~n27736 ;
  assign n29693 = ~n13291 & n29692 ;
  assign n29694 = n8084 & ~n19757 ;
  assign n29695 = n29694 ^ n5745 ^ 1'b0 ;
  assign n29696 = n29695 ^ n16163 ^ 1'b0 ;
  assign n29697 = ~n6679 & n13593 ;
  assign n29698 = ~n10075 & n29697 ;
  assign n29699 = n13531 ^ n7475 ^ 1'b0 ;
  assign n29700 = n11837 | n29699 ;
  assign n29701 = ( n22050 & ~n29698 ) | ( n22050 & n29700 ) | ( ~n29698 & n29700 ) ;
  assign n29702 = n10720 | n28939 ;
  assign n29703 = ~n10498 & n15275 ;
  assign n29704 = n16064 ^ n15648 ^ 1'b0 ;
  assign n29705 = n1600 & ~n4941 ;
  assign n29706 = n2022 | n29705 ;
  assign n29707 = n20010 | n29706 ;
  assign n29708 = n29707 ^ n13405 ^ 1'b0 ;
  assign n29709 = n29704 & n29708 ;
  assign n29710 = n10791 ^ n6357 ^ n5892 ;
  assign n29711 = n29710 ^ n8533 ^ 1'b0 ;
  assign n29712 = ~n861 & n11163 ;
  assign n29713 = n29712 ^ n22162 ^ n17633 ;
  assign n29714 = n11801 ^ n3849 ^ 1'b0 ;
  assign n29715 = n15063 | n29714 ;
  assign n29716 = n7841 & ~n29715 ;
  assign n29717 = n11469 & n29716 ;
  assign n29718 = n3126 & n6441 ;
  assign n29719 = n11535 & n12910 ;
  assign n29720 = ~x104 & n29719 ;
  assign n29721 = n13068 & n27646 ;
  assign n29722 = n1402 & ~n16444 ;
  assign n29723 = n9714 & n29722 ;
  assign n29724 = n6447 ^ n2314 ^ 1'b0 ;
  assign n29725 = ~n29723 & n29724 ;
  assign n29726 = ~n4469 & n29725 ;
  assign n29727 = n29721 & n29726 ;
  assign n29728 = n16109 | n29727 ;
  assign n29729 = n27328 ^ n8541 ^ 1'b0 ;
  assign n29730 = n10413 | n29729 ;
  assign n29731 = ( x73 & n368 ) | ( x73 & ~n29730 ) | ( n368 & ~n29730 ) ;
  assign n29732 = n8038 & ~n19353 ;
  assign n29733 = ~n5606 & n29732 ;
  assign n29734 = n29090 | n29733 ;
  assign n29735 = ( n2082 & n20631 ) | ( n2082 & n28444 ) | ( n20631 & n28444 ) ;
  assign n29736 = n18409 | n25690 ;
  assign n29737 = n29736 ^ n10942 ^ 1'b0 ;
  assign n29738 = ~n9419 & n22035 ;
  assign n29739 = n6162 & ~n29738 ;
  assign n29740 = n29739 ^ n15966 ^ 1'b0 ;
  assign n29741 = n7939 | n10380 ;
  assign n29742 = n11533 & n29741 ;
  assign n29743 = ~n20932 & n29742 ;
  assign n29744 = n29743 ^ n20811 ^ 1'b0 ;
  assign n29745 = n862 & n13698 ;
  assign n29746 = n2984 & ~n10411 ;
  assign n29747 = ~n3948 & n29746 ;
  assign n29748 = n29747 ^ n6436 ^ 1'b0 ;
  assign n29749 = n29748 ^ n25849 ^ n25629 ;
  assign n29750 = n8508 ^ n7039 ^ 1'b0 ;
  assign n29751 = ( n5071 & n11593 ) | ( n5071 & ~n29750 ) | ( n11593 & ~n29750 ) ;
  assign n29752 = n10117 ^ n260 ^ 1'b0 ;
  assign n29753 = n11187 ^ n1757 ^ 1'b0 ;
  assign n29754 = ~n29752 & n29753 ;
  assign n29755 = ~n22989 & n28280 ;
  assign n29756 = n14988 & n29755 ;
  assign n29757 = n13236 & ~n17337 ;
  assign n29758 = ~n8716 & n25465 ;
  assign n29759 = ~n1106 & n1628 ;
  assign n29760 = n29759 ^ n29736 ^ 1'b0 ;
  assign n29762 = n9824 | n15303 ;
  assign n29761 = n3658 & ~n20342 ;
  assign n29763 = n29762 ^ n29761 ^ 1'b0 ;
  assign n29764 = ~n26645 & n29763 ;
  assign n29765 = n13429 & n29764 ;
  assign n29766 = n15486 ^ n3351 ^ 1'b0 ;
  assign n29767 = ~n9988 & n26564 ;
  assign n29768 = n10992 & ~n12290 ;
  assign n29769 = ~n4083 & n29768 ;
  assign n29770 = n29769 ^ n6597 ^ 1'b0 ;
  assign n29771 = n29770 ^ n29007 ^ n17971 ;
  assign n29772 = n28133 ^ n21530 ^ n9611 ;
  assign n29773 = n562 & ~n9752 ;
  assign n29774 = n29773 ^ n9521 ^ 1'b0 ;
  assign n29775 = x186 & ~n4154 ;
  assign n29776 = n29775 ^ n10371 ^ n3526 ;
  assign n29777 = n12026 & ~n29776 ;
  assign n29778 = ~n29774 & n29777 ;
  assign n29779 = n19619 ^ n2119 ^ 1'b0 ;
  assign n29780 = n7064 | n10340 ;
  assign n29781 = n10845 & n15686 ;
  assign n29782 = n15451 & n29781 ;
  assign n29783 = ( n16100 & ~n26520 ) | ( n16100 & n29782 ) | ( ~n26520 & n29782 ) ;
  assign n29784 = ~n5894 & n16977 ;
  assign n29785 = ~n21310 & n29784 ;
  assign n29786 = n3477 & ~n9002 ;
  assign n29787 = n10117 ^ n3790 ^ 1'b0 ;
  assign n29788 = n29787 ^ n18557 ^ 1'b0 ;
  assign n29789 = ( n11823 & n17206 ) | ( n11823 & n29788 ) | ( n17206 & n29788 ) ;
  assign n29790 = ~n14172 & n29600 ;
  assign n29791 = n16571 & ~n29790 ;
  assign n29792 = n20917 ^ n16687 ^ 1'b0 ;
  assign n29793 = n12344 & ~n29792 ;
  assign n29794 = n4389 & n8551 ;
  assign n29795 = ~n6476 & n29794 ;
  assign n29796 = n4818 | n8659 ;
  assign n29797 = n29796 ^ n7876 ^ 1'b0 ;
  assign n29798 = n29797 ^ n8646 ^ 1'b0 ;
  assign n29799 = n2828 & n29798 ;
  assign n29800 = n29795 & n29799 ;
  assign n29801 = ~n10065 & n20703 ;
  assign n29802 = n12350 ^ n5197 ^ x103 ;
  assign n29803 = n4992 & ~n7385 ;
  assign n29804 = n29803 ^ n14322 ^ 1'b0 ;
  assign n29805 = n29802 | n29804 ;
  assign n29806 = n29805 ^ n4067 ^ 1'b0 ;
  assign n29807 = n3047 ^ n2126 ^ 1'b0 ;
  assign n29808 = n26572 & n29807 ;
  assign n29809 = n13112 & n29808 ;
  assign n29810 = n1069 & ~n20846 ;
  assign n29811 = n14598 | n29810 ;
  assign n29812 = n14580 & ~n29811 ;
  assign n29813 = n29812 ^ n23110 ^ 1'b0 ;
  assign n29814 = n29809 & n29813 ;
  assign n29815 = n10116 | n24354 ;
  assign n29816 = n29815 ^ n5197 ^ 1'b0 ;
  assign n29817 = ( ~n6531 & n26470 ) | ( ~n6531 & n29816 ) | ( n26470 & n29816 ) ;
  assign n29818 = n11578 & ~n29817 ;
  assign n29819 = ~n783 & n4207 ;
  assign n29820 = ~n22004 & n29819 ;
  assign n29821 = n2334 & ~n15771 ;
  assign n29822 = ~n2678 & n29821 ;
  assign n29823 = n29640 | n29822 ;
  assign n29824 = n18977 | n29823 ;
  assign n29825 = ~n857 & n23729 ;
  assign n29826 = ( ~n28045 & n29824 ) | ( ~n28045 & n29825 ) | ( n29824 & n29825 ) ;
  assign n29827 = ~n8009 & n23162 ;
  assign n29828 = ( n20443 & ~n29826 ) | ( n20443 & n29827 ) | ( ~n29826 & n29827 ) ;
  assign n29829 = n3717 & n29399 ;
  assign n29830 = n27313 ^ n13017 ^ 1'b0 ;
  assign n29831 = ( ~n6345 & n8688 ) | ( ~n6345 & n11015 ) | ( n8688 & n11015 ) ;
  assign n29832 = n21106 ^ n332 ^ 1'b0 ;
  assign n29833 = n29832 ^ n16443 ^ 1'b0 ;
  assign n29834 = n29831 & ~n29833 ;
  assign n29835 = ( n8754 & n15185 ) | ( n8754 & n29834 ) | ( n15185 & n29834 ) ;
  assign n29836 = n29835 ^ n27302 ^ 1'b0 ;
  assign n29838 = n5899 | n14145 ;
  assign n29839 = n29838 ^ n5881 ^ 1'b0 ;
  assign n29840 = n2892 & n29839 ;
  assign n29841 = n29840 ^ n10106 ^ 1'b0 ;
  assign n29837 = n17780 ^ n6684 ^ 1'b0 ;
  assign n29842 = n29841 ^ n29837 ^ n2231 ;
  assign n29843 = n7040 | n24237 ;
  assign n29844 = ( x87 & ~n3264 ) | ( x87 & n8930 ) | ( ~n3264 & n8930 ) ;
  assign n29845 = n22952 & n29844 ;
  assign n29846 = ( ~n12321 & n13084 ) | ( ~n12321 & n16717 ) | ( n13084 & n16717 ) ;
  assign n29847 = n29846 ^ n3905 ^ 1'b0 ;
  assign n29848 = x173 & ~n1853 ;
  assign n29849 = ~n4090 & n29848 ;
  assign n29850 = n29849 ^ n23729 ^ 1'b0 ;
  assign n29851 = n26301 & ~n29850 ;
  assign n29852 = ( ~n1197 & n3540 ) | ( ~n1197 & n14023 ) | ( n3540 & n14023 ) ;
  assign n29853 = n15221 ^ n7822 ^ 1'b0 ;
  assign n29854 = n29852 | n29853 ;
  assign n29855 = n28036 & ~n29854 ;
  assign n29856 = n12194 & ~n28967 ;
  assign n29857 = n29856 ^ n15101 ^ 1'b0 ;
  assign n29858 = n9478 & ~n21370 ;
  assign n29859 = n10168 ^ n1755 ^ 1'b0 ;
  assign n29860 = n1080 & ~n26385 ;
  assign n29861 = n29860 ^ n25498 ^ 1'b0 ;
  assign n29862 = n5828 | n13740 ;
  assign n29863 = n29862 ^ n7891 ^ 1'b0 ;
  assign n29864 = n10142 ^ n7231 ^ 1'b0 ;
  assign n29865 = ~n29863 & n29864 ;
  assign n29866 = n29865 ^ n22873 ^ n4690 ;
  assign n29867 = n8902 | n10549 ;
  assign n29868 = n29867 ^ n16455 ^ 1'b0 ;
  assign n29869 = n1168 | n15738 ;
  assign n29870 = n29869 ^ n26578 ^ 1'b0 ;
  assign n29871 = n15788 ^ n14577 ^ 1'b0 ;
  assign n29872 = n28889 ^ n8697 ^ n4529 ;
  assign n29873 = n29872 ^ n14318 ^ n671 ;
  assign n29874 = ( n471 & ~n3997 ) | ( n471 & n29873 ) | ( ~n3997 & n29873 ) ;
  assign n29875 = n7223 | n22687 ;
  assign n29876 = ( n2645 & n27084 ) | ( n2645 & ~n29875 ) | ( n27084 & ~n29875 ) ;
  assign n29877 = n19406 ^ n11013 ^ 1'b0 ;
  assign n29878 = ~n29876 & n29877 ;
  assign n29879 = n18560 ^ n11389 ^ 1'b0 ;
  assign n29880 = ~n6357 & n29879 ;
  assign n29881 = ( n15690 & n29878 ) | ( n15690 & ~n29880 ) | ( n29878 & ~n29880 ) ;
  assign n29882 = n8072 & ~n24293 ;
  assign n29883 = ( n10982 & ~n14489 ) | ( n10982 & n21855 ) | ( ~n14489 & n21855 ) ;
  assign n29884 = ~n5174 & n6030 ;
  assign n29885 = ~n29883 & n29884 ;
  assign n29886 = n19300 & ~n26197 ;
  assign n29887 = n16573 & n29886 ;
  assign n29888 = ( n2529 & ~n3588 ) | ( n2529 & n5341 ) | ( ~n3588 & n5341 ) ;
  assign n29889 = n29888 ^ n14102 ^ n8001 ;
  assign n29890 = ( n13310 & ~n24196 ) | ( n13310 & n26369 ) | ( ~n24196 & n26369 ) ;
  assign n29891 = n23212 ^ n5347 ^ n2389 ;
  assign n29892 = n10593 ^ n8504 ^ 1'b0 ;
  assign n29893 = n4935 & n11078 ;
  assign n29894 = ~n9874 & n29893 ;
  assign n29895 = n29892 & ~n29894 ;
  assign n29896 = n18235 & n29895 ;
  assign n29897 = n23417 | n29896 ;
  assign n29898 = n29897 ^ n4308 ^ 1'b0 ;
  assign n29899 = n29891 & n29898 ;
  assign n29900 = n17799 ^ n1476 ^ 1'b0 ;
  assign n29901 = n5573 & ~n15943 ;
  assign n29902 = n29901 ^ n21635 ^ 1'b0 ;
  assign n29903 = n16521 ^ n14965 ^ 1'b0 ;
  assign n29904 = n26075 ^ n17063 ^ n8668 ;
  assign n29905 = n29904 ^ n25893 ^ n24334 ;
  assign n29906 = n27263 & ~n29905 ;
  assign n29907 = n29906 ^ n20983 ^ 1'b0 ;
  assign n29908 = n26704 ^ n24605 ^ 1'b0 ;
  assign n29909 = n29908 ^ n22095 ^ n19380 ;
  assign n29910 = ~n20524 & n29909 ;
  assign n29911 = n26550 & n29910 ;
  assign n29914 = n5522 ^ n5316 ^ n968 ;
  assign n29912 = n15486 & n21833 ;
  assign n29913 = n29912 ^ n5246 ^ 1'b0 ;
  assign n29915 = n29914 ^ n29913 ^ n18983 ;
  assign n29916 = ( n6253 & n8996 ) | ( n6253 & n16812 ) | ( n8996 & n16812 ) ;
  assign n29917 = n29916 ^ n16425 ^ n9750 ;
  assign n29918 = n29917 ^ n7851 ^ 1'b0 ;
  assign n29919 = n5307 & ~n16898 ;
  assign n29920 = ( ~n13809 & n22326 ) | ( ~n13809 & n29919 ) | ( n22326 & n29919 ) ;
  assign n29921 = n2137 | n8735 ;
  assign n29922 = n4729 | n8624 ;
  assign n29923 = n29922 ^ n28021 ^ 1'b0 ;
  assign n29924 = ~n29921 & n29923 ;
  assign n29925 = n3564 ^ n1354 ^ 1'b0 ;
  assign n29926 = ~n20115 & n29925 ;
  assign n29927 = n29926 ^ n22521 ^ 1'b0 ;
  assign n29929 = n2359 | n3792 ;
  assign n29928 = n10525 | n13806 ;
  assign n29930 = n29929 ^ n29928 ^ 1'b0 ;
  assign n29931 = n9406 ^ n2744 ^ n1869 ;
  assign n29932 = ~n9101 & n29931 ;
  assign n29933 = n29429 ^ n11741 ^ n887 ;
  assign n29934 = ( n7780 & ~n13183 ) | ( n7780 & n15107 ) | ( ~n13183 & n15107 ) ;
  assign n29935 = n1980 & ~n2847 ;
  assign n29936 = ~n18575 & n29935 ;
  assign n29937 = n27679 ^ n15450 ^ 1'b0 ;
  assign n29939 = n25592 ^ n18623 ^ 1'b0 ;
  assign n29938 = n8721 | n20825 ;
  assign n29940 = n29939 ^ n29938 ^ 1'b0 ;
  assign n29941 = n28217 ^ n5287 ^ 1'b0 ;
  assign n29942 = n23810 ^ n19696 ^ n16499 ;
  assign n29943 = ~n1519 & n29942 ;
  assign n29944 = n11970 ^ n6654 ^ 1'b0 ;
  assign n29945 = ( n763 & ~n10025 ) | ( n763 & n11279 ) | ( ~n10025 & n11279 ) ;
  assign n29946 = n23844 ^ n19058 ^ n6788 ;
  assign n29947 = ( n12259 & ~n12674 ) | ( n12259 & n29946 ) | ( ~n12674 & n29946 ) ;
  assign n29948 = n29945 & ~n29947 ;
  assign n29949 = n2109 & ~n8621 ;
  assign n29950 = n7077 ^ n3532 ^ 1'b0 ;
  assign n29951 = n29949 & ~n29950 ;
  assign n29952 = ~n25568 & n29951 ;
  assign n29953 = n29952 ^ n24709 ^ 1'b0 ;
  assign n29956 = n12050 ^ n11301 ^ 1'b0 ;
  assign n29957 = n29956 ^ n6085 ^ x6 ;
  assign n29955 = n1698 & n2531 ;
  assign n29954 = ~n14177 & n25877 ;
  assign n29958 = n29957 ^ n29955 ^ n29954 ;
  assign n29959 = ( ~n15305 & n29953 ) | ( ~n15305 & n29958 ) | ( n29953 & n29958 ) ;
  assign n29960 = n3816 ^ n1231 ^ 1'b0 ;
  assign n29961 = n2263 | n29960 ;
  assign n29962 = n27263 | n29961 ;
  assign n29965 = n20384 ^ n7262 ^ 1'b0 ;
  assign n29963 = n7617 ^ n2662 ^ 1'b0 ;
  assign n29964 = n11722 & n29963 ;
  assign n29966 = n29965 ^ n29964 ^ 1'b0 ;
  assign n29967 = n4197 ^ n1002 ^ 1'b0 ;
  assign n29968 = n28245 ^ n10096 ^ n9485 ;
  assign n29969 = n22617 & n29968 ;
  assign n29970 = n29969 ^ n10042 ^ 1'b0 ;
  assign n29971 = ( n1366 & n29967 ) | ( n1366 & ~n29970 ) | ( n29967 & ~n29970 ) ;
  assign n29972 = n9437 & n25718 ;
  assign n29973 = ( n3955 & n29971 ) | ( n3955 & n29972 ) | ( n29971 & n29972 ) ;
  assign n29974 = n20280 ^ n9897 ^ 1'b0 ;
  assign n29975 = n26675 ^ n14210 ^ 1'b0 ;
  assign n29976 = n1187 & n4639 ;
  assign n29977 = n17541 ^ n13459 ^ 1'b0 ;
  assign n29978 = ~n6174 & n29977 ;
  assign n29979 = ~n14805 & n27889 ;
  assign n29980 = n29979 ^ n8185 ^ 1'b0 ;
  assign n29981 = n11125 ^ n5109 ^ 1'b0 ;
  assign n29982 = n29981 ^ n23306 ^ n12750 ;
  assign n29983 = ( ~n15721 & n19911 ) | ( ~n15721 & n20015 ) | ( n19911 & n20015 ) ;
  assign n29984 = n29983 ^ n2779 ^ 1'b0 ;
  assign n29988 = n23468 ^ n14787 ^ n4881 ;
  assign n29989 = ~n3802 & n8221 ;
  assign n29990 = ~n29988 & n29989 ;
  assign n29985 = ( n2359 & ~n6098 ) | ( n2359 & n14603 ) | ( ~n6098 & n14603 ) ;
  assign n29986 = n23757 ^ n11572 ^ n10432 ;
  assign n29987 = n29985 & n29986 ;
  assign n29991 = n29990 ^ n29987 ^ n11505 ;
  assign n29992 = n3087 & n5497 ;
  assign n29993 = n29992 ^ n1869 ^ 1'b0 ;
  assign n29994 = ~n2895 & n29993 ;
  assign n29995 = n17083 & n29994 ;
  assign n29996 = n1780 & ~n29995 ;
  assign n29997 = n29991 & n29996 ;
  assign n30005 = n19240 ^ n18857 ^ n4063 ;
  assign n29998 = ( n620 & n2016 ) | ( n620 & ~n15063 ) | ( n2016 & ~n15063 ) ;
  assign n29999 = n23137 & ~n29998 ;
  assign n30000 = n2518 ^ x175 ^ 1'b0 ;
  assign n30001 = n29999 | n30000 ;
  assign n30002 = n5868 | n17968 ;
  assign n30003 = n30001 & ~n30002 ;
  assign n30004 = n7800 & ~n30003 ;
  assign n30006 = n30005 ^ n30004 ^ 1'b0 ;
  assign n30007 = n18822 ^ n16313 ^ 1'b0 ;
  assign n30008 = n17892 ^ n5484 ^ 1'b0 ;
  assign n30009 = n23037 ^ n16757 ^ n6368 ;
  assign n30010 = n10523 & ~n30009 ;
  assign n30011 = n28944 ^ n25796 ^ 1'b0 ;
  assign n30012 = n4441 | n14704 ;
  assign n30013 = ~n5860 & n29661 ;
  assign n30014 = n20699 & n30013 ;
  assign n30015 = ~n30012 & n30014 ;
  assign n30016 = n21655 ^ n1476 ^ 1'b0 ;
  assign n30017 = n9705 & ~n30016 ;
  assign n30018 = ~n13701 & n30017 ;
  assign n30019 = n9097 ^ n3526 ^ n3408 ;
  assign n30020 = n802 & ~n8833 ;
  assign n30021 = n21000 ^ n18683 ^ 1'b0 ;
  assign n30022 = ( n30019 & n30020 ) | ( n30019 & n30021 ) | ( n30020 & n30021 ) ;
  assign n30023 = n11279 & n13313 ;
  assign n30024 = n30023 ^ n25309 ^ n1429 ;
  assign n30025 = n23434 ^ n11910 ^ 1'b0 ;
  assign n30026 = n621 & ~n8287 ;
  assign n30027 = n30026 ^ n25783 ^ 1'b0 ;
  assign n30028 = ~n1298 & n30027 ;
  assign n30029 = n2348 | n7841 ;
  assign n30030 = n6597 | n28178 ;
  assign n30031 = n28178 & ~n30030 ;
  assign n30032 = n6896 & ~n30031 ;
  assign n30033 = n30031 & n30032 ;
  assign n30034 = n20216 & ~n30033 ;
  assign n30035 = n30034 ^ n1941 ^ 1'b0 ;
  assign n30036 = ~n10196 & n14531 ;
  assign n30037 = n30036 ^ n3341 ^ 1'b0 ;
  assign n30038 = n9118 | n13326 ;
  assign n30039 = n11728 | n30038 ;
  assign n30040 = ( n26675 & n26712 ) | ( n26675 & ~n30039 ) | ( n26712 & ~n30039 ) ;
  assign n30041 = n26973 ^ n19068 ^ n1301 ;
  assign n30042 = ( ~n30037 & n30040 ) | ( ~n30037 & n30041 ) | ( n30040 & n30041 ) ;
  assign n30043 = n1536 | n5736 ;
  assign n30044 = n2085 | n30043 ;
  assign n30045 = ~n7412 & n30044 ;
  assign n30046 = n30045 ^ n7195 ^ n6626 ;
  assign n30047 = n16706 ^ n14321 ^ n537 ;
  assign n30048 = n3292 | n10327 ;
  assign n30049 = n5718 & ~n19036 ;
  assign n30050 = ~n5961 & n30049 ;
  assign n30051 = n27166 ^ n15721 ^ n13048 ;
  assign n30052 = n30051 ^ n21767 ^ n5173 ;
  assign n30053 = n6675 & ~n12981 ;
  assign n30054 = ( ~n7468 & n18359 ) | ( ~n7468 & n30053 ) | ( n18359 & n30053 ) ;
  assign n30057 = n13925 | n17841 ;
  assign n30058 = n7376 & ~n30057 ;
  assign n30055 = n12926 ^ n11105 ^ n5298 ;
  assign n30056 = ~n14056 & n30055 ;
  assign n30059 = n30058 ^ n30056 ^ n19552 ;
  assign n30060 = n15001 | n17094 ;
  assign n30061 = n23635 ^ n19677 ^ n16710 ;
  assign n30062 = n30061 ^ n14150 ^ n2219 ;
  assign n30063 = n30062 ^ n3525 ^ 1'b0 ;
  assign n30064 = n18456 ^ n3804 ^ 1'b0 ;
  assign n30065 = n12887 & n20605 ;
  assign n30066 = n22917 & n30065 ;
  assign n30067 = n30066 ^ n7655 ^ 1'b0 ;
  assign n30068 = ~n7526 & n30067 ;
  assign n30069 = ( n20643 & n30064 ) | ( n20643 & n30068 ) | ( n30064 & n30068 ) ;
  assign n30070 = n14984 ^ n5664 ^ n1538 ;
  assign n30071 = n17773 ^ n1158 ^ 1'b0 ;
  assign n30072 = n4985 & ~n24651 ;
  assign n30073 = ~n30071 & n30072 ;
  assign n30074 = n3207 & ~n7934 ;
  assign n30075 = n21656 ^ n13721 ^ n12818 ;
  assign n30076 = n30075 ^ n14920 ^ 1'b0 ;
  assign n30077 = n15147 | n19137 ;
  assign n30078 = n19704 ^ n18753 ^ 1'b0 ;
  assign n30079 = n3936 ^ n835 ^ x141 ;
  assign n30080 = n28926 ^ n2317 ^ 1'b0 ;
  assign n30081 = n30079 | n30080 ;
  assign n30082 = ( n30077 & n30078 ) | ( n30077 & n30081 ) | ( n30078 & n30081 ) ;
  assign n30083 = n12923 | n18370 ;
  assign n30084 = n11839 | n30083 ;
  assign n30085 = n22382 ^ n5021 ^ 1'b0 ;
  assign n30086 = n1328 & n29017 ;
  assign n30087 = n30086 ^ n8431 ^ 1'b0 ;
  assign n30088 = n9314 & n15022 ;
  assign n30089 = n30088 ^ n10940 ^ 1'b0 ;
  assign n30090 = n7806 ^ n2551 ^ 1'b0 ;
  assign n30091 = n28939 ^ n10687 ^ 1'b0 ;
  assign n30092 = ~n5781 & n30091 ;
  assign n30093 = n4243 & n10926 ;
  assign n30094 = ~n30092 & n30093 ;
  assign n30095 = ( n29859 & n30090 ) | ( n29859 & n30094 ) | ( n30090 & n30094 ) ;
  assign n30096 = n24350 ^ n21949 ^ 1'b0 ;
  assign n30097 = n630 | n19164 ;
  assign n30098 = n20369 | n30097 ;
  assign n30099 = ( n1204 & n5091 ) | ( n1204 & ~n11054 ) | ( n5091 & ~n11054 ) ;
  assign n30100 = ~n2356 & n21030 ;
  assign n30106 = ( n11842 & n23065 ) | ( n11842 & n26073 ) | ( n23065 & n26073 ) ;
  assign n30104 = n902 & n16783 ;
  assign n30101 = n442 & n22380 ;
  assign n30102 = n30101 ^ n14835 ^ 1'b0 ;
  assign n30103 = n4493 & n30102 ;
  assign n30105 = n30104 ^ n30103 ^ n945 ;
  assign n30107 = n30106 ^ n30105 ^ 1'b0 ;
  assign n30108 = n13862 | n29231 ;
  assign n30109 = n25045 & ~n30108 ;
  assign n30110 = n2137 | n30109 ;
  assign n30111 = n4995 | n23293 ;
  assign n30112 = n19456 | n30111 ;
  assign n30113 = n5203 & n27473 ;
  assign n30114 = ~n30112 & n30113 ;
  assign n30115 = n7644 ^ n460 ^ 1'b0 ;
  assign n30116 = n30115 ^ n8681 ^ 1'b0 ;
  assign n30117 = n4598 & n30116 ;
  assign n30118 = n30117 ^ n5264 ^ 1'b0 ;
  assign n30119 = ( n371 & ~n2465 ) | ( n371 & n2990 ) | ( ~n2465 & n2990 ) ;
  assign n30120 = ~n8361 & n12118 ;
  assign n30121 = n5039 ^ n3430 ^ n2811 ;
  assign n30122 = ( n2994 & ~n12362 ) | ( n2994 & n30121 ) | ( ~n12362 & n30121 ) ;
  assign n30123 = ~n1701 & n30122 ;
  assign n30124 = ~n30120 & n30123 ;
  assign n30125 = n30119 & ~n30124 ;
  assign n30126 = ~n30118 & n30125 ;
  assign n30127 = n7338 & n9364 ;
  assign n30128 = ( n4004 & n8116 ) | ( n4004 & ~n30127 ) | ( n8116 & ~n30127 ) ;
  assign n30130 = n5011 ^ n2758 ^ n1750 ;
  assign n30129 = n9842 ^ n6903 ^ n845 ;
  assign n30131 = n30130 ^ n30129 ^ 1'b0 ;
  assign n30132 = ~n697 & n30131 ;
  assign n30133 = n30132 ^ n9434 ^ 1'b0 ;
  assign n30134 = n6619 ^ n733 ^ 1'b0 ;
  assign n30135 = n30134 ^ n5245 ^ 1'b0 ;
  assign n30136 = ~n30133 & n30135 ;
  assign n30137 = n4141 & ~n25404 ;
  assign n30138 = n5095 & n30137 ;
  assign n30139 = n30138 ^ n29540 ^ 1'b0 ;
  assign n30140 = n30139 ^ n23936 ^ 1'b0 ;
  assign n30141 = n25605 ^ n12346 ^ 1'b0 ;
  assign n30142 = ( n1291 & ~n2915 ) | ( n1291 & n21560 ) | ( ~n2915 & n21560 ) ;
  assign n30143 = n9423 ^ n6255 ^ 1'b0 ;
  assign n30144 = n9635 | n30143 ;
  assign n30145 = n8306 & n30144 ;
  assign n30146 = n30145 ^ n17412 ^ 1'b0 ;
  assign n30147 = n30146 ^ n12407 ^ 1'b0 ;
  assign n30148 = n24420 ^ n4760 ^ 1'b0 ;
  assign n30149 = n25450 ^ n19444 ^ n17589 ;
  assign n30150 = n5254 | n12925 ;
  assign n30151 = n8960 | n30150 ;
  assign n30152 = n15184 ^ n13218 ^ n5548 ;
  assign n30153 = n30152 ^ n26944 ^ 1'b0 ;
  assign n30154 = ( x166 & x251 ) | ( x166 & ~n4874 ) | ( x251 & ~n4874 ) ;
  assign n30155 = n3054 & n4141 ;
  assign n30156 = n30154 & n30155 ;
  assign n30157 = n30156 ^ n9539 ^ n8025 ;
  assign n30158 = n18723 ^ n11731 ^ 1'b0 ;
  assign n30159 = n27169 ^ n943 ^ 1'b0 ;
  assign n30160 = ~n30158 & n30159 ;
  assign n30161 = n30160 ^ n4842 ^ 1'b0 ;
  assign n30162 = n30161 ^ n8948 ^ 1'b0 ;
  assign n30163 = n30157 & n30162 ;
  assign n30164 = n19178 ^ n3750 ^ 1'b0 ;
  assign n30165 = ( n3030 & ~n17381 ) | ( n3030 & n18864 ) | ( ~n17381 & n18864 ) ;
  assign n30166 = n24630 & ~n30165 ;
  assign n30167 = n4927 | n10509 ;
  assign n30168 = n24887 ^ n9631 ^ 1'b0 ;
  assign n30169 = ( ~n7193 & n7650 ) | ( ~n7193 & n15500 ) | ( n7650 & n15500 ) ;
  assign n30170 = n14943 | n30169 ;
  assign n30171 = n30170 ^ n23131 ^ 1'b0 ;
  assign n30172 = ~n3640 & n13186 ;
  assign n30173 = n30172 ^ n2822 ^ 1'b0 ;
  assign n30174 = n2243 & ~n20317 ;
  assign n30175 = n15171 ^ n4977 ^ n3660 ;
  assign n30176 = n28112 ^ n12812 ^ 1'b0 ;
  assign n30177 = n25726 ^ n7733 ^ n7540 ;
  assign n30178 = n23587 ^ n14044 ^ 1'b0 ;
  assign n30179 = n23616 & n30178 ;
  assign n30180 = n3810 | n18306 ;
  assign n30183 = n8180 ^ n259 ^ 1'b0 ;
  assign n30184 = n2539 & n30183 ;
  assign n30181 = n12401 ^ n4453 ^ n2995 ;
  assign n30182 = ( n3286 & n13881 ) | ( n3286 & n30181 ) | ( n13881 & n30181 ) ;
  assign n30185 = n30184 ^ n30182 ^ 1'b0 ;
  assign n30186 = n30185 ^ n6110 ^ 1'b0 ;
  assign n30187 = ~n30180 & n30186 ;
  assign n30188 = n9483 & n10707 ;
  assign n30189 = n15621 & n30188 ;
  assign n30190 = ~n5814 & n8230 ;
  assign n30191 = n30190 ^ n859 ^ 1'b0 ;
  assign n30192 = ~n6815 & n13667 ;
  assign n30193 = ~n6228 & n30192 ;
  assign n30194 = n13226 ^ n9997 ^ 1'b0 ;
  assign n30195 = ~n1463 & n30194 ;
  assign n30196 = n30195 ^ n4016 ^ 1'b0 ;
  assign n30197 = n30196 ^ n5290 ^ 1'b0 ;
  assign n30198 = n29796 & n30197 ;
  assign n30200 = n22252 ^ n6632 ^ n4341 ;
  assign n30201 = n30200 ^ n13865 ^ n9948 ;
  assign n30202 = n30201 ^ n11992 ^ 1'b0 ;
  assign n30199 = ~n6904 & n19370 ;
  assign n30203 = n30202 ^ n30199 ^ 1'b0 ;
  assign n30205 = n16081 & n20943 ;
  assign n30206 = n2435 & n30205 ;
  assign n30204 = n4980 & ~n17332 ;
  assign n30207 = n30206 ^ n30204 ^ 1'b0 ;
  assign n30208 = n23965 ^ n18043 ^ n6218 ;
  assign n30209 = x165 & n30208 ;
  assign n30210 = n9519 ^ n2580 ^ 1'b0 ;
  assign n30214 = ( ~n10112 & n10242 ) | ( ~n10112 & n13189 ) | ( n10242 & n13189 ) ;
  assign n30211 = n9337 ^ n9177 ^ 1'b0 ;
  assign n30212 = ~n22152 & n30211 ;
  assign n30213 = n30212 ^ n29007 ^ n27935 ;
  assign n30215 = n30214 ^ n30213 ^ n5134 ;
  assign n30219 = n7788 & n10034 ;
  assign n30220 = n18512 ^ n1364 ^ 1'b0 ;
  assign n30221 = ( n27727 & n30219 ) | ( n27727 & n30220 ) | ( n30219 & n30220 ) ;
  assign n30216 = n11758 ^ n1430 ^ 1'b0 ;
  assign n30217 = n30216 ^ n26856 ^ n12515 ;
  assign n30218 = n30217 ^ n19181 ^ 1'b0 ;
  assign n30222 = n30221 ^ n30218 ^ n16066 ;
  assign n30223 = ~n19036 & n30222 ;
  assign n30224 = n17489 & n30223 ;
  assign n30225 = n7608 | n22636 ;
  assign n30226 = n12959 ^ n7957 ^ 1'b0 ;
  assign n30227 = ~n6156 & n30226 ;
  assign n30228 = ~n1653 & n4525 ;
  assign n30229 = n8233 & n10287 ;
  assign n30230 = ~n4367 & n30229 ;
  assign n30231 = ~n26704 & n30230 ;
  assign n30232 = ~n1908 & n30231 ;
  assign n30233 = n30228 & n30232 ;
  assign n30234 = n1050 & n15133 ;
  assign n30235 = n30234 ^ n6851 ^ 1'b0 ;
  assign n30236 = ~n27172 & n28189 ;
  assign n30237 = ~n8331 & n30236 ;
  assign n30238 = n19404 ^ n5239 ^ 1'b0 ;
  assign n30239 = n29444 | n30238 ;
  assign n30240 = n22610 ^ n4423 ^ 1'b0 ;
  assign n30241 = n20977 & ~n30240 ;
  assign n30242 = n5972 ^ n612 ^ 1'b0 ;
  assign n30243 = n25942 ^ n19636 ^ n11750 ;
  assign n30244 = n30243 ^ n16032 ^ n2012 ;
  assign n30245 = ( ~n702 & n11762 ) | ( ~n702 & n21545 ) | ( n11762 & n21545 ) ;
  assign n30246 = n7578 & n30245 ;
  assign n30247 = ~n19720 & n30246 ;
  assign n30248 = n18066 & ~n30247 ;
  assign n30249 = n30248 ^ n23046 ^ n1655 ;
  assign n30250 = ( ~n15971 & n16647 ) | ( ~n15971 & n23351 ) | ( n16647 & n23351 ) ;
  assign n30251 = n9327 ^ n3910 ^ 1'b0 ;
  assign n30252 = n9872 & ~n19317 ;
  assign n30253 = n1216 | n13446 ;
  assign n30254 = n30252 | n30253 ;
  assign n30255 = ( n30250 & n30251 ) | ( n30250 & n30254 ) | ( n30251 & n30254 ) ;
  assign n30256 = n30255 ^ n15941 ^ n3858 ;
  assign n30257 = n18920 ^ n15991 ^ n3184 ;
  assign n30258 = ~n4609 & n23312 ;
  assign n30259 = n10272 | n25647 ;
  assign n30260 = n17716 & n30259 ;
  assign n30261 = n30260 ^ n4227 ^ 1'b0 ;
  assign n30262 = n1630 & n30261 ;
  assign n30263 = n1454 & n7739 ;
  assign n30264 = n21421 ^ n4578 ^ 1'b0 ;
  assign n30265 = ~n1869 & n30264 ;
  assign n30266 = n30263 | n30265 ;
  assign n30267 = n22661 ^ n10056 ^ x128 ;
  assign n30268 = n4068 | n28423 ;
  assign n30269 = n30268 ^ n4849 ^ 1'b0 ;
  assign n30270 = ~n3158 & n30269 ;
  assign n30271 = n30270 ^ n11493 ^ 1'b0 ;
  assign n30272 = n22128 & ~n30271 ;
  assign n30273 = ~n2638 & n30272 ;
  assign n30274 = n14969 ^ n9159 ^ n1010 ;
  assign n30275 = n30274 ^ n10194 ^ 1'b0 ;
  assign n30276 = n14366 & ~n30275 ;
  assign n30277 = n18997 ^ n16383 ^ 1'b0 ;
  assign n30278 = n30276 & n30277 ;
  assign n30279 = n675 | n8976 ;
  assign n30280 = n22499 ^ n6934 ^ 1'b0 ;
  assign n30281 = n20965 & ~n30280 ;
  assign n30282 = n30279 & n30281 ;
  assign n30283 = n13478 & n30282 ;
  assign n30286 = n9889 ^ n2585 ^ 1'b0 ;
  assign n30287 = n22713 & n30286 ;
  assign n30288 = n9223 | n15877 ;
  assign n30289 = n30287 | n30288 ;
  assign n30284 = n3624 & ~n13127 ;
  assign n30285 = n20543 & n30284 ;
  assign n30290 = n30289 ^ n30285 ^ 1'b0 ;
  assign n30295 = n8300 & ~n11160 ;
  assign n30291 = n3034 & ~n5254 ;
  assign n30292 = n2892 & n30291 ;
  assign n30293 = n21004 ^ n642 ^ 1'b0 ;
  assign n30294 = ( ~n8948 & n30292 ) | ( ~n8948 & n30293 ) | ( n30292 & n30293 ) ;
  assign n30296 = n30295 ^ n30294 ^ n5376 ;
  assign n30297 = n740 | n30296 ;
  assign n30298 = n1766 & n4306 ;
  assign n30299 = n30298 ^ n13793 ^ 1'b0 ;
  assign n30300 = n30299 ^ n1583 ^ 1'b0 ;
  assign n30301 = n22824 | n30300 ;
  assign n30302 = ( n335 & n7582 ) | ( n335 & n15278 ) | ( n7582 & n15278 ) ;
  assign n30303 = n4683 & n24685 ;
  assign n30304 = n8185 & ~n22310 ;
  assign n30305 = n18512 | n30304 ;
  assign n30306 = n15493 | n30305 ;
  assign n30307 = n27573 ^ n2136 ^ 1'b0 ;
  assign n30308 = n10614 & ~n10699 ;
  assign n30309 = n7850 & ~n11035 ;
  assign n30310 = n18960 ^ n11283 ^ n5207 ;
  assign n30311 = n8993 ^ n5144 ^ 1'b0 ;
  assign n30312 = n30310 | n30311 ;
  assign n30313 = n15701 ^ n4533 ^ 1'b0 ;
  assign n30314 = n16215 ^ n7006 ^ 1'b0 ;
  assign n30315 = n17568 & n24667 ;
  assign n30316 = n30315 ^ n25461 ^ n25377 ;
  assign n30317 = n8628 | n15904 ;
  assign n30318 = ( n8765 & n29176 ) | ( n8765 & n30317 ) | ( n29176 & n30317 ) ;
  assign n30319 = n9451 | n20747 ;
  assign n30320 = n10613 ^ n1341 ^ 1'b0 ;
  assign n30321 = n8496 & ~n30320 ;
  assign n30322 = n7734 & n13150 ;
  assign n30323 = ( n519 & n3722 ) | ( n519 & ~n30322 ) | ( n3722 & ~n30322 ) ;
  assign n30324 = n30323 ^ n24638 ^ n2194 ;
  assign n30325 = n7167 ^ n3705 ^ n2796 ;
  assign n30326 = n30325 ^ n17957 ^ n5793 ;
  assign n30327 = n12917 ^ x126 ^ 1'b0 ;
  assign n30328 = n21669 ^ n7302 ^ 1'b0 ;
  assign n30329 = n30327 & ~n30328 ;
  assign n30330 = n30326 | n30329 ;
  assign n30331 = ( ~n18006 & n24619 ) | ( ~n18006 & n30330 ) | ( n24619 & n30330 ) ;
  assign n30334 = n5877 & n17731 ;
  assign n30335 = n30334 ^ n23676 ^ 1'b0 ;
  assign n30336 = n30335 ^ n17789 ^ n2771 ;
  assign n30332 = n17340 ^ n12259 ^ 1'b0 ;
  assign n30333 = ( n729 & ~n4493 ) | ( n729 & n30332 ) | ( ~n4493 & n30332 ) ;
  assign n30337 = n30336 ^ n30333 ^ 1'b0 ;
  assign n30339 = n15107 ^ n5610 ^ x41 ;
  assign n30340 = ~n7602 & n30339 ;
  assign n30341 = n30340 ^ n9268 ^ 1'b0 ;
  assign n30338 = n835 & ~n27894 ;
  assign n30342 = n30341 ^ n30338 ^ 1'b0 ;
  assign n30343 = n24032 ^ n17161 ^ 1'b0 ;
  assign n30344 = n4083 & ~n30343 ;
  assign n30345 = n19421 ^ n10339 ^ 1'b0 ;
  assign n30346 = n7066 & n7669 ;
  assign n30347 = n13061 | n16063 ;
  assign n30348 = n30347 ^ n23559 ^ 1'b0 ;
  assign n30349 = n378 | n24808 ;
  assign n30350 = n10001 | n30349 ;
  assign n30351 = n30350 ^ n16096 ^ 1'b0 ;
  assign n30352 = ~n30348 & n30351 ;
  assign n30353 = n1489 & ~n14835 ;
  assign n30354 = n10754 ^ n4780 ^ 1'b0 ;
  assign n30355 = ( ~x198 & n2849 ) | ( ~x198 & n30354 ) | ( n2849 & n30354 ) ;
  assign n30356 = ( n27712 & ~n30353 ) | ( n27712 & n30355 ) | ( ~n30353 & n30355 ) ;
  assign n30357 = n30356 ^ n20739 ^ n947 ;
  assign n30358 = n19955 & ~n30357 ;
  assign n30359 = ~n12346 & n30358 ;
  assign n30360 = ~n857 & n28190 ;
  assign n30361 = n27879 ^ n20002 ^ n17405 ;
  assign n30362 = n30361 ^ n20438 ^ n4959 ;
  assign n30363 = n28042 ^ n27942 ^ n19159 ;
  assign n30365 = ( n6510 & n8526 ) | ( n6510 & n9789 ) | ( n8526 & n9789 ) ;
  assign n30366 = ( n1998 & n3307 ) | ( n1998 & ~n30365 ) | ( n3307 & ~n30365 ) ;
  assign n30367 = n1262 & n4752 ;
  assign n30368 = n14758 & n30367 ;
  assign n30369 = n30366 & n30368 ;
  assign n30364 = n2886 & n15098 ;
  assign n30370 = n30369 ^ n30364 ^ 1'b0 ;
  assign n30371 = ~n7980 & n23673 ;
  assign n30372 = n16779 & n30371 ;
  assign n30373 = n9025 & ~n24543 ;
  assign n30374 = n30373 ^ n19032 ^ n8533 ;
  assign n30375 = n30374 ^ n2270 ^ 1'b0 ;
  assign n30376 = n8335 | n10968 ;
  assign n30377 = n30376 ^ n25549 ^ n3237 ;
  assign n30378 = n25518 ^ n18683 ^ n5827 ;
  assign n30379 = ~n19181 & n30378 ;
  assign n30380 = n30379 ^ n6962 ^ 1'b0 ;
  assign n30381 = n5381 | n11796 ;
  assign n30382 = n30381 ^ x244 ^ 1'b0 ;
  assign n30383 = ~n21003 & n30382 ;
  assign n30384 = n18726 ^ n16270 ^ n8252 ;
  assign n30385 = ( ~n2253 & n9576 ) | ( ~n2253 & n30384 ) | ( n9576 & n30384 ) ;
  assign n30386 = ( n5283 & n19146 ) | ( n5283 & ~n30385 ) | ( n19146 & ~n30385 ) ;
  assign n30387 = n18808 ^ n7909 ^ 1'b0 ;
  assign n30388 = n29589 & ~n30387 ;
  assign n30389 = ~n21198 & n27666 ;
  assign n30390 = ~n18856 & n30389 ;
  assign n30391 = n30390 ^ n28545 ^ 1'b0 ;
  assign n30392 = n10261 | n30391 ;
  assign n30393 = n17696 ^ n5768 ^ 1'b0 ;
  assign n30394 = n11152 & ~n30393 ;
  assign n30395 = n12234 ^ n11837 ^ 1'b0 ;
  assign n30396 = ( ~n2453 & n5528 ) | ( ~n2453 & n14575 ) | ( n5528 & n14575 ) ;
  assign n30397 = ( n6723 & ~n18142 ) | ( n6723 & n30396 ) | ( ~n18142 & n30396 ) ;
  assign n30398 = ( x149 & n3775 ) | ( x149 & n5554 ) | ( n3775 & n5554 ) ;
  assign n30399 = n945 & n30398 ;
  assign n30400 = ~n30397 & n30399 ;
  assign n30401 = n10545 & ~n30400 ;
  assign n30402 = n30401 ^ n30124 ^ 1'b0 ;
  assign n30405 = n11934 ^ n8907 ^ 1'b0 ;
  assign n30404 = n18394 ^ n5042 ^ 1'b0 ;
  assign n30406 = n30405 ^ n30404 ^ n3016 ;
  assign n30407 = n8114 ^ n3869 ^ 1'b0 ;
  assign n30408 = n30406 & n30407 ;
  assign n30403 = n13680 | n15313 ;
  assign n30409 = n30408 ^ n30403 ^ 1'b0 ;
  assign n30410 = n2950 | n23374 ;
  assign n30411 = n27115 ^ n24605 ^ 1'b0 ;
  assign n30414 = n4132 & ~n20159 ;
  assign n30415 = ~n3831 & n30414 ;
  assign n30412 = n5862 ^ n4460 ^ 1'b0 ;
  assign n30413 = ( n5166 & n9587 ) | ( n5166 & n30412 ) | ( n9587 & n30412 ) ;
  assign n30416 = n30415 ^ n30413 ^ 1'b0 ;
  assign n30417 = n2106 & n2362 ;
  assign n30418 = ~n5800 & n30417 ;
  assign n30422 = ( ~n2616 & n3961 ) | ( ~n2616 & n15327 ) | ( n3961 & n15327 ) ;
  assign n30423 = n30422 ^ n19041 ^ 1'b0 ;
  assign n30419 = n12524 ^ n5879 ^ 1'b0 ;
  assign n30420 = n30419 ^ n18466 ^ n13578 ;
  assign n30421 = n30420 ^ n19689 ^ 1'b0 ;
  assign n30424 = n30423 ^ n30421 ^ 1'b0 ;
  assign n30425 = n6152 ^ n938 ^ 1'b0 ;
  assign n30426 = n29294 & n30425 ;
  assign n30427 = n1284 & ~n2469 ;
  assign n30428 = n24168 | n30427 ;
  assign n30429 = n20521 ^ n8642 ^ 1'b0 ;
  assign n30430 = ~n5289 & n30429 ;
  assign n30431 = n1312 & ~n1734 ;
  assign n30432 = n13768 & ~n30431 ;
  assign n30433 = n11035 ^ n1339 ^ 1'b0 ;
  assign n30434 = n14017 ^ x211 ^ 1'b0 ;
  assign n30435 = n30434 ^ n15156 ^ 1'b0 ;
  assign n30436 = n2301 & n25220 ;
  assign n30437 = n30436 ^ n12508 ^ 1'b0 ;
  assign n30438 = n5842 ^ n1209 ^ 1'b0 ;
  assign n30439 = n23239 ^ n7788 ^ 1'b0 ;
  assign n30440 = n13356 & ~n30439 ;
  assign n30441 = n30440 ^ n18238 ^ n4540 ;
  assign n30442 = n11291 ^ n4611 ^ 1'b0 ;
  assign n30443 = n3608 & n30442 ;
  assign n30444 = ~n490 & n30443 ;
  assign n30445 = n1025 | n27064 ;
  assign n30451 = n4306 & n25912 ;
  assign n30452 = n12671 & n30451 ;
  assign n30447 = n9581 & n23256 ;
  assign n30448 = n14358 & n30447 ;
  assign n30449 = n30448 ^ n8810 ^ 1'b0 ;
  assign n30450 = n11377 | n30449 ;
  assign n30446 = n21549 ^ n608 ^ 1'b0 ;
  assign n30453 = n30452 ^ n30450 ^ n30446 ;
  assign n30454 = n8757 | n16201 ;
  assign n30455 = ( n11522 & n30119 ) | ( n11522 & n30454 ) | ( n30119 & n30454 ) ;
  assign n30456 = n22906 & ~n30455 ;
  assign n30457 = ~n6569 & n14049 ;
  assign n30458 = n30457 ^ n9299 ^ 1'b0 ;
  assign n30459 = n30458 ^ n10436 ^ n6174 ;
  assign n30460 = ~n9788 & n30459 ;
  assign n30461 = n2005 ^ x175 ^ 1'b0 ;
  assign n30462 = n14246 & n30461 ;
  assign n30463 = n4043 & n15382 ;
  assign n30464 = n20233 ^ n7386 ^ n5042 ;
  assign n30465 = n30464 ^ n29807 ^ 1'b0 ;
  assign n30466 = n30465 ^ n10055 ^ n5483 ;
  assign n30467 = ~n1689 & n27225 ;
  assign n30468 = n22009 ^ n10680 ^ 1'b0 ;
  assign n30469 = n8702 & n30468 ;
  assign n30470 = n30467 | n30469 ;
  assign n30471 = ( ~n1653 & n5361 ) | ( ~n1653 & n17583 ) | ( n5361 & n17583 ) ;
  assign n30472 = n2119 & ~n30471 ;
  assign n30475 = n10713 ^ n3191 ^ 1'b0 ;
  assign n30476 = n30040 | n30475 ;
  assign n30473 = x205 | n3318 ;
  assign n30474 = n30473 ^ n2054 ^ n1506 ;
  assign n30477 = n30476 ^ n30474 ^ n12396 ;
  assign n30478 = n9337 ^ n7525 ^ 1'b0 ;
  assign n30479 = n7900 ^ n4662 ^ 1'b0 ;
  assign n30480 = n17343 & ~n23905 ;
  assign n30481 = ~n30479 & n30480 ;
  assign n30482 = n14801 ^ n4618 ^ 1'b0 ;
  assign n30483 = n22759 & n30482 ;
  assign n30484 = ( ~n5163 & n13341 ) | ( ~n5163 & n29443 ) | ( n13341 & n29443 ) ;
  assign n30485 = n12191 & ~n21862 ;
  assign n30486 = n30485 ^ n16327 ^ 1'b0 ;
  assign n30487 = n30486 ^ n2061 ^ 1'b0 ;
  assign n30488 = n19424 ^ n12792 ^ 1'b0 ;
  assign n30489 = ~n19873 & n30488 ;
  assign n30490 = ( x97 & n15654 ) | ( x97 & ~n30489 ) | ( n15654 & ~n30489 ) ;
  assign n30491 = n12423 & ~n28397 ;
  assign n30492 = ( n4130 & ~n14257 ) | ( n4130 & n21213 ) | ( ~n14257 & n21213 ) ;
  assign n30493 = n2937 | n30492 ;
  assign n30494 = n1374 & ~n30493 ;
  assign n30495 = n30494 ^ n16783 ^ 1'b0 ;
  assign n30496 = n16132 & ~n30495 ;
  assign n30497 = n9660 & ~n10200 ;
  assign n30498 = n30497 ^ n29958 ^ 1'b0 ;
  assign n30499 = n15876 | n30498 ;
  assign n30500 = n1064 | n30499 ;
  assign n30501 = n8684 & ~n24213 ;
  assign n30502 = n16232 | n30501 ;
  assign n30503 = n30502 ^ n6062 ^ 1'b0 ;
  assign n30504 = ~n1309 & n2769 ;
  assign n30505 = n30504 ^ n8253 ^ 1'b0 ;
  assign n30506 = n5789 ^ n574 ^ 1'b0 ;
  assign n30507 = ( n4039 & n8684 ) | ( n4039 & n30506 ) | ( n8684 & n30506 ) ;
  assign n30508 = n24463 ^ n20995 ^ n14316 ;
  assign n30509 = n5726 & ~n30508 ;
  assign n30510 = n5170 & n30509 ;
  assign n30511 = ~n19624 & n21371 ;
  assign n30512 = n2821 & n30511 ;
  assign n30513 = n13652 ^ n12212 ^ n7294 ;
  assign n30514 = n17045 ^ n4579 ^ 1'b0 ;
  assign n30515 = ( ~n615 & n4220 ) | ( ~n615 & n11384 ) | ( n4220 & n11384 ) ;
  assign n30516 = ( ~n6534 & n7618 ) | ( ~n6534 & n30515 ) | ( n7618 & n30515 ) ;
  assign n30517 = n3995 & ~n30516 ;
  assign n30518 = n10449 ^ n5821 ^ 1'b0 ;
  assign n30519 = ~n7132 & n30518 ;
  assign n30520 = n3855 & n9607 ;
  assign n30521 = n30519 & n30520 ;
  assign n30522 = n6252 & n8461 ;
  assign n30523 = n3296 & n30522 ;
  assign n30524 = n30523 ^ n29982 ^ 1'b0 ;
  assign n30525 = n3198 | n14050 ;
  assign n30526 = n6730 & ~n30525 ;
  assign n30527 = n5634 | n12246 ;
  assign n30528 = n30527 ^ n10609 ^ 1'b0 ;
  assign n30529 = n30528 ^ n22930 ^ n2169 ;
  assign n30530 = n2500 & ~n12341 ;
  assign n30531 = ( ~n1183 & n7990 ) | ( ~n1183 & n11320 ) | ( n7990 & n11320 ) ;
  assign n30532 = n16689 & n30531 ;
  assign n30533 = x158 & ~n13340 ;
  assign n30534 = n30533 ^ n4585 ^ 1'b0 ;
  assign n30535 = n2015 & ~n30534 ;
  assign n30536 = n30535 ^ n3820 ^ 1'b0 ;
  assign n30537 = n17146 ^ n3510 ^ 1'b0 ;
  assign n30538 = n14895 | n30537 ;
  assign n30539 = n22627 | n30538 ;
  assign n30540 = ~n2675 & n3768 ;
  assign n30541 = n30540 ^ n9103 ^ 1'b0 ;
  assign n30542 = ( ~n13378 & n30012 ) | ( ~n13378 & n30541 ) | ( n30012 & n30541 ) ;
  assign n30543 = n26437 ^ n3327 ^ 1'b0 ;
  assign n30544 = ( n6280 & n7758 ) | ( n6280 & ~n13515 ) | ( n7758 & ~n13515 ) ;
  assign n30545 = n7195 | n10134 ;
  assign n30546 = n30545 ^ n5417 ^ 1'b0 ;
  assign n30547 = n30546 ^ n7599 ^ 1'b0 ;
  assign n30548 = n30547 ^ n14887 ^ n13497 ;
  assign n30549 = n12412 & n30548 ;
  assign n30550 = n30549 ^ n21859 ^ 1'b0 ;
  assign n30551 = n7298 | n7691 ;
  assign n30552 = n30551 ^ n3100 ^ 1'b0 ;
  assign n30553 = n30552 ^ n7284 ^ n5516 ;
  assign n30554 = n841 & n30553 ;
  assign n30555 = n30554 ^ n5920 ^ 1'b0 ;
  assign n30556 = ( n1669 & n15272 ) | ( n1669 & n17427 ) | ( n15272 & n17427 ) ;
  assign n30557 = n30556 ^ n23771 ^ 1'b0 ;
  assign n30558 = n12209 & ~n30557 ;
  assign n30559 = n17843 ^ n11804 ^ 1'b0 ;
  assign n30560 = n7184 & n24787 ;
  assign n30561 = ~n30559 & n30560 ;
  assign n30562 = n25461 ^ n4838 ^ 1'b0 ;
  assign n30563 = ( n28643 & n30561 ) | ( n28643 & ~n30562 ) | ( n30561 & ~n30562 ) ;
  assign n30564 = ( n1084 & n2582 ) | ( n1084 & ~n5305 ) | ( n2582 & ~n5305 ) ;
  assign n30565 = n21377 | n25577 ;
  assign n30566 = n30564 | n30565 ;
  assign n30567 = x120 | n16120 ;
  assign n30568 = n6999 | n15965 ;
  assign n30569 = n30568 ^ n5573 ^ 1'b0 ;
  assign n30570 = n4904 & ~n15933 ;
  assign n30571 = ~n4334 & n30570 ;
  assign n30572 = n5500 & ~n12648 ;
  assign n30573 = n30572 ^ n5888 ^ n2702 ;
  assign n30574 = n30571 | n30573 ;
  assign n30575 = n14302 & ~n30574 ;
  assign n30576 = n30575 ^ n22184 ^ n15897 ;
  assign n30577 = n30576 ^ n11665 ^ 1'b0 ;
  assign n30578 = ~n9238 & n11135 ;
  assign n30579 = n30578 ^ n12371 ^ 1'b0 ;
  assign n30582 = ~n6251 & n12370 ;
  assign n30580 = n18882 | n23099 ;
  assign n30581 = n30580 ^ n13721 ^ 1'b0 ;
  assign n30583 = n30582 ^ n30581 ^ n23782 ;
  assign n30584 = ( n15727 & n16337 ) | ( n15727 & n29816 ) | ( n16337 & n29816 ) ;
  assign n30585 = n1848 & n5905 ;
  assign n30586 = n5539 | n10145 ;
  assign n30587 = n30586 ^ n11786 ^ 1'b0 ;
  assign n30588 = n2114 & ~n30587 ;
  assign n30589 = n30588 ^ n23765 ^ 1'b0 ;
  assign n30590 = n27105 ^ n4465 ^ 1'b0 ;
  assign n30591 = n16659 ^ n684 ^ 1'b0 ;
  assign n30592 = ~n15826 & n18602 ;
  assign n30593 = n17841 & ~n30592 ;
  assign n30594 = n5379 | n8631 ;
  assign n30595 = n30594 ^ n14515 ^ 1'b0 ;
  assign n30596 = n30595 ^ n21270 ^ n2615 ;
  assign n30597 = ( n1343 & ~n7145 ) | ( n1343 & n26509 ) | ( ~n7145 & n26509 ) ;
  assign n30599 = n9806 | n15604 ;
  assign n30600 = n8365 | n30599 ;
  assign n30601 = n19457 | n30600 ;
  assign n30598 = ~n12899 & n25287 ;
  assign n30602 = n30601 ^ n30598 ^ 1'b0 ;
  assign n30603 = n8387 | n23518 ;
  assign n30604 = n27273 | n30603 ;
  assign n30605 = n8024 | n23963 ;
  assign n30606 = n30605 ^ n410 ^ 1'b0 ;
  assign n30607 = n16860 & n21784 ;
  assign n30608 = n8983 ^ n854 ^ 1'b0 ;
  assign n30609 = n20531 & n30608 ;
  assign n30610 = n11409 ^ x209 ^ 1'b0 ;
  assign n30611 = x230 & n30610 ;
  assign n30612 = n30611 ^ n19690 ^ 1'b0 ;
  assign n30613 = n30609 & ~n30612 ;
  assign n30614 = n25781 ^ n6817 ^ 1'b0 ;
  assign n30615 = ( n11126 & n14993 ) | ( n11126 & ~n19113 ) | ( n14993 & ~n19113 ) ;
  assign n30616 = n30614 & n30615 ;
  assign n30617 = n30616 ^ n12206 ^ 1'b0 ;
  assign n30618 = n17133 ^ n4239 ^ 1'b0 ;
  assign n30619 = n21357 & n30618 ;
  assign n30620 = ~n9467 & n19655 ;
  assign n30621 = n8244 | n30620 ;
  assign n30622 = n19104 | n30621 ;
  assign n30623 = n16662 & ~n19435 ;
  assign n30624 = n1234 & n30623 ;
  assign n30625 = n30624 ^ n7210 ^ 1'b0 ;
  assign n30626 = n13952 ^ n10828 ^ n9331 ;
  assign n30627 = n24513 ^ n341 ^ x233 ;
  assign n30628 = n5102 & n13716 ;
  assign n30629 = ~n13322 & n30628 ;
  assign n30630 = n20142 ^ n7646 ^ 1'b0 ;
  assign n30631 = n30629 | n30630 ;
  assign n30632 = n13998 | n17420 ;
  assign n30633 = n30632 ^ n17296 ^ 1'b0 ;
  assign n30634 = n21018 & n30633 ;
  assign n30635 = ~n26105 & n30634 ;
  assign n30636 = n28700 ^ n22354 ^ 1'b0 ;
  assign n30637 = ( n8600 & ~n8924 ) | ( n8600 & n27015 ) | ( ~n8924 & n27015 ) ;
  assign n30638 = n24691 ^ n5065 ^ 1'b0 ;
  assign n30639 = ~n1930 & n11364 ;
  assign n30640 = n12502 & n30639 ;
  assign n30641 = n26370 ^ n7144 ^ n4592 ;
  assign n30642 = ~n13729 & n15921 ;
  assign n30643 = n30642 ^ n1140 ^ 1'b0 ;
  assign n30644 = n30643 ^ n7570 ^ 1'b0 ;
  assign n30645 = n30641 & n30644 ;
  assign n30646 = ~n21962 & n30645 ;
  assign n30647 = n30646 ^ n25217 ^ 1'b0 ;
  assign n30648 = n15854 ^ n13197 ^ n3979 ;
  assign n30649 = n6283 | n30648 ;
  assign n30650 = n30649 ^ n12459 ^ 1'b0 ;
  assign n30651 = ~n30647 & n30650 ;
  assign n30652 = n6082 | n26566 ;
  assign n30653 = n30652 ^ n6294 ^ n1468 ;
  assign n30654 = n11273 ^ n8332 ^ 1'b0 ;
  assign n30655 = ( ~n3344 & n10018 ) | ( ~n3344 & n21465 ) | ( n10018 & n21465 ) ;
  assign n30656 = n30655 ^ n2173 ^ 1'b0 ;
  assign n30657 = n15704 ^ n7538 ^ 1'b0 ;
  assign n30658 = n10528 | n30657 ;
  assign n30659 = ~n18305 & n30658 ;
  assign n30660 = ( ~n13346 & n14617 ) | ( ~n13346 & n21230 ) | ( n14617 & n21230 ) ;
  assign n30661 = n23249 & ~n30660 ;
  assign n30662 = ( ~n4070 & n7339 ) | ( ~n4070 & n8622 ) | ( n7339 & n8622 ) ;
  assign n30663 = n982 | n30662 ;
  assign n30664 = n3727 & ~n3985 ;
  assign n30665 = n19666 ^ n15224 ^ 1'b0 ;
  assign n30666 = n2665 | n30665 ;
  assign n30667 = n30666 ^ n4618 ^ 1'b0 ;
  assign n30668 = n30667 ^ n8454 ^ 1'b0 ;
  assign n30669 = n5846 & ~n30668 ;
  assign n30670 = ( n21379 & n30664 ) | ( n21379 & ~n30669 ) | ( n30664 & ~n30669 ) ;
  assign n30672 = n8258 ^ n1444 ^ 1'b0 ;
  assign n30673 = n4003 & ~n30672 ;
  assign n30674 = ~n9460 & n30673 ;
  assign n30675 = n9071 & n30674 ;
  assign n30671 = n15294 | n22710 ;
  assign n30676 = n30675 ^ n30671 ^ 1'b0 ;
  assign n30677 = ~n8783 & n16286 ;
  assign n30678 = n5237 & n30677 ;
  assign n30679 = n21071 | n27438 ;
  assign n30680 = n5027 & ~n30679 ;
  assign n30681 = n12051 & ~n15838 ;
  assign n30682 = ~n25757 & n29602 ;
  assign n30683 = n30682 ^ n5261 ^ 1'b0 ;
  assign n30684 = n2036 | n26073 ;
  assign n30685 = n24057 | n30684 ;
  assign n30686 = ( n7068 & n9002 ) | ( n7068 & ~n30685 ) | ( n9002 & ~n30685 ) ;
  assign n30687 = ( n28625 & n29730 ) | ( n28625 & ~n30686 ) | ( n29730 & ~n30686 ) ;
  assign n30690 = n16643 & ~n19356 ;
  assign n30688 = x130 & ~n21424 ;
  assign n30689 = n30688 ^ n18602 ^ 1'b0 ;
  assign n30691 = n30690 ^ n30689 ^ 1'b0 ;
  assign n30694 = n8029 & n11147 ;
  assign n30695 = ~n6021 & n30694 ;
  assign n30692 = n21463 ^ n7660 ^ 1'b0 ;
  assign n30693 = n10892 & ~n30692 ;
  assign n30696 = n30695 ^ n30693 ^ n385 ;
  assign n30697 = n25490 ^ n1103 ^ 1'b0 ;
  assign n30698 = ~n2769 & n30697 ;
  assign n30699 = ( ~n9711 & n11252 ) | ( ~n9711 & n20866 ) | ( n11252 & n20866 ) ;
  assign n30700 = n30699 ^ n2748 ^ 1'b0 ;
  assign n30701 = n7393 & n30700 ;
  assign n30702 = ~n5984 & n30701 ;
  assign n30703 = n14004 ^ n3747 ^ 1'b0 ;
  assign n30704 = n16915 | n30703 ;
  assign n30705 = ~n6717 & n11457 ;
  assign n30706 = n26638 ^ n14081 ^ 1'b0 ;
  assign n30707 = ~n6783 & n30706 ;
  assign n30708 = ( n3329 & n24039 ) | ( n3329 & n30707 ) | ( n24039 & n30707 ) ;
  assign n30710 = n2642 ^ n1816 ^ 1'b0 ;
  assign n30709 = n13921 | n14690 ;
  assign n30711 = n30710 ^ n30709 ^ 1'b0 ;
  assign n30712 = ~n3877 & n4661 ;
  assign n30713 = n30712 ^ n28172 ^ 1'b0 ;
  assign n30714 = n4703 & n25773 ;
  assign n30715 = n29642 & n30714 ;
  assign n30716 = n4090 ^ x184 ^ 1'b0 ;
  assign n30717 = n2690 & n30716 ;
  assign n30718 = n679 & ~n10566 ;
  assign n30719 = n30718 ^ n4114 ^ 1'b0 ;
  assign n30720 = n30719 ^ n1576 ^ 1'b0 ;
  assign n30721 = n5948 ^ n4326 ^ 1'b0 ;
  assign n30724 = n14717 & n27122 ;
  assign n30722 = n26718 ^ n14711 ^ n6810 ;
  assign n30723 = n7850 & ~n30722 ;
  assign n30725 = n30724 ^ n30723 ^ 1'b0 ;
  assign n30726 = n23785 | n30725 ;
  assign n30727 = n4693 | n22001 ;
  assign n30728 = n30727 ^ n6869 ^ 1'b0 ;
  assign n30729 = n1970 ^ n290 ^ 1'b0 ;
  assign n30730 = ~n7723 & n30729 ;
  assign n30731 = ( n14071 & n22831 ) | ( n14071 & ~n30730 ) | ( n22831 & ~n30730 ) ;
  assign n30732 = n30731 ^ n29413 ^ 1'b0 ;
  assign n30733 = n30728 | n30732 ;
  assign n30734 = n4910 & ~n9560 ;
  assign n30735 = ~n7929 & n30734 ;
  assign n30736 = n30735 ^ n8391 ^ 1'b0 ;
  assign n30737 = n19685 ^ n8424 ^ 1'b0 ;
  assign n30738 = n30736 | n30737 ;
  assign n30739 = ~n9860 & n12986 ;
  assign n30740 = n29543 ^ n9586 ^ n8374 ;
  assign n30748 = ~n5257 & n7867 ;
  assign n30741 = n13099 ^ n6129 ^ 1'b0 ;
  assign n30742 = ~n14172 & n30741 ;
  assign n30743 = n30742 ^ n14704 ^ n7579 ;
  assign n30744 = n30743 ^ n29649 ^ 1'b0 ;
  assign n30745 = ~n16062 & n30744 ;
  assign n30746 = ( n13229 & ~n19121 ) | ( n13229 & n30745 ) | ( ~n19121 & n30745 ) ;
  assign n30747 = n12898 & n30746 ;
  assign n30749 = n30748 ^ n30747 ^ 1'b0 ;
  assign n30750 = n30749 ^ n9562 ^ 1'b0 ;
  assign n30751 = n30740 & n30750 ;
  assign n30752 = n30751 ^ n10387 ^ 1'b0 ;
  assign n30753 = n9698 ^ n1206 ^ 1'b0 ;
  assign n30754 = n21299 | n30753 ;
  assign n30755 = n30754 ^ n27160 ^ 1'b0 ;
  assign n30756 = n4514 & n18656 ;
  assign n30757 = n30756 ^ n1452 ^ 1'b0 ;
  assign n30758 = n30757 ^ n28007 ^ n8605 ;
  assign n30759 = n3387 & ~n17089 ;
  assign n30760 = n5816 & n19920 ;
  assign n30761 = n2268 ^ n702 ^ 1'b0 ;
  assign n30762 = n17011 ^ n4274 ^ 1'b0 ;
  assign n30763 = ~n13350 & n30762 ;
  assign n30764 = n7231 ^ n6264 ^ n1898 ;
  assign n30765 = n30764 ^ n3328 ^ 1'b0 ;
  assign n30766 = n30763 & ~n30765 ;
  assign n30767 = n20879 & n30766 ;
  assign n30768 = n5071 | n16525 ;
  assign n30769 = ~n9297 & n30768 ;
  assign n30770 = n5990 ^ n792 ^ 1'b0 ;
  assign n30771 = n23909 ^ n17057 ^ 1'b0 ;
  assign n30772 = n28444 ^ n8172 ^ 1'b0 ;
  assign n30773 = n11270 & n30772 ;
  assign n30774 = ~n2280 & n3555 ;
  assign n30775 = n28807 ^ n18700 ^ 1'b0 ;
  assign n30776 = n4654 & n30775 ;
  assign n30777 = ~n1665 & n5601 ;
  assign n30778 = n30777 ^ n21508 ^ n19844 ;
  assign n30779 = ( n4115 & ~n21692 ) | ( n4115 & n30778 ) | ( ~n21692 & n30778 ) ;
  assign n30780 = n13495 ^ x238 ^ 1'b0 ;
  assign n30781 = n11518 | n30780 ;
  assign n30782 = n15730 | n30781 ;
  assign n30783 = ~n1385 & n30782 ;
  assign n30784 = n4979 & n18649 ;
  assign n30785 = n30784 ^ n1028 ^ 1'b0 ;
  assign n30786 = n10667 & ~n25223 ;
  assign n30787 = ~n30785 & n30786 ;
  assign n30788 = n30787 ^ n23587 ^ n9873 ;
  assign n30789 = n30788 ^ n18159 ^ n11357 ;
  assign n30790 = n30789 ^ n15331 ^ n2953 ;
  assign n30791 = n7841 & n11076 ;
  assign n30792 = n30791 ^ n7324 ^ 1'b0 ;
  assign n30793 = ~n18086 & n30792 ;
  assign n30794 = n22773 & n30793 ;
  assign n30800 = n14480 ^ n12471 ^ 1'b0 ;
  assign n30795 = n6620 ^ n829 ^ x238 ;
  assign n30796 = n30795 ^ x17 ^ 1'b0 ;
  assign n30797 = n5426 | n30796 ;
  assign n30798 = ~n7447 & n11418 ;
  assign n30799 = n30797 & n30798 ;
  assign n30801 = n30800 ^ n30799 ^ 1'b0 ;
  assign n30802 = n4896 & ~n30801 ;
  assign n30803 = n8444 & n10446 ;
  assign n30804 = ~n18722 & n30803 ;
  assign n30805 = n30804 ^ n7644 ^ 1'b0 ;
  assign n30806 = n17345 & n30012 ;
  assign n30807 = n15000 ^ n10532 ^ 1'b0 ;
  assign n30808 = n22627 & n30807 ;
  assign n30809 = ( n9654 & n18329 ) | ( n9654 & ~n30808 ) | ( n18329 & ~n30808 ) ;
  assign n30810 = n735 | n5884 ;
  assign n30811 = n16845 & ~n30810 ;
  assign n30812 = n1895 & n30811 ;
  assign n30813 = n5846 & ~n18938 ;
  assign n30814 = n30813 ^ n16495 ^ 1'b0 ;
  assign n30815 = ~n13350 & n30814 ;
  assign n30816 = n30815 ^ n7358 ^ 1'b0 ;
  assign n30817 = n18492 | n18758 ;
  assign n30818 = n6100 & ~n30817 ;
  assign n30819 = n30818 ^ n11631 ^ 1'b0 ;
  assign n30820 = ~n28229 & n30819 ;
  assign n30821 = ( ~x252 & n10782 ) | ( ~x252 & n10791 ) | ( n10782 & n10791 ) ;
  assign n30822 = ~n4093 & n25632 ;
  assign n30823 = ~n30821 & n30822 ;
  assign n30824 = n4600 ^ n4003 ^ n572 ;
  assign n30825 = n30824 ^ n1626 ^ 1'b0 ;
  assign n30826 = n15704 ^ n12362 ^ n5270 ;
  assign n30827 = n26180 & ~n30826 ;
  assign n30828 = ~n1958 & n30827 ;
  assign n30829 = n1196 & n15774 ;
  assign n30830 = n30829 ^ n19938 ^ 1'b0 ;
  assign n30831 = n3304 | n6458 ;
  assign n30832 = n30831 ^ n7338 ^ 1'b0 ;
  assign n30833 = ~n5642 & n30832 ;
  assign n30834 = n12788 & n30833 ;
  assign n30835 = n904 | n30834 ;
  assign n30836 = n30835 ^ n3175 ^ 1'b0 ;
  assign n30837 = n29136 & ~n30836 ;
  assign n30838 = n30837 ^ n1985 ^ 1'b0 ;
  assign n30839 = n30830 & n30838 ;
  assign n30840 = ( n3660 & ~n12052 ) | ( n3660 & n14779 ) | ( ~n12052 & n14779 ) ;
  assign n30841 = n30840 ^ n4693 ^ 1'b0 ;
  assign n30842 = n4592 ^ x70 ^ 1'b0 ;
  assign n30843 = ~n5760 & n23974 ;
  assign n30844 = n30842 & ~n30843 ;
  assign n30845 = n4221 ^ n625 ^ 1'b0 ;
  assign n30846 = n30845 ^ n1862 ^ 1'b0 ;
  assign n30847 = n15534 & n30846 ;
  assign n30848 = n13961 & ~n19078 ;
  assign n30849 = n30848 ^ n26878 ^ 1'b0 ;
  assign n30850 = n4154 & ~n30849 ;
  assign n30851 = n11531 & ~n28420 ;
  assign n30852 = ~n30440 & n30851 ;
  assign n30853 = n25720 | n30852 ;
  assign n30854 = n30853 ^ n25011 ^ 1'b0 ;
  assign n30855 = n275 | n10208 ;
  assign n30856 = n9193 ^ n4013 ^ n2670 ;
  assign n30857 = ( ~n8603 & n16341 ) | ( ~n8603 & n30856 ) | ( n16341 & n30856 ) ;
  assign n30859 = n26463 ^ n22178 ^ n12548 ;
  assign n30858 = n6546 ^ n1727 ^ n845 ;
  assign n30860 = n30859 ^ n30858 ^ n21967 ;
  assign n30861 = n17754 ^ n9050 ^ 1'b0 ;
  assign n30862 = n12053 & n27123 ;
  assign n30863 = ~n8888 & n30800 ;
  assign n30864 = n30863 ^ n17923 ^ 1'b0 ;
  assign n30866 = ~n2478 & n6820 ;
  assign n30867 = n30866 ^ n19780 ^ 1'b0 ;
  assign n30865 = n7298 | n16855 ;
  assign n30868 = n30867 ^ n30865 ^ n5134 ;
  assign n30869 = n30868 ^ n25329 ^ 1'b0 ;
  assign n30870 = n18586 ^ n17761 ^ n6945 ;
  assign n30871 = n4228 & n5535 ;
  assign n30872 = n30553 ^ n1211 ^ 1'b0 ;
  assign n30873 = ( n6069 & n27887 ) | ( n6069 & ~n30872 ) | ( n27887 & ~n30872 ) ;
  assign n30874 = ( n876 & ~n3328 ) | ( n876 & n16409 ) | ( ~n3328 & n16409 ) ;
  assign n30875 = n30874 ^ n5880 ^ 1'b0 ;
  assign n30876 = n23292 & ~n30875 ;
  assign n30877 = n9958 ^ n8286 ^ 1'b0 ;
  assign n30878 = n9044 & n30877 ;
  assign n30879 = n13986 & n17796 ;
  assign n30880 = n30879 ^ n11583 ^ 1'b0 ;
  assign n30881 = n1667 & n30880 ;
  assign n30882 = n30881 ^ n3862 ^ 1'b0 ;
  assign n30883 = n30882 ^ n6153 ^ 1'b0 ;
  assign n30884 = n2723 | n6253 ;
  assign n30885 = n30884 ^ n2183 ^ 1'b0 ;
  assign n30886 = n22030 ^ n14157 ^ 1'b0 ;
  assign n30887 = ( n21989 & ~n30885 ) | ( n21989 & n30886 ) | ( ~n30885 & n30886 ) ;
  assign n30888 = n14562 & n30785 ;
  assign n30889 = n30888 ^ n1733 ^ 1'b0 ;
  assign n30890 = n2831 & n19939 ;
  assign n30891 = ~n11691 & n30890 ;
  assign n30892 = n9083 | n25654 ;
  assign n30893 = n3945 ^ n884 ^ 1'b0 ;
  assign n30894 = n30892 & n30893 ;
  assign n30895 = ( ~n25446 & n30891 ) | ( ~n25446 & n30894 ) | ( n30891 & n30894 ) ;
  assign n30896 = ( ~n19058 & n30889 ) | ( ~n19058 & n30895 ) | ( n30889 & n30895 ) ;
  assign n30897 = n20697 ^ n3633 ^ 1'b0 ;
  assign n30898 = n22870 | n30897 ;
  assign n30899 = n2342 & n9311 ;
  assign n30900 = n7016 | n30899 ;
  assign n30901 = n30900 ^ n16788 ^ 1'b0 ;
  assign n30902 = n30898 | n30901 ;
  assign n30903 = n3196 & n10706 ;
  assign n30904 = n30902 & ~n30903 ;
  assign n30905 = ~n12812 & n26989 ;
  assign n30906 = ~n28479 & n30905 ;
  assign n30907 = n810 | n27530 ;
  assign n30908 = n4203 & ~n25185 ;
  assign n30909 = n1088 | n6967 ;
  assign n30910 = n5285 & ~n30909 ;
  assign n30911 = n30910 ^ n522 ^ 1'b0 ;
  assign n30912 = n30908 | n30911 ;
  assign n30913 = n4739 ^ n2909 ^ 1'b0 ;
  assign n30914 = n7263 & ~n30913 ;
  assign n30915 = n7736 & n11741 ;
  assign n30916 = n1204 | n30915 ;
  assign n30917 = n935 | n19479 ;
  assign n30918 = ~n2541 & n16970 ;
  assign n30919 = ~n300 & n30918 ;
  assign n30921 = n1558 | n16036 ;
  assign n30922 = n30921 ^ n8986 ^ 1'b0 ;
  assign n30920 = ~n552 & n18791 ;
  assign n30923 = n30922 ^ n30920 ^ 1'b0 ;
  assign n30924 = n27007 | n30923 ;
  assign n30925 = n30924 ^ n13066 ^ 1'b0 ;
  assign n30926 = n402 & ~n14217 ;
  assign n30927 = n30926 ^ n7464 ^ 1'b0 ;
  assign n30928 = ~n16874 & n30927 ;
  assign n30929 = n4557 & ~n30928 ;
  assign n30930 = n19940 | n30929 ;
  assign n30931 = ~n10087 & n30930 ;
  assign n30932 = n17661 ^ n8181 ^ 1'b0 ;
  assign n30933 = n14827 & n30932 ;
  assign n30934 = n25328 ^ n16258 ^ 1'b0 ;
  assign n30935 = n30933 & n30934 ;
  assign n30937 = n23539 ^ n17530 ^ 1'b0 ;
  assign n30938 = ~n6668 & n30937 ;
  assign n30936 = n12175 ^ n8079 ^ 1'b0 ;
  assign n30939 = n30938 ^ n30936 ^ 1'b0 ;
  assign n30940 = n14250 ^ n7881 ^ 1'b0 ;
  assign n30941 = n22792 & n30940 ;
  assign n30942 = n17782 & n30941 ;
  assign n30943 = n10644 & ~n12723 ;
  assign n30944 = n30943 ^ n9294 ^ 1'b0 ;
  assign n30945 = n13135 | n30944 ;
  assign n30946 = n5645 ^ n516 ^ 1'b0 ;
  assign n30947 = n21198 ^ n8438 ^ 1'b0 ;
  assign n30948 = n7554 & ~n30947 ;
  assign n30949 = n30948 ^ n7085 ^ 1'b0 ;
  assign n30950 = ~n19469 & n30949 ;
  assign n30951 = ~n15957 & n30950 ;
  assign n30952 = ~n26192 & n30951 ;
  assign n30953 = n30952 ^ n29063 ^ n5860 ;
  assign n30954 = ( n12197 & ~n30946 ) | ( n12197 & n30953 ) | ( ~n30946 & n30953 ) ;
  assign n30956 = ( n12486 & n13975 ) | ( n12486 & ~n17041 ) | ( n13975 & ~n17041 ) ;
  assign n30957 = n12120 ^ n2258 ^ 1'b0 ;
  assign n30958 = ( n1024 & n30956 ) | ( n1024 & n30957 ) | ( n30956 & n30957 ) ;
  assign n30955 = n7988 | n20804 ;
  assign n30959 = n30958 ^ n30955 ^ 1'b0 ;
  assign n30960 = n11946 ^ n8001 ^ 1'b0 ;
  assign n30961 = ~n29990 & n30960 ;
  assign n30962 = n30961 ^ n29916 ^ 1'b0 ;
  assign n30963 = n25745 ^ n9757 ^ 1'b0 ;
  assign n30964 = n6856 & ~n23254 ;
  assign n30965 = ~n30963 & n30964 ;
  assign n30966 = n30965 ^ n24928 ^ 1'b0 ;
  assign n30971 = n16138 & ~n21567 ;
  assign n30972 = n30971 ^ n25798 ^ 1'b0 ;
  assign n30967 = n16572 ^ n5827 ^ 1'b0 ;
  assign n30968 = n16101 & ~n30967 ;
  assign n30969 = n13443 ^ n12610 ^ 1'b0 ;
  assign n30970 = n30968 & ~n30969 ;
  assign n30973 = n30972 ^ n30970 ^ 1'b0 ;
  assign n30974 = n10301 ^ n3837 ^ 1'b0 ;
  assign n30975 = n20504 & ~n30974 ;
  assign n30976 = n9824 & n30975 ;
  assign n30977 = ( n16540 & ~n26175 ) | ( n16540 & n30976 ) | ( ~n26175 & n30976 ) ;
  assign n30978 = n16496 ^ n4432 ^ 1'b0 ;
  assign n30979 = ~n17130 & n30978 ;
  assign n30980 = n6001 | n6782 ;
  assign n30981 = n5992 & ~n30980 ;
  assign n30983 = n29558 ^ n28600 ^ n20497 ;
  assign n30982 = n20803 ^ n5961 ^ 1'b0 ;
  assign n30984 = n30983 ^ n30982 ^ 1'b0 ;
  assign n30985 = n22682 & ~n30984 ;
  assign n30987 = n5596 | n16917 ;
  assign n30988 = n17924 & n30987 ;
  assign n30986 = n12839 & n24222 ;
  assign n30989 = n30988 ^ n30986 ^ 1'b0 ;
  assign n30990 = ( ~n7912 & n9223 ) | ( ~n7912 & n25189 ) | ( n9223 & n25189 ) ;
  assign n30991 = n13756 & ~n20634 ;
  assign n30992 = n25618 ^ n7678 ^ 1'b0 ;
  assign n30993 = n30546 | n30992 ;
  assign n30994 = ( n6018 & n22462 ) | ( n6018 & n30993 ) | ( n22462 & n30993 ) ;
  assign n30995 = n30994 ^ n24005 ^ n1401 ;
  assign n30996 = n14934 ^ n7313 ^ 1'b0 ;
  assign n30997 = n30995 & ~n30996 ;
  assign n30998 = ( ~n30990 & n30991 ) | ( ~n30990 & n30997 ) | ( n30991 & n30997 ) ;
  assign n30999 = ( n9509 & ~n11388 ) | ( n9509 & n17188 ) | ( ~n11388 & n17188 ) ;
  assign n31000 = n5397 & ~n26071 ;
  assign n31001 = n2680 & n31000 ;
  assign n31002 = n9414 ^ n4882 ^ 1'b0 ;
  assign n31003 = n18791 ^ n9173 ^ 1'b0 ;
  assign n31004 = ~n5047 & n31003 ;
  assign n31005 = ~n31002 & n31004 ;
  assign n31006 = n13592 | n31005 ;
  assign n31007 = n31001 & ~n31006 ;
  assign n31008 = ~n18534 & n21080 ;
  assign n31009 = ~n14100 & n31008 ;
  assign n31010 = n4542 & ~n25155 ;
  assign n31011 = n17612 & n31010 ;
  assign n31012 = n16969 ^ n9948 ^ n8585 ;
  assign n31013 = ( n4465 & ~n4981 ) | ( n4465 & n7325 ) | ( ~n4981 & n7325 ) ;
  assign n31014 = n31013 ^ n26408 ^ n6606 ;
  assign n31015 = ( n11506 & n22739 ) | ( n11506 & n31014 ) | ( n22739 & n31014 ) ;
  assign n31016 = n1376 | n26108 ;
  assign n31017 = n3321 & n31016 ;
  assign n31018 = n31017 ^ n25250 ^ n13403 ;
  assign n31019 = ~n3317 & n10179 ;
  assign n31020 = n1865 & n31019 ;
  assign n31021 = n31020 ^ n12094 ^ n2061 ;
  assign n31022 = n27950 ^ n23306 ^ n18450 ;
  assign n31023 = n22427 & n31022 ;
  assign n31024 = ~n17471 & n18223 ;
  assign n31025 = n19631 & n31024 ;
  assign n31026 = n31025 ^ n30636 ^ 1'b0 ;
  assign n31027 = n16094 ^ n7252 ^ 1'b0 ;
  assign n31028 = n7427 & n31027 ;
  assign n31029 = n12500 & n16042 ;
  assign n31030 = ( ~n26878 & n31028 ) | ( ~n26878 & n31029 ) | ( n31028 & n31029 ) ;
  assign n31031 = ( n2831 & n11926 ) | ( n2831 & n11956 ) | ( n11926 & n11956 ) ;
  assign n31032 = n10194 ^ n6260 ^ 1'b0 ;
  assign n31033 = n4448 | n31032 ;
  assign n31034 = n4184 | n31033 ;
  assign n31035 = ~n7691 & n26434 ;
  assign n31036 = n31035 ^ n23522 ^ 1'b0 ;
  assign n31037 = n5739 & n31036 ;
  assign n31038 = n31037 ^ n5503 ^ 1'b0 ;
  assign n31039 = n10039 ^ n284 ^ 1'b0 ;
  assign n31040 = ~n31005 & n31039 ;
  assign n31042 = ~n1524 & n8454 ;
  assign n31043 = ~n4842 & n31042 ;
  assign n31044 = ~n5860 & n31043 ;
  assign n31045 = n509 | n31044 ;
  assign n31041 = n10804 & n19648 ;
  assign n31046 = n31045 ^ n31041 ^ 1'b0 ;
  assign n31047 = n11377 ^ n5760 ^ n1694 ;
  assign n31048 = n22127 | n31047 ;
  assign n31049 = ( ~n12912 & n16358 ) | ( ~n12912 & n18916 ) | ( n16358 & n18916 ) ;
  assign n31050 = n6284 ^ n1682 ^ 1'b0 ;
  assign n31051 = n5798 | n31050 ;
  assign n31052 = n7772 & ~n30421 ;
  assign n31058 = n7184 & ~n18182 ;
  assign n31059 = ( n8888 & n27279 ) | ( n8888 & ~n31058 ) | ( n27279 & ~n31058 ) ;
  assign n31060 = ~n10255 & n31059 ;
  assign n31061 = n7777 & n31060 ;
  assign n31053 = n4365 ^ n2845 ^ 1'b0 ;
  assign n31054 = n4461 | n31053 ;
  assign n31055 = n31054 ^ n4874 ^ 1'b0 ;
  assign n31056 = ( n4815 & n5611 ) | ( n4815 & ~n31055 ) | ( n5611 & ~n31055 ) ;
  assign n31057 = n24213 & ~n31056 ;
  assign n31062 = n31061 ^ n31057 ^ 1'b0 ;
  assign n31063 = n31062 ^ n16408 ^ 1'b0 ;
  assign n31064 = ( n10285 & n16246 ) | ( n10285 & n19004 ) | ( n16246 & n19004 ) ;
  assign n31065 = n10891 ^ n5174 ^ 1'b0 ;
  assign n31066 = ~n1971 & n31065 ;
  assign n31067 = ( n11931 & n22982 ) | ( n11931 & ~n31066 ) | ( n22982 & ~n31066 ) ;
  assign n31068 = n31067 ^ n16628 ^ 1'b0 ;
  assign n31069 = n16340 ^ n9755 ^ n517 ;
  assign n31070 = n24219 ^ n17976 ^ 1'b0 ;
  assign n31071 = n29949 ^ n843 ^ 1'b0 ;
  assign n31072 = ~n15058 & n31071 ;
  assign n31073 = n6141 & ~n31072 ;
  assign n31074 = n22959 ^ n12716 ^ 1'b0 ;
  assign n31075 = ( n8767 & n8939 ) | ( n8767 & ~n28287 ) | ( n8939 & ~n28287 ) ;
  assign n31076 = n31074 & ~n31075 ;
  assign n31077 = n31076 ^ n25793 ^ 1'b0 ;
  assign n31078 = ~n31073 & n31077 ;
  assign n31079 = n4115 & ~n23945 ;
  assign n31080 = n12301 | n14270 ;
  assign n31081 = n14119 | n31080 ;
  assign n31082 = n17123 ^ n2613 ^ 1'b0 ;
  assign n31083 = n7754 ^ n3160 ^ 1'b0 ;
  assign n31084 = ( n11463 & n16232 ) | ( n11463 & ~n31083 ) | ( n16232 & ~n31083 ) ;
  assign n31085 = n14227 ^ n13800 ^ n11973 ;
  assign n31086 = n31084 & ~n31085 ;
  assign n31087 = ( ~n8942 & n10661 ) | ( ~n8942 & n31086 ) | ( n10661 & n31086 ) ;
  assign n31088 = n1719 | n2062 ;
  assign n31089 = n1555 & ~n31088 ;
  assign n31090 = n12160 & ~n31089 ;
  assign n31091 = n31090 ^ n4200 ^ 1'b0 ;
  assign n31092 = n31091 ^ n16254 ^ 1'b0 ;
  assign n31093 = ( n4795 & n10226 ) | ( n4795 & n18983 ) | ( n10226 & n18983 ) ;
  assign n31094 = n11575 & ~n31093 ;
  assign n31095 = ( n20034 & n31092 ) | ( n20034 & ~n31094 ) | ( n31092 & ~n31094 ) ;
  assign n31096 = n6484 ^ n1271 ^ 1'b0 ;
  assign n31097 = n9948 | n31096 ;
  assign n31098 = n9095 & ~n31097 ;
  assign n31099 = ~n6484 & n11931 ;
  assign n31100 = n5973 | n6406 ;
  assign n31101 = n2016 & ~n31100 ;
  assign n31102 = ( n4112 & ~n31099 ) | ( n4112 & n31101 ) | ( ~n31099 & n31101 ) ;
  assign n31103 = n24048 & ~n31102 ;
  assign n31104 = n15859 ^ n4933 ^ 1'b0 ;
  assign n31105 = ~n31103 & n31104 ;
  assign n31106 = n21797 ^ n2680 ^ n1717 ;
  assign n31107 = n9075 | n10209 ;
  assign n31108 = n31107 ^ n10587 ^ 1'b0 ;
  assign n31109 = n5076 | n31108 ;
  assign n31110 = n23702 & ~n31109 ;
  assign n31111 = n2278 & ~n14696 ;
  assign n31114 = n9251 ^ n3775 ^ 1'b0 ;
  assign n31112 = n10044 & ~n21717 ;
  assign n31113 = n31112 ^ n29654 ^ 1'b0 ;
  assign n31115 = n31114 ^ n31113 ^ n436 ;
  assign n31116 = n2448 & ~n19532 ;
  assign n31118 = n2996 & ~n5276 ;
  assign n31119 = n31118 ^ n2708 ^ 1'b0 ;
  assign n31120 = ( n6835 & n13378 ) | ( n6835 & n31119 ) | ( n13378 & n31119 ) ;
  assign n31117 = n2854 & ~n2983 ;
  assign n31121 = n31120 ^ n31117 ^ n4460 ;
  assign n31122 = n31116 | n31121 ;
  assign n31123 = n19252 ^ n16338 ^ 1'b0 ;
  assign n31124 = n26928 ^ n15909 ^ 1'b0 ;
  assign n31125 = n22351 & n31124 ;
  assign n31126 = n2005 & ~n25084 ;
  assign n31127 = n19897 & n31126 ;
  assign n31128 = n2907 & n22236 ;
  assign n31129 = ( ~x167 & n6536 ) | ( ~x167 & n28243 ) | ( n6536 & n28243 ) ;
  assign n31130 = n31129 ^ n25512 ^ 1'b0 ;
  assign n31131 = n12313 ^ n7998 ^ 1'b0 ;
  assign n31132 = n18027 ^ n7927 ^ 1'b0 ;
  assign n31133 = n31131 | n31132 ;
  assign n31134 = n23801 & n31133 ;
  assign n31140 = n3559 & n5672 ;
  assign n31141 = n11586 & n31140 ;
  assign n31135 = n23858 ^ n834 ^ 1'b0 ;
  assign n31136 = n22070 ^ n9939 ^ 1'b0 ;
  assign n31137 = n31135 & n31136 ;
  assign n31138 = n19031 & n31137 ;
  assign n31139 = n13213 | n31138 ;
  assign n31142 = n31141 ^ n31139 ^ 1'b0 ;
  assign n31143 = ~n787 & n2054 ;
  assign n31144 = n17562 | n27626 ;
  assign n31145 = n24335 ^ n15285 ^ 1'b0 ;
  assign n31146 = n8225 | n31145 ;
  assign n31147 = n16857 & ~n28143 ;
  assign n31148 = ~n20239 & n31147 ;
  assign n31149 = n25231 ^ n24416 ^ 1'b0 ;
  assign n31150 = n10928 | n21831 ;
  assign n31151 = ( n9467 & ~n10272 ) | ( n9467 & n18310 ) | ( ~n10272 & n18310 ) ;
  assign n31152 = ( n24618 & n27540 ) | ( n24618 & ~n31151 ) | ( n27540 & ~n31151 ) ;
  assign n31153 = n31150 & ~n31152 ;
  assign n31154 = n6068 ^ n2138 ^ 1'b0 ;
  assign n31155 = ~n2481 & n31154 ;
  assign n31156 = ( n4234 & ~n10381 ) | ( n4234 & n31155 ) | ( ~n10381 & n31155 ) ;
  assign n31157 = n5014 & ~n17428 ;
  assign n31158 = n31157 ^ n16172 ^ 1'b0 ;
  assign n31159 = n2643 | n12843 ;
  assign n31160 = n20772 ^ n3148 ^ 1'b0 ;
  assign n31161 = n14243 ^ n8281 ^ 1'b0 ;
  assign n31162 = ~n30908 & n31161 ;
  assign n31163 = n3223 | n12826 ;
  assign n31164 = n31163 ^ n29029 ^ 1'b0 ;
  assign n31165 = n6213 & ~n31164 ;
  assign n31166 = n369 & n31165 ;
  assign n31167 = n22089 ^ n6547 ^ 1'b0 ;
  assign n31168 = n4764 & ~n25403 ;
  assign n31169 = n11838 & ~n27327 ;
  assign n31170 = n31169 ^ n2028 ^ 1'b0 ;
  assign n31171 = ( n8896 & n17270 ) | ( n8896 & n23091 ) | ( n17270 & n23091 ) ;
  assign n31172 = ( n8922 & ~n12621 ) | ( n8922 & n22986 ) | ( ~n12621 & n22986 ) ;
  assign n31173 = n31172 ^ n30757 ^ 1'b0 ;
  assign n31174 = n31173 ^ n10900 ^ 1'b0 ;
  assign n31175 = ~n31171 & n31174 ;
  assign n31176 = ~n5170 & n13129 ;
  assign n31177 = ~n14242 & n31176 ;
  assign n31178 = n500 | n14234 ;
  assign n31179 = ( n5416 & n6703 ) | ( n5416 & ~n31178 ) | ( n6703 & ~n31178 ) ;
  assign n31180 = n31179 ^ n6124 ^ n587 ;
  assign n31181 = n5060 | n12677 ;
  assign n31182 = n20252 & n31181 ;
  assign n31183 = n31180 & ~n31182 ;
  assign n31184 = n15493 & n25516 ;
  assign n31185 = n28133 ^ n7569 ^ n369 ;
  assign n31186 = ~n26615 & n31185 ;
  assign n31187 = n31186 ^ n21331 ^ 1'b0 ;
  assign n31188 = n27912 | n31187 ;
  assign n31189 = n31188 ^ n14721 ^ 1'b0 ;
  assign n31190 = ~n10885 & n22896 ;
  assign n31191 = n13297 ^ n4024 ^ 1'b0 ;
  assign n31192 = n5753 | n31191 ;
  assign n31193 = n5741 | n22287 ;
  assign n31194 = n31192 | n31193 ;
  assign n31195 = n31194 ^ n23952 ^ 1'b0 ;
  assign n31196 = n10777 ^ n5984 ^ 1'b0 ;
  assign n31197 = ~n8878 & n31196 ;
  assign n31198 = n16987 & ~n25657 ;
  assign n31199 = n7789 | n31198 ;
  assign n31200 = n9874 ^ n8191 ^ 1'b0 ;
  assign n31201 = n19915 & ~n31200 ;
  assign n31202 = n31201 ^ n16749 ^ 1'b0 ;
  assign n31203 = n6645 ^ n2283 ^ 1'b0 ;
  assign n31204 = ~n2445 & n31203 ;
  assign n31205 = ( n5376 & n27752 ) | ( n5376 & n31204 ) | ( n27752 & n31204 ) ;
  assign n31207 = n9719 ^ n2209 ^ n686 ;
  assign n31208 = n31207 ^ n18079 ^ 1'b0 ;
  assign n31209 = ( n10558 & n28727 ) | ( n10558 & ~n31208 ) | ( n28727 & ~n31208 ) ;
  assign n31210 = n1176 | n31209 ;
  assign n31206 = ~n11420 & n23359 ;
  assign n31211 = n31210 ^ n31206 ^ 1'b0 ;
  assign n31212 = n7529 & n31211 ;
  assign n31213 = x250 & ~n11376 ;
  assign n31214 = n31213 ^ n14597 ^ 1'b0 ;
  assign n31215 = ( n920 & n14691 ) | ( n920 & n28614 ) | ( n14691 & n28614 ) ;
  assign n31216 = ( ~n644 & n2449 ) | ( ~n644 & n9678 ) | ( n2449 & n9678 ) ;
  assign n31217 = n20806 | n31216 ;
  assign n31218 = n31217 ^ n16175 ^ 1'b0 ;
  assign n31219 = n20678 ^ n6585 ^ 1'b0 ;
  assign n31220 = n17131 & n31219 ;
  assign n31221 = ~n14810 & n31220 ;
  assign n31222 = n26604 & ~n31221 ;
  assign n31225 = n8515 ^ n7585 ^ 1'b0 ;
  assign n31226 = n17912 & ~n31225 ;
  assign n31223 = n5206 & n12962 ;
  assign n31224 = n31223 ^ n19775 ^ 1'b0 ;
  assign n31227 = n31226 ^ n31224 ^ 1'b0 ;
  assign n31228 = n8697 & ~n16826 ;
  assign n31229 = n30995 & n31228 ;
  assign n31230 = n9217 & ~n13079 ;
  assign n31231 = n15696 & n22917 ;
  assign n31232 = ~n16751 & n17654 ;
  assign n31233 = ~n4975 & n31232 ;
  assign n31234 = x128 & ~n10902 ;
  assign n31235 = n31234 ^ n12471 ^ 1'b0 ;
  assign n31236 = ~n1450 & n19281 ;
  assign n31237 = n2645 | n8851 ;
  assign n31238 = n6468 | n17652 ;
  assign n31239 = n8029 | n31238 ;
  assign n31240 = n936 & n14606 ;
  assign n31241 = ( n27817 & ~n31239 ) | ( n27817 & n31240 ) | ( ~n31239 & n31240 ) ;
  assign n31242 = n790 & ~n16104 ;
  assign n31243 = n24179 ^ n3568 ^ 1'b0 ;
  assign n31244 = n23631 & ~n31243 ;
  assign n31245 = n4410 & n31244 ;
  assign n31246 = n25710 ^ n12677 ^ 1'b0 ;
  assign n31247 = ( n2056 & ~n2202 ) | ( n2056 & n31246 ) | ( ~n2202 & n31246 ) ;
  assign n31248 = n4761 ^ n2637 ^ 1'b0 ;
  assign n31249 = ( n2469 & n3621 ) | ( n2469 & n17414 ) | ( n3621 & n17414 ) ;
  assign n31250 = n21689 & n31249 ;
  assign n31251 = n31250 ^ n16740 ^ 1'b0 ;
  assign n31252 = ( ~n5033 & n16187 ) | ( ~n5033 & n23427 ) | ( n16187 & n23427 ) ;
  assign n31253 = ~n8964 & n31252 ;
  assign n31254 = ~n14626 & n26236 ;
  assign n31255 = n31254 ^ n25784 ^ 1'b0 ;
  assign n31256 = n28046 ^ n18674 ^ n13158 ;
  assign n31257 = ( n9881 & ~n25135 ) | ( n9881 & n29890 ) | ( ~n25135 & n29890 ) ;
  assign n31258 = n21369 ^ n12340 ^ n2994 ;
  assign n31259 = ~n5536 & n31258 ;
  assign n31260 = n10687 ^ n2613 ^ 1'b0 ;
  assign n31263 = n17371 ^ n7329 ^ 1'b0 ;
  assign n31264 = n31263 ^ n28889 ^ n18926 ;
  assign n31265 = n13669 ^ n12812 ^ 1'b0 ;
  assign n31266 = ~n19802 & n31265 ;
  assign n31267 = n31266 ^ n17250 ^ n14850 ;
  assign n31268 = ( ~n27426 & n31264 ) | ( ~n27426 & n31267 ) | ( n31264 & n31267 ) ;
  assign n31261 = n9345 & n9548 ;
  assign n31262 = n31261 ^ n6156 ^ 1'b0 ;
  assign n31269 = n31268 ^ n31262 ^ 1'b0 ;
  assign n31270 = n9044 ^ n7684 ^ 1'b0 ;
  assign n31271 = ~n20280 & n27384 ;
  assign n31272 = n31271 ^ n15614 ^ 1'b0 ;
  assign n31273 = n20899 ^ n16462 ^ n14869 ;
  assign n31274 = ~n11364 & n22146 ;
  assign n31275 = ( n15590 & n24839 ) | ( n15590 & ~n31274 ) | ( n24839 & ~n31274 ) ;
  assign n31276 = n31275 ^ n19228 ^ n10127 ;
  assign n31277 = ~n18017 & n29386 ;
  assign n31278 = n2178 & n7499 ;
  assign n31279 = n23905 ^ n7091 ^ 1'b0 ;
  assign n31280 = ~n31278 & n31279 ;
  assign n31281 = n30669 & ~n31280 ;
  assign n31282 = n14955 & n15506 ;
  assign n31283 = n31282 ^ n16847 ^ 1'b0 ;
  assign n31284 = n31283 ^ n1283 ^ 1'b0 ;
  assign n31285 = n17180 & n31284 ;
  assign n31286 = n16094 ^ n5296 ^ 1'b0 ;
  assign n31287 = ( ~n5071 & n15766 ) | ( ~n5071 & n23936 ) | ( n15766 & n23936 ) ;
  assign n31288 = ( n29017 & n31286 ) | ( n29017 & n31287 ) | ( n31286 & n31287 ) ;
  assign n31289 = n25932 ^ n18208 ^ n4432 ;
  assign n31290 = n20363 & n31158 ;
  assign n31291 = n31290 ^ n5425 ^ 1'b0 ;
  assign n31292 = n17661 ^ n12624 ^ 1'b0 ;
  assign n31293 = n4084 & n16996 ;
  assign n31294 = ~n31292 & n31293 ;
  assign n31295 = n31294 ^ n25198 ^ 1'b0 ;
  assign n31296 = n1366 & n31295 ;
  assign n31297 = n9154 & n22326 ;
  assign n31298 = n31297 ^ n6403 ^ n1239 ;
  assign n31299 = n3073 & ~n7522 ;
  assign n31300 = n31299 ^ n15524 ^ n1754 ;
  assign n31302 = n360 & n789 ;
  assign n31303 = ~x99 & n31302 ;
  assign n31301 = n13774 ^ n9944 ^ x184 ;
  assign n31304 = n31303 ^ n31301 ^ n2171 ;
  assign n31305 = ( ~n8777 & n31300 ) | ( ~n8777 & n31304 ) | ( n31300 & n31304 ) ;
  assign n31306 = ( n2204 & ~n14324 ) | ( n2204 & n19929 ) | ( ~n14324 & n19929 ) ;
  assign n31307 = ( n459 & n8963 ) | ( n459 & n22269 ) | ( n8963 & n22269 ) ;
  assign n31308 = n21654 ^ n13583 ^ 1'b0 ;
  assign n31309 = ~n7057 & n31308 ;
  assign n31310 = n10704 | n31309 ;
  assign n31311 = ~n2208 & n24024 ;
  assign n31312 = n31311 ^ n14805 ^ 1'b0 ;
  assign n31313 = ~n13503 & n31312 ;
  assign n31314 = n17570 ^ n5798 ^ 1'b0 ;
  assign n31315 = n792 & n31314 ;
  assign n31316 = n31315 ^ n19299 ^ 1'b0 ;
  assign n31317 = n31313 & ~n31316 ;
  assign n31318 = n25177 & ~n26928 ;
  assign n31319 = n3136 | n7814 ;
  assign n31320 = n31319 ^ n7840 ^ 1'b0 ;
  assign n31321 = n22905 ^ n18844 ^ 1'b0 ;
  assign n31322 = ~n4609 & n31321 ;
  assign n31323 = ~n13516 & n31322 ;
  assign n31324 = ~n30087 & n31323 ;
  assign n31325 = n31320 & n31324 ;
  assign n31326 = n10318 & ~n17826 ;
  assign n31327 = n20009 ^ n366 ^ 1'b0 ;
  assign n31328 = n256 & n945 ;
  assign n31329 = n30972 & n31328 ;
  assign n31330 = ( ~n8949 & n9815 ) | ( ~n8949 & n18255 ) | ( n9815 & n18255 ) ;
  assign n31331 = n31330 ^ n5317 ^ 1'b0 ;
  assign n31332 = ~n16083 & n31331 ;
  assign n31333 = ( n20517 & n27754 ) | ( n20517 & n31332 ) | ( n27754 & n31332 ) ;
  assign n31334 = n14172 ^ n1155 ^ 1'b0 ;
  assign n31335 = n31334 ^ n11093 ^ n11087 ;
  assign n31336 = ~n841 & n31335 ;
  assign n31337 = n10205 & n31336 ;
  assign n31338 = n24634 ^ n18158 ^ 1'b0 ;
  assign n31339 = ~n15487 & n31338 ;
  assign n31340 = n13010 | n31339 ;
  assign n31341 = ( n6717 & ~n8251 ) | ( n6717 & n31340 ) | ( ~n8251 & n31340 ) ;
  assign n31342 = n12194 & n12244 ;
  assign n31343 = ~n1307 & n14658 ;
  assign n31344 = ~n31342 & n31343 ;
  assign n31345 = n1893 ^ n801 ^ 1'b0 ;
  assign n31346 = ~n13831 & n16901 ;
  assign n31347 = ~n31345 & n31346 ;
  assign n31348 = n17033 | n17991 ;
  assign n31349 = n4351 & ~n31348 ;
  assign n31350 = n31349 ^ n15931 ^ n9472 ;
  assign n31351 = ~n1769 & n31350 ;
  assign n31352 = n23338 ^ n21780 ^ 1'b0 ;
  assign n31353 = n20731 | n31352 ;
  assign n31358 = ~n4791 & n8149 ;
  assign n31359 = n31358 ^ n18711 ^ n4707 ;
  assign n31354 = n16095 ^ n7331 ^ n1558 ;
  assign n31355 = n31354 ^ n9221 ^ n8927 ;
  assign n31356 = ~n27993 & n31355 ;
  assign n31357 = ~n14603 & n31356 ;
  assign n31360 = n31359 ^ n31357 ^ n12619 ;
  assign n31361 = n20645 & ~n26421 ;
  assign n31362 = n31361 ^ n16550 ^ 1'b0 ;
  assign n31363 = n2189 & n29568 ;
  assign n31364 = n1349 & ~n4806 ;
  assign n31365 = n31364 ^ n19873 ^ n14085 ;
  assign n31366 = n12676 & n31365 ;
  assign n31367 = ~n26993 & n31366 ;
  assign n31368 = n3088 & ~n14517 ;
  assign n31369 = n31367 & n31368 ;
  assign n31370 = n4270 | n16075 ;
  assign n31371 = n31370 ^ n14886 ^ 1'b0 ;
  assign n31372 = n17056 & n31371 ;
  assign n31373 = n10661 ^ n390 ^ 1'b0 ;
  assign n31374 = n27816 & n31373 ;
  assign n31375 = n20530 & ~n31374 ;
  assign n31376 = n18084 ^ n11622 ^ 1'b0 ;
  assign n31377 = ( n4686 & n9548 ) | ( n4686 & ~n16232 ) | ( n9548 & ~n16232 ) ;
  assign n31378 = n31377 ^ n24914 ^ n10661 ;
  assign n31379 = n8200 & n19066 ;
  assign n31380 = n31379 ^ n15782 ^ 1'b0 ;
  assign n31381 = n3518 | n17589 ;
  assign n31382 = n10503 | n31381 ;
  assign n31383 = n10301 | n15451 ;
  assign n31384 = n27752 & ~n31383 ;
  assign n31385 = ( n14097 & n21834 ) | ( n14097 & n21875 ) | ( n21834 & n21875 ) ;
  assign n31386 = ~n10247 & n26566 ;
  assign n31387 = ~n10194 & n31386 ;
  assign n31388 = n31387 ^ n20389 ^ 1'b0 ;
  assign n31389 = n4505 & n24438 ;
  assign n31390 = n31388 & ~n31389 ;
  assign n31391 = n31385 & n31390 ;
  assign n31392 = n3637 | n9721 ;
  assign n31393 = n31392 ^ n9373 ^ 1'b0 ;
  assign n31394 = n15411 & n31393 ;
  assign n31395 = n6829 & ~n27703 ;
  assign n31396 = ~n31394 & n31395 ;
  assign n31397 = ( ~n5386 & n12671 ) | ( ~n5386 & n18913 ) | ( n12671 & n18913 ) ;
  assign n31398 = ( n9880 & ~n11388 ) | ( n9880 & n20293 ) | ( ~n11388 & n20293 ) ;
  assign n31399 = ~n6232 & n31398 ;
  assign n31401 = n16202 ^ n9967 ^ n7519 ;
  assign n31402 = ~n1964 & n15035 ;
  assign n31403 = ( n4827 & n31401 ) | ( n4827 & ~n31402 ) | ( n31401 & ~n31402 ) ;
  assign n31400 = n14694 | n25269 ;
  assign n31404 = n31403 ^ n31400 ^ 1'b0 ;
  assign n31405 = n8244 | n31404 ;
  assign n31406 = n13618 ^ n7342 ^ 1'b0 ;
  assign n31407 = n1300 & ~n31406 ;
  assign n31408 = ( n12282 & ~n17116 ) | ( n12282 & n22771 ) | ( ~n17116 & n22771 ) ;
  assign n31410 = n7878 | n16187 ;
  assign n31409 = n14542 ^ n11510 ^ 1'b0 ;
  assign n31411 = n31410 ^ n31409 ^ n29839 ;
  assign n31412 = n30310 ^ n9454 ^ n7675 ;
  assign n31413 = n9995 ^ n6487 ^ 1'b0 ;
  assign n31414 = n21381 & n31413 ;
  assign n31415 = ~n18983 & n31414 ;
  assign n31416 = ~n4107 & n31415 ;
  assign n31417 = n18697 ^ n16638 ^ 1'b0 ;
  assign n31418 = n13267 ^ n9447 ^ n2680 ;
  assign n31419 = n11428 | n11923 ;
  assign n31420 = n31418 | n31419 ;
  assign n31421 = n14381 & ~n31420 ;
  assign n31422 = n6665 & n31421 ;
  assign n31423 = ~n31417 & n31422 ;
  assign n31424 = n15989 ^ n14538 ^ 1'b0 ;
  assign n31425 = n23073 ^ n1211 ^ 1'b0 ;
  assign n31426 = n13716 & ~n31425 ;
  assign n31427 = ~n28998 & n31426 ;
  assign n31428 = ~n6074 & n31427 ;
  assign n31429 = n20155 ^ n4763 ^ 1'b0 ;
  assign n31430 = n5688 & ~n31429 ;
  assign n31431 = n4789 & n31430 ;
  assign n31432 = n23617 ^ n20862 ^ n14863 ;
  assign n31433 = n31432 ^ n7339 ^ x251 ;
  assign n31434 = n18758 | n31433 ;
  assign n31435 = n23991 | n31434 ;
  assign n31436 = ( n19319 & n27875 ) | ( n19319 & ~n28627 ) | ( n27875 & ~n28627 ) ;
  assign n31437 = n9461 ^ n7699 ^ 1'b0 ;
  assign n31438 = n23503 | n31437 ;
  assign n31440 = ~n1636 & n7649 ;
  assign n31441 = ~n27049 & n31440 ;
  assign n31439 = n7575 | n13519 ;
  assign n31442 = n31441 ^ n31439 ^ 1'b0 ;
  assign n31443 = ( n6850 & ~n13250 ) | ( n6850 & n16193 ) | ( ~n13250 & n16193 ) ;
  assign n31444 = ~n2827 & n6981 ;
  assign n31445 = n743 & ~n31444 ;
  assign n31446 = ~n31443 & n31445 ;
  assign n31447 = n6735 | n17626 ;
  assign n31451 = n12787 ^ n12579 ^ n3023 ;
  assign n31450 = n7370 | n9853 ;
  assign n31448 = n21259 ^ n16609 ^ 1'b0 ;
  assign n31449 = n4046 | n31448 ;
  assign n31452 = n31451 ^ n31450 ^ n31449 ;
  assign n31453 = n11095 & n28158 ;
  assign n31454 = n22773 ^ n16085 ^ 1'b0 ;
  assign n31455 = ~n11361 & n14102 ;
  assign n31456 = n31455 ^ n21997 ^ 1'b0 ;
  assign n31457 = n1904 & ~n31456 ;
  assign n31458 = ~n19042 & n31457 ;
  assign n31459 = n1559 & n5535 ;
  assign n31460 = n31459 ^ n21640 ^ 1'b0 ;
  assign n31465 = n11230 ^ n944 ^ 1'b0 ;
  assign n31466 = ~n14366 & n31465 ;
  assign n31461 = n22839 & n25678 ;
  assign n31462 = n31461 ^ n19074 ^ 1'b0 ;
  assign n31463 = ( n4455 & n10165 ) | ( n4455 & ~n31462 ) | ( n10165 & ~n31462 ) ;
  assign n31464 = n31028 & n31463 ;
  assign n31467 = n31466 ^ n31464 ^ 1'b0 ;
  assign n31468 = ( n6483 & n11370 ) | ( n6483 & n18336 ) | ( n11370 & n18336 ) ;
  assign n31469 = n21755 & ~n31468 ;
  assign n31470 = n5675 ^ n5447 ^ 1'b0 ;
  assign n31471 = ( x162 & n12985 ) | ( x162 & n26488 ) | ( n12985 & n26488 ) ;
  assign n31472 = n22801 ^ n4985 ^ 1'b0 ;
  assign n31473 = n31471 & ~n31472 ;
  assign n31474 = n9802 ^ n9076 ^ 1'b0 ;
  assign n31475 = n2022 | n7186 ;
  assign n31476 = ( ~n2908 & n24691 ) | ( ~n2908 & n31475 ) | ( n24691 & n31475 ) ;
  assign n31477 = ~n29183 & n31476 ;
  assign n31478 = n17259 & n31477 ;
  assign n31479 = ~n3556 & n22799 ;
  assign n31480 = n23391 | n26181 ;
  assign n31482 = ( ~n5097 & n5712 ) | ( ~n5097 & n21203 ) | ( n5712 & n21203 ) ;
  assign n31481 = n14867 ^ n5137 ^ n282 ;
  assign n31483 = n31482 ^ n31481 ^ 1'b0 ;
  assign n31484 = n6896 & n21343 ;
  assign n31485 = n13620 & n18780 ;
  assign n31486 = n31485 ^ n19195 ^ 1'b0 ;
  assign n31487 = n15156 & ~n31486 ;
  assign n31488 = n16349 ^ n12353 ^ n7282 ;
  assign n31489 = n18416 & ~n31488 ;
  assign n31490 = n4476 | n23374 ;
  assign n31491 = n31490 ^ n14588 ^ 1'b0 ;
  assign n31492 = n14026 & ~n14138 ;
  assign n31493 = n14831 & n31492 ;
  assign n31494 = n31493 ^ n8155 ^ 1'b0 ;
  assign n31500 = n2893 ^ n2527 ^ 1'b0 ;
  assign n31501 = n2150 & ~n31500 ;
  assign n31502 = ( ~n13295 & n18275 ) | ( ~n13295 & n31501 ) | ( n18275 & n31501 ) ;
  assign n31495 = n4447 & n7413 ;
  assign n31496 = ~n23795 & n24487 ;
  assign n31497 = n31495 & n31496 ;
  assign n31498 = n15838 | n22802 ;
  assign n31499 = n31497 & ~n31498 ;
  assign n31503 = n31502 ^ n31499 ^ n14881 ;
  assign n31504 = n7823 & n9141 ;
  assign n31505 = ~n3361 & n31504 ;
  assign n31506 = n21272 & n30689 ;
  assign n31507 = n31506 ^ n10473 ^ 1'b0 ;
  assign n31508 = n393 & n31507 ;
  assign n31509 = n27068 & n31508 ;
  assign n31510 = ~n9742 & n28970 ;
  assign n31511 = n8523 & n31510 ;
  assign n31512 = n19669 | n19728 ;
  assign n31513 = n27199 ^ n26566 ^ n1140 ;
  assign n31514 = n31513 ^ n24445 ^ n17348 ;
  assign n31515 = n5741 | n7952 ;
  assign n31516 = n10381 | n31515 ;
  assign n31517 = n8589 & n21222 ;
  assign n31518 = ~n31516 & n31517 ;
  assign n31519 = n6547 & n11007 ;
  assign n31520 = n13640 ^ n10220 ^ x79 ;
  assign n31521 = n16693 & n16781 ;
  assign n31522 = ~n31520 & n31521 ;
  assign n31523 = n31522 ^ n14387 ^ 1'b0 ;
  assign n31524 = ~n15707 & n19674 ;
  assign n31525 = n31524 ^ n10076 ^ 1'b0 ;
  assign n31526 = n701 & n31525 ;
  assign n31527 = n21625 ^ n9155 ^ 1'b0 ;
  assign n31528 = n6292 & ~n21919 ;
  assign n31529 = n31528 ^ n25577 ^ n1944 ;
  assign n31530 = ( n10527 & ~n25274 ) | ( n10527 & n27160 ) | ( ~n25274 & n27160 ) ;
  assign n31531 = n3102 & ~n6606 ;
  assign n31532 = n5449 & n11900 ;
  assign n31533 = ~n16104 & n31532 ;
  assign n31534 = ~n3719 & n26612 ;
  assign n31535 = n31533 & n31534 ;
  assign n31538 = n15664 ^ n12812 ^ n12275 ;
  assign n31539 = n31538 ^ n10230 ^ 1'b0 ;
  assign n31536 = n11187 & ~n28535 ;
  assign n31537 = n9944 & n31536 ;
  assign n31540 = n31539 ^ n31537 ^ n16761 ;
  assign n31541 = n31540 ^ n6775 ^ 1'b0 ;
  assign n31542 = n20021 & n31541 ;
  assign n31543 = n7208 | n19302 ;
  assign n31544 = ( n21709 & ~n30766 ) | ( n21709 & n31543 ) | ( ~n30766 & n31543 ) ;
  assign n31545 = n23898 ^ n21003 ^ n16325 ;
  assign n31546 = ( ~n17639 & n17987 ) | ( ~n17639 & n31545 ) | ( n17987 & n31545 ) ;
  assign n31547 = n519 ^ x246 ^ 1'b0 ;
  assign n31548 = n31547 ^ n23287 ^ n18794 ;
  assign n31549 = n8026 ^ n1832 ^ 1'b0 ;
  assign n31550 = ~n5134 & n31549 ;
  assign n31551 = n31550 ^ n19690 ^ 1'b0 ;
  assign n31552 = n10654 ^ n9575 ^ n2135 ;
  assign n31553 = n31552 ^ n4698 ^ 1'b0 ;
  assign n31560 = n17603 ^ n4260 ^ 1'b0 ;
  assign n31561 = n14909 & n31560 ;
  assign n31562 = n31561 ^ n19858 ^ n16911 ;
  assign n31555 = ~n4641 & n7037 ;
  assign n31556 = n31555 ^ n3556 ^ 1'b0 ;
  assign n31554 = ~n5235 & n11839 ;
  assign n31557 = n31556 ^ n31554 ^ 1'b0 ;
  assign n31558 = n932 | n31557 ;
  assign n31559 = n9078 & ~n31558 ;
  assign n31563 = n31562 ^ n31559 ^ 1'b0 ;
  assign n31564 = ~n10221 & n11920 ;
  assign n31565 = n31564 ^ n9548 ^ 1'b0 ;
  assign n31566 = n26930 ^ n12589 ^ n743 ;
  assign n31567 = ~n16874 & n30874 ;
  assign n31568 = ~n4007 & n12114 ;
  assign n31569 = n9164 & n31568 ;
  assign n31570 = ~n260 & n5185 ;
  assign n31571 = n19421 & n31570 ;
  assign n31572 = n9399 | n22827 ;
  assign n31573 = n18460 ^ n13675 ^ 1'b0 ;
  assign n31574 = ~n2511 & n31573 ;
  assign n31575 = n31574 ^ n15713 ^ n12322 ;
  assign n31576 = n15733 ^ n11370 ^ 1'b0 ;
  assign n31577 = n797 & n31576 ;
  assign n31578 = n21826 & ~n24223 ;
  assign n31579 = n31577 | n31578 ;
  assign n31580 = n8633 | n30028 ;
  assign n31581 = n1034 & ~n31580 ;
  assign n31582 = ~n5819 & n24986 ;
  assign n31583 = n13837 & n25853 ;
  assign n31584 = ~n6231 & n31583 ;
  assign n31585 = n31584 ^ n17262 ^ 1'b0 ;
  assign n31586 = ( n19092 & n31582 ) | ( n19092 & ~n31585 ) | ( n31582 & ~n31585 ) ;
  assign n31587 = ~n12315 & n15962 ;
  assign n31588 = ~n7639 & n31587 ;
  assign n31589 = ~n3190 & n31588 ;
  assign n31590 = n13140 ^ n5761 ^ 1'b0 ;
  assign n31591 = ( n10770 & n10937 ) | ( n10770 & n21574 ) | ( n10937 & n21574 ) ;
  assign n31592 = n31591 ^ n9217 ^ 1'b0 ;
  assign n31593 = n31590 & n31592 ;
  assign n31594 = n6114 & ~n12920 ;
  assign n31595 = n22860 ^ n268 ^ 1'b0 ;
  assign n31596 = n7389 & n31595 ;
  assign n31597 = n3057 & n7339 ;
  assign n31598 = n31597 ^ n18636 ^ 1'b0 ;
  assign n31599 = n31598 ^ n13578 ^ 1'b0 ;
  assign n31600 = ( n3770 & n24211 ) | ( n3770 & n31285 ) | ( n24211 & n31285 ) ;
  assign n31601 = n18145 & ~n18329 ;
  assign n31602 = n2730 & n31601 ;
  assign n31603 = x162 & ~n15771 ;
  assign n31604 = n31603 ^ n15373 ^ 1'b0 ;
  assign n31605 = n22016 & ~n31604 ;
  assign n31606 = n31605 ^ n31249 ^ 1'b0 ;
  assign n31607 = n4952 & ~n11231 ;
  assign n31608 = n31607 ^ n29048 ^ n10261 ;
  assign n31609 = n18894 ^ n11380 ^ n3274 ;
  assign n31610 = n27411 | n31609 ;
  assign n31611 = n2722 | n4327 ;
  assign n31612 = n15486 & ~n20665 ;
  assign n31613 = ~n31611 & n31612 ;
  assign n31614 = n31182 ^ n22549 ^ 1'b0 ;
  assign n31615 = n5681 & ~n11336 ;
  assign n31616 = n21181 & ~n25081 ;
  assign n31617 = n17015 & n31616 ;
  assign n31618 = n16491 & ~n16876 ;
  assign n31619 = n25372 ^ n3147 ^ 1'b0 ;
  assign n31620 = n31619 ^ n4242 ^ 1'b0 ;
  assign n31621 = ~n31618 & n31620 ;
  assign n31622 = n10138 & ~n11221 ;
  assign n31623 = ~n2750 & n26470 ;
  assign n31624 = ( ~n5519 & n11047 ) | ( ~n5519 & n31623 ) | ( n11047 & n31623 ) ;
  assign n31625 = n31624 ^ n5813 ^ n629 ;
  assign n31626 = n8515 & ~n24474 ;
  assign n31629 = ~n4556 & n8837 ;
  assign n31630 = ~n6207 & n31629 ;
  assign n31627 = n3088 & ~n20219 ;
  assign n31628 = n3675 & n31627 ;
  assign n31631 = n31630 ^ n31628 ^ n5402 ;
  assign n31632 = ~n3403 & n14057 ;
  assign n31633 = ( n19821 & ~n31631 ) | ( n19821 & n31632 ) | ( ~n31631 & n31632 ) ;
  assign n31634 = n5721 | n7378 ;
  assign n31635 = n20821 | n31634 ;
  assign n31636 = n22798 | n31635 ;
  assign n31637 = n7003 | n13327 ;
  assign n31638 = n31637 ^ n27209 ^ 1'b0 ;
  assign n31639 = n20459 | n31638 ;
  assign n31640 = n3464 | n31639 ;
  assign n31641 = ~n2524 & n8556 ;
  assign n31642 = n7578 ^ n6756 ^ 1'b0 ;
  assign n31643 = n31642 ^ n29027 ^ n602 ;
  assign n31648 = n8542 | n13503 ;
  assign n31649 = n3508 & ~n31648 ;
  assign n31650 = ~n31029 & n31649 ;
  assign n31644 = n23845 ^ n6006 ^ n692 ;
  assign n31645 = n8299 ^ n6606 ^ 1'b0 ;
  assign n31646 = n31644 & ~n31645 ;
  assign n31647 = n12766 & n31646 ;
  assign n31651 = n31650 ^ n31647 ^ 1'b0 ;
  assign n31652 = n1479 & n5532 ;
  assign n31653 = n31652 ^ n18253 ^ 1'b0 ;
  assign n31654 = n22917 | n31653 ;
  assign n31655 = n7065 ^ n3980 ^ 1'b0 ;
  assign n31656 = n2736 & n31655 ;
  assign n31657 = n7620 ^ n7488 ^ 1'b0 ;
  assign n31658 = n31657 ^ n13218 ^ 1'b0 ;
  assign n31659 = ~n17916 & n31658 ;
  assign n31660 = n12904 ^ n697 ^ 1'b0 ;
  assign n31661 = n7099 & n31660 ;
  assign n31662 = ~n15969 & n25286 ;
  assign n31663 = n31662 ^ n27044 ^ n2873 ;
  assign n31664 = n4788 & n8129 ;
  assign n31665 = n15577 & ~n31664 ;
  assign n31666 = ~n5331 & n31665 ;
  assign n31667 = n31666 ^ n10825 ^ 1'b0 ;
  assign n31668 = n23887 | n31667 ;
  assign n31669 = ( n7088 & n21756 ) | ( n7088 & n31168 ) | ( n21756 & n31168 ) ;
  assign n31670 = n4467 ^ n1002 ^ 1'b0 ;
  assign n31671 = ( n19499 & n27166 ) | ( n19499 & ~n31670 ) | ( n27166 & ~n31670 ) ;
  assign n31672 = ( n26206 & ~n29325 ) | ( n26206 & n31671 ) | ( ~n29325 & n31671 ) ;
  assign n31673 = n16280 ^ n5177 ^ n3821 ;
  assign n31674 = n31673 ^ n8346 ^ 1'b0 ;
  assign n31675 = n28632 ^ n6402 ^ 1'b0 ;
  assign n31676 = n31675 ^ n29957 ^ 1'b0 ;
  assign n31677 = n2313 & n10832 ;
  assign n31678 = n13273 ^ n970 ^ 1'b0 ;
  assign n31679 = n27035 | n31678 ;
  assign n31680 = n1495 & ~n7805 ;
  assign n31684 = n3917 & n9163 ;
  assign n31685 = n31684 ^ n17233 ^ n13933 ;
  assign n31686 = n31685 ^ n17821 ^ 1'b0 ;
  assign n31687 = n25943 & n31686 ;
  assign n31681 = n28567 ^ n27166 ^ n23808 ;
  assign n31682 = n31681 ^ n14353 ^ n2907 ;
  assign n31683 = n28018 & ~n31682 ;
  assign n31688 = n31687 ^ n31683 ^ 1'b0 ;
  assign n31689 = n31688 ^ n15477 ^ n2210 ;
  assign n31690 = n21567 ^ n20566 ^ n8609 ;
  assign n31691 = n10471 | n23274 ;
  assign n31692 = n1055 | n7137 ;
  assign n31693 = n26665 | n31692 ;
  assign n31694 = n31693 ^ n14677 ^ 1'b0 ;
  assign n31695 = ~n1382 & n5118 ;
  assign n31696 = n31695 ^ n8314 ^ 1'b0 ;
  assign n31697 = n3692 | n31696 ;
  assign n31698 = n9516 & ~n31697 ;
  assign n31699 = n3492 & ~n31698 ;
  assign n31700 = n13498 & n31699 ;
  assign n31701 = n31700 ^ n14335 ^ n11504 ;
  assign n31702 = ( n30202 & n31694 ) | ( n30202 & n31701 ) | ( n31694 & n31701 ) ;
  assign n31703 = n31702 ^ n27509 ^ 1'b0 ;
  assign n31704 = ~n26650 & n31703 ;
  assign n31705 = n10120 & ~n18524 ;
  assign n31706 = n25237 ^ n6344 ^ 1'b0 ;
  assign n31707 = n25687 ^ n6241 ^ n3532 ;
  assign n31708 = n1688 & ~n15186 ;
  assign n31709 = n15096 & n31708 ;
  assign n31710 = n17306 | n18865 ;
  assign n31711 = n8457 & ~n31710 ;
  assign n31712 = n31709 & n31711 ;
  assign n31713 = n17221 | n31712 ;
  assign n31714 = n31707 | n31713 ;
  assign n31715 = n17614 ^ n6861 ^ 1'b0 ;
  assign n31716 = n31715 ^ n29206 ^ n6398 ;
  assign n31717 = n1545 | n6962 ;
  assign n31718 = n19268 ^ n14217 ^ 1'b0 ;
  assign n31719 = n23820 | n31718 ;
  assign n31720 = n22960 & ~n31719 ;
  assign n31721 = ~x172 & n31720 ;
  assign n31723 = n7851 & ~n8311 ;
  assign n31724 = n25891 & ~n31723 ;
  assign n31722 = n19503 & ~n21142 ;
  assign n31725 = n31724 ^ n31722 ^ 1'b0 ;
  assign n31726 = ( n22047 & n24566 ) | ( n22047 & n30382 ) | ( n24566 & n30382 ) ;
  assign n31727 = n7402 ^ n7315 ^ 1'b0 ;
  assign n31728 = n13380 ^ n1702 ^ 1'b0 ;
  assign n31729 = x157 | n31728 ;
  assign n31730 = x46 & ~n31729 ;
  assign n31731 = n25630 & n31730 ;
  assign n31732 = n16686 ^ n13898 ^ 1'b0 ;
  assign n31733 = n21142 ^ n7611 ^ 1'b0 ;
  assign n31734 = n26078 ^ n8327 ^ 1'b0 ;
  assign n31735 = n8527 & n31734 ;
  assign n31736 = ~n31733 & n31735 ;
  assign n31737 = n10130 & ~n24258 ;
  assign n31738 = ~n27290 & n31737 ;
  assign n31739 = n11953 | n13259 ;
  assign n31740 = n11649 | n12118 ;
  assign n31741 = n31740 ^ n5319 ^ 1'b0 ;
  assign n31742 = n31741 ^ n24164 ^ n7801 ;
  assign n31743 = n9491 ^ n7803 ^ 1'b0 ;
  assign n31744 = n20283 & n31743 ;
  assign n31745 = ( n6776 & n13263 ) | ( n6776 & ~n31744 ) | ( n13263 & ~n31744 ) ;
  assign n31746 = n27449 ^ n536 ^ 1'b0 ;
  assign n31747 = n1996 & n31746 ;
  assign n31748 = n8733 & n31747 ;
  assign n31749 = ~n9255 & n31748 ;
  assign n31750 = n4809 | n5330 ;
  assign n31751 = n31750 ^ n10038 ^ 1'b0 ;
  assign n31752 = n31751 ^ n27206 ^ 1'b0 ;
  assign n31753 = n26633 & ~n31752 ;
  assign n31754 = n18202 ^ n11664 ^ 1'b0 ;
  assign n31755 = n16199 | n31754 ;
  assign n31756 = ( n15026 & n26319 ) | ( n15026 & ~n31755 ) | ( n26319 & ~n31755 ) ;
  assign n31757 = n30452 ^ n25471 ^ n4128 ;
  assign n31761 = n17029 ^ n7769 ^ n7513 ;
  assign n31758 = ~n10405 & n24184 ;
  assign n31759 = ~n27839 & n31758 ;
  assign n31760 = n31759 ^ n26569 ^ 1'b0 ;
  assign n31762 = n31761 ^ n31760 ^ n5535 ;
  assign n31763 = n11781 ^ n6353 ^ 1'b0 ;
  assign n31764 = n4347 & n31763 ;
  assign n31765 = ~n4579 & n7856 ;
  assign n31766 = n31765 ^ n7557 ^ 1'b0 ;
  assign n31767 = ( n12326 & ~n31764 ) | ( n12326 & n31766 ) | ( ~n31764 & n31766 ) ;
  assign n31768 = n31767 ^ n27561 ^ n7904 ;
  assign n31769 = ~n3153 & n13967 ;
  assign n31770 = n31769 ^ n22716 ^ n11741 ;
  assign n31771 = n4598 & n17999 ;
  assign n31772 = n31771 ^ n7669 ^ 1'b0 ;
  assign n31773 = n30946 ^ n17562 ^ 1'b0 ;
  assign n31774 = ~n31772 & n31773 ;
  assign n31775 = n4876 & n7598 ;
  assign n31776 = ( ~n3344 & n10550 ) | ( ~n3344 & n21168 ) | ( n10550 & n21168 ) ;
  assign n31777 = n28412 ^ n6986 ^ n4317 ;
  assign n31778 = n26704 ^ n1453 ^ n952 ;
  assign n31779 = n12722 & n31778 ;
  assign n31780 = n11043 & ~n26370 ;
  assign n31781 = ( n3585 & n6488 ) | ( n3585 & n31780 ) | ( n6488 & n31780 ) ;
  assign n31782 = n12139 | n31781 ;
  assign n31783 = ( ~n15562 & n19356 ) | ( ~n15562 & n31782 ) | ( n19356 & n31782 ) ;
  assign n31784 = n31779 & n31783 ;
  assign n31785 = n15085 & ~n19391 ;
  assign n31786 = ~n15703 & n26431 ;
  assign n31787 = n31786 ^ n10555 ^ 1'b0 ;
  assign n31788 = n4162 | n7062 ;
  assign n31789 = n31788 ^ n27147 ^ 1'b0 ;
  assign n31790 = ~n22538 & n31462 ;
  assign n31791 = n30156 & n31790 ;
  assign n31792 = ( n16895 & n31789 ) | ( n16895 & ~n31791 ) | ( n31789 & ~n31791 ) ;
  assign n31793 = n26808 ^ n25618 ^ n6184 ;
  assign n31794 = n31793 ^ n8167 ^ 1'b0 ;
  assign n31795 = n5670 | n14756 ;
  assign n31796 = n2660 & ~n31795 ;
  assign n31797 = n4052 & n31796 ;
  assign n31798 = ( ~n27068 & n31794 ) | ( ~n27068 & n31797 ) | ( n31794 & n31797 ) ;
  assign n31800 = n1786 | n8869 ;
  assign n31801 = n6305 | n31800 ;
  assign n31802 = n31801 ^ n30970 ^ n23240 ;
  assign n31803 = n18405 | n31802 ;
  assign n31799 = n15827 | n28531 ;
  assign n31804 = n31803 ^ n31799 ^ 1'b0 ;
  assign n31805 = n25383 ^ n22783 ^ 1'b0 ;
  assign n31806 = n10165 & ~n31805 ;
  assign n31807 = ~n2931 & n31806 ;
  assign n31808 = n9421 & n31807 ;
  assign n31809 = n15838 ^ x24 ^ 1'b0 ;
  assign n31810 = n19865 ^ n7810 ^ 1'b0 ;
  assign n31811 = n1325 & n31810 ;
  assign n31812 = n11457 ^ n4723 ^ 1'b0 ;
  assign n31813 = ~n3581 & n31812 ;
  assign n31814 = ~n16800 & n31813 ;
  assign n31815 = n13662 ^ n5771 ^ 1'b0 ;
  assign n31816 = n19886 ^ n5042 ^ 1'b0 ;
  assign n31817 = ( ~n6348 & n9759 ) | ( ~n6348 & n12027 ) | ( n9759 & n12027 ) ;
  assign n31818 = ( n7599 & n10960 ) | ( n7599 & n31817 ) | ( n10960 & n31817 ) ;
  assign n31819 = n31818 ^ n31550 ^ 1'b0 ;
  assign n31820 = ( n797 & ~n10072 ) | ( n797 & n10953 ) | ( ~n10072 & n10953 ) ;
  assign n31821 = n8161 & n26301 ;
  assign n31822 = n31820 & n31821 ;
  assign n31823 = n5593 & n9522 ;
  assign n31824 = n2085 | n17672 ;
  assign n31825 = n21380 ^ n10373 ^ 1'b0 ;
  assign n31826 = ~n31824 & n31825 ;
  assign n31827 = n13962 & n31826 ;
  assign n31828 = ~n15110 & n20617 ;
  assign n31829 = n18217 ^ n6732 ^ n515 ;
  assign n31830 = n13066 ^ n6754 ^ 1'b0 ;
  assign n31831 = n31829 & n31830 ;
  assign n31832 = n1680 ^ n1241 ^ 1'b0 ;
  assign n31833 = n31831 & n31832 ;
  assign n31834 = ( ~n14960 & n21542 ) | ( ~n14960 & n31833 ) | ( n21542 & n31833 ) ;
  assign n31835 = n5139 ^ n302 ^ 1'b0 ;
  assign n31836 = n11245 ^ n10164 ^ 1'b0 ;
  assign n31837 = n4079 & ~n31836 ;
  assign n31838 = n19303 & n31837 ;
  assign n31839 = n17450 | n26628 ;
  assign n31840 = n31838 | n31839 ;
  assign n31841 = n19206 & ~n20230 ;
  assign n31842 = ( n4373 & ~n18830 ) | ( n4373 & n31486 ) | ( ~n18830 & n31486 ) ;
  assign n31843 = n18971 ^ n5911 ^ 1'b0 ;
  assign n31844 = n19364 | n31843 ;
  assign n31845 = n31844 ^ n10830 ^ n8248 ;
  assign n31846 = n24085 | n25117 ;
  assign n31847 = n12082 & n30385 ;
  assign n31848 = n18732 ^ n7285 ^ 1'b0 ;
  assign n31849 = n9351 | n31848 ;
  assign n31850 = n15722 | n26641 ;
  assign n31851 = n31849 & ~n31850 ;
  assign n31852 = n16547 ^ n13662 ^ n6351 ;
  assign n31853 = n4435 & ~n27176 ;
  assign n31854 = ( n6682 & n31852 ) | ( n6682 & ~n31853 ) | ( n31852 & ~n31853 ) ;
  assign n31855 = n11634 & ~n15927 ;
  assign n31856 = n31855 ^ n15839 ^ 1'b0 ;
  assign n31858 = n16001 ^ n15357 ^ n3188 ;
  assign n31857 = n3085 & n21018 ;
  assign n31859 = n31858 ^ n31857 ^ 1'b0 ;
  assign n31860 = n31859 ^ n23423 ^ 1'b0 ;
  assign n31862 = n11778 ^ n3990 ^ 1'b0 ;
  assign n31863 = n27879 | n31862 ;
  assign n31861 = n11651 & n17516 ;
  assign n31864 = n31863 ^ n31861 ^ 1'b0 ;
  assign n31865 = n16827 & n27050 ;
  assign n31866 = ~n31864 & n31865 ;
  assign n31867 = n18496 ^ n14234 ^ x193 ;
  assign n31868 = n30249 ^ n7780 ^ 1'b0 ;
  assign n31869 = ~n5789 & n31868 ;
  assign n31870 = n15169 & n17924 ;
  assign n31871 = ~n15502 & n31870 ;
  assign n31872 = n3237 & ~n12664 ;
  assign n31873 = n28243 & n31872 ;
  assign n31874 = n14439 ^ n7163 ^ 1'b0 ;
  assign n31875 = n2580 | n31874 ;
  assign n31876 = n2493 & n27612 ;
  assign n31877 = n10497 ^ n3732 ^ n2197 ;
  assign n31878 = ~n2223 & n31877 ;
  assign n31879 = ~n5956 & n31878 ;
  assign n31880 = ~x144 & n2469 ;
  assign n31881 = n22309 & n31880 ;
  assign n31882 = n7484 | n8465 ;
  assign n31883 = n813 & ~n31882 ;
  assign n31884 = n31883 ^ n12021 ^ 1'b0 ;
  assign n31885 = ~n3281 & n31884 ;
  assign n31886 = ~n12049 & n12145 ;
  assign n31887 = n31886 ^ n22903 ^ 1'b0 ;
  assign n31888 = n30019 ^ n15965 ^ 1'b0 ;
  assign n31889 = n31888 ^ n12207 ^ 1'b0 ;
  assign n31890 = ~n2842 & n9430 ;
  assign n31891 = n28937 ^ n23784 ^ n518 ;
  assign n31892 = n2236 & n6011 ;
  assign n31893 = n11652 & ~n31892 ;
  assign n31894 = n24927 ^ n16337 ^ n1318 ;
  assign n31895 = n28191 ^ n22796 ^ 1'b0 ;
  assign n31897 = n8420 | n12062 ;
  assign n31896 = n27426 | n29740 ;
  assign n31898 = n31897 ^ n31896 ^ 1'b0 ;
  assign n31899 = n31072 ^ n18468 ^ n8387 ;
  assign n31900 = n9711 & ~n31899 ;
  assign n31901 = n31900 ^ n14230 ^ 1'b0 ;
  assign n31902 = n28676 ^ n17341 ^ x21 ;
  assign n31903 = n31783 ^ n31670 ^ n26575 ;
  assign n31904 = ~n6698 & n10244 ;
  assign n31905 = n31904 ^ n4223 ^ 1'b0 ;
  assign n31906 = ~n25249 & n31905 ;
  assign n31907 = n18334 ^ n3932 ^ 1'b0 ;
  assign n31908 = n26712 ^ n1882 ^ 1'b0 ;
  assign n31909 = n31907 | n31908 ;
  assign n31910 = n15732 | n23447 ;
  assign n31911 = n26564 ^ n19742 ^ 1'b0 ;
  assign n31913 = n19534 ^ n17519 ^ 1'b0 ;
  assign n31912 = ( n19766 & n25270 ) | ( n19766 & n27573 ) | ( n25270 & n27573 ) ;
  assign n31914 = n31913 ^ n31912 ^ n22678 ;
  assign n31915 = n2746 & n23766 ;
  assign n31916 = n31915 ^ n29125 ^ 1'b0 ;
  assign n31917 = ( x87 & n3737 ) | ( x87 & n31916 ) | ( n3737 & n31916 ) ;
  assign n31918 = n2506 | n3277 ;
  assign n31919 = n21888 ^ n2386 ^ 1'b0 ;
  assign n31920 = n31918 & n31919 ;
  assign n31921 = n19865 ^ n18483 ^ 1'b0 ;
  assign n31922 = ( n10764 & n13026 ) | ( n10764 & ~n14150 ) | ( n13026 & ~n14150 ) ;
  assign n31923 = n7210 & ~n18637 ;
  assign n31924 = n27935 & n31923 ;
  assign n31925 = n4449 & ~n10320 ;
  assign n31926 = n14416 ^ n14128 ^ n8384 ;
  assign n31927 = n31926 ^ n1807 ^ 1'b0 ;
  assign n31928 = n31925 | n31927 ;
  assign n31929 = n31924 & ~n31928 ;
  assign n31930 = n6971 | n31929 ;
  assign n31931 = n31922 | n31930 ;
  assign n31932 = n21100 ^ n15509 ^ n7475 ;
  assign n31933 = n31932 ^ n28722 ^ n2133 ;
  assign n31934 = n18390 ^ n16363 ^ 1'b0 ;
  assign n31935 = n6512 | n24038 ;
  assign n31936 = n10863 ^ x158 ^ 1'b0 ;
  assign n31937 = n1754 & ~n31936 ;
  assign n31938 = n31937 ^ n29559 ^ n20115 ;
  assign n31939 = ( n1120 & ~n9925 ) | ( n1120 & n29956 ) | ( ~n9925 & n29956 ) ;
  assign n31940 = n31939 ^ n23222 ^ 1'b0 ;
  assign n31941 = ~n4419 & n31940 ;
  assign n31942 = ( ~n6580 & n12198 ) | ( ~n6580 & n31941 ) | ( n12198 & n31941 ) ;
  assign n31943 = n6268 & n7322 ;
  assign n31944 = n4280 & ~n24219 ;
  assign n31945 = ~n16012 & n31944 ;
  assign n31946 = n12443 ^ n5544 ^ 1'b0 ;
  assign n31947 = n29712 ^ n15729 ^ 1'b0 ;
  assign n31948 = n31946 | n31947 ;
  assign n31949 = n18386 ^ n4699 ^ 1'b0 ;
  assign n31950 = n29700 ^ n9563 ^ 1'b0 ;
  assign n31951 = n31949 & n31950 ;
  assign n31952 = n31951 ^ n21093 ^ n14212 ;
  assign n31953 = ( ~n483 & n1579 ) | ( ~n483 & n30119 ) | ( n1579 & n30119 ) ;
  assign n31954 = n31953 ^ n31618 ^ n27130 ;
  assign n31955 = n2983 & ~n14984 ;
  assign n31956 = ~n7504 & n31955 ;
  assign n31957 = ~n2799 & n14947 ;
  assign n31958 = n31957 ^ n2405 ^ 1'b0 ;
  assign n31959 = ( n18880 & n31956 ) | ( n18880 & ~n31958 ) | ( n31956 & ~n31958 ) ;
  assign n31960 = n18896 | n19701 ;
  assign n31961 = n15515 ^ n6597 ^ 1'b0 ;
  assign n31962 = n21624 & ~n31961 ;
  assign n31963 = n8815 & n31962 ;
  assign n31964 = n30627 ^ n6118 ^ 1'b0 ;
  assign n31965 = n22209 ^ n8492 ^ n5842 ;
  assign n31966 = n2774 & n2899 ;
  assign n31967 = n5426 & n31966 ;
  assign n31968 = n31965 & ~n31967 ;
  assign n31969 = n31968 ^ n4480 ^ 1'b0 ;
  assign n31970 = n21583 ^ n17504 ^ n3796 ;
  assign n31971 = n31970 ^ n8683 ^ 1'b0 ;
  assign n31972 = n19531 ^ n9303 ^ n2588 ;
  assign n31973 = n15316 ^ n10095 ^ 1'b0 ;
  assign n31974 = n31973 ^ n18374 ^ 1'b0 ;
  assign n31975 = ~n31972 & n31974 ;
  assign n31976 = ( n7649 & ~n28813 ) | ( n7649 & n31975 ) | ( ~n28813 & n31975 ) ;
  assign n31977 = n23636 & n24161 ;
  assign n31978 = ( ~n5203 & n8942 ) | ( ~n5203 & n31977 ) | ( n8942 & n31977 ) ;
  assign n31979 = n11113 | n14230 ;
  assign n31980 = n12852 | n31979 ;
  assign n31981 = ~n3095 & n31980 ;
  assign n31982 = ~n2722 & n5800 ;
  assign n31983 = n31982 ^ n11211 ^ 1'b0 ;
  assign n31984 = n14762 | n31983 ;
  assign n31985 = ( ~n3440 & n11022 ) | ( ~n3440 & n15428 ) | ( n11022 & n15428 ) ;
  assign n31986 = n7430 | n31985 ;
  assign n31987 = n24025 & n25099 ;
  assign n31989 = n7055 | n13994 ;
  assign n31988 = n15073 & n16277 ;
  assign n31990 = n31989 ^ n31988 ^ 1'b0 ;
  assign n31991 = n13451 ^ n9251 ^ 1'b0 ;
  assign n31992 = ~n11450 & n31991 ;
  assign n31993 = n31992 ^ n6616 ^ n4355 ;
  assign n31994 = ~n260 & n6010 ;
  assign n31995 = n31993 & n31994 ;
  assign n31996 = n28416 | n31995 ;
  assign n31997 = n11992 ^ n1500 ^ 1'b0 ;
  assign n31998 = n17881 ^ n3274 ^ 1'b0 ;
  assign n31999 = n16261 ^ n7561 ^ 1'b0 ;
  assign n32000 = n6445 & n31999 ;
  assign n32001 = n32000 ^ n8222 ^ 1'b0 ;
  assign n32002 = ( n2616 & n8447 ) | ( n2616 & ~n20098 ) | ( n8447 & ~n20098 ) ;
  assign n32008 = n15671 ^ n10744 ^ n1329 ;
  assign n32009 = ( n24397 & n30926 ) | ( n24397 & n32008 ) | ( n30926 & n32008 ) ;
  assign n32004 = n10315 ^ n3430 ^ 1'b0 ;
  assign n32005 = n3949 | n13058 ;
  assign n32006 = n32005 ^ n26317 ^ 1'b0 ;
  assign n32007 = n32004 & ~n32006 ;
  assign n32010 = n32009 ^ n32007 ^ n4055 ;
  assign n32003 = n7057 | n20093 ;
  assign n32011 = n32010 ^ n32003 ^ 1'b0 ;
  assign n32012 = n21251 ^ n20949 ^ 1'b0 ;
  assign n32013 = n32012 ^ n3696 ^ n1899 ;
  assign n32014 = n8315 ^ x60 ^ 1'b0 ;
  assign n32015 = ( n4189 & n7145 ) | ( n4189 & n10317 ) | ( n7145 & n10317 ) ;
  assign n32016 = n17061 & ~n32015 ;
  assign n32020 = n14443 | n17363 ;
  assign n32017 = ~n11655 & n14587 ;
  assign n32018 = n32017 ^ n14989 ^ 1'b0 ;
  assign n32019 = n15976 | n32018 ;
  assign n32021 = n32020 ^ n32019 ^ 1'b0 ;
  assign n32022 = n7521 ^ n673 ^ 1'b0 ;
  assign n32023 = n14239 & ~n29386 ;
  assign n32024 = ( n11581 & n32022 ) | ( n11581 & ~n32023 ) | ( n32022 & ~n32023 ) ;
  assign n32025 = ~n12035 & n32024 ;
  assign n32026 = n32025 ^ n12972 ^ n5323 ;
  assign n32027 = n26637 ^ n13079 ^ n4884 ;
  assign n32028 = n6989 | n32027 ;
  assign n32029 = n32028 ^ x116 ^ 1'b0 ;
  assign n32030 = n7055 | n16964 ;
  assign n32031 = n32030 ^ n8160 ^ 1'b0 ;
  assign n32032 = n32031 ^ n10451 ^ n10255 ;
  assign n32033 = ( n8735 & ~n32029 ) | ( n8735 & n32032 ) | ( ~n32029 & n32032 ) ;
  assign n32034 = n31198 ^ n2700 ^ 1'b0 ;
  assign n32035 = n3957 ^ n3386 ^ 1'b0 ;
  assign n32037 = n1444 ^ x176 ^ 1'b0 ;
  assign n32038 = n6640 & n32037 ;
  assign n32036 = ~n13099 & n31486 ;
  assign n32039 = n32038 ^ n32036 ^ 1'b0 ;
  assign n32040 = n2136 & n6938 ;
  assign n32041 = ~n19819 & n32040 ;
  assign n32042 = ( ~n27573 & n28072 ) | ( ~n27573 & n32041 ) | ( n28072 & n32041 ) ;
  assign n32043 = n10245 ^ n3889 ^ 1'b0 ;
  assign n32044 = n6296 | n32043 ;
  assign n32045 = n19328 | n32044 ;
  assign n32046 = n10662 ^ n2937 ^ 1'b0 ;
  assign n32047 = n28308 & n32046 ;
  assign n32048 = n398 | n21493 ;
  assign n32049 = n20643 & ~n32048 ;
  assign n32050 = n19518 ^ x31 ^ 1'b0 ;
  assign n32051 = n32049 | n32050 ;
  assign n32052 = n31349 ^ n3896 ^ 1'b0 ;
  assign n32053 = n18837 & n18844 ;
  assign n32054 = n9336 & ~n11652 ;
  assign n32055 = x247 & n2313 ;
  assign n32056 = n32055 ^ n15359 ^ n13278 ;
  assign n32057 = n30630 ^ n8685 ^ 1'b0 ;
  assign n32058 = n28824 ^ n25071 ^ n19078 ;
  assign n32059 = n21848 ^ n14412 ^ 1'b0 ;
  assign n32060 = n2958 ^ n335 ^ 1'b0 ;
  assign n32061 = n7512 | n8045 ;
  assign n32062 = n32061 ^ n17535 ^ 1'b0 ;
  assign n32063 = ~n10709 & n11066 ;
  assign n32064 = n32063 ^ n22410 ^ 1'b0 ;
  assign n32065 = n32062 & n32064 ;
  assign n32066 = n26224 ^ n18470 ^ n15861 ;
  assign n32067 = n6448 | n19154 ;
  assign n32068 = n16679 & ~n32067 ;
  assign n32069 = n32068 ^ n30367 ^ n22296 ;
  assign n32070 = n2313 & ~n3239 ;
  assign n32071 = n32070 ^ n9586 ^ 1'b0 ;
  assign n32072 = n3178 & n32071 ;
  assign n32073 = ~n9852 & n13493 ;
  assign n32074 = n32073 ^ n658 ^ 1'b0 ;
  assign n32075 = n7741 | n8024 ;
  assign n32076 = n3564 | n12644 ;
  assign n32080 = n12929 ^ n8761 ^ 1'b0 ;
  assign n32081 = n32080 ^ n31185 ^ n7986 ;
  assign n32077 = ~n20991 & n30867 ;
  assign n32078 = n1596 & n32077 ;
  assign n32079 = n32078 ^ n23845 ^ 1'b0 ;
  assign n32082 = n32081 ^ n32079 ^ n5722 ;
  assign n32083 = ~n14800 & n21527 ;
  assign n32084 = ~n12239 & n32083 ;
  assign n32085 = n32084 ^ n12854 ^ 1'b0 ;
  assign n32086 = n31783 & n32085 ;
  assign n32087 = n2268 & n6256 ;
  assign n32088 = n3821 | n12686 ;
  assign n32089 = n32088 ^ n26244 ^ 1'b0 ;
  assign n32090 = n32089 ^ n29432 ^ n4226 ;
  assign n32091 = n11837 ^ n873 ^ 1'b0 ;
  assign n32092 = n5803 & ~n32091 ;
  assign n32093 = n3667 & n20801 ;
  assign n32094 = n13680 & n32093 ;
  assign n32095 = n1707 ^ x24 ^ 1'b0 ;
  assign n32096 = n32095 ^ n14486 ^ 1'b0 ;
  assign n32097 = n32094 | n32096 ;
  assign n32098 = ( n18011 & ~n32092 ) | ( n18011 & n32097 ) | ( ~n32092 & n32097 ) ;
  assign n32099 = n1859 | n12118 ;
  assign n32100 = n27655 & ~n32099 ;
  assign n32101 = ~n18377 & n32100 ;
  assign n32102 = n17697 & n26828 ;
  assign n32103 = n32102 ^ n7880 ^ 1'b0 ;
  assign n32105 = n4090 ^ n3821 ^ 1'b0 ;
  assign n32104 = ~n9949 & n16394 ;
  assign n32106 = n32105 ^ n32104 ^ 1'b0 ;
  assign n32107 = ( n1553 & n2903 ) | ( n1553 & n5335 ) | ( n2903 & n5335 ) ;
  assign n32108 = n30836 & n32107 ;
  assign n32109 = x222 & ~n1722 ;
  assign n32110 = n22856 ^ n19261 ^ n9347 ;
  assign n32111 = n22631 | n26348 ;
  assign n32112 = n32111 ^ n27520 ^ n24767 ;
  assign n32113 = n17668 & ~n32112 ;
  assign n32114 = ( ~n10072 & n18160 ) | ( ~n10072 & n31554 ) | ( n18160 & n31554 ) ;
  assign n32115 = n7780 & ~n26522 ;
  assign n32116 = n19765 ^ n6094 ^ 1'b0 ;
  assign n32117 = n23130 & ~n32116 ;
  assign n32118 = n17431 & n32117 ;
  assign n32119 = ~n4468 & n8481 ;
  assign n32120 = n32119 ^ n10221 ^ 1'b0 ;
  assign n32121 = ( n11666 & n13148 ) | ( n11666 & n20727 ) | ( n13148 & n20727 ) ;
  assign n32122 = n9457 & ~n32121 ;
  assign n32123 = n18801 & n32122 ;
  assign n32124 = ~n32120 & n32123 ;
  assign n32125 = n25006 ^ n932 ^ 1'b0 ;
  assign n32126 = ~n22150 & n32125 ;
  assign n32127 = n32126 ^ n10726 ^ 1'b0 ;
  assign n32128 = n1605 & ~n4490 ;
  assign n32129 = n29329 ^ n24055 ^ 1'b0 ;
  assign n32130 = n32128 & ~n32129 ;
  assign n32131 = n28617 ^ n9013 ^ 1'b0 ;
  assign n32132 = ~n9702 & n32131 ;
  assign n32133 = n24438 ^ n10229 ^ n3402 ;
  assign n32134 = n15539 & ~n32133 ;
  assign n32135 = ~n32132 & n32134 ;
  assign n32136 = n32135 ^ n28455 ^ 1'b0 ;
  assign n32140 = ~n19328 & n19646 ;
  assign n32141 = n15040 & n32140 ;
  assign n32142 = n2422 & ~n26949 ;
  assign n32143 = n32141 & ~n32142 ;
  assign n32137 = ~n3583 & n9164 ;
  assign n32138 = ~n28635 & n32137 ;
  assign n32139 = ~n7089 & n32138 ;
  assign n32144 = n32143 ^ n32139 ^ n7186 ;
  assign n32145 = n1838 & n22440 ;
  assign n32146 = n32145 ^ n11721 ^ 1'b0 ;
  assign n32147 = n27737 ^ n12916 ^ n11015 ;
  assign n32148 = n10112 ^ n2536 ^ 1'b0 ;
  assign n32149 = n10259 ^ n8314 ^ 1'b0 ;
  assign n32150 = ( n7260 & n8794 ) | ( n7260 & n17076 ) | ( n8794 & n17076 ) ;
  assign n32151 = n32150 ^ n3781 ^ 1'b0 ;
  assign n32152 = n32149 | n32151 ;
  assign n32153 = n12837 & ~n23202 ;
  assign n32154 = n1789 | n13698 ;
  assign n32155 = n32154 ^ n1604 ^ n678 ;
  assign n32156 = n32155 ^ n22199 ^ 1'b0 ;
  assign n32157 = n5618 | n19191 ;
  assign n32158 = n16062 ^ n14397 ^ n3471 ;
  assign n32159 = n32158 ^ n29236 ^ n1291 ;
  assign n32160 = n633 & ~n3172 ;
  assign n32161 = n8794 | n23720 ;
  assign n32162 = n5149 | n32161 ;
  assign n32163 = n2927 & n11381 ;
  assign n32164 = ~n13916 & n32163 ;
  assign n32165 = n25021 ^ n24090 ^ 1'b0 ;
  assign n32171 = n12726 & ~n16923 ;
  assign n32166 = n8696 & n10498 ;
  assign n32167 = n8578 ^ n3483 ^ 1'b0 ;
  assign n32168 = ( ~n16075 & n25911 ) | ( ~n16075 & n32167 ) | ( n25911 & n32167 ) ;
  assign n32169 = ~n26403 & n32168 ;
  assign n32170 = n32166 & n32169 ;
  assign n32172 = n32171 ^ n32170 ^ n17554 ;
  assign n32173 = ~n10778 & n12678 ;
  assign n32174 = n13187 ^ n7486 ^ 1'b0 ;
  assign n32175 = ( n8640 & n9326 ) | ( n8640 & n15029 ) | ( n9326 & n15029 ) ;
  assign n32176 = n32175 ^ n16462 ^ n4809 ;
  assign n32177 = n22502 & ~n32176 ;
  assign n32178 = n32177 ^ n21716 ^ 1'b0 ;
  assign n32179 = n12126 ^ n11888 ^ 1'b0 ;
  assign n32180 = n18138 ^ n1641 ^ n710 ;
  assign n32181 = ~n7009 & n18481 ;
  assign n32182 = n30609 ^ n4869 ^ n787 ;
  assign n32183 = n32182 ^ n15518 ^ 1'b0 ;
  assign n32184 = n32183 ^ n30814 ^ n19804 ;
  assign n32185 = ( n16474 & n27629 ) | ( n16474 & ~n30700 ) | ( n27629 & ~n30700 ) ;
  assign n32186 = n7015 & ~n11447 ;
  assign n32187 = ( n2889 & ~n11551 ) | ( n2889 & n12674 ) | ( ~n11551 & n12674 ) ;
  assign n32188 = ~n2295 & n32187 ;
  assign n32189 = n6370 & n32188 ;
  assign n32190 = n14076 ^ n12287 ^ n5090 ;
  assign n32191 = n32190 ^ n9724 ^ 1'b0 ;
  assign n32192 = n3389 | n32191 ;
  assign n32193 = n15778 & n26567 ;
  assign n32194 = n32193 ^ n945 ^ 1'b0 ;
  assign n32195 = ~n30518 & n32194 ;
  assign n32196 = n9998 | n24511 ;
  assign n32197 = n32196 ^ n22021 ^ 1'b0 ;
  assign n32200 = n7963 & ~n26137 ;
  assign n32198 = n28357 ^ n11445 ^ 1'b0 ;
  assign n32199 = n11393 | n32198 ;
  assign n32201 = n32200 ^ n32199 ^ 1'b0 ;
  assign n32202 = ( n11240 & n13925 ) | ( n11240 & n22755 ) | ( n13925 & n22755 ) ;
  assign n32203 = n1110 | n26386 ;
  assign n32204 = n32203 ^ n29521 ^ 1'b0 ;
  assign n32205 = n32204 ^ n23724 ^ 1'b0 ;
  assign n32206 = n21981 ^ n20418 ^ 1'b0 ;
  assign n32207 = n23991 ^ n932 ^ 1'b0 ;
  assign n32208 = n32207 ^ n30850 ^ 1'b0 ;
  assign n32209 = n23567 ^ n3037 ^ 1'b0 ;
  assign n32210 = n26887 ^ n3773 ^ 1'b0 ;
  assign n32211 = n32209 | n32210 ;
  assign n32212 = n21337 ^ n18753 ^ n9631 ;
  assign n32213 = n21663 & n32212 ;
  assign n32214 = ( n13320 & n23897 ) | ( n13320 & n32213 ) | ( n23897 & n32213 ) ;
  assign n32215 = ( n5429 & n6018 ) | ( n5429 & ~n20429 ) | ( n6018 & ~n20429 ) ;
  assign n32216 = n2435 | n5935 ;
  assign n32217 = n9058 & ~n16286 ;
  assign n32218 = ( n10667 & ~n22190 ) | ( n10667 & n32217 ) | ( ~n22190 & n32217 ) ;
  assign n32219 = n6062 & n32218 ;
  assign n32220 = n32216 & n32219 ;
  assign n32221 = n3100 & n3144 ;
  assign n32222 = n32221 ^ n3335 ^ 1'b0 ;
  assign n32223 = ( n1247 & n18008 ) | ( n1247 & ~n32222 ) | ( n18008 & ~n32222 ) ;
  assign n32224 = n27153 | n32223 ;
  assign n32225 = n2055 & ~n25354 ;
  assign n32226 = ( n4159 & n5646 ) | ( n4159 & ~n8129 ) | ( n5646 & ~n8129 ) ;
  assign n32227 = n32226 ^ n26181 ^ 1'b0 ;
  assign n32228 = n32227 ^ n1729 ^ 1'b0 ;
  assign n32229 = n8393 & ~n12010 ;
  assign n32230 = n2919 ^ n1452 ^ n837 ;
  assign n32231 = n32230 ^ n21926 ^ n1647 ;
  assign n32232 = n25680 ^ n19553 ^ n8020 ;
  assign n32233 = ~n2212 & n4711 ;
  assign n32234 = ( ~n10314 & n15383 ) | ( ~n10314 & n32233 ) | ( n15383 & n32233 ) ;
  assign n32235 = ( n11270 & ~n19490 ) | ( n11270 & n32234 ) | ( ~n19490 & n32234 ) ;
  assign n32236 = n6413 & ~n15859 ;
  assign n32237 = ~n23845 & n32236 ;
  assign n32238 = ~n14920 & n17902 ;
  assign n32239 = n32237 & n32238 ;
  assign n32240 = n2344 | n32239 ;
  assign n32241 = n32235 | n32240 ;
  assign n32242 = n5575 & n19197 ;
  assign n32243 = n3883 | n12768 ;
  assign n32244 = n32243 ^ n27166 ^ 1'b0 ;
  assign n32245 = n10094 & n22361 ;
  assign n32246 = n14805 & n32245 ;
  assign n32247 = ( ~n1028 & n23769 ) | ( ~n1028 & n32246 ) | ( n23769 & n32246 ) ;
  assign n32248 = n15986 ^ n15938 ^ 1'b0 ;
  assign n32249 = n14528 & ~n32248 ;
  assign n32250 = ( ~n12291 & n16613 ) | ( ~n12291 & n32249 ) | ( n16613 & n32249 ) ;
  assign n32251 = n6306 | n15813 ;
  assign n32252 = n32251 ^ n18683 ^ 1'b0 ;
  assign n32253 = n10181 ^ n8507 ^ x167 ;
  assign n32254 = ~n31101 & n32253 ;
  assign n32255 = n1327 & ~n32254 ;
  assign n32256 = n17661 | n27861 ;
  assign n32257 = n2119 & n5311 ;
  assign n32258 = ( ~n12788 & n14172 ) | ( ~n12788 & n19321 ) | ( n14172 & n19321 ) ;
  assign n32259 = n22152 & ~n28554 ;
  assign n32260 = ~n32258 & n32259 ;
  assign n32261 = n22484 ^ n6457 ^ 1'b0 ;
  assign n32262 = ~n32260 & n32261 ;
  assign n32263 = ( n5682 & n19507 ) | ( n5682 & n19814 ) | ( n19507 & n19814 ) ;
  assign n32264 = ( n6915 & n25119 ) | ( n6915 & n32263 ) | ( n25119 & n32263 ) ;
  assign n32265 = n16740 ^ n2983 ^ 1'b0 ;
  assign n32266 = n17464 & n32265 ;
  assign n32267 = n32266 ^ n16615 ^ 1'b0 ;
  assign n32268 = n32267 ^ n16020 ^ 1'b0 ;
  assign n32271 = n3073 & ~n6782 ;
  assign n32269 = n7104 & n16417 ;
  assign n32270 = n32269 ^ n31226 ^ 1'b0 ;
  assign n32272 = n32271 ^ n32270 ^ n25674 ;
  assign n32273 = n1294 & n17946 ;
  assign n32274 = ~n14866 & n32273 ;
  assign n32275 = n9587 | n32274 ;
  assign n32276 = n32275 ^ n18403 ^ 1'b0 ;
  assign n32277 = n21346 ^ n8193 ^ 1'b0 ;
  assign n32278 = n32276 & ~n32277 ;
  assign n32279 = n614 & ~n28177 ;
  assign n32280 = ~n4327 & n32279 ;
  assign n32281 = n345 | n18001 ;
  assign n32282 = n14869 | n32281 ;
  assign n32283 = n21508 & ~n21944 ;
  assign n32284 = ( ~n31244 & n32282 ) | ( ~n31244 & n32283 ) | ( n32282 & n32283 ) ;
  assign n32285 = ( n1134 & n23942 ) | ( n1134 & n26908 ) | ( n23942 & n26908 ) ;
  assign n32286 = n3958 ^ n1079 ^ 1'b0 ;
  assign n32287 = n20449 & ~n29231 ;
  assign n32288 = ( ~n1588 & n12708 ) | ( ~n1588 & n15699 ) | ( n12708 & n15699 ) ;
  assign n32289 = n17718 & n32288 ;
  assign n32290 = n12668 ^ n5112 ^ 1'b0 ;
  assign n32291 = n2009 | n9363 ;
  assign n32292 = n32291 ^ n20047 ^ 1'b0 ;
  assign n32293 = n32292 ^ n1034 ^ 1'b0 ;
  assign n32294 = n32290 & ~n32293 ;
  assign n32302 = ( n1673 & ~n5628 ) | ( n1673 & n15287 ) | ( ~n5628 & n15287 ) ;
  assign n32303 = ~n8244 & n20323 ;
  assign n32304 = n32302 & n32303 ;
  assign n32296 = ( n4760 & n6738 ) | ( n4760 & n9421 ) | ( n6738 & n9421 ) ;
  assign n32295 = ~n2154 & n6772 ;
  assign n32297 = n32296 ^ n32295 ^ 1'b0 ;
  assign n32298 = ( n3433 & n14840 ) | ( n3433 & n32297 ) | ( n14840 & n32297 ) ;
  assign n32299 = n10164 & n32298 ;
  assign n32300 = ~n17541 & n32299 ;
  assign n32301 = n26320 | n32300 ;
  assign n32305 = n32304 ^ n32301 ^ 1'b0 ;
  assign n32306 = ~n23191 & n26605 ;
  assign n32308 = n12888 ^ n7812 ^ n3831 ;
  assign n32309 = ( x249 & n28500 ) | ( x249 & ~n32308 ) | ( n28500 & ~n32308 ) ;
  assign n32307 = n451 & ~n14789 ;
  assign n32310 = n32309 ^ n32307 ^ 1'b0 ;
  assign n32311 = n23093 ^ n20618 ^ 1'b0 ;
  assign n32312 = ( n15208 & ~n20544 ) | ( n15208 & n25438 ) | ( ~n20544 & n25438 ) ;
  assign n32313 = n2386 | n12554 ;
  assign n32314 = n11304 | n32313 ;
  assign n32315 = n28269 & n32314 ;
  assign n32316 = n24314 ^ n7862 ^ 1'b0 ;
  assign n32317 = n17129 ^ n12575 ^ 1'b0 ;
  assign n32318 = n7413 | n10971 ;
  assign n32319 = n987 & n15335 ;
  assign n32320 = n32319 ^ n3910 ^ n2390 ;
  assign n32321 = n3133 & ~n7400 ;
  assign n32322 = n19379 | n32321 ;
  assign n32323 = n32322 ^ n25023 ^ 1'b0 ;
  assign n32324 = n3755 & ~n32323 ;
  assign n32325 = n1007 & ~n1611 ;
  assign n32326 = n1611 & n32325 ;
  assign n32327 = n3242 & ~n32326 ;
  assign n32328 = n32326 & n32327 ;
  assign n32329 = n11203 | n32328 ;
  assign n32330 = n10092 & ~n32329 ;
  assign n32331 = n32330 ^ n13744 ^ 1'b0 ;
  assign n32332 = ( x97 & n8323 ) | ( x97 & n21138 ) | ( n8323 & n21138 ) ;
  assign n32333 = n32332 ^ n25654 ^ n8784 ;
  assign n32334 = n7619 & n20588 ;
  assign n32335 = n32334 ^ n19806 ^ 1'b0 ;
  assign n32336 = n11951 ^ n3529 ^ 1'b0 ;
  assign n32337 = n32336 ^ n28317 ^ 1'b0 ;
  assign n32338 = n7912 ^ n6551 ^ 1'b0 ;
  assign n32339 = n15371 & ~n32338 ;
  assign n32340 = ( n1781 & ~n4068 ) | ( n1781 & n14068 ) | ( ~n4068 & n14068 ) ;
  assign n32341 = n3009 | n32340 ;
  assign n32342 = n16209 ^ n14927 ^ 1'b0 ;
  assign n32343 = n32342 ^ n27643 ^ 1'b0 ;
  assign n32344 = n6406 ^ n831 ^ 1'b0 ;
  assign n32345 = n32344 ^ n1031 ^ 1'b0 ;
  assign n32346 = n23470 & n32345 ;
  assign n32347 = ~n29956 & n32346 ;
  assign n32348 = ~n3994 & n32347 ;
  assign n32349 = n729 | n10046 ;
  assign n32350 = n32349 ^ n20749 ^ n14750 ;
  assign n32351 = n8288 & n32350 ;
  assign n32352 = n32351 ^ n9350 ^ 1'b0 ;
  assign n32353 = n19404 ^ n2197 ^ 1'b0 ;
  assign n32354 = n1673 | n9540 ;
  assign n32355 = n15528 & ~n32354 ;
  assign n32356 = n4574 & ~n32355 ;
  assign n32357 = ~n31877 & n32356 ;
  assign n32358 = n1266 & ~n6917 ;
  assign n32359 = n6195 | n21780 ;
  assign n32360 = n32359 ^ x26 ^ 1'b0 ;
  assign n32361 = ~n17325 & n32360 ;
  assign n32362 = n32358 & n32361 ;
  assign n32363 = n21756 ^ n12050 ^ n897 ;
  assign n32364 = n21421 ^ n12147 ^ n1768 ;
  assign n32365 = n32364 ^ n32304 ^ n961 ;
  assign n32366 = n30317 ^ n5263 ^ 1'b0 ;
  assign n32367 = n12532 ^ n11908 ^ 1'b0 ;
  assign n32368 = n18234 & n32367 ;
  assign n32369 = n32368 ^ n17371 ^ 1'b0 ;
  assign n32370 = n2575 & n23915 ;
  assign n32371 = ~n12591 & n32370 ;
  assign n32372 = n6445 & n32314 ;
  assign n32373 = n32372 ^ x183 ^ 1'b0 ;
  assign n32374 = ( ~n11601 & n30103 ) | ( ~n11601 & n32373 ) | ( n30103 & n32373 ) ;
  assign n32375 = n10652 ^ n8609 ^ n4489 ;
  assign n32376 = n6002 ^ n2038 ^ x91 ;
  assign n32377 = n18121 & n32376 ;
  assign n32378 = ~n5445 & n18158 ;
  assign n32379 = ( n32375 & n32377 ) | ( n32375 & ~n32378 ) | ( n32377 & ~n32378 ) ;
  assign n32385 = n764 & ~n9241 ;
  assign n32386 = ~n9635 & n32385 ;
  assign n32384 = n14752 ^ n9835 ^ 1'b0 ;
  assign n32380 = n2912 & ~n21656 ;
  assign n32381 = ~n12116 & n32380 ;
  assign n32382 = n18348 | n32381 ;
  assign n32383 = n1273 & ~n32382 ;
  assign n32387 = n32386 ^ n32384 ^ n32383 ;
  assign n32388 = n1962 | n18850 ;
  assign n32389 = n32388 ^ n8477 ^ 1'b0 ;
  assign n32390 = n28190 ^ n9806 ^ 1'b0 ;
  assign n32392 = n1684 & ~n8046 ;
  assign n32391 = x184 & n4226 ;
  assign n32393 = n32392 ^ n32391 ^ 1'b0 ;
  assign n32394 = n32393 ^ n13967 ^ 1'b0 ;
  assign n32395 = n32390 & n32394 ;
  assign n32396 = n9068 ^ n3523 ^ 1'b0 ;
  assign n32397 = n16981 | n32396 ;
  assign n32398 = n32397 ^ n21151 ^ 1'b0 ;
  assign n32399 = n7384 & ~n32398 ;
  assign n32400 = n32399 ^ x103 ^ 1'b0 ;
  assign n32401 = n1553 & n5394 ;
  assign n32402 = n5447 & n32401 ;
  assign n32403 = n440 | n11661 ;
  assign n32404 = n32403 ^ n7929 ^ 1'b0 ;
  assign n32405 = n32404 ^ n19109 ^ 1'b0 ;
  assign n32410 = ( n2078 & n5054 ) | ( n2078 & ~n8074 ) | ( n5054 & ~n8074 ) ;
  assign n32406 = n14489 ^ n10497 ^ n294 ;
  assign n32407 = n32406 ^ n30038 ^ 1'b0 ;
  assign n32408 = ~n26141 & n32407 ;
  assign n32409 = n32408 ^ n10977 ^ 1'b0 ;
  assign n32411 = n32410 ^ n32409 ^ 1'b0 ;
  assign n32412 = ( n4326 & n5004 ) | ( n4326 & ~n19742 ) | ( n5004 & ~n19742 ) ;
  assign n32413 = n22481 | n32412 ;
  assign n32414 = n20703 | n32413 ;
  assign n32415 = ~n7043 & n16351 ;
  assign n32416 = n1247 & ~n5776 ;
  assign n32417 = n20958 ^ n17367 ^ n4067 ;
  assign n32418 = ( n9586 & n12823 ) | ( n9586 & n32417 ) | ( n12823 & n32417 ) ;
  assign n32419 = n8352 ^ n5905 ^ 1'b0 ;
  assign n32420 = n31981 ^ n9192 ^ 1'b0 ;
  assign n32421 = n10244 ^ n8169 ^ 1'b0 ;
  assign n32422 = ~n31928 & n32421 ;
  assign n32423 = n14041 ^ n2135 ^ 1'b0 ;
  assign n32424 = n10984 & ~n32423 ;
  assign n32425 = n2614 & ~n6376 ;
  assign n32426 = n32425 ^ n12188 ^ n10451 ;
  assign n32427 = n32426 ^ n28866 ^ n22896 ;
  assign n32428 = n6791 & ~n31538 ;
  assign n32429 = n25045 & ~n32428 ;
  assign n32430 = n9937 ^ n2191 ^ n1666 ;
  assign n32431 = n18558 & n27333 ;
  assign n32432 = n2577 & n32431 ;
  assign n32433 = n16267 ^ n8613 ^ 1'b0 ;
  assign n32434 = n32433 ^ n16558 ^ 1'b0 ;
  assign n32435 = n660 & ~n32434 ;
  assign n32436 = n24488 | n29432 ;
  assign n32437 = n471 | n4345 ;
  assign n32438 = n10454 ^ n3014 ^ 1'b0 ;
  assign n32439 = n32437 & n32438 ;
  assign n32440 = ~n15826 & n32439 ;
  assign n32441 = ~n4959 & n32440 ;
  assign n32442 = n32441 ^ n8257 ^ 1'b0 ;
  assign n32443 = ~n21879 & n32442 ;
  assign n32444 = n32443 ^ n10613 ^ 1'b0 ;
  assign n32445 = n1511 & n9021 ;
  assign n32446 = n6669 & n15870 ;
  assign n32447 = ~n32445 & n32446 ;
  assign n32448 = n12709 ^ n2449 ^ 1'b0 ;
  assign n32449 = ( n19213 & ~n21989 ) | ( n19213 & n31978 ) | ( ~n21989 & n31978 ) ;
  assign n32450 = n28444 ^ n9054 ^ 1'b0 ;
  assign n32451 = ~n12118 & n32450 ;
  assign n32452 = n2006 & n6253 ;
  assign n32453 = n32452 ^ n32263 ^ 1'b0 ;
  assign n32454 = ~n7225 & n32453 ;
  assign n32455 = n21364 | n32454 ;
  assign n32456 = ~n9290 & n26097 ;
  assign n32457 = n2980 ^ x196 ^ 1'b0 ;
  assign n32458 = n32456 & ~n32457 ;
  assign n32459 = n593 & ~n9414 ;
  assign n32460 = ~n17853 & n32459 ;
  assign n32461 = n10563 & ~n32460 ;
  assign n32462 = ~n6320 & n6990 ;
  assign n32463 = n21048 ^ n514 ^ 1'b0 ;
  assign n32464 = ( ~n1037 & n32462 ) | ( ~n1037 & n32463 ) | ( n32462 & n32463 ) ;
  assign n32465 = n16301 ^ n6248 ^ 1'b0 ;
  assign n32466 = n18362 & ~n32465 ;
  assign n32467 = n32466 ^ n11844 ^ 1'b0 ;
  assign n32468 = n16400 ^ n13017 ^ n2505 ;
  assign n32469 = ~n8160 & n32468 ;
  assign n32470 = ~n390 & n32469 ;
  assign n32471 = n32470 ^ n16433 ^ 1'b0 ;
  assign n32473 = n5089 & n15494 ;
  assign n32472 = n16907 & n23874 ;
  assign n32474 = n32473 ^ n32472 ^ 1'b0 ;
  assign n32475 = n9063 & n17630 ;
  assign n32476 = n1405 & ~n8676 ;
  assign n32477 = ~n15712 & n32476 ;
  assign n32478 = n32477 ^ n3575 ^ 1'b0 ;
  assign n32479 = n14888 ^ n12105 ^ n2932 ;
  assign n32480 = n3093 & ~n7319 ;
  assign n32481 = n32479 & n32480 ;
  assign n32483 = n12526 ^ n4830 ^ 1'b0 ;
  assign n32484 = ~n12581 & n32483 ;
  assign n32482 = n7189 | n17481 ;
  assign n32485 = n32484 ^ n32482 ^ 1'b0 ;
  assign n32486 = n2691 & n13711 ;
  assign n32487 = n21486 ^ n3053 ^ 1'b0 ;
  assign n32488 = n11966 & n13603 ;
  assign n32489 = ~n32487 & n32488 ;
  assign n32490 = n12794 ^ n5364 ^ 1'b0 ;
  assign n32491 = n11691 & n31231 ;
  assign n32492 = ~n20819 & n32491 ;
  assign n32493 = n2147 & ~n8743 ;
  assign n32494 = n32493 ^ n30587 ^ 1'b0 ;
  assign n32495 = n22325 ^ n10754 ^ n8418 ;
  assign n32496 = ~n857 & n8246 ;
  assign n32497 = n32496 ^ n13326 ^ 1'b0 ;
  assign n32498 = n13885 | n32497 ;
  assign n32499 = ( n424 & ~n7473 ) | ( n424 & n32498 ) | ( ~n7473 & n32498 ) ;
  assign n32500 = n17906 | n32499 ;
  assign n32501 = n9652 | n32500 ;
  assign n32502 = ~n4648 & n18106 ;
  assign n32503 = ( n1476 & ~n4133 ) | ( n1476 & n17429 ) | ( ~n4133 & n17429 ) ;
  assign n32504 = n19669 | n32503 ;
  assign n32505 = n2962 | n32504 ;
  assign n32506 = n8639 & ~n12032 ;
  assign n32507 = n32506 ^ n12929 ^ 1'b0 ;
  assign n32508 = ( n1592 & n15818 ) | ( n1592 & ~n16826 ) | ( n15818 & ~n16826 ) ;
  assign n32509 = n32508 ^ n23218 ^ n485 ;
  assign n32510 = n9605 & n32509 ;
  assign n32511 = n18291 & n32510 ;
  assign n32512 = ~n10599 & n18723 ;
  assign n32513 = ~n19189 & n32512 ;
  assign n32514 = n19244 ^ n16809 ^ 1'b0 ;
  assign n32515 = n8343 & n32514 ;
  assign n32516 = n15526 | n27664 ;
  assign n32517 = n32516 ^ n21951 ^ 1'b0 ;
  assign n32520 = n13542 ^ n12598 ^ 1'b0 ;
  assign n32518 = n8683 | n9008 ;
  assign n32519 = n24713 | n32518 ;
  assign n32521 = n32520 ^ n32519 ^ 1'b0 ;
  assign n32522 = ~n3217 & n13770 ;
  assign n32523 = n32522 ^ n4646 ^ 1'b0 ;
  assign n32524 = n32523 ^ n29982 ^ n1476 ;
  assign n32525 = ( n5149 & ~n18448 ) | ( n5149 & n18874 ) | ( ~n18448 & n18874 ) ;
  assign n32526 = ( n3589 & ~n17724 ) | ( n3589 & n32525 ) | ( ~n17724 & n32525 ) ;
  assign n32527 = n9226 & ~n12709 ;
  assign n32528 = n4311 & n32527 ;
  assign n32529 = n8294 & ~n22254 ;
  assign n32530 = n32529 ^ n31837 ^ n3679 ;
  assign n32531 = n27297 & ~n32530 ;
  assign n32532 = ~n27147 & n28411 ;
  assign n32533 = ~n14655 & n32532 ;
  assign n32534 = ~n1357 & n9880 ;
  assign n32535 = n32534 ^ n28927 ^ 1'b0 ;
  assign n32536 = ~n1930 & n32390 ;
  assign n32537 = n9342 & n32536 ;
  assign n32538 = ( ~n13618 & n28611 ) | ( ~n13618 & n32537 ) | ( n28611 & n32537 ) ;
  assign n32539 = n6001 ^ n1271 ^ 1'b0 ;
  assign n32540 = ( ~n10617 & n20895 ) | ( ~n10617 & n29562 ) | ( n20895 & n29562 ) ;
  assign n32541 = n19256 ^ n9335 ^ 1'b0 ;
  assign n32542 = n11503 & n32541 ;
  assign n32545 = ( ~n4739 & n5241 ) | ( ~n4739 & n32089 ) | ( n5241 & n32089 ) ;
  assign n32543 = n29348 ^ n14529 ^ 1'b0 ;
  assign n32544 = n3255 | n32543 ;
  assign n32546 = n32545 ^ n32544 ^ n1573 ;
  assign n32547 = ~n4383 & n11562 ;
  assign n32548 = n28554 ^ n21495 ^ n1899 ;
  assign n32549 = n390 & ~n23057 ;
  assign n32550 = ~n7875 & n32549 ;
  assign n32551 = ( n14498 & ~n16697 ) | ( n14498 & n26102 ) | ( ~n16697 & n26102 ) ;
  assign n32552 = n22269 ^ n14476 ^ n6946 ;
  assign n32553 = n3282 | n32552 ;
  assign n32554 = n32553 ^ n16040 ^ 1'b0 ;
  assign n32555 = n32554 ^ n424 ^ 1'b0 ;
  assign n32556 = n32551 | n32555 ;
  assign n32557 = ( n1682 & ~n17337 ) | ( n1682 & n23580 ) | ( ~n17337 & n23580 ) ;
  assign n32558 = ( ~n12333 & n20738 ) | ( ~n12333 & n32557 ) | ( n20738 & n32557 ) ;
  assign n32559 = n7821 & n27151 ;
  assign n32560 = n32559 ^ n13783 ^ 1'b0 ;
  assign n32561 = ~n10794 & n32560 ;
  assign n32562 = n32561 ^ n2293 ^ 1'b0 ;
  assign n32563 = n32562 ^ n25458 ^ 1'b0 ;
  assign n32564 = n11529 & ~n21363 ;
  assign n32565 = n32564 ^ n32107 ^ 1'b0 ;
  assign n32566 = n451 & n589 ;
  assign n32567 = n5128 & n32566 ;
  assign n32569 = n4271 & ~n9745 ;
  assign n32570 = ( n19311 & n19888 ) | ( n19311 & ~n32569 ) | ( n19888 & ~n32569 ) ;
  assign n32568 = n2746 ^ n2680 ^ 1'b0 ;
  assign n32571 = n32570 ^ n32568 ^ n4129 ;
  assign n32578 = ( n2818 & n6195 ) | ( n2818 & n11680 ) | ( n6195 & n11680 ) ;
  assign n32575 = n14544 ^ n12315 ^ n3257 ;
  assign n32576 = n32575 ^ n15414 ^ 1'b0 ;
  assign n32577 = ~n8437 & n32576 ;
  assign n32572 = n3090 & ~n28190 ;
  assign n32573 = n5043 ^ n4502 ^ 1'b0 ;
  assign n32574 = ( n2744 & ~n32572 ) | ( n2744 & n32573 ) | ( ~n32572 & n32573 ) ;
  assign n32579 = n32578 ^ n32577 ^ n32574 ;
  assign n32580 = n2263 | n10463 ;
  assign n32581 = x157 & n32580 ;
  assign n32582 = n17690 & ~n24356 ;
  assign n32583 = n32582 ^ n28997 ^ 1'b0 ;
  assign n32584 = ( n5038 & n6367 ) | ( n5038 & ~n8676 ) | ( n6367 & ~n8676 ) ;
  assign n32585 = ( n1413 & n3837 ) | ( n1413 & ~n17355 ) | ( n3837 & ~n17355 ) ;
  assign n32586 = n16491 ^ n11043 ^ 1'b0 ;
  assign n32587 = n3561 | n32586 ;
  assign n32588 = ( n2389 & n9752 ) | ( n2389 & n32587 ) | ( n9752 & n32587 ) ;
  assign n32589 = n9103 & ~n32588 ;
  assign n32590 = ~n32585 & n32589 ;
  assign n32591 = n32584 | n32590 ;
  assign n32592 = n18345 | n32591 ;
  assign n32593 = ~n4332 & n12169 ;
  assign n32594 = n20021 & n32226 ;
  assign n32595 = n32593 & n32594 ;
  assign n32596 = n4310 & n19356 ;
  assign n32597 = n3835 & ~n32596 ;
  assign n32598 = n7851 & n12744 ;
  assign n32599 = n32598 ^ n3972 ^ 1'b0 ;
  assign n32600 = ~n28722 & n32599 ;
  assign n32601 = n23556 & ~n32600 ;
  assign n32602 = ( n5233 & ~n20630 ) | ( n5233 & n20747 ) | ( ~n20630 & n20747 ) ;
  assign n32603 = ( n9660 & ~n18009 ) | ( n9660 & n32013 ) | ( ~n18009 & n32013 ) ;
  assign n32604 = n6826 & ~n14559 ;
  assign n32605 = n32604 ^ n3693 ^ 1'b0 ;
  assign n32606 = n32605 ^ n14364 ^ n13005 ;
  assign n32607 = ~n14953 & n19779 ;
  assign n32608 = n3483 & n7634 ;
  assign n32609 = ~x17 & n32608 ;
  assign n32610 = n5923 ^ n5345 ^ 1'b0 ;
  assign n32611 = n13090 | n32610 ;
  assign n32612 = n3819 & ~n4543 ;
  assign n32613 = n1178 & ~n18762 ;
  assign n32614 = ~n32612 & n32613 ;
  assign n32615 = n32614 ^ n12622 ^ 1'b0 ;
  assign n32617 = n27294 ^ n13803 ^ 1'b0 ;
  assign n32616 = n14725 & n26287 ;
  assign n32618 = n32617 ^ n32616 ^ 1'b0 ;
  assign n32619 = n30519 ^ n15843 ^ 1'b0 ;
  assign n32620 = n24781 ^ n2685 ^ 1'b0 ;
  assign n32621 = n28094 ^ n27411 ^ 1'b0 ;
  assign n32622 = n32620 | n32621 ;
  assign n32623 = n10822 | n32622 ;
  assign n32624 = n32623 ^ n18561 ^ 1'b0 ;
  assign n32625 = n8331 ^ n7916 ^ 1'b0 ;
  assign n32626 = n18783 & n32625 ;
  assign n32627 = n3188 & ~n32626 ;
  assign n32628 = ~n32094 & n32627 ;
  assign n32629 = n17918 ^ n14046 ^ n10899 ;
  assign n32630 = n32629 ^ n7480 ^ n5834 ;
  assign n32631 = n32628 & n32630 ;
  assign n32632 = ( ~n17703 & n17944 ) | ( ~n17703 & n23837 ) | ( n17944 & n23837 ) ;
  assign n32633 = n11285 ^ n9157 ^ n6669 ;
  assign n32634 = n32633 ^ n21336 ^ n12057 ;
  assign n32635 = n32634 ^ n10964 ^ n2310 ;
  assign n32636 = ~n13041 & n32635 ;
  assign n32637 = n5368 | n18868 ;
  assign n32638 = n8208 | n13061 ;
  assign n32639 = n32638 ^ n18439 ^ 1'b0 ;
  assign n32640 = n20261 & ~n32639 ;
  assign n32641 = n4756 & ~n5850 ;
  assign n32642 = n3227 | n5245 ;
  assign n32643 = n32642 ^ n32514 ^ 1'b0 ;
  assign n32644 = n32641 & n32643 ;
  assign n32645 = ~n1022 & n16640 ;
  assign n32646 = n22783 ^ n284 ^ 1'b0 ;
  assign n32647 = ~n2051 & n23437 ;
  assign n32648 = n4114 | n17589 ;
  assign n32649 = n6888 | n32648 ;
  assign n32650 = n16366 & n32649 ;
  assign n32651 = n21605 & n32650 ;
  assign n32652 = n10661 & n13615 ;
  assign n32653 = ( ~x6 & n24327 ) | ( ~x6 & n26818 ) | ( n24327 & n26818 ) ;
  assign n32654 = n7655 ^ n1285 ^ 1'b0 ;
  assign n32655 = n424 | n29186 ;
  assign n32656 = ( ~n17106 & n32654 ) | ( ~n17106 & n32655 ) | ( n32654 & n32655 ) ;
  assign n32657 = n11802 & ~n15086 ;
  assign n32658 = n27230 ^ n722 ^ 1'b0 ;
  assign n32659 = n32658 ^ n23795 ^ n20136 ;
  assign n32660 = ~n8821 & n32659 ;
  assign n32661 = n32657 & n32660 ;
  assign n32662 = n11116 | n23614 ;
  assign n32663 = n2144 | n15760 ;
  assign n32664 = n22065 | n32663 ;
  assign n32665 = n32249 ^ n21206 ^ n4326 ;
  assign n32666 = n32665 ^ n24948 ^ n5466 ;
  assign n32667 = ~n25620 & n32666 ;
  assign n32668 = n32667 ^ n15033 ^ 1'b0 ;
  assign n32669 = ( n4600 & n25059 ) | ( n4600 & n26995 ) | ( n25059 & n26995 ) ;
  assign n32670 = n28813 ^ n25362 ^ n19810 ;
  assign n32673 = n9064 ^ n7598 ^ 1'b0 ;
  assign n32672 = ~n6077 & n14946 ;
  assign n32674 = n32673 ^ n32672 ^ 1'b0 ;
  assign n32671 = n3923 | n5767 ;
  assign n32675 = n32674 ^ n32671 ^ n2769 ;
  assign n32676 = ( n6606 & n12418 ) | ( n6606 & ~n25189 ) | ( n12418 & ~n25189 ) ;
  assign n32677 = n16366 & ~n32676 ;
  assign n32678 = n32677 ^ n7966 ^ 1'b0 ;
  assign n32679 = n11703 ^ n10784 ^ 1'b0 ;
  assign n32680 = n20117 | n32679 ;
  assign n32682 = ( n7256 & ~n7560 ) | ( n7256 & n11384 ) | ( ~n7560 & n11384 ) ;
  assign n32681 = x177 & n9235 ;
  assign n32683 = n32682 ^ n32681 ^ 1'b0 ;
  assign n32684 = n10380 & ~n32683 ;
  assign n32685 = ~n495 & n6326 ;
  assign n32686 = n32685 ^ n10728 ^ 1'b0 ;
  assign n32687 = ~n29084 & n32686 ;
  assign n32691 = n9818 | n10398 ;
  assign n32692 = n32691 ^ n17979 ^ 1'b0 ;
  assign n32693 = n3587 | n32692 ;
  assign n32688 = n4112 & n9434 ;
  assign n32689 = n32688 ^ n1749 ^ 1'b0 ;
  assign n32690 = n16012 & ~n32689 ;
  assign n32694 = n32693 ^ n32690 ^ 1'b0 ;
  assign n32695 = n15304 ^ n3440 ^ x244 ;
  assign n32696 = n32695 ^ n21870 ^ 1'b0 ;
  assign n32697 = n32696 ^ n13809 ^ n8268 ;
  assign n32698 = n10038 & ~n17098 ;
  assign n32699 = n24419 | n32698 ;
  assign n32700 = n1415 & ~n23012 ;
  assign n32701 = n16439 | n32700 ;
  assign n32702 = n32699 | n32701 ;
  assign n32703 = n10850 ^ n1542 ^ n913 ;
  assign n32704 = n25446 ^ n21144 ^ 1'b0 ;
  assign n32705 = ~n7814 & n21827 ;
  assign n32706 = ~n12941 & n32705 ;
  assign n32707 = n6585 & n32706 ;
  assign n32708 = ( n24629 & n31056 ) | ( n24629 & n32707 ) | ( n31056 & n32707 ) ;
  assign n32709 = n10005 ^ n7550 ^ 1'b0 ;
  assign n32710 = n13407 ^ n6858 ^ n3190 ;
  assign n32711 = n11984 & n32710 ;
  assign n32712 = n32709 & ~n32711 ;
  assign n32713 = ~n10045 & n18785 ;
  assign n32714 = n24387 & n32713 ;
  assign n32715 = n6385 | n32714 ;
  assign n32716 = n6341 & ~n32715 ;
  assign n32717 = n853 & ~n1434 ;
  assign n32718 = n32706 ^ n8315 ^ n3674 ;
  assign n32719 = ~n8290 & n32718 ;
  assign n32720 = n3521 & n8957 ;
  assign n32721 = n12760 & ~n15008 ;
  assign n32722 = n11097 & n12039 ;
  assign n32723 = n9296 & n32722 ;
  assign n32724 = n3433 & n20957 ;
  assign n32725 = n32723 & n32724 ;
  assign n32726 = n32725 ^ n26029 ^ n22991 ;
  assign n32727 = n19936 ^ n16150 ^ n9296 ;
  assign n32728 = n1494 | n32727 ;
  assign n32729 = n32728 ^ n10259 ^ 1'b0 ;
  assign n32730 = n32729 ^ n11857 ^ n4935 ;
  assign n32731 = n5949 ^ n1773 ^ 1'b0 ;
  assign n32732 = n3869 | n32731 ;
  assign n32733 = n22541 ^ n6379 ^ 1'b0 ;
  assign n32734 = n32732 | n32733 ;
  assign n32735 = n30066 ^ n22155 ^ n5135 ;
  assign n32736 = n32735 ^ n5108 ^ n5071 ;
  assign n32737 = n10990 | n31654 ;
  assign n32738 = n32736 | n32737 ;
  assign n32739 = n10464 | n13067 ;
  assign n32740 = ( n10865 & n26298 ) | ( n10865 & n29684 ) | ( n26298 & n29684 ) ;
  assign n32743 = n6094 & ~n23941 ;
  assign n32744 = n8631 & n32743 ;
  assign n32741 = n3854 ^ n2006 ^ 1'b0 ;
  assign n32742 = n19273 & ~n32741 ;
  assign n32745 = n32744 ^ n32742 ^ 1'b0 ;
  assign n32746 = n9658 & ~n19239 ;
  assign n32747 = ( ~n2294 & n23541 ) | ( ~n2294 & n32746 ) | ( n23541 & n32746 ) ;
  assign n32748 = n32747 ^ n21456 ^ n5994 ;
  assign n32749 = n32748 ^ n16474 ^ 1'b0 ;
  assign n32750 = n32745 & n32749 ;
  assign n32751 = n6606 & n25707 ;
  assign n32757 = ( n4593 & n5203 ) | ( n4593 & ~n12092 ) | ( n5203 & ~n12092 ) ;
  assign n32752 = ~n9927 & n14528 ;
  assign n32753 = n5792 & n32752 ;
  assign n32754 = n18409 | n32753 ;
  assign n32755 = n13212 | n32754 ;
  assign n32756 = n13418 & n32755 ;
  assign n32758 = n32757 ^ n32756 ^ 1'b0 ;
  assign n32759 = ~n6562 & n18700 ;
  assign n32760 = n26281 ^ n22519 ^ n9641 ;
  assign n32761 = n30700 ^ n20201 ^ 1'b0 ;
  assign n32762 = n31747 ^ n13944 ^ 1'b0 ;
  assign n32763 = n14641 & n32762 ;
  assign n32764 = ( ~n10475 & n16495 ) | ( ~n10475 & n32763 ) | ( n16495 & n32763 ) ;
  assign n32766 = n23795 ^ n5527 ^ 1'b0 ;
  assign n32767 = n7140 & n32766 ;
  assign n32768 = n32767 ^ n22386 ^ n1715 ;
  assign n32769 = ( n1554 & n23418 ) | ( n1554 & n32768 ) | ( n23418 & n32768 ) ;
  assign n32765 = n7867 | n13494 ;
  assign n32770 = n32769 ^ n32765 ^ 1'b0 ;
  assign n32771 = ~n15780 & n18579 ;
  assign n32772 = ~n2904 & n32771 ;
  assign n32773 = n10776 ^ n5881 ^ 1'b0 ;
  assign n32774 = n17073 | n32773 ;
  assign n32775 = n1403 & ~n2906 ;
  assign n32776 = n32775 ^ n16581 ^ 1'b0 ;
  assign n32777 = ( n23064 & n27215 ) | ( n23064 & n32776 ) | ( n27215 & n32776 ) ;
  assign n32778 = ( n1639 & n20406 ) | ( n1639 & ~n31812 ) | ( n20406 & ~n31812 ) ;
  assign n32779 = n18454 ^ n8614 ^ 1'b0 ;
  assign n32780 = n32779 ^ n3200 ^ 1'b0 ;
  assign n32781 = n32780 ^ n13593 ^ x26 ;
  assign n32782 = ~n22498 & n32781 ;
  assign n32783 = n32782 ^ n15126 ^ 1'b0 ;
  assign n32787 = n7370 ^ n1271 ^ 1'b0 ;
  assign n32784 = ( n1034 & n7100 ) | ( n1034 & n16583 ) | ( n7100 & n16583 ) ;
  assign n32785 = n18716 ^ n1553 ^ 1'b0 ;
  assign n32786 = n32784 & ~n32785 ;
  assign n32788 = n32787 ^ n32786 ^ 1'b0 ;
  assign n32789 = ( n6001 & n17558 ) | ( n6001 & ~n32788 ) | ( n17558 & ~n32788 ) ;
  assign n32792 = n23412 ^ n10736 ^ 1'b0 ;
  assign n32791 = x236 & n22101 ;
  assign n32790 = n18928 ^ n17916 ^ 1'b0 ;
  assign n32793 = n32792 ^ n32791 ^ n32790 ;
  assign n32794 = ( n24094 & ~n24394 ) | ( n24094 & n28416 ) | ( ~n24394 & n28416 ) ;
  assign n32795 = n13009 ^ n7988 ^ 1'b0 ;
  assign n32796 = n32795 ^ n24996 ^ 1'b0 ;
  assign n32797 = n6783 ^ n857 ^ 1'b0 ;
  assign n32798 = n22059 | n32797 ;
  assign n32799 = n10959 ^ n1548 ^ n316 ;
  assign n32800 = n32799 ^ n17401 ^ 1'b0 ;
  assign n32801 = ~n8047 & n30315 ;
  assign n32802 = n12263 ^ n7988 ^ 1'b0 ;
  assign n32803 = n13407 & n32802 ;
  assign n32804 = ( n1463 & n21354 ) | ( n1463 & n29651 ) | ( n21354 & n29651 ) ;
  assign n32805 = n1789 | n11480 ;
  assign n32806 = n32805 ^ n8678 ^ 1'b0 ;
  assign n32807 = n9835 & n32806 ;
  assign n32808 = ( n1521 & ~n6847 ) | ( n1521 & n9336 ) | ( ~n6847 & n9336 ) ;
  assign n32809 = n20323 & n29507 ;
  assign n32810 = n32809 ^ n4280 ^ 1'b0 ;
  assign n32811 = n1684 & n8891 ;
  assign n32812 = n19737 & n32811 ;
  assign n32813 = n3934 & ~n6558 ;
  assign n32814 = ~n15996 & n32813 ;
  assign n32815 = n24639 ^ n2878 ^ 1'b0 ;
  assign n32816 = ( n4512 & n26730 ) | ( n4512 & ~n32815 ) | ( n26730 & ~n32815 ) ;
  assign n32817 = ~n1205 & n13251 ;
  assign n32818 = ~n10515 & n32817 ;
  assign n32819 = n19192 & ~n32818 ;
  assign n32820 = n11516 & n32819 ;
  assign n32821 = n17620 & ~n21597 ;
  assign n32822 = ~n21530 & n32821 ;
  assign n32823 = ( n4835 & ~n32820 ) | ( n4835 & n32822 ) | ( ~n32820 & n32822 ) ;
  assign n32824 = n4351 & ~n7484 ;
  assign n32825 = ~n1736 & n6708 ;
  assign n32826 = n22190 & n32825 ;
  assign n32829 = n17773 ^ n15239 ^ 1'b0 ;
  assign n32827 = n17357 ^ n5264 ^ 1'b0 ;
  assign n32828 = n12716 & n32827 ;
  assign n32830 = n32829 ^ n32828 ^ 1'b0 ;
  assign n32831 = ( ~x144 & n5624 ) | ( ~x144 & n18413 ) | ( n5624 & n18413 ) ;
  assign n32832 = n2391 & n32831 ;
  assign n32833 = n31292 ^ n14246 ^ 1'b0 ;
  assign n32834 = ( n5214 & n8056 ) | ( n5214 & ~n26556 ) | ( n8056 & ~n26556 ) ;
  assign n32835 = n32834 ^ n28825 ^ 1'b0 ;
  assign n32836 = x168 & n15613 ;
  assign n32837 = n32836 ^ n22784 ^ n8079 ;
  assign n32838 = n18720 & ~n29112 ;
  assign n32839 = ~n19072 & n32838 ;
  assign n32840 = n32839 ^ n20086 ^ 1'b0 ;
  assign n32841 = n23758 & ~n32840 ;
  assign n32842 = ( n9778 & n11807 ) | ( n9778 & n29057 ) | ( n11807 & n29057 ) ;
  assign n32843 = n31281 & ~n32842 ;
  assign n32844 = n28575 & n32843 ;
  assign n32845 = n973 & n22254 ;
  assign n32846 = n10799 & n12160 ;
  assign n32847 = n32846 ^ n10157 ^ 1'b0 ;
  assign n32848 = n32847 ^ n9919 ^ 1'b0 ;
  assign n32849 = n32848 ^ n27140 ^ 1'b0 ;
  assign n32851 = n12301 ^ n9640 ^ 1'b0 ;
  assign n32852 = ~n13393 & n32851 ;
  assign n32853 = n28309 & n32852 ;
  assign n32854 = n32853 ^ n21430 ^ 1'b0 ;
  assign n32850 = n12344 & n27387 ;
  assign n32855 = n32854 ^ n32850 ^ 1'b0 ;
  assign n32856 = ~n3342 & n32855 ;
  assign n32857 = n32856 ^ n24588 ^ 1'b0 ;
  assign n32858 = ~n6302 & n8947 ;
  assign n32859 = n9990 & ~n28718 ;
  assign n32860 = n10017 & n32859 ;
  assign n32861 = ~n9250 & n17562 ;
  assign n32862 = n1563 & n32861 ;
  assign n32863 = n32862 ^ n2843 ^ 1'b0 ;
  assign n32864 = n808 & ~n32863 ;
  assign n32865 = n32864 ^ n16783 ^ 1'b0 ;
  assign n32866 = ~n16083 & n23298 ;
  assign n32867 = ~n2314 & n10052 ;
  assign n32868 = ( n3235 & n14975 ) | ( n3235 & ~n22292 ) | ( n14975 & ~n22292 ) ;
  assign n32869 = n3959 & n28281 ;
  assign n32870 = n32868 & n32869 ;
  assign n32871 = n11446 | n11506 ;
  assign n32872 = n7043 ^ n669 ^ 1'b0 ;
  assign n32873 = ~n12929 & n32872 ;
  assign n32874 = n32873 ^ n26172 ^ 1'b0 ;
  assign n32875 = ( ~x84 & n1548 ) | ( ~x84 & n2958 ) | ( n1548 & n2958 ) ;
  assign n32876 = n32875 ^ n9014 ^ 1'b0 ;
  assign n32877 = n17448 & n32876 ;
  assign n32878 = n32874 & n32877 ;
  assign n32879 = ( n23012 & n27495 ) | ( n23012 & n30464 ) | ( n27495 & n30464 ) ;
  assign n32880 = ~n2723 & n5758 ;
  assign n32881 = n32880 ^ n1972 ^ 1'b0 ;
  assign n32882 = n10757 & n32881 ;
  assign n32883 = n32882 ^ n9030 ^ n5934 ;
  assign n32884 = n2199 & n15788 ;
  assign n32885 = ( n3056 & n10643 ) | ( n3056 & ~n18197 ) | ( n10643 & ~n18197 ) ;
  assign n32886 = n32885 ^ n10287 ^ n7288 ;
  assign n32887 = n10179 | n32886 ;
  assign n32888 = n14895 ^ n10656 ^ 1'b0 ;
  assign n32889 = n19296 ^ n6606 ^ 1'b0 ;
  assign n32890 = ~n11085 & n32889 ;
  assign n32893 = n20039 & n27368 ;
  assign n32891 = n4287 & n19399 ;
  assign n32892 = n32891 ^ n11502 ^ 1'b0 ;
  assign n32894 = n32893 ^ n32892 ^ n13140 ;
  assign n32895 = n28686 ^ n13758 ^ 1'b0 ;
  assign n32896 = n4431 & ~n32895 ;
  assign n32897 = n15614 ^ n2505 ^ 1'b0 ;
  assign n32898 = n4140 & ~n32897 ;
  assign n32899 = n32898 ^ n2769 ^ 1'b0 ;
  assign n32900 = n10688 & n32899 ;
  assign n32903 = n1451 & n10768 ;
  assign n32904 = ~n26856 & n32903 ;
  assign n32905 = x36 & ~n32904 ;
  assign n32906 = ~n5879 & n32905 ;
  assign n32907 = n32906 ^ n14527 ^ n337 ;
  assign n32901 = n411 | n24565 ;
  assign n32902 = n15343 | n32901 ;
  assign n32908 = n32907 ^ n32902 ^ 1'b0 ;
  assign n32909 = n17532 | n32908 ;
  assign n32911 = ~n1931 & n4411 ;
  assign n32910 = n1653 | n19560 ;
  assign n32912 = n32911 ^ n32910 ^ 1'b0 ;
  assign n32913 = n6969 & n7741 ;
  assign n32914 = n16337 & ~n32913 ;
  assign n32915 = n2476 ^ n2050 ^ 1'b0 ;
  assign n32916 = n15476 ^ n8481 ^ 1'b0 ;
  assign n32917 = n26232 ^ n4411 ^ 1'b0 ;
  assign n32918 = n17631 ^ n12715 ^ 1'b0 ;
  assign n32919 = n24429 & n32918 ;
  assign n32920 = n27075 ^ n2204 ^ 1'b0 ;
  assign n32921 = n12920 & ~n16142 ;
  assign n32922 = n32921 ^ n19992 ^ n5458 ;
  assign n32923 = ~n29243 & n32922 ;
  assign n32924 = ( ~n7416 & n10402 ) | ( ~n7416 & n32923 ) | ( n10402 & n32923 ) ;
  assign n32925 = n675 | n17749 ;
  assign n32926 = n32925 ^ n997 ^ 1'b0 ;
  assign n32927 = n32297 & n32926 ;
  assign n32928 = n17306 ^ n5676 ^ 1'b0 ;
  assign n32929 = n32927 | n32928 ;
  assign n32930 = ( n2427 & n4120 ) | ( n2427 & n5737 ) | ( n4120 & n5737 ) ;
  assign n32931 = n32930 ^ n6710 ^ n3203 ;
  assign n32932 = n32931 ^ n9101 ^ 1'b0 ;
  assign n32933 = n13587 & ~n32932 ;
  assign n32934 = n13951 | n29891 ;
  assign n32935 = n9085 & ~n32934 ;
  assign n32936 = n22833 & n32935 ;
  assign n32937 = ( n4257 & n11897 ) | ( n4257 & ~n12522 ) | ( n11897 & ~n12522 ) ;
  assign n32938 = ~n6393 & n23677 ;
  assign n32939 = ~n945 & n32938 ;
  assign n32940 = ( n22918 & ~n32937 ) | ( n22918 & n32939 ) | ( ~n32937 & n32939 ) ;
  assign n32941 = ( n10058 & n29867 ) | ( n10058 & n32940 ) | ( n29867 & n32940 ) ;
  assign n32942 = ( ~n3689 & n25635 ) | ( ~n3689 & n32941 ) | ( n25635 & n32941 ) ;
  assign n32943 = n6094 ^ n5897 ^ n5611 ;
  assign n32944 = n32943 ^ n20776 ^ n3707 ;
  assign n32945 = n29688 ^ n591 ^ 1'b0 ;
  assign n32946 = n10326 & ~n32945 ;
  assign n32947 = n29154 ^ n4065 ^ 1'b0 ;
  assign n32948 = ~n2003 & n3260 ;
  assign n32949 = n16553 & n32948 ;
  assign n32950 = n2950 & ~n32949 ;
  assign n32951 = n7085 & ~n32950 ;
  assign n32952 = ~n32947 & n32951 ;
  assign n32953 = n10476 & ~n30650 ;
  assign n32954 = n4879 & n23699 ;
  assign n32955 = n32954 ^ n2931 ^ 1'b0 ;
  assign n32956 = ( n7690 & n9656 ) | ( n7690 & n13540 ) | ( n9656 & n13540 ) ;
  assign n32957 = n2351 & n2466 ;
  assign n32958 = n19780 ^ n14978 ^ 1'b0 ;
  assign n32959 = ~n32957 & n32958 ;
  assign n32960 = n22699 ^ n14496 ^ 1'b0 ;
  assign n32961 = n32959 & ~n32960 ;
  assign n32962 = n32961 ^ n17407 ^ n2997 ;
  assign n32963 = n21392 ^ n21343 ^ 1'b0 ;
  assign n32964 = n8815 & ~n23541 ;
  assign n32965 = ( n32962 & ~n32963 ) | ( n32962 & n32964 ) | ( ~n32963 & n32964 ) ;
  assign n32966 = n31450 ^ n24184 ^ n19694 ;
  assign n32967 = n32966 ^ n22773 ^ x159 ;
  assign n32968 = n12400 & n32230 ;
  assign n32969 = n15835 & n32968 ;
  assign n32970 = n14393 ^ n8206 ^ 1'b0 ;
  assign n32974 = n8017 & ~n29769 ;
  assign n32975 = n9885 & n32974 ;
  assign n32976 = n32975 ^ n32015 ^ n15132 ;
  assign n32971 = ~n15257 & n16698 ;
  assign n32972 = ~n25798 & n27473 ;
  assign n32973 = n32971 & ~n32972 ;
  assign n32977 = n32976 ^ n32973 ^ n27520 ;
  assign n32979 = n15743 | n25165 ;
  assign n32980 = n32979 ^ n15433 ^ 1'b0 ;
  assign n32978 = n6504 ^ n2962 ^ 1'b0 ;
  assign n32981 = n32980 ^ n32978 ^ 1'b0 ;
  assign n32982 = n32981 ^ n20752 ^ n15865 ;
  assign n32983 = n4039 | n29059 ;
  assign n32984 = ~n23901 & n31096 ;
  assign n32985 = ~n1955 & n2613 ;
  assign n32986 = n22170 & n32985 ;
  assign n32987 = n29600 ^ n6272 ^ 1'b0 ;
  assign n32988 = n6194 | n32987 ;
  assign n32989 = n32988 ^ n7113 ^ 1'b0 ;
  assign n32990 = n14758 & n32989 ;
  assign n32991 = n32990 ^ n2857 ^ 1'b0 ;
  assign n32992 = ~n6192 & n32991 ;
  assign n32995 = n10132 & ~n14628 ;
  assign n32996 = n32995 ^ n9080 ^ 1'b0 ;
  assign n32993 = n2099 & n32757 ;
  assign n32994 = n32993 ^ n21785 ^ 1'b0 ;
  assign n32997 = n32996 ^ n32994 ^ n8201 ;
  assign n32998 = n32997 ^ n21304 ^ n17984 ;
  assign n32999 = n923 | n9540 ;
  assign n33000 = n15525 | n32999 ;
  assign n33001 = n33000 ^ n32829 ^ n9308 ;
  assign n33002 = n11817 ^ n5779 ^ n3803 ;
  assign n33003 = n6113 ^ n3819 ^ n3039 ;
  assign n33004 = ( n12410 & ~n33002 ) | ( n12410 & n33003 ) | ( ~n33002 & n33003 ) ;
  assign n33005 = ( n12730 & n26369 ) | ( n12730 & ~n33004 ) | ( n26369 & ~n33004 ) ;
  assign n33006 = n23651 ^ n2165 ^ 1'b0 ;
  assign n33007 = ~n1106 & n10830 ;
  assign n33008 = n17507 & n33007 ;
  assign n33009 = n11381 & ~n33008 ;
  assign n33010 = n33009 ^ n14639 ^ n1516 ;
  assign n33011 = n33010 ^ n15664 ^ 1'b0 ;
  assign n33012 = n19709 ^ n4179 ^ 1'b0 ;
  assign n33013 = ( x59 & n5235 ) | ( x59 & n8630 ) | ( n5235 & n8630 ) ;
  assign n33014 = ~n1286 & n33013 ;
  assign n33015 = ~n33012 & n33014 ;
  assign n33016 = ( n2856 & n11268 ) | ( n2856 & ~n29088 ) | ( n11268 & ~n29088 ) ;
  assign n33017 = n15038 ^ n5873 ^ 1'b0 ;
  assign n33018 = ( ~n6117 & n16276 ) | ( ~n6117 & n33017 ) | ( n16276 & n33017 ) ;
  assign n33019 = n11106 | n19329 ;
  assign n33020 = n24314 | n33019 ;
  assign n33021 = n2171 | n24706 ;
  assign n33022 = n18227 & ~n33021 ;
  assign n33023 = ~n4108 & n4554 ;
  assign n33024 = n6103 ^ n1705 ^ 1'b0 ;
  assign n33025 = ( ~n3347 & n33023 ) | ( ~n3347 & n33024 ) | ( n33023 & n33024 ) ;
  assign n33026 = n15969 ^ n12567 ^ n992 ;
  assign n33027 = ( n7798 & ~n11502 ) | ( n7798 & n33026 ) | ( ~n11502 & n33026 ) ;
  assign n33028 = n33027 ^ n5715 ^ 1'b0 ;
  assign n33029 = n13119 | n32886 ;
  assign n33030 = n33029 ^ n21414 ^ 1'b0 ;
  assign n33031 = n23963 ^ n6542 ^ n4683 ;
  assign n33032 = n33031 ^ n27115 ^ n9732 ;
  assign n33033 = ~n32031 & n33032 ;
  assign n33034 = n33033 ^ n18711 ^ 1'b0 ;
  assign n33035 = n11804 & ~n27436 ;
  assign n33036 = ~n9529 & n33035 ;
  assign n33037 = n19115 | n33036 ;
  assign n33038 = n33037 ^ n26208 ^ 1'b0 ;
  assign n33039 = n839 & n15996 ;
  assign n33040 = n33039 ^ n5841 ^ 1'b0 ;
  assign n33041 = x12 & ~n5573 ;
  assign n33042 = n33041 ^ n3142 ^ 1'b0 ;
  assign n33043 = ( n11663 & n33040 ) | ( n11663 & ~n33042 ) | ( n33040 & ~n33042 ) ;
  assign n33044 = ~n9723 & n31682 ;
  assign n33045 = n33044 ^ n22822 ^ n16345 ;
  assign n33046 = n29570 ^ n17159 ^ n7611 ;
  assign n33047 = n4237 | n6357 ;
  assign n33048 = n12766 | n13120 ;
  assign n33049 = n33047 | n33048 ;
  assign n33050 = n8279 ^ n3793 ^ n2771 ;
  assign n33051 = n33050 ^ n3085 ^ 1'b0 ;
  assign n33052 = n25583 & ~n33051 ;
  assign n33053 = n902 | n3619 ;
  assign n33054 = n33053 ^ n3104 ^ 1'b0 ;
  assign n33055 = n22278 ^ n21736 ^ n7031 ;
  assign n33056 = ( n3034 & ~n19051 ) | ( n3034 & n33055 ) | ( ~n19051 & n33055 ) ;
  assign n33057 = ( n18647 & n25988 ) | ( n18647 & ~n26613 ) | ( n25988 & ~n26613 ) ;
  assign n33058 = n953 & ~n22943 ;
  assign n33059 = ( n18920 & n33057 ) | ( n18920 & n33058 ) | ( n33057 & n33058 ) ;
  assign n33060 = ( n6402 & n8345 ) | ( n6402 & n15838 ) | ( n8345 & n15838 ) ;
  assign n33061 = n12109 ^ n6860 ^ 1'b0 ;
  assign n33062 = n33060 | n33061 ;
  assign n33063 = n15803 & n33062 ;
  assign n33064 = n4209 & n18569 ;
  assign n33065 = n15686 | n33064 ;
  assign n33066 = n17075 & n23630 ;
  assign n33067 = ~n31182 & n33066 ;
  assign n33068 = ( n1104 & n1637 ) | ( n1104 & n14533 ) | ( n1637 & n14533 ) ;
  assign n33069 = ( n1174 & n17624 ) | ( n1174 & ~n25316 ) | ( n17624 & ~n25316 ) ;
  assign n33070 = n12550 ^ n4784 ^ 1'b0 ;
  assign n33071 = ( n1064 & n18953 ) | ( n1064 & n33070 ) | ( n18953 & n33070 ) ;
  assign n33072 = n7912 ^ n6074 ^ 1'b0 ;
  assign n33073 = ~n28305 & n33072 ;
  assign n33074 = n4615 & ~n5478 ;
  assign n33075 = n33074 ^ n2385 ^ 1'b0 ;
  assign n33076 = n33075 ^ n26706 ^ n26693 ;
  assign n33077 = n3899 & n10695 ;
  assign n33078 = n33077 ^ n23852 ^ 1'b0 ;
  assign n33079 = n15447 ^ n7710 ^ 1'b0 ;
  assign n33080 = ~x48 & n33079 ;
  assign n33081 = n11113 ^ n7515 ^ 1'b0 ;
  assign n33082 = n30339 & ~n33081 ;
  assign n33083 = n27479 ^ n14102 ^ 1'b0 ;
  assign n33084 = n4427 & ~n10350 ;
  assign n33085 = n33084 ^ n30310 ^ 1'b0 ;
  assign n33086 = n33085 ^ n30867 ^ 1'b0 ;
  assign n33087 = n19883 ^ n5715 ^ 1'b0 ;
  assign n33088 = n29590 ^ n9068 ^ n2722 ;
  assign n33089 = n33088 ^ n8496 ^ 1'b0 ;
  assign n33090 = n6196 & n28925 ;
  assign n33091 = n1048 & n33090 ;
  assign n33092 = n33091 ^ n19551 ^ 1'b0 ;
  assign n33093 = n33092 ^ n30810 ^ 1'b0 ;
  assign n33094 = ( n8716 & n13721 ) | ( n8716 & ~n16540 ) | ( n13721 & ~n16540 ) ;
  assign n33095 = n33094 ^ n28133 ^ n12598 ;
  assign n33096 = ~n33093 & n33095 ;
  assign n33097 = n9641 & n10044 ;
  assign n33098 = n1209 & n33097 ;
  assign n33099 = ( ~n3222 & n3768 ) | ( ~n3222 & n33098 ) | ( n3768 & n33098 ) ;
  assign n33100 = n14178 & n33099 ;
  assign n33101 = n8343 & ~n22284 ;
  assign n33102 = n33101 ^ n25793 ^ 1'b0 ;
  assign n33103 = n3514 | n33102 ;
  assign n33104 = ( n1409 & n2106 ) | ( n1409 & n3943 ) | ( n2106 & n3943 ) ;
  assign n33105 = n21794 ^ n7001 ^ 1'b0 ;
  assign n33106 = n8328 & ~n14713 ;
  assign n33107 = n33106 ^ n25799 ^ 1'b0 ;
  assign n33108 = n19070 ^ n11104 ^ 1'b0 ;
  assign n33109 = n10734 ^ n8629 ^ n507 ;
  assign n33110 = ( n6425 & ~n8670 ) | ( n6425 & n11128 ) | ( ~n8670 & n11128 ) ;
  assign n33111 = ~n33109 & n33110 ;
  assign n33112 = ( n10555 & ~n18841 ) | ( n10555 & n32990 ) | ( ~n18841 & n32990 ) ;
  assign n33113 = n26566 & ~n33112 ;
  assign n33114 = ~n14014 & n33113 ;
  assign n33115 = n11025 ^ n7011 ^ 1'b0 ;
  assign n33116 = n3640 | n33115 ;
  assign n33117 = ( n4395 & n13478 ) | ( n4395 & n17394 ) | ( n13478 & n17394 ) ;
  assign n33118 = n23364 & n33117 ;
  assign n33119 = n33116 & n33118 ;
  assign n33120 = n9061 ^ n3247 ^ 1'b0 ;
  assign n33121 = n17129 ^ n10342 ^ 1'b0 ;
  assign n33122 = ( n9937 & n33120 ) | ( n9937 & ~n33121 ) | ( n33120 & ~n33121 ) ;
  assign n33123 = n16736 ^ n8930 ^ 1'b0 ;
  assign n33124 = n816 & n2339 ;
  assign n33125 = ~n15921 & n33124 ;
  assign n33126 = n8512 & ~n11219 ;
  assign n33127 = n32681 & n33126 ;
  assign n33128 = n32961 ^ n20635 ^ 1'b0 ;
  assign n33129 = n5781 & n17179 ;
  assign n33130 = n5773 | n5942 ;
  assign n33131 = n1693 & ~n33130 ;
  assign n33132 = n17631 & ~n25026 ;
  assign n33133 = ( ~n21139 & n33131 ) | ( ~n21139 & n33132 ) | ( n33131 & n33132 ) ;
  assign n33134 = ( n2445 & n5919 ) | ( n2445 & ~n8674 ) | ( n5919 & ~n8674 ) ;
  assign n33135 = n9351 | n33134 ;
  assign n33136 = n33135 ^ n30515 ^ 1'b0 ;
  assign n33137 = n15686 & n26381 ;
  assign n33138 = ~n23893 & n33137 ;
  assign n33139 = n18435 | n23096 ;
  assign n33140 = n33139 ^ n24250 ^ 1'b0 ;
  assign n33141 = n6251 ^ n4394 ^ n1993 ;
  assign n33142 = ( n4909 & n6393 ) | ( n4909 & n28230 ) | ( n6393 & n28230 ) ;
  assign n33143 = n6960 & n10106 ;
  assign n33144 = ( n9665 & n33142 ) | ( n9665 & ~n33143 ) | ( n33142 & ~n33143 ) ;
  assign n33145 = n9064 ^ n4795 ^ 1'b0 ;
  assign n33146 = ( n5188 & n10356 ) | ( n5188 & ~n33145 ) | ( n10356 & ~n33145 ) ;
  assign n33147 = n14353 & n33146 ;
  assign n33148 = n31221 & n33147 ;
  assign n33150 = n14912 ^ n12969 ^ 1'b0 ;
  assign n33151 = n9108 & n33150 ;
  assign n33152 = n33151 ^ n18248 ^ 1'b0 ;
  assign n33153 = n6538 | n33152 ;
  assign n33149 = n7295 & n18041 ;
  assign n33154 = n33153 ^ n33149 ^ 1'b0 ;
  assign n33155 = n8579 ^ n2453 ^ 1'b0 ;
  assign n33156 = n31945 ^ n29543 ^ n8043 ;
  assign n33157 = n1659 & n4711 ;
  assign n33158 = n7051 ^ n615 ^ 1'b0 ;
  assign n33159 = ~n33157 & n33158 ;
  assign n33160 = n27587 & ~n33159 ;
  assign n33161 = ~n6893 & n31392 ;
  assign n33162 = n33161 ^ n26109 ^ n10122 ;
  assign n33165 = n13354 ^ n12000 ^ 1'b0 ;
  assign n33166 = n17773 & ~n33165 ;
  assign n33163 = ( n2914 & n6121 ) | ( n2914 & n32412 ) | ( n6121 & n32412 ) ;
  assign n33164 = n10646 & ~n33163 ;
  assign n33167 = n33166 ^ n33164 ^ 1'b0 ;
  assign n33168 = n18958 ^ n343 ^ 1'b0 ;
  assign n33169 = ~n326 & n7006 ;
  assign n33170 = n33169 ^ n5859 ^ 1'b0 ;
  assign n33171 = n17554 ^ n6102 ^ 1'b0 ;
  assign n33172 = ( n6960 & ~n10171 ) | ( n6960 & n16933 ) | ( ~n10171 & n16933 ) ;
  assign n33173 = n9177 ^ n8964 ^ 1'b0 ;
  assign n33174 = n18102 & ~n33173 ;
  assign n33175 = n12714 ^ n2621 ^ n947 ;
  assign n33176 = n33172 & ~n33175 ;
  assign n33177 = n10290 ^ n2822 ^ n588 ;
  assign n33178 = n3773 & n10403 ;
  assign n33179 = n33178 ^ n9408 ^ n6266 ;
  assign n33180 = n33179 ^ n19171 ^ n4502 ;
  assign n33181 = n33180 ^ n8683 ^ 1'b0 ;
  assign n33182 = n33177 & n33181 ;
  assign n33183 = n28755 ^ n3012 ^ 1'b0 ;
  assign n33184 = n4187 & ~n33183 ;
  assign n33185 = n9738 ^ n5934 ^ 1'b0 ;
  assign n33186 = n1185 & n33185 ;
  assign n33187 = n3212 | n15273 ;
  assign n33188 = n1938 | n33187 ;
  assign n33189 = ~n14748 & n33188 ;
  assign n33190 = n33186 & n33189 ;
  assign n33191 = n11550 ^ n7499 ^ 1'b0 ;
  assign n33192 = n3302 & ~n33191 ;
  assign n33193 = n33192 ^ n9345 ^ n7026 ;
  assign n33194 = n31207 ^ n18138 ^ 1'b0 ;
  assign n33195 = n33193 & ~n33194 ;
  assign n33199 = n3404 & n4402 ;
  assign n33200 = n33199 ^ n16293 ^ n8760 ;
  assign n33196 = n24200 ^ n22542 ^ n4617 ;
  assign n33197 = n15410 & ~n33196 ;
  assign n33198 = n33197 ^ n21566 ^ 1'b0 ;
  assign n33201 = n33200 ^ n33198 ^ n18976 ;
  assign n33202 = n3669 ^ n3075 ^ 1'b0 ;
  assign n33203 = n26677 | n33202 ;
  assign n33204 = ~n28373 & n30438 ;
  assign n33205 = n16413 & n33204 ;
  assign n33206 = n787 | n11301 ;
  assign n33207 = x129 & n22190 ;
  assign n33208 = n17838 & ~n19324 ;
  assign n33209 = n20987 ^ n9318 ^ 1'b0 ;
  assign n33210 = n490 & n33209 ;
  assign n33211 = n1862 & n33210 ;
  assign n33212 = ( n11085 & n33208 ) | ( n11085 & n33211 ) | ( n33208 & n33211 ) ;
  assign n33213 = n16429 & n19567 ;
  assign n33214 = n22691 & n33213 ;
  assign n33215 = n26380 & ~n33214 ;
  assign n33216 = n16961 | n19358 ;
  assign n33217 = n24545 ^ n16521 ^ n4699 ;
  assign n33218 = ( n14669 & n16087 ) | ( n14669 & ~n33217 ) | ( n16087 & ~n33217 ) ;
  assign n33219 = n15228 ^ n7179 ^ n2511 ;
  assign n33220 = n32571 ^ n15929 ^ 1'b0 ;
  assign n33221 = n18934 & n33220 ;
  assign n33222 = ~n12126 & n21310 ;
  assign n33223 = ( ~n2505 & n2777 ) | ( ~n2505 & n32018 ) | ( n2777 & n32018 ) ;
  assign n33224 = n32957 ^ n2754 ^ 1'b0 ;
  assign n33225 = n33224 ^ n21771 ^ 1'b0 ;
  assign n33226 = n13285 & ~n13467 ;
  assign n33227 = n33226 ^ n13017 ^ n8073 ;
  assign n33228 = n9145 | n33227 ;
  assign n33229 = n22835 & ~n31313 ;
  assign n33230 = n14685 & ~n33229 ;
  assign n33231 = ~n1566 & n27164 ;
  assign n33232 = ~n12703 & n33231 ;
  assign n33233 = n7942 ^ n4479 ^ 1'b0 ;
  assign n33234 = ~n302 & n12451 ;
  assign n33235 = n26328 & n33234 ;
  assign n33236 = n8821 | n33235 ;
  assign n33237 = n33236 ^ n21396 ^ 1'b0 ;
  assign n33238 = ( n16293 & n25453 ) | ( n16293 & ~n28166 ) | ( n25453 & ~n28166 ) ;
  assign n33239 = n19004 & n26841 ;
  assign n33240 = ( n3466 & n17753 ) | ( n3466 & n33239 ) | ( n17753 & n33239 ) ;
  assign n33241 = n33240 ^ n15469 ^ n11455 ;
  assign n33243 = n20808 ^ n6853 ^ 1'b0 ;
  assign n33244 = n20982 & ~n33243 ;
  assign n33242 = n10829 ^ n1804 ^ 1'b0 ;
  assign n33245 = n33244 ^ n33242 ^ 1'b0 ;
  assign n33246 = ~n22992 & n33245 ;
  assign n33247 = n2766 | n17049 ;
  assign n33248 = n24005 & ~n33247 ;
  assign n33249 = n16997 ^ n7607 ^ 1'b0 ;
  assign n33250 = n33249 ^ n27438 ^ 1'b0 ;
  assign n33251 = n26527 & n33250 ;
  assign n33252 = n18556 ^ n17969 ^ 1'b0 ;
  assign n33253 = n3449 ^ n1613 ^ 1'b0 ;
  assign n33254 = n9506 | n33253 ;
  assign n33255 = ~n7952 & n33254 ;
  assign n33256 = ( n25914 & n33252 ) | ( n25914 & ~n33255 ) | ( n33252 & ~n33255 ) ;
  assign n33257 = n32933 ^ n20927 ^ 1'b0 ;
  assign n33258 = ~n33256 & n33257 ;
  assign n33259 = n22427 ^ n10659 ^ n9457 ;
  assign n33260 = n11655 | n33259 ;
  assign n33261 = n26844 | n33260 ;
  assign n33262 = n25803 ^ n8940 ^ 1'b0 ;
  assign n33263 = n2111 & n33262 ;
  assign n33264 = n16346 ^ x73 ^ 1'b0 ;
  assign n33265 = n33263 & n33264 ;
  assign n33266 = n33265 ^ n2493 ^ 1'b0 ;
  assign n33267 = ( n5070 & n13866 ) | ( n5070 & ~n33266 ) | ( n13866 & ~n33266 ) ;
  assign n33268 = n31507 ^ n8100 ^ 1'b0 ;
  assign n33269 = n15715 ^ n3237 ^ 1'b0 ;
  assign n33270 = n23744 | n33269 ;
  assign n33271 = n820 | n20458 ;
  assign n33272 = n29232 ^ n22351 ^ 1'b0 ;
  assign n33273 = n33271 & n33272 ;
  assign n33274 = n4948 & n25557 ;
  assign n33275 = n26074 ^ n14068 ^ 1'b0 ;
  assign n33276 = n11545 & ~n33275 ;
  assign n33281 = n29914 ^ n9861 ^ n9523 ;
  assign n33282 = ( ~x129 & n14179 ) | ( ~x129 & n33281 ) | ( n14179 & n33281 ) ;
  assign n33277 = n16337 ^ n13081 ^ 1'b0 ;
  assign n33278 = n1170 | n33277 ;
  assign n33279 = ( n7854 & n28948 ) | ( n7854 & ~n33278 ) | ( n28948 & ~n33278 ) ;
  assign n33280 = ~n9775 & n33279 ;
  assign n33283 = n33282 ^ n33280 ^ 1'b0 ;
  assign n33284 = n30861 ^ n15534 ^ 1'b0 ;
  assign n33285 = ( n8632 & ~n14124 ) | ( n8632 & n24843 ) | ( ~n14124 & n24843 ) ;
  assign n33286 = ~n655 & n6351 ;
  assign n33287 = n2233 & ~n13041 ;
  assign n33288 = ~n6756 & n7303 ;
  assign n33289 = n3975 & n33288 ;
  assign n33290 = n1273 | n33289 ;
  assign n33291 = n33287 | n33290 ;
  assign n33292 = n23288 ^ n7766 ^ 1'b0 ;
  assign n33293 = n6879 & n33292 ;
  assign n33294 = n4991 | n5208 ;
  assign n33295 = n33294 ^ n2452 ^ 1'b0 ;
  assign n33296 = ( n1757 & n2764 ) | ( n1757 & n33295 ) | ( n2764 & n33295 ) ;
  assign n33297 = n20384 ^ n5057 ^ x24 ;
  assign n33298 = n33296 | n33297 ;
  assign n33299 = n33298 ^ n14153 ^ 1'b0 ;
  assign n33300 = n32175 ^ n21133 ^ 1'b0 ;
  assign n33301 = n19993 | n33300 ;
  assign n33302 = ~n16795 & n28129 ;
  assign n33303 = n6170 ^ n1382 ^ 1'b0 ;
  assign n33304 = n16558 & ~n33303 ;
  assign n33307 = n10805 ^ n3385 ^ 1'b0 ;
  assign n33308 = n17403 & ~n33307 ;
  assign n33309 = n33308 ^ n2551 ^ x128 ;
  assign n33310 = n33309 ^ n9037 ^ 1'b0 ;
  assign n33305 = n16505 ^ n10351 ^ 1'b0 ;
  assign n33306 = n17621 | n33305 ;
  assign n33311 = n33310 ^ n33306 ^ n7339 ;
  assign n33312 = n2064 & ~n20479 ;
  assign n33314 = n2700 | n27810 ;
  assign n33315 = n24146 | n33314 ;
  assign n33313 = n32587 ^ n11089 ^ 1'b0 ;
  assign n33316 = n33315 ^ n33313 ^ 1'b0 ;
  assign n33317 = ~n16596 & n30989 ;
  assign n33318 = n1000 & n33317 ;
  assign n33319 = n8298 ^ n3738 ^ 1'b0 ;
  assign n33320 = n2162 & ~n33319 ;
  assign n33321 = n27071 & n33320 ;
  assign n33322 = n1474 & ~n2738 ;
  assign n33323 = n33322 ^ x13 ^ 1'b0 ;
  assign n33324 = n26248 ^ n6260 ^ x158 ;
  assign n33325 = n17334 ^ n362 ^ 1'b0 ;
  assign n33326 = n33325 ^ n10313 ^ 1'b0 ;
  assign n33327 = ~n33324 & n33326 ;
  assign n33328 = n33327 ^ n4767 ^ 1'b0 ;
  assign n33329 = n4692 & n20864 ;
  assign n33330 = ( n4935 & n24668 ) | ( n4935 & n25915 ) | ( n24668 & n25915 ) ;
  assign n33331 = ( n29707 & ~n33329 ) | ( n29707 & n33330 ) | ( ~n33329 & n33330 ) ;
  assign n33332 = n1626 | n9516 ;
  assign n33333 = x243 | n33332 ;
  assign n33334 = n33333 ^ n31209 ^ 1'b0 ;
  assign n33335 = ~n7988 & n11228 ;
  assign n33336 = n12738 | n33335 ;
  assign n33337 = n8284 & n14881 ;
  assign n33338 = ~n31013 & n33337 ;
  assign n33339 = ~n7242 & n33338 ;
  assign n33340 = n30012 & ~n33339 ;
  assign n33341 = n932 | n9738 ;
  assign n33342 = n27453 ^ n7637 ^ 1'b0 ;
  assign n33343 = n1696 & ~n33342 ;
  assign n33344 = n33341 & n33343 ;
  assign n33345 = n11412 & ~n25103 ;
  assign n33346 = n33345 ^ x98 ^ 1'b0 ;
  assign n33347 = n8644 & ~n13531 ;
  assign n33348 = n5818 & n33347 ;
  assign n33349 = n33346 & n33348 ;
  assign n33350 = ~n1002 & n4230 ;
  assign n33351 = n33350 ^ n1110 ^ 1'b0 ;
  assign n33352 = n19724 | n33351 ;
  assign n33353 = n10949 | n20067 ;
  assign n33354 = n33353 ^ n12486 ^ 1'b0 ;
  assign n33355 = n20263 | n21864 ;
  assign n33356 = n2209 | n16553 ;
  assign n33357 = n17411 ^ n17111 ^ 1'b0 ;
  assign n33358 = ( n5002 & ~n13726 ) | ( n5002 & n33357 ) | ( ~n13726 & n33357 ) ;
  assign n33359 = ~n8633 & n16700 ;
  assign n33360 = n33359 ^ n24230 ^ 1'b0 ;
  assign n33361 = ~n17871 & n25681 ;
  assign n33362 = n18933 & n21597 ;
  assign n33363 = n3595 | n33362 ;
  assign n33364 = n33361 | n33363 ;
  assign n33365 = n2155 & ~n29603 ;
  assign n33366 = ( n10785 & ~n12362 ) | ( n10785 & n33365 ) | ( ~n12362 & n33365 ) ;
  assign n33367 = ( ~n6914 & n10370 ) | ( ~n6914 & n12933 ) | ( n10370 & n12933 ) ;
  assign n33368 = n22792 ^ n10509 ^ 1'b0 ;
  assign n33369 = n4215 | n33368 ;
  assign n33371 = n4623 ^ n1853 ^ 1'b0 ;
  assign n33372 = n8722 & n33371 ;
  assign n33370 = n10131 ^ n5400 ^ 1'b0 ;
  assign n33373 = n33372 ^ n33370 ^ 1'b0 ;
  assign n33374 = ~n888 & n5251 ;
  assign n33375 = n26744 ^ n22839 ^ 1'b0 ;
  assign n33376 = n17694 & ~n33375 ;
  assign n33377 = n17620 ^ n14415 ^ 1'b0 ;
  assign n33378 = n23835 ^ n8991 ^ 1'b0 ;
  assign n33379 = n8048 | n33378 ;
  assign n33380 = ( ~n7319 & n16172 ) | ( ~n7319 & n17426 ) | ( n16172 & n17426 ) ;
  assign n33381 = n3830 & n16461 ;
  assign n33382 = n16556 | n33381 ;
  assign n33383 = n16004 | n16841 ;
  assign n33384 = n4145 | n33383 ;
  assign n33385 = ( n1809 & n33382 ) | ( n1809 & ~n33384 ) | ( n33382 & ~n33384 ) ;
  assign n33386 = ~n9518 & n23377 ;
  assign n33387 = n28481 | n33386 ;
  assign n33388 = n21309 & n28625 ;
  assign n33389 = n33388 ^ n32926 ^ 1'b0 ;
  assign n33390 = n9349 & n17379 ;
  assign n33391 = n15294 & n33390 ;
  assign n33392 = n18280 | n33391 ;
  assign n33393 = n25872 & ~n33392 ;
  assign n33394 = n33016 ^ n28919 ^ 1'b0 ;
  assign n33395 = n27840 & ~n33394 ;
  assign n33396 = ~n4638 & n22699 ;
  assign n33397 = n33396 ^ n2897 ^ 1'b0 ;
  assign n33398 = n17632 | n25355 ;
  assign n33399 = n33398 ^ n19765 ^ 1'b0 ;
  assign n33400 = n21105 & ~n33399 ;
  assign n33402 = n4944 & ~n7871 ;
  assign n33401 = ~n30296 & n30899 ;
  assign n33403 = n33402 ^ n33401 ^ n3604 ;
  assign n33404 = n20292 ^ n11706 ^ 1'b0 ;
  assign n33405 = n20819 & ~n33404 ;
  assign n33406 = n23212 ^ n22330 ^ n15526 ;
  assign n33407 = n7184 ^ n6011 ^ 1'b0 ;
  assign n33408 = ~n33406 & n33407 ;
  assign n33409 = n11914 & n33408 ;
  assign n33410 = n12315 & n33409 ;
  assign n33411 = n15632 ^ n12922 ^ 1'b0 ;
  assign n33412 = n2994 & ~n24168 ;
  assign n33413 = n6612 & n33412 ;
  assign n33414 = ( n9052 & n25647 ) | ( n9052 & n33413 ) | ( n25647 & n33413 ) ;
  assign n33415 = n1963 & n32639 ;
  assign n33416 = n33414 | n33415 ;
  assign n33421 = n738 & n18250 ;
  assign n33417 = ( ~x13 & n16864 ) | ( ~x13 & n23584 ) | ( n16864 & n23584 ) ;
  assign n33418 = n12710 ^ n9916 ^ n4316 ;
  assign n33419 = n20265 | n33418 ;
  assign n33420 = n33417 & ~n33419 ;
  assign n33422 = n33421 ^ n33420 ^ n13241 ;
  assign n33423 = n2216 & n14565 ;
  assign n33424 = ~n18837 & n33423 ;
  assign n33425 = n33424 ^ n2061 ^ 1'b0 ;
  assign n33426 = n2763 & n15447 ;
  assign n33427 = n33426 ^ n30161 ^ 1'b0 ;
  assign n33428 = n24663 ^ n23201 ^ n16443 ;
  assign n33429 = n19622 ^ n3519 ^ 1'b0 ;
  assign n33430 = n9866 & ~n33429 ;
  assign n33431 = ~n3759 & n33430 ;
  assign n33432 = ~n33428 & n33431 ;
  assign n33434 = n24189 ^ n15331 ^ n10486 ;
  assign n33433 = n28939 ^ n6846 ^ 1'b0 ;
  assign n33435 = n33434 ^ n33433 ^ 1'b0 ;
  assign n33436 = n16796 ^ n8103 ^ 1'b0 ;
  assign n33437 = n29498 ^ n23029 ^ n8062 ;
  assign n33438 = n15321 | n25249 ;
  assign n33439 = n33438 ^ n2097 ^ 1'b0 ;
  assign n33440 = n23163 ^ n5197 ^ 1'b0 ;
  assign n33441 = n2192 | n3255 ;
  assign n33442 = n3667 & n33441 ;
  assign n33443 = n13391 & n33442 ;
  assign n33444 = n3404 & n10603 ;
  assign n33445 = n19302 & n33444 ;
  assign n33446 = n9897 | n17030 ;
  assign n33447 = n6734 & ~n33446 ;
  assign n33448 = n33445 & n33447 ;
  assign n33449 = n8544 & n13275 ;
  assign n33450 = n33449 ^ n12883 ^ n9024 ;
  assign n33451 = n33450 ^ n26495 ^ 1'b0 ;
  assign n33452 = n33448 & ~n33451 ;
  assign n33453 = n17059 & ~n19650 ;
  assign n33454 = n33453 ^ n8057 ^ n2547 ;
  assign n33455 = n3093 & n5522 ;
  assign n33456 = n5929 & n33455 ;
  assign n33457 = ( n26349 & n30867 ) | ( n26349 & n33456 ) | ( n30867 & n33456 ) ;
  assign n33458 = n3848 ^ n1613 ^ 1'b0 ;
  assign n33459 = n20934 | n26997 ;
  assign n33460 = n6854 ^ n3423 ^ 1'b0 ;
  assign n33461 = n14546 & n33460 ;
  assign n33462 = n33461 ^ n913 ^ 1'b0 ;
  assign n33463 = n33462 ^ n14566 ^ 1'b0 ;
  assign n33464 = n16473 ^ n15808 ^ n11425 ;
  assign n33465 = ( n12065 & n31397 ) | ( n12065 & ~n33464 ) | ( n31397 & ~n33464 ) ;
  assign n33466 = n26128 ^ n21004 ^ 1'b0 ;
  assign n33469 = ~n1042 & n4815 ;
  assign n33470 = n33469 ^ n310 ^ 1'b0 ;
  assign n33467 = ( n2222 & n5525 ) | ( n2222 & n16993 ) | ( n5525 & n16993 ) ;
  assign n33468 = n8603 | n33467 ;
  assign n33471 = n33470 ^ n33468 ^ 1'b0 ;
  assign n33472 = n14328 ^ n10527 ^ 1'b0 ;
  assign n33473 = ~n15266 & n33472 ;
  assign n33474 = n1110 & n7277 ;
  assign n33475 = ~n33473 & n33474 ;
  assign n33476 = n19738 ^ n14274 ^ 1'b0 ;
  assign n33477 = ~n19621 & n33476 ;
  assign n33478 = n495 & n6261 ;
  assign n33479 = n33478 ^ n26639 ^ n19915 ;
  assign n33480 = ( n3424 & n26241 ) | ( n3424 & n26256 ) | ( n26241 & n26256 ) ;
  assign n33481 = n11053 ^ n2086 ^ 1'b0 ;
  assign n33482 = n28370 | n33481 ;
  assign n33483 = n23981 ^ n393 ^ 1'b0 ;
  assign n33484 = n5057 & ~n33483 ;
  assign n33485 = n668 | n3931 ;
  assign n33486 = n668 & ~n33485 ;
  assign n33487 = n1995 & n4625 ;
  assign n33488 = ~n1995 & n33487 ;
  assign n33489 = n14938 | n33488 ;
  assign n33490 = n33486 & ~n33489 ;
  assign n33491 = ~n4227 & n8647 ;
  assign n33492 = n33490 & n33491 ;
  assign n33493 = n951 & n19709 ;
  assign n33494 = n33492 | n33493 ;
  assign n33495 = n33492 & ~n33494 ;
  assign n33496 = n33495 ^ n4437 ^ 1'b0 ;
  assign n33497 = ~n1457 & n33496 ;
  assign n33498 = n6640 ^ n5085 ^ 1'b0 ;
  assign n33499 = ~n8971 & n33498 ;
  assign n33500 = ~n5365 & n33499 ;
  assign n33501 = n29163 ^ n6915 ^ 1'b0 ;
  assign n33502 = n19823 | n33501 ;
  assign n33503 = n33502 ^ n6646 ^ n4053 ;
  assign n33504 = ( n2041 & n33500 ) | ( n2041 & ~n33503 ) | ( n33500 & ~n33503 ) ;
  assign n33505 = ( n19675 & n33497 ) | ( n19675 & ~n33504 ) | ( n33497 & ~n33504 ) ;
  assign n33506 = n33484 & n33505 ;
  assign n33507 = n33506 ^ n3292 ^ 1'b0 ;
  assign n33508 = ~n8023 & n12037 ;
  assign n33509 = n33508 ^ n17999 ^ n11796 ;
  assign n33510 = n16275 ^ n1804 ^ 1'b0 ;
  assign n33511 = n33510 ^ n19393 ^ n11977 ;
  assign n33512 = n24002 ^ n9530 ^ 1'b0 ;
  assign n33513 = ( ~n15401 & n29694 ) | ( ~n15401 & n33512 ) | ( n29694 & n33512 ) ;
  assign n33514 = n32671 & ~n33513 ;
  assign n33515 = n33514 ^ n3638 ^ 1'b0 ;
  assign n33516 = n21217 ^ n17851 ^ n5914 ;
  assign n33517 = n33516 ^ n20040 ^ 1'b0 ;
  assign n33518 = n4544 & ~n7761 ;
  assign n33519 = n33518 ^ n16014 ^ 1'b0 ;
  assign n33520 = n17542 | n33519 ;
  assign n33521 = n33517 & ~n33520 ;
  assign n33522 = n1634 & ~n26224 ;
  assign n33523 = ~n11715 & n33522 ;
  assign n33524 = n31721 ^ n2488 ^ 1'b0 ;
  assign n33525 = n5190 & n33524 ;
  assign n33526 = n12315 | n30895 ;
  assign n33527 = n24848 ^ n6981 ^ n2080 ;
  assign n33528 = n7066 & ~n19874 ;
  assign n33529 = n1250 & ~n6125 ;
  assign n33530 = n1979 & n33529 ;
  assign n33531 = n29227 ^ n25442 ^ 1'b0 ;
  assign n33532 = n25819 & ~n33531 ;
  assign n33533 = n15744 ^ n13793 ^ 1'b0 ;
  assign n33534 = n33532 & n33533 ;
  assign n33535 = n33530 | n33534 ;
  assign n33536 = n12971 ^ n4243 ^ 1'b0 ;
  assign n33537 = n18656 & n33536 ;
  assign n33538 = ~n9139 & n11139 ;
  assign n33539 = ~n4496 & n33538 ;
  assign n33540 = n31129 ^ n1281 ^ 1'b0 ;
  assign n33541 = n292 | n14460 ;
  assign n33542 = n12450 & ~n25613 ;
  assign n33543 = n33542 ^ n7584 ^ 1'b0 ;
  assign n33544 = ( n17663 & ~n33541 ) | ( n17663 & n33543 ) | ( ~n33541 & n33543 ) ;
  assign n33545 = n5775 | n14452 ;
  assign n33546 = n24629 & ~n33545 ;
  assign n33547 = n33546 ^ n21417 ^ 1'b0 ;
  assign n33548 = n5412 ^ n4304 ^ 1'b0 ;
  assign n33549 = ( n8303 & n20119 ) | ( n8303 & ~n29490 ) | ( n20119 & ~n29490 ) ;
  assign n33550 = n33549 ^ n2259 ^ 1'b0 ;
  assign n33551 = n3794 ^ n2892 ^ 1'b0 ;
  assign n33552 = n7425 | n33551 ;
  assign n33553 = n5905 | n26872 ;
  assign n33554 = n33552 & ~n33553 ;
  assign n33555 = n2354 | n12744 ;
  assign n33556 = n3197 & n33555 ;
  assign n33557 = n6204 & n33556 ;
  assign n33558 = n8089 & n12711 ;
  assign n33559 = ( n3156 & n10419 ) | ( n3156 & ~n23884 ) | ( n10419 & ~n23884 ) ;
  assign n33560 = n13338 & ~n33559 ;
  assign n33563 = n4132 ^ n1844 ^ 1'b0 ;
  assign n33564 = n3953 & n19645 ;
  assign n33565 = n33563 & n33564 ;
  assign n33561 = n1766 | n13545 ;
  assign n33562 = ~n18693 & n33561 ;
  assign n33566 = n33565 ^ n33562 ^ 1'b0 ;
  assign n33567 = ( n10968 & n16580 ) | ( n10968 & ~n33566 ) | ( n16580 & ~n33566 ) ;
  assign n33568 = n19761 ^ n3093 ^ 1'b0 ;
  assign n33569 = n33568 ^ n12137 ^ 1'b0 ;
  assign n33570 = n20938 | n33569 ;
  assign n33571 = n16750 ^ n16101 ^ 1'b0 ;
  assign n33572 = ~n1709 & n4617 ;
  assign n33573 = n33572 ^ n13170 ^ n10234 ;
  assign n33574 = ~n32098 & n33573 ;
  assign n33575 = ~n25258 & n33574 ;
  assign n33576 = n18894 & ~n31961 ;
  assign n33577 = n7720 | n20080 ;
  assign n33578 = n33577 ^ n15382 ^ 1'b0 ;
  assign n33579 = n19709 ^ n13017 ^ n10117 ;
  assign n33580 = n33579 ^ n30733 ^ 1'b0 ;
  assign n33581 = n12657 ^ n1430 ^ 1'b0 ;
  assign n33582 = ~n4091 & n33581 ;
  assign n33583 = ~n18174 & n33582 ;
  assign n33584 = ( ~x12 & n11963 ) | ( ~x12 & n23862 ) | ( n11963 & n23862 ) ;
  assign n33585 = n33584 ^ n3005 ^ n2903 ;
  assign n33586 = n25853 ^ n2970 ^ 1'b0 ;
  assign n33587 = n3928 & n33586 ;
  assign n33588 = n33587 ^ n13152 ^ n3196 ;
  assign n33589 = n33585 & n33588 ;
  assign n33590 = n6962 ^ n5901 ^ 1'b0 ;
  assign n33591 = n21694 ^ n9525 ^ 1'b0 ;
  assign n33592 = ( ~n652 & n33590 ) | ( ~n652 & n33591 ) | ( n33590 & n33591 ) ;
  assign n33593 = n9944 | n33592 ;
  assign n33594 = n33593 ^ n1933 ^ 1'b0 ;
  assign n33595 = n4426 & ~n33594 ;
  assign n33596 = n31543 ^ n6209 ^ n1602 ;
  assign n33597 = n9073 ^ n3865 ^ 1'b0 ;
  assign n33598 = ~n19154 & n33597 ;
  assign n33599 = n33598 ^ n20723 ^ n9333 ;
  assign n33600 = n7570 ^ n5875 ^ 1'b0 ;
  assign n33601 = ~n15934 & n33600 ;
  assign n33602 = n15689 ^ n6623 ^ 1'b0 ;
  assign n33603 = ( n33599 & n33601 ) | ( n33599 & ~n33602 ) | ( n33601 & ~n33602 ) ;
  assign n33604 = n33603 ^ n21013 ^ 1'b0 ;
  assign n33605 = n3203 & ~n11973 ;
  assign n33606 = n11788 | n31729 ;
  assign n33607 = n3914 & ~n33606 ;
  assign n33608 = n21567 ^ n11631 ^ n3506 ;
  assign n33609 = n2272 | n3053 ;
  assign n33610 = ~n33608 & n33609 ;
  assign n33611 = ~n25052 & n33610 ;
  assign n33612 = n33167 ^ n27798 ^ 1'b0 ;
  assign n33613 = ~n33611 & n33612 ;
  assign n33614 = ( n600 & n5486 ) | ( n600 & n17091 ) | ( n5486 & n17091 ) ;
  assign n33615 = n16303 & n33614 ;
  assign n33616 = n33615 ^ x59 ^ 1'b0 ;
  assign n33618 = n17907 ^ n6557 ^ 1'b0 ;
  assign n33619 = n12370 & n33618 ;
  assign n33617 = n8163 & ~n12865 ;
  assign n33620 = n33619 ^ n33617 ^ n21404 ;
  assign n33621 = n28393 ^ x90 ^ 1'b0 ;
  assign n33624 = n14953 ^ n7622 ^ n365 ;
  assign n33625 = n3061 & n33624 ;
  assign n33622 = n32682 ^ n14761 ^ 1'b0 ;
  assign n33623 = ( ~n3056 & n18568 ) | ( ~n3056 & n33622 ) | ( n18568 & n33622 ) ;
  assign n33626 = n33625 ^ n33623 ^ n12849 ;
  assign n33627 = ( ~n2340 & n3345 ) | ( ~n2340 & n10900 ) | ( n3345 & n10900 ) ;
  assign n33628 = n20814 ^ n15686 ^ n12004 ;
  assign n33629 = n33627 & ~n33628 ;
  assign n33630 = n3191 & ~n33629 ;
  assign n33631 = n5441 & ~n23728 ;
  assign n33632 = ~n2405 & n33631 ;
  assign n33633 = n21833 ^ n9159 ^ 1'b0 ;
  assign n33634 = n26793 & n33633 ;
  assign n33637 = n22923 ^ n1201 ^ 1'b0 ;
  assign n33635 = ~n7055 & n13591 ;
  assign n33636 = n33635 ^ n18807 ^ 1'b0 ;
  assign n33638 = n33637 ^ n33636 ^ n6413 ;
  assign n33639 = ( ~n8183 & n17494 ) | ( ~n8183 & n22788 ) | ( n17494 & n22788 ) ;
  assign n33640 = n4644 ^ n4089 ^ 1'b0 ;
  assign n33641 = n6710 & n23914 ;
  assign n33642 = ~n33640 & n33641 ;
  assign n33643 = n31723 ^ n27950 ^ 1'b0 ;
  assign n33644 = n33643 ^ n3705 ^ 1'b0 ;
  assign n33645 = n14528 & ~n33644 ;
  assign n33647 = ( n8069 & n8398 ) | ( n8069 & n18454 ) | ( n8398 & n18454 ) ;
  assign n33646 = ~n4712 & n10243 ;
  assign n33648 = n33647 ^ n33646 ^ 1'b0 ;
  assign n33649 = ~n17630 & n26974 ;
  assign n33650 = n5073 ^ n1728 ^ 1'b0 ;
  assign n33651 = n33650 ^ n28167 ^ n2724 ;
  assign n33652 = n33651 ^ n6792 ^ 1'b0 ;
  assign n33653 = n14966 & ~n24086 ;
  assign n33654 = n29849 | n33653 ;
  assign n33655 = n33654 ^ n20936 ^ 1'b0 ;
  assign n33656 = n17429 & ~n33655 ;
  assign n33657 = n21314 ^ n17894 ^ n7825 ;
  assign n33658 = n19960 ^ n3379 ^ 1'b0 ;
  assign n33659 = n17607 ^ n12234 ^ n10628 ;
  assign n33660 = n11500 & n20043 ;
  assign n33661 = n33660 ^ n29534 ^ 1'b0 ;
  assign n33662 = n25317 ^ n17835 ^ 1'b0 ;
  assign n33663 = n4402 | n33662 ;
  assign n33664 = n13527 & ~n33663 ;
  assign n33665 = ~n33661 & n33664 ;
  assign n33666 = n7437 ^ n2763 ^ 1'b0 ;
  assign n33667 = n33666 ^ n9423 ^ 1'b0 ;
  assign n33668 = n6938 & ~n33667 ;
  assign n33669 = n9381 ^ n7078 ^ 1'b0 ;
  assign n33670 = n33669 ^ n29922 ^ n21661 ;
  assign n33671 = ~n2997 & n33670 ;
  assign n33672 = ~n13659 & n33671 ;
  assign n33673 = ~n15794 & n23505 ;
  assign n33674 = n26704 ^ n9266 ^ n7488 ;
  assign n33675 = ( n7769 & n25424 ) | ( n7769 & n33674 ) | ( n25424 & n33674 ) ;
  assign n33676 = n18280 | n25677 ;
  assign n33677 = n10150 | n33676 ;
  assign n33678 = ( n3300 & n16601 ) | ( n3300 & ~n33677 ) | ( n16601 & ~n33677 ) ;
  assign n33679 = n33678 ^ n33293 ^ 1'b0 ;
  assign n33680 = ~n8993 & n33679 ;
  assign n33681 = n4203 & n4700 ;
  assign n33682 = n33681 ^ n24266 ^ 1'b0 ;
  assign n33683 = n29179 & ~n33622 ;
  assign n33684 = n15063 | n20170 ;
  assign n33685 = ~n5660 & n10826 ;
  assign n33686 = n28142 | n33685 ;
  assign n33687 = n459 & n13582 ;
  assign n33688 = n17159 & n21951 ;
  assign n33689 = n33688 ^ n12202 ^ 1'b0 ;
  assign n33690 = ( n1758 & ~n3139 ) | ( n1758 & n20273 ) | ( ~n3139 & n20273 ) ;
  assign n33691 = n11967 & n33690 ;
  assign n33692 = n33691 ^ n20403 ^ 1'b0 ;
  assign n33694 = n4685 & n13609 ;
  assign n33695 = n10781 ^ n9957 ^ 1'b0 ;
  assign n33696 = n33694 & ~n33695 ;
  assign n33693 = n19629 & n30434 ;
  assign n33697 = n33696 ^ n33693 ^ 1'b0 ;
  assign n33698 = n32344 ^ n826 ^ 1'b0 ;
  assign n33699 = n33698 ^ n27664 ^ n15625 ;
  assign n33700 = n28373 ^ n5935 ^ 1'b0 ;
  assign n33701 = ~n19792 & n29909 ;
  assign n33702 = ~n10961 & n33701 ;
  assign n33703 = n7592 & ~n29353 ;
  assign n33704 = n33703 ^ n1946 ^ 1'b0 ;
  assign n33705 = ~n14407 & n33704 ;
  assign n33706 = ~n27622 & n33705 ;
  assign n33707 = n28271 & ~n28598 ;
  assign n33708 = n11187 & n33707 ;
  assign n33709 = ( x235 & ~n300 ) | ( x235 & n26499 ) | ( ~n300 & n26499 ) ;
  assign n33710 = ~n2464 & n12003 ;
  assign n33711 = n2754 & n33710 ;
  assign n33712 = n22117 & ~n33711 ;
  assign n33714 = n655 & ~n5305 ;
  assign n33715 = n33714 ^ x69 ^ 1'b0 ;
  assign n33716 = n15431 | n33715 ;
  assign n33717 = n33716 ^ n21565 ^ 1'b0 ;
  assign n33713 = ~n9642 & n14146 ;
  assign n33718 = n33717 ^ n33713 ^ 1'b0 ;
  assign n33719 = n4838 & n10628 ;
  assign n33720 = n8958 & n33719 ;
  assign n33721 = n33720 ^ n19196 ^ n5588 ;
  assign n33722 = ~n4177 & n28359 ;
  assign n33723 = ( n690 & n9931 ) | ( n690 & ~n22420 ) | ( n9931 & ~n22420 ) ;
  assign n33724 = n451 & n33723 ;
  assign n33725 = n33724 ^ n29209 ^ n5979 ;
  assign n33726 = ~n8013 & n25010 ;
  assign n33727 = n10661 & n33726 ;
  assign n33728 = n4282 | n33727 ;
  assign n33729 = n30161 & ~n33728 ;
  assign n33730 = n2219 & n20328 ;
  assign n33731 = n5054 | n12206 ;
  assign n33732 = n33730 | n33731 ;
  assign n33733 = ( n12985 & n33729 ) | ( n12985 & n33732 ) | ( n33729 & n33732 ) ;
  assign n33737 = n14328 ^ n14252 ^ 1'b0 ;
  assign n33738 = ~n14781 & n33737 ;
  assign n33739 = ~n4995 & n33738 ;
  assign n33740 = n33739 ^ n19503 ^ 1'b0 ;
  assign n33741 = n7470 & ~n33740 ;
  assign n33742 = n33741 ^ n835 ^ 1'b0 ;
  assign n33734 = n13795 ^ n1655 ^ n1377 ;
  assign n33735 = n33734 ^ n12136 ^ n2439 ;
  assign n33736 = n24862 & ~n33735 ;
  assign n33743 = n33742 ^ n33736 ^ 1'b0 ;
  assign n33744 = n1462 & ~n16173 ;
  assign n33745 = n33744 ^ n2589 ^ 1'b0 ;
  assign n33746 = n4364 | n33745 ;
  assign n33747 = n33746 ^ n25732 ^ 1'b0 ;
  assign n33748 = n7678 ^ n4512 ^ 1'b0 ;
  assign n33749 = n29057 & n33748 ;
  assign n33750 = ( ~n6240 & n6580 ) | ( ~n6240 & n21840 ) | ( n6580 & n21840 ) ;
  assign n33751 = n19919 ^ n4679 ^ n2445 ;
  assign n33752 = n33751 ^ n31444 ^ 1'b0 ;
  assign n33753 = n22226 & n29040 ;
  assign n33754 = n17059 ^ n7068 ^ 1'b0 ;
  assign n33755 = n33753 & ~n33754 ;
  assign n33756 = n1357 | n14789 ;
  assign n33757 = n10459 & n33756 ;
  assign n33758 = n22665 ^ n2549 ^ 1'b0 ;
  assign n33759 = ~n6191 & n14227 ;
  assign n33760 = ~n21266 & n33759 ;
  assign n33761 = n5364 & ~n21183 ;
  assign n33762 = n10794 | n14635 ;
  assign n33763 = n33762 ^ n10124 ^ 1'b0 ;
  assign n33764 = n33763 ^ n20484 ^ 1'b0 ;
  assign n33765 = n10170 & n24965 ;
  assign n33766 = n33765 ^ n15389 ^ 1'b0 ;
  assign n33767 = ( ~n8651 & n9005 ) | ( ~n8651 & n13209 ) | ( n9005 & n13209 ) ;
  assign n33768 = n10974 ^ n6580 ^ 1'b0 ;
  assign n33769 = n33767 & n33768 ;
  assign n33770 = ~n2355 & n16163 ;
  assign n33771 = ( ~n1487 & n20898 ) | ( ~n1487 & n21762 ) | ( n20898 & n21762 ) ;
  assign n33772 = n22165 | n33771 ;
  assign n33773 = ~n5094 & n18163 ;
  assign n33774 = ( n5368 & n12865 ) | ( n5368 & n27917 ) | ( n12865 & n27917 ) ;
  assign n33775 = ( n18997 & ~n33773 ) | ( n18997 & n33774 ) | ( ~n33773 & n33774 ) ;
  assign n33780 = n21365 ^ n8582 ^ n5479 ;
  assign n33779 = n22208 ^ n5366 ^ n4341 ;
  assign n33781 = n33780 ^ n33779 ^ n19345 ;
  assign n33776 = ( n9879 & ~n13231 ) | ( n9879 & n16736 ) | ( ~n13231 & n16736 ) ;
  assign n33777 = n33776 ^ n24603 ^ 1'b0 ;
  assign n33778 = n33777 ^ n15331 ^ n11332 ;
  assign n33782 = n33781 ^ n33778 ^ n1353 ;
  assign n33783 = n341 & ~n17537 ;
  assign n33784 = n33783 ^ n21477 ^ 1'b0 ;
  assign n33785 = ~n12829 & n21463 ;
  assign n33786 = n19923 ^ n1508 ^ 1'b0 ;
  assign n33787 = n33785 | n33786 ;
  assign n33788 = n33787 ^ n4694 ^ 1'b0 ;
  assign n33789 = n33784 & n33788 ;
  assign n33790 = ~n23785 & n24263 ;
  assign n33791 = n33790 ^ n15530 ^ 1'b0 ;
  assign n33792 = n12746 | n16668 ;
  assign n33793 = n33792 ^ n5611 ^ 1'b0 ;
  assign n33794 = ( n15177 & ~n24418 ) | ( n15177 & n33793 ) | ( ~n24418 & n33793 ) ;
  assign n33795 = n21287 & n33794 ;
  assign n33796 = n33795 ^ n31418 ^ 1'b0 ;
  assign n33797 = n10046 | n14275 ;
  assign n33798 = n4425 | n33797 ;
  assign n33799 = n7875 & n19600 ;
  assign n33800 = n26483 | n33799 ;
  assign n33801 = n33800 ^ n29257 ^ n11611 ;
  assign n33802 = n21782 ^ n10326 ^ n2871 ;
  assign n33803 = ~n9776 & n16286 ;
  assign n33804 = n4229 ^ n2102 ^ 1'b0 ;
  assign n33805 = n13060 ^ n12129 ^ 1'b0 ;
  assign n33806 = n33804 & n33805 ;
  assign n33807 = n27652 | n33806 ;
  assign n33808 = ~n3023 & n33807 ;
  assign n33809 = n26759 ^ n7718 ^ 1'b0 ;
  assign n33810 = n17858 & n33809 ;
  assign n33811 = ( n565 & n2362 ) | ( n565 & ~n5830 ) | ( n2362 & ~n5830 ) ;
  assign n33812 = ~n17303 & n33811 ;
  assign n33813 = ( x120 & n12664 ) | ( x120 & ~n33812 ) | ( n12664 & ~n33812 ) ;
  assign n33814 = n33813 ^ n10431 ^ 1'b0 ;
  assign n33815 = n33810 & ~n33814 ;
  assign n33816 = n4468 | n10582 ;
  assign n33817 = n3821 & ~n33816 ;
  assign n33818 = n31890 ^ n21904 ^ 1'b0 ;
  assign n33819 = n402 | n33818 ;
  assign n33820 = n21048 ^ n2972 ^ 1'b0 ;
  assign n33821 = n20116 & n33820 ;
  assign n33822 = n20282 & ~n21957 ;
  assign n33823 = n6968 | n33822 ;
  assign n33824 = n28866 ^ n16349 ^ 1'b0 ;
  assign n33825 = ( n25769 & n30845 ) | ( n25769 & ~n33824 ) | ( n30845 & ~n33824 ) ;
  assign n33826 = n21637 & n30148 ;
  assign n33827 = n18243 & n33826 ;
  assign n33828 = n14274 | n30898 ;
  assign n33829 = n18070 ^ n16444 ^ 1'b0 ;
  assign n33830 = ~n33828 & n33829 ;
  assign n33831 = n33830 ^ n517 ^ 1'b0 ;
  assign n33832 = n19180 ^ n8984 ^ n390 ;
  assign n33833 = n15525 & ~n17614 ;
  assign n33834 = ~n8614 & n19629 ;
  assign n33835 = ~n21691 & n33834 ;
  assign n33836 = n33835 ^ n31224 ^ n19072 ;
  assign n33837 = ( n1423 & n2111 ) | ( n1423 & n11034 ) | ( n2111 & n11034 ) ;
  assign n33838 = n2598 & n33837 ;
  assign n33839 = n12483 & ~n33838 ;
  assign n33840 = n19695 ^ n11714 ^ 1'b0 ;
  assign n33841 = n1781 | n33840 ;
  assign n33842 = n795 & n27018 ;
  assign n33849 = ~n2172 & n20737 ;
  assign n33850 = n32915 & n33849 ;
  assign n33843 = n11357 | n15257 ;
  assign n33844 = n25237 ^ n1999 ^ 1'b0 ;
  assign n33845 = ~n33843 & n33844 ;
  assign n33846 = n8025 ^ x222 ^ 1'b0 ;
  assign n33847 = n33845 & n33846 ;
  assign n33848 = ( n14212 & ~n26349 ) | ( n14212 & n33847 ) | ( ~n26349 & n33847 ) ;
  assign n33851 = n33850 ^ n33848 ^ n21900 ;
  assign n33852 = n3999 | n21555 ;
  assign n33853 = n33852 ^ n6922 ^ 1'b0 ;
  assign n33854 = ( ~n3885 & n11934 ) | ( ~n3885 & n25942 ) | ( n11934 & n25942 ) ;
  assign n33855 = n19875 | n25396 ;
  assign n33856 = ( n2822 & n33854 ) | ( n2822 & ~n33855 ) | ( n33854 & ~n33855 ) ;
  assign n33857 = n2524 & n33856 ;
  assign n33858 = n20175 & n33857 ;
  assign n33859 = n23970 | n25277 ;
  assign n33860 = n33859 ^ n8812 ^ 1'b0 ;
  assign n33861 = ~n1359 & n6119 ;
  assign n33862 = ~n8278 & n33861 ;
  assign n33863 = n33862 ^ n32926 ^ n21344 ;
  assign n33864 = n13248 | n24915 ;
  assign n33865 = n33864 ^ n24058 ^ n8276 ;
  assign n33866 = n1867 & n21297 ;
  assign n33867 = ~n22982 & n33866 ;
  assign n33868 = n6777 ^ n6692 ^ 1'b0 ;
  assign n33869 = n20456 ^ n14321 ^ 1'b0 ;
  assign n33870 = ( n829 & n11905 ) | ( n829 & ~n33869 ) | ( n11905 & ~n33869 ) ;
  assign n33871 = n13896 & ~n23869 ;
  assign n33872 = n30873 ^ n4154 ^ 1'b0 ;
  assign n33873 = ~n4725 & n33872 ;
  assign n33874 = n18120 ^ n3445 ^ 1'b0 ;
  assign n33875 = n18238 ^ n5014 ^ 1'b0 ;
  assign n33876 = n16488 ^ n4462 ^ 1'b0 ;
  assign n33877 = ~n16427 & n33876 ;
  assign n33878 = n33875 & n33877 ;
  assign n33879 = ~n6670 & n24678 ;
  assign n33880 = n4184 | n5355 ;
  assign n33881 = ~n493 & n33880 ;
  assign n33882 = n22868 ^ n11844 ^ n7968 ;
  assign n33883 = n15250 ^ n8389 ^ 1'b0 ;
  assign n33884 = ~n8430 & n33883 ;
  assign n33885 = ~n18270 & n33884 ;
  assign n33886 = n11615 ^ n7336 ^ 1'b0 ;
  assign n33887 = n3467 & ~n30392 ;
  assign n33888 = ~n663 & n33887 ;
  assign n33890 = n29273 ^ n14186 ^ 1'b0 ;
  assign n33891 = n19575 ^ n10763 ^ n482 ;
  assign n33892 = n33890 & n33891 ;
  assign n33889 = n24226 ^ n22302 ^ 1'b0 ;
  assign n33893 = n33892 ^ n33889 ^ n32058 ;
  assign n33894 = n33893 ^ n13706 ^ 1'b0 ;
  assign n33895 = n19557 & n33894 ;
  assign n33896 = n24265 ^ n604 ^ 1'b0 ;
  assign n33897 = n15074 & n33896 ;
  assign n33898 = n33897 ^ n7792 ^ 1'b0 ;
  assign n33899 = n33898 ^ n12617 ^ 1'b0 ;
  assign n33900 = n19037 ^ n6597 ^ n3231 ;
  assign n33901 = n1963 & ~n12939 ;
  assign n33902 = ( ~n3637 & n21285 ) | ( ~n3637 & n33901 ) | ( n21285 & n33901 ) ;
  assign n33905 = n14651 ^ n4768 ^ 1'b0 ;
  assign n33903 = n9485 | n13592 ;
  assign n33904 = n23089 & ~n33903 ;
  assign n33906 = n33905 ^ n33904 ^ 1'b0 ;
  assign n33907 = n25512 & ~n32758 ;
  assign n33908 = n33907 ^ n17146 ^ 1'b0 ;
  assign n33909 = n530 | n14145 ;
  assign n33910 = n22296 | n33909 ;
  assign n33911 = ( ~n5237 & n6031 ) | ( ~n5237 & n7120 ) | ( n6031 & n7120 ) ;
  assign n33912 = ( ~n3755 & n7569 ) | ( ~n3755 & n9062 ) | ( n7569 & n9062 ) ;
  assign n33913 = ~n33911 & n33912 ;
  assign n33914 = n5472 & n13749 ;
  assign n33915 = n33914 ^ n4390 ^ 1'b0 ;
  assign n33916 = ~n31470 & n33915 ;
  assign n33917 = n33916 ^ n29797 ^ 1'b0 ;
  assign n33918 = ( n3958 & n8853 ) | ( n3958 & ~n33917 ) | ( n8853 & ~n33917 ) ;
  assign n33919 = n9240 & n24420 ;
  assign n33920 = n33919 ^ n26759 ^ n22208 ;
  assign n33921 = n4812 & ~n6135 ;
  assign n33922 = n33921 ^ n25662 ^ 1'b0 ;
  assign n33923 = n292 & ~n15941 ;
  assign n33924 = n953 & n19656 ;
  assign n33929 = n6254 & ~n20303 ;
  assign n33925 = n30845 ^ n28970 ^ 1'b0 ;
  assign n33926 = n25646 & n33925 ;
  assign n33927 = n15629 & ~n33926 ;
  assign n33928 = n26946 & ~n33927 ;
  assign n33930 = n33929 ^ n33928 ^ 1'b0 ;
  assign n33931 = n4461 ^ n2032 ^ n1434 ;
  assign n33932 = ~n28379 & n33931 ;
  assign n33933 = ~n3352 & n33932 ;
  assign n33934 = n5674 & n27158 ;
  assign n33935 = n33934 ^ n9787 ^ 1'b0 ;
  assign n33936 = n33935 ^ n20606 ^ n1499 ;
  assign n33937 = n2259 & ~n3644 ;
  assign n33938 = n15677 ^ n8433 ^ 1'b0 ;
  assign n33939 = ~n20471 & n33938 ;
  assign n33940 = ~n9035 & n30153 ;
  assign n33941 = n13728 | n29822 ;
  assign n33942 = n26718 | n33941 ;
  assign n33943 = n14071 & n33942 ;
  assign n33944 = ~n24079 & n33943 ;
  assign n33946 = n1510 & n6404 ;
  assign n33947 = ~n31831 & n33946 ;
  assign n33945 = ~n7493 & n23212 ;
  assign n33948 = n33947 ^ n33945 ^ 1'b0 ;
  assign n33949 = n8920 & n13712 ;
  assign n33950 = n7275 | n33949 ;
  assign n33951 = n12512 & ~n27602 ;
  assign n33952 = ~n1630 & n33951 ;
  assign n33953 = n33952 ^ n32698 ^ n2338 ;
  assign n33954 = x163 & n14352 ;
  assign n33955 = ~n18362 & n33954 ;
  assign n33956 = n20031 ^ n5367 ^ 1'b0 ;
  assign n33957 = ~n17825 & n33956 ;
  assign n33958 = n33957 ^ n12306 ^ n4783 ;
  assign n33959 = ( n20021 & n33955 ) | ( n20021 & ~n33958 ) | ( n33955 & ~n33958 ) ;
  assign n33960 = n21900 & n25037 ;
  assign n33961 = n33960 ^ n1156 ^ 1'b0 ;
  assign n33962 = n4919 | n13614 ;
  assign n33963 = n33962 ^ n4824 ^ 1'b0 ;
  assign n33964 = n11491 & ~n33963 ;
  assign n33965 = n7996 & n16139 ;
  assign n33966 = n33965 ^ n6855 ^ 1'b0 ;
  assign n33967 = n7189 | n33966 ;
  assign n33968 = n33964 & n33967 ;
  assign n33969 = ~n7622 & n25444 ;
  assign n33970 = n33969 ^ n18394 ^ 1'b0 ;
  assign n33971 = n22703 ^ n11504 ^ 1'b0 ;
  assign n33972 = n29199 ^ n4661 ^ 1'b0 ;
  assign n33973 = n6319 & n33972 ;
  assign n33974 = n20080 ^ n11279 ^ 1'b0 ;
  assign n33975 = n11719 ^ n5296 ^ n4378 ;
  assign n33976 = n22849 ^ n943 ^ 1'b0 ;
  assign n33977 = ( ~n7619 & n19066 ) | ( ~n7619 & n33976 ) | ( n19066 & n33976 ) ;
  assign n33978 = n33977 ^ n26098 ^ n1640 ;
  assign n33979 = n20402 | n29890 ;
  assign n33980 = n18822 & ~n31932 ;
  assign n33981 = n1863 & n5710 ;
  assign n33983 = n782 | n2685 ;
  assign n33984 = n2230 | n33983 ;
  assign n33982 = ~n10287 & n14322 ;
  assign n33985 = n33984 ^ n33982 ^ n4959 ;
  assign n33986 = n1923 ^ n1542 ^ 1'b0 ;
  assign n33987 = ( ~n11389 & n19241 ) | ( ~n11389 & n33986 ) | ( n19241 & n33986 ) ;
  assign n33988 = ( x159 & n19727 ) | ( x159 & ~n33987 ) | ( n19727 & ~n33987 ) ;
  assign n33989 = n5672 & ~n29073 ;
  assign n33990 = n3455 & ~n6393 ;
  assign n33991 = ~n7349 & n33990 ;
  assign n33992 = ( n9823 & n13933 ) | ( n9823 & ~n33991 ) | ( n13933 & ~n33991 ) ;
  assign n33993 = n33992 ^ n19909 ^ 1'b0 ;
  assign n33994 = ~n15168 & n33993 ;
  assign n33995 = n1685 & n33994 ;
  assign n33996 = n21561 ^ n17572 ^ 1'b0 ;
  assign n33997 = n22710 ^ n1000 ^ 1'b0 ;
  assign n33998 = ~n33996 & n33997 ;
  assign n33999 = n1813 & n16682 ;
  assign n34000 = n9010 & n33999 ;
  assign n34001 = n34000 ^ n3185 ^ 1'b0 ;
  assign n34003 = n15370 ^ n1170 ^ 1'b0 ;
  assign n34002 = ( n1918 & n8018 ) | ( n1918 & ~n11472 ) | ( n8018 & ~n11472 ) ;
  assign n34004 = n34003 ^ n34002 ^ n7322 ;
  assign n34005 = n30707 ^ n21911 ^ n2092 ;
  assign n34006 = n31275 | n34005 ;
  assign n34007 = n20883 ^ n15030 ^ 1'b0 ;
  assign n34008 = n11562 & ~n34007 ;
  assign n34009 = n3547 & n34008 ;
  assign n34010 = ~n15635 & n34009 ;
  assign n34011 = n11070 & ~n13854 ;
  assign n34012 = n13835 & n34011 ;
  assign n34013 = n5443 | n26818 ;
  assign n34014 = ( n1995 & n15544 ) | ( n1995 & n21941 ) | ( n15544 & n21941 ) ;
  assign n34015 = n34014 ^ n11451 ^ n292 ;
  assign n34016 = n19698 & n21485 ;
  assign n34025 = n1664 & ~n16209 ;
  assign n34017 = n764 & n2311 ;
  assign n34018 = n34017 ^ n6754 ^ 1'b0 ;
  assign n34019 = x84 & ~n34018 ;
  assign n34020 = n34019 ^ n8211 ^ 1'b0 ;
  assign n34021 = n17626 ^ n8429 ^ 1'b0 ;
  assign n34022 = n9059 & n9844 ;
  assign n34023 = ~n34021 & n34022 ;
  assign n34024 = n34020 | n34023 ;
  assign n34026 = n34025 ^ n34024 ^ 1'b0 ;
  assign n34027 = ~n4469 & n33599 ;
  assign n34028 = n34027 ^ n7873 ^ 1'b0 ;
  assign n34029 = n24914 & ~n30028 ;
  assign n34030 = ( n6365 & ~n12720 ) | ( n6365 & n27215 ) | ( ~n12720 & n27215 ) ;
  assign n34031 = ~n2856 & n5203 ;
  assign n34032 = n34031 ^ n3368 ^ 1'b0 ;
  assign n34033 = ( ~n9379 & n24166 ) | ( ~n9379 & n34032 ) | ( n24166 & n34032 ) ;
  assign n34034 = ~n20596 & n30361 ;
  assign n34035 = ~n8448 & n29796 ;
  assign n34036 = n30523 & n34035 ;
  assign n34037 = n1322 & ~n7547 ;
  assign n34038 = n34037 ^ n7940 ^ n3749 ;
  assign n34039 = n34038 ^ n19796 ^ 1'b0 ;
  assign n34040 = n7342 & n29214 ;
  assign n34041 = n22020 & ~n22330 ;
  assign n34042 = ~n4334 & n20142 ;
  assign n34043 = n11108 | n21780 ;
  assign n34044 = ( n16777 & ~n27669 ) | ( n16777 & n34043 ) | ( ~n27669 & n34043 ) ;
  assign n34045 = ~n9832 & n24445 ;
  assign n34046 = n27149 ^ n12957 ^ n10562 ;
  assign n34047 = ~n11687 & n27622 ;
  assign n34048 = n26809 & n34047 ;
  assign n34049 = n15869 ^ n14692 ^ 1'b0 ;
  assign n34050 = n15338 & n34049 ;
  assign n34051 = n8935 ^ x38 ^ 1'b0 ;
  assign n34052 = ~n1257 & n34051 ;
  assign n34053 = ~n10449 & n34052 ;
  assign n34054 = n7004 | n7604 ;
  assign n34055 = n34054 ^ n15180 ^ 1'b0 ;
  assign n34056 = ~n34053 & n34055 ;
  assign n34057 = ~n5405 & n34056 ;
  assign n34058 = n34057 ^ n13633 ^ 1'b0 ;
  assign n34059 = n20645 & ~n34058 ;
  assign n34060 = n9222 & n24327 ;
  assign n34061 = n13124 & n34060 ;
  assign n34062 = n22201 ^ n20627 ^ 1'b0 ;
  assign n34063 = n15003 ^ n3078 ^ 1'b0 ;
  assign n34064 = n34062 & n34063 ;
  assign n34065 = n8523 | n32957 ;
  assign n34066 = n32895 ^ n2755 ^ 1'b0 ;
  assign n34067 = ( n14787 & ~n16022 ) | ( n14787 & n28222 ) | ( ~n16022 & n28222 ) ;
  assign n34068 = n356 & ~n11880 ;
  assign n34069 = n5472 & n34068 ;
  assign n34070 = n34067 & n34069 ;
  assign n34071 = n17949 & ~n34070 ;
  assign n34072 = n34071 ^ n29163 ^ 1'b0 ;
  assign n34073 = n8391 ^ n3091 ^ 1'b0 ;
  assign n34074 = n16967 ^ n1265 ^ 1'b0 ;
  assign n34075 = n34073 & n34074 ;
  assign n34076 = n9907 ^ n4484 ^ n3557 ;
  assign n34077 = n27449 ^ n6060 ^ 1'b0 ;
  assign n34078 = ~n34076 & n34077 ;
  assign n34079 = ( n27074 & ~n34075 ) | ( n27074 & n34078 ) | ( ~n34075 & n34078 ) ;
  assign n34080 = n11714 ^ n6201 ^ n907 ;
  assign n34081 = n9724 ^ n412 ^ 1'b0 ;
  assign n34082 = n34080 & ~n34081 ;
  assign n34083 = ( n4690 & n13249 ) | ( n4690 & n34082 ) | ( n13249 & n34082 ) ;
  assign n34084 = n34083 ^ n11348 ^ 1'b0 ;
  assign n34085 = ~n16718 & n34084 ;
  assign n34090 = n24551 ^ n22051 ^ 1'b0 ;
  assign n34091 = n11351 & ~n34090 ;
  assign n34087 = n5706 ^ n1328 ^ 1'b0 ;
  assign n34088 = ~n5165 & n34087 ;
  assign n34086 = ~n16933 & n19840 ;
  assign n34089 = n34088 ^ n34086 ^ 1'b0 ;
  assign n34092 = n34091 ^ n34089 ^ 1'b0 ;
  assign n34093 = n28130 ^ n11367 ^ 1'b0 ;
  assign n34094 = n8858 ^ n4801 ^ 1'b0 ;
  assign n34095 = n7586 & ~n14182 ;
  assign n34096 = n34095 ^ n17403 ^ 1'b0 ;
  assign n34097 = n34096 ^ n12521 ^ n11160 ;
  assign n34098 = ( ~n22306 & n34094 ) | ( ~n22306 & n34097 ) | ( n34094 & n34097 ) ;
  assign n34099 = ( n5360 & n11518 ) | ( n5360 & n12521 ) | ( n11518 & n12521 ) ;
  assign n34100 = ( n23107 & ~n33041 ) | ( n23107 & n34099 ) | ( ~n33041 & n34099 ) ;
  assign n34101 = n6176 ^ n1247 ^ 1'b0 ;
  assign n34102 = n33617 ^ n16168 ^ n3763 ;
  assign n34103 = n34101 & ~n34102 ;
  assign n34104 = n34103 ^ n13187 ^ 1'b0 ;
  assign n34105 = n24281 ^ n18082 ^ 1'b0 ;
  assign n34106 = n26271 | n34105 ;
  assign n34107 = ~n15268 & n16581 ;
  assign n34108 = ~n2007 & n2150 ;
  assign n34109 = n16518 & n34108 ;
  assign n34110 = n15116 & ~n34109 ;
  assign n34111 = ~n34107 & n34110 ;
  assign n34112 = n19353 | n29451 ;
  assign n34113 = n457 | n34112 ;
  assign n34114 = n4395 ^ n576 ^ 1'b0 ;
  assign n34115 = ~n3173 & n34114 ;
  assign n34116 = n34115 ^ n24002 ^ n6865 ;
  assign n34117 = n10794 ^ n9739 ^ n3481 ;
  assign n34118 = n1265 & n12570 ;
  assign n34119 = n34118 ^ n31182 ^ 1'b0 ;
  assign n34120 = n34119 ^ n13147 ^ 1'b0 ;
  assign n34121 = n4101 & ~n34120 ;
  assign n34122 = n22380 | n31777 ;
  assign n34123 = n34122 ^ n18588 ^ 1'b0 ;
  assign n34124 = n19399 ^ n1454 ^ 1'b0 ;
  assign n34125 = n34124 ^ n27975 ^ 1'b0 ;
  assign n34126 = ( x1 & ~n13092 ) | ( x1 & n21962 ) | ( ~n13092 & n21962 ) ;
  assign n34127 = n12240 & n18404 ;
  assign n34128 = ~n2016 & n34127 ;
  assign n34129 = n34128 ^ n12499 ^ 1'b0 ;
  assign n34130 = n34129 ^ n3985 ^ 1'b0 ;
  assign n34131 = n3630 & ~n34130 ;
  assign n34132 = n28740 & ~n34131 ;
  assign n34133 = n16439 & ~n34132 ;
  assign n34134 = n29476 ^ n26982 ^ n12102 ;
  assign n34135 = ( n20680 & ~n32876 ) | ( n20680 & n34134 ) | ( ~n32876 & n34134 ) ;
  assign n34136 = n27131 ^ n5011 ^ 1'b0 ;
  assign n34137 = ~n9388 & n34136 ;
  assign n34138 = n34137 ^ n9475 ^ 1'b0 ;
  assign n34139 = n26316 ^ n9897 ^ 1'b0 ;
  assign n34140 = n12796 | n14360 ;
  assign n34141 = ( ~n8850 & n9433 ) | ( ~n8850 & n30629 ) | ( n9433 & n30629 ) ;
  assign n34142 = n8875 ^ n4669 ^ 1'b0 ;
  assign n34143 = ~n34141 & n34142 ;
  assign n34144 = n21321 & n34143 ;
  assign n34145 = n10427 | n26515 ;
  assign n34146 = n14306 | n34145 ;
  assign n34147 = n34146 ^ n9433 ^ 1'b0 ;
  assign n34148 = n22819 | n34147 ;
  assign n34149 = n1486 ^ n854 ^ 1'b0 ;
  assign n34150 = n15988 & ~n22317 ;
  assign n34151 = n34149 & n34150 ;
  assign n34152 = n21985 ^ n17497 ^ 1'b0 ;
  assign n34153 = n5556 ^ n3133 ^ 1'b0 ;
  assign n34154 = n34153 ^ n475 ^ 1'b0 ;
  assign n34155 = n12153 & ~n34154 ;
  assign n34156 = n24540 ^ n1204 ^ 1'b0 ;
  assign n34157 = n14851 & ~n25959 ;
  assign n34158 = n34157 ^ n4787 ^ 1'b0 ;
  assign n34159 = ( n14690 & n32190 ) | ( n14690 & ~n34158 ) | ( n32190 & ~n34158 ) ;
  assign n34160 = n34159 ^ n3880 ^ 1'b0 ;
  assign n34161 = n34156 | n34160 ;
  assign n34162 = n34161 ^ n10781 ^ 1'b0 ;
  assign n34163 = n4219 & n23246 ;
  assign n34164 = n19250 ^ n14084 ^ n8151 ;
  assign n34165 = ( n28210 & n34163 ) | ( n28210 & ~n34164 ) | ( n34163 & ~n34164 ) ;
  assign n34166 = n5329 | n17983 ;
  assign n34167 = n1797 & n19909 ;
  assign n34168 = n12418 & n34167 ;
  assign n34169 = n4989 & n34168 ;
  assign n34170 = n9503 & n16440 ;
  assign n34171 = n34170 ^ n9890 ^ 1'b0 ;
  assign n34172 = n5625 & n14789 ;
  assign n34173 = n14743 ^ n10966 ^ 1'b0 ;
  assign n34174 = n34172 | n34173 ;
  assign n34175 = ( n28547 & n34171 ) | ( n28547 & n34174 ) | ( n34171 & n34174 ) ;
  assign n34176 = n1185 & ~n26759 ;
  assign n34177 = n11628 & n34176 ;
  assign n34178 = ( n34169 & n34175 ) | ( n34169 & ~n34177 ) | ( n34175 & ~n34177 ) ;
  assign n34179 = n9896 | n12644 ;
  assign n34180 = n30976 & ~n34179 ;
  assign n34181 = n2001 & ~n32552 ;
  assign n34182 = ( n5166 & n13182 ) | ( n5166 & ~n32233 ) | ( n13182 & ~n32233 ) ;
  assign n34183 = n34182 ^ n16357 ^ n2221 ;
  assign n34185 = ~n7678 & n14003 ;
  assign n34186 = n6501 & n34185 ;
  assign n34184 = ~n10339 & n17377 ;
  assign n34187 = n34186 ^ n34184 ^ 1'b0 ;
  assign n34188 = n34187 ^ n10025 ^ 1'b0 ;
  assign n34189 = n9148 & n30200 ;
  assign n34190 = ~n9156 & n34189 ;
  assign n34191 = n22784 ^ n17763 ^ n9509 ;
  assign n34192 = n34191 ^ n19976 ^ n10832 ;
  assign n34193 = ~n34190 & n34192 ;
  assign n34194 = ~n2028 & n9828 ;
  assign n34195 = n9602 ^ n7160 ^ 1'b0 ;
  assign n34196 = n4855 | n34195 ;
  assign n34197 = n34196 ^ n23884 ^ 1'b0 ;
  assign n34198 = n34197 ^ n10960 ^ n9304 ;
  assign n34199 = n34198 ^ n8078 ^ 1'b0 ;
  assign n34200 = ~n28051 & n34199 ;
  assign n34201 = n34200 ^ n3939 ^ 1'b0 ;
  assign n34202 = n34194 & ~n34201 ;
  assign n34203 = ~n10688 & n34202 ;
  assign n34204 = ~n3285 & n26885 ;
  assign n34205 = n13681 | n14880 ;
  assign n34206 = n34205 ^ n1383 ^ 1'b0 ;
  assign n34207 = n34206 ^ n10644 ^ 1'b0 ;
  assign n34208 = n34207 ^ n31995 ^ 1'b0 ;
  assign n34209 = n9282 ^ n5610 ^ 1'b0 ;
  assign n34210 = n23516 & ~n34209 ;
  assign n34213 = n5929 | n8179 ;
  assign n34214 = n34213 ^ n19907 ^ 1'b0 ;
  assign n34211 = n10884 ^ n5795 ^ n1655 ;
  assign n34212 = n21483 | n34211 ;
  assign n34215 = n34214 ^ n34212 ^ 1'b0 ;
  assign n34220 = ~n16826 & n30826 ;
  assign n34219 = n32848 ^ n20332 ^ n18516 ;
  assign n34216 = n9379 ^ n5485 ^ 1'b0 ;
  assign n34217 = n19581 & ~n34216 ;
  assign n34218 = n16757 & n34217 ;
  assign n34221 = n34220 ^ n34219 ^ n34218 ;
  assign n34222 = n11703 ^ n7279 ^ 1'b0 ;
  assign n34223 = n34222 ^ n471 ^ x38 ;
  assign n34224 = ( n7142 & n7998 ) | ( n7142 & n34223 ) | ( n7998 & n34223 ) ;
  assign n34225 = n8709 ^ n2107 ^ 1'b0 ;
  assign n34226 = n34225 ^ n9794 ^ 1'b0 ;
  assign n34227 = n6784 & ~n12671 ;
  assign n34228 = n19182 | n26583 ;
  assign n34229 = n7559 & ~n34228 ;
  assign n34230 = ~n24611 & n34229 ;
  assign n34231 = n33546 ^ n12281 ^ n660 ;
  assign n34232 = n18331 ^ n15761 ^ n7113 ;
  assign n34233 = n2688 & n18753 ;
  assign n34234 = n28516 | n29965 ;
  assign n34240 = n14724 ^ n2339 ^ 1'b0 ;
  assign n34241 = n9773 | n34240 ;
  assign n34235 = ~n4439 & n22260 ;
  assign n34236 = n9491 ^ x146 ^ 1'b0 ;
  assign n34237 = n4278 & ~n34236 ;
  assign n34238 = n34235 & ~n34237 ;
  assign n34239 = n33354 & ~n34238 ;
  assign n34242 = n34241 ^ n34239 ^ 1'b0 ;
  assign n34243 = ~n14108 & n26495 ;
  assign n34244 = ( n2955 & ~n17011 ) | ( n2955 & n17754 ) | ( ~n17011 & n17754 ) ;
  assign n34245 = n33609 ^ n9333 ^ n5776 ;
  assign n34246 = ( n4034 & n6944 ) | ( n4034 & ~n34245 ) | ( n6944 & ~n34245 ) ;
  assign n34247 = ~n7900 & n18928 ;
  assign n34248 = n14510 ^ n5637 ^ 1'b0 ;
  assign n34249 = n34247 & n34248 ;
  assign n34250 = ~n3019 & n15761 ;
  assign n34253 = ~n804 & n11232 ;
  assign n34254 = n34253 ^ n9010 ^ 1'b0 ;
  assign n34255 = n34254 ^ n22950 ^ n8361 ;
  assign n34251 = n33189 ^ n30307 ^ 1'b0 ;
  assign n34252 = ~n18394 & n34251 ;
  assign n34256 = n34255 ^ n34252 ^ 1'b0 ;
  assign n34257 = n29277 ^ n18466 ^ 1'b0 ;
  assign n34258 = n34257 ^ n17836 ^ n259 ;
  assign n34259 = n12230 ^ n11361 ^ 1'b0 ;
  assign n34260 = n22192 | n34259 ;
  assign n34261 = n34260 ^ n27318 ^ 1'b0 ;
  assign n34262 = n12656 ^ n7759 ^ n608 ;
  assign n34263 = n6998 & n7381 ;
  assign n34264 = n11884 & n34263 ;
  assign n34265 = n29314 | n34264 ;
  assign n34266 = n34262 & ~n34265 ;
  assign n34267 = n22317 | n34266 ;
  assign n34273 = ( n1472 & ~n7104 ) | ( n1472 & n8287 ) | ( ~n7104 & n8287 ) ;
  assign n34268 = n853 & n9260 ;
  assign n34269 = n17587 & n34268 ;
  assign n34270 = n34269 ^ n25930 ^ 1'b0 ;
  assign n34271 = n31883 | n34270 ;
  assign n34272 = n15881 & n34271 ;
  assign n34274 = n34273 ^ n34272 ^ 1'b0 ;
  assign n34275 = n8181 & ~n34211 ;
  assign n34276 = n11443 & n31219 ;
  assign n34277 = n32038 ^ n14998 ^ 1'b0 ;
  assign n34278 = n13530 & n34277 ;
  assign n34279 = ~n4394 & n33186 ;
  assign n34280 = n34279 ^ n19765 ^ 1'b0 ;
  assign n34281 = n4310 & ~n8228 ;
  assign n34282 = n19736 & n34281 ;
  assign n34283 = n808 & ~n34282 ;
  assign n34284 = n34283 ^ n21664 ^ 1'b0 ;
  assign n34285 = n34284 ^ n23795 ^ n11000 ;
  assign n34286 = n17520 | n19911 ;
  assign n34287 = n5909 | n34286 ;
  assign n34288 = n34287 ^ n14785 ^ 1'b0 ;
  assign n34289 = n25912 ^ n3033 ^ 1'b0 ;
  assign n34290 = n2639 | n18732 ;
  assign n34291 = n34290 ^ n2476 ^ x182 ;
  assign n34292 = n14741 ^ n1937 ^ 1'b0 ;
  assign n34293 = ~n19031 & n34292 ;
  assign n34294 = n34293 ^ n23388 ^ n6543 ;
  assign n34295 = ~n14439 & n19649 ;
  assign n34296 = ~n4438 & n34295 ;
  assign n34297 = n34296 ^ n33417 ^ n26412 ;
  assign n34298 = x185 & n18448 ;
  assign n34299 = n12893 & n34298 ;
  assign n34300 = n7824 & n34299 ;
  assign n34301 = n10046 ^ n3212 ^ 1'b0 ;
  assign n34302 = ~n34300 & n34301 ;
  assign n34303 = n34302 ^ n12480 ^ 1'b0 ;
  assign n34304 = n8746 | n34303 ;
  assign n34308 = n5975 & n17661 ;
  assign n34309 = n34308 ^ n5475 ^ 1'b0 ;
  assign n34310 = n6870 & n34309 ;
  assign n34311 = ~n20403 & n34310 ;
  assign n34305 = n18465 ^ n11566 ^ 1'b0 ;
  assign n34306 = n3049 ^ n2294 ^ 1'b0 ;
  assign n34307 = n34305 & ~n34306 ;
  assign n34312 = n34311 ^ n34307 ^ n17519 ;
  assign n34313 = n22716 | n34312 ;
  assign n34314 = n34313 ^ n9242 ^ 1'b0 ;
  assign n34315 = n12353 | n17508 ;
  assign n34316 = n34315 ^ n3878 ^ 1'b0 ;
  assign n34317 = ( x97 & n7630 ) | ( x97 & ~n9717 ) | ( n7630 & ~n9717 ) ;
  assign n34318 = n24707 ^ n5334 ^ n2993 ;
  assign n34319 = ( n5070 & n34317 ) | ( n5070 & n34318 ) | ( n34317 & n34318 ) ;
  assign n34322 = n256 | n343 ;
  assign n34323 = n343 & ~n34322 ;
  assign n34320 = n5702 & ~n6899 ;
  assign n34321 = n6899 & n34320 ;
  assign n34324 = n34323 ^ n34321 ^ n7515 ;
  assign n34325 = n6710 & n12779 ;
  assign n34326 = n34325 ^ n21311 ^ n14981 ;
  assign n34327 = n31061 & n34326 ;
  assign n34328 = n12874 & n27906 ;
  assign n34329 = n34328 ^ n27716 ^ 1'b0 ;
  assign n34330 = ~x87 & n21277 ;
  assign n34331 = n33929 ^ n27678 ^ 1'b0 ;
  assign n34332 = n31787 & n34331 ;
  assign n34333 = n34330 & n34332 ;
  assign n34334 = n4501 | n17646 ;
  assign n34335 = n16478 & ~n34334 ;
  assign n34336 = n34335 ^ n19866 ^ 1'b0 ;
  assign n34337 = n26545 ^ n10803 ^ n8930 ;
  assign n34338 = ( ~n9277 & n12036 ) | ( ~n9277 & n34337 ) | ( n12036 & n34337 ) ;
  assign n34339 = n34338 ^ n20713 ^ 1'b0 ;
  assign n34340 = n34336 & n34339 ;
  assign n34341 = n21768 | n27010 ;
  assign n34342 = n16897 | n34341 ;
  assign n34343 = n34342 ^ n4454 ^ n3299 ;
  assign n34344 = n1928 & ~n12986 ;
  assign n34345 = n34344 ^ n2978 ^ 1'b0 ;
  assign n34346 = ( ~n25892 & n33362 ) | ( ~n25892 & n34345 ) | ( n33362 & n34345 ) ;
  assign n34347 = n34346 ^ n20925 ^ n8017 ;
  assign n34348 = n375 & n4441 ;
  assign n34349 = n20501 & ~n23306 ;
  assign n34350 = n11005 & n34349 ;
  assign n34351 = n3262 & ~n18554 ;
  assign n34352 = n33858 ^ n28764 ^ 1'b0 ;
  assign n34353 = n14018 & n34352 ;
  assign n34356 = n10105 ^ n3145 ^ n2094 ;
  assign n34354 = ( ~n6362 & n6681 ) | ( ~n6362 & n6940 ) | ( n6681 & n6940 ) ;
  assign n34355 = ( n21898 & n22617 ) | ( n21898 & n34354 ) | ( n22617 & n34354 ) ;
  assign n34357 = n34356 ^ n34355 ^ 1'b0 ;
  assign n34358 = n34357 ^ n19303 ^ 1'b0 ;
  assign n34359 = ( ~x247 & n4888 ) | ( ~x247 & n15963 ) | ( n4888 & n15963 ) ;
  assign n34360 = n4763 ^ n994 ^ 1'b0 ;
  assign n34361 = n22451 & ~n34360 ;
  assign n34362 = ~n17098 & n34361 ;
  assign n34363 = ( n3810 & ~n13968 ) | ( n3810 & n34362 ) | ( ~n13968 & n34362 ) ;
  assign n34364 = n1285 | n7994 ;
  assign n34365 = ~n19584 & n34364 ;
  assign n34366 = n34365 ^ n9897 ^ 1'b0 ;
  assign n34367 = ( n12597 & n13545 ) | ( n12597 & ~n34366 ) | ( n13545 & ~n34366 ) ;
  assign n34368 = n17796 & ~n18048 ;
  assign n34369 = ( ~n2769 & n3007 ) | ( ~n2769 & n34368 ) | ( n3007 & n34368 ) ;
  assign n34370 = n12726 & ~n24270 ;
  assign n34371 = n16681 & ~n28191 ;
  assign n34372 = ~n8343 & n34371 ;
  assign n34374 = n13788 ^ n2349 ^ 1'b0 ;
  assign n34373 = n12962 ^ n1899 ^ 1'b0 ;
  assign n34375 = n34374 ^ n34373 ^ n5105 ;
  assign n34376 = n34375 ^ n21132 ^ 1'b0 ;
  assign n34377 = ( ~n2543 & n14016 ) | ( ~n2543 & n33822 ) | ( n14016 & n33822 ) ;
  assign n34378 = n8835 ^ n3191 ^ 1'b0 ;
  assign n34379 = n18406 & n34378 ;
  assign n34380 = n17647 ^ n9121 ^ 1'b0 ;
  assign n34381 = n8507 ^ n5195 ^ 1'b0 ;
  assign n34382 = ( x92 & ~n7520 ) | ( x92 & n34381 ) | ( ~n7520 & n34381 ) ;
  assign n34383 = ~n8841 & n9333 ;
  assign n34384 = ~n34382 & n34383 ;
  assign n34385 = n26724 ^ n9146 ^ 1'b0 ;
  assign n34386 = ~n26097 & n34385 ;
  assign n34387 = n9986 | n19524 ;
  assign n34388 = n1725 | n34387 ;
  assign n34389 = n21243 & n34388 ;
  assign n34390 = n10767 & ~n26865 ;
  assign n34391 = n23213 & n34390 ;
  assign n34392 = n20927 & n34391 ;
  assign n34393 = x65 & ~n19575 ;
  assign n34394 = ~n8372 & n34393 ;
  assign n34395 = n34394 ^ n34273 ^ n2349 ;
  assign n34397 = ( ~n2835 & n25722 ) | ( ~n2835 & n26712 ) | ( n25722 & n26712 ) ;
  assign n34396 = n14859 | n24003 ;
  assign n34398 = n34397 ^ n34396 ^ n9772 ;
  assign n34399 = n34398 ^ n15151 ^ n14242 ;
  assign n34400 = n30101 ^ n704 ^ 1'b0 ;
  assign n34401 = n29277 ^ n25396 ^ n17023 ;
  assign n34402 = n27774 ^ n23292 ^ 1'b0 ;
  assign n34403 = n1362 & ~n34402 ;
  assign n34405 = ( x194 & n8778 ) | ( x194 & n21573 ) | ( n8778 & n21573 ) ;
  assign n34406 = n4104 | n16002 ;
  assign n34407 = n34405 | n34406 ;
  assign n34408 = n34407 ^ n3896 ^ 1'b0 ;
  assign n34404 = n2389 & ~n6001 ;
  assign n34409 = n34408 ^ n34404 ^ 1'b0 ;
  assign n34410 = n10879 | n27725 ;
  assign n34411 = n18160 | n30046 ;
  assign n34412 = n34410 | n34411 ;
  assign n34413 = n7865 | n26770 ;
  assign n34414 = n9628 ^ n8460 ^ 1'b0 ;
  assign n34415 = n3197 & n34414 ;
  assign n34416 = n31928 ^ n20436 ^ n1593 ;
  assign n34417 = n34416 ^ n2164 ^ 1'b0 ;
  assign n34418 = n14923 ^ n10629 ^ 1'b0 ;
  assign n34419 = n12437 ^ n10537 ^ n2850 ;
  assign n34420 = n29816 ^ n6318 ^ 1'b0 ;
  assign n34421 = n9569 | n34420 ;
  assign n34422 = n16276 ^ n3010 ^ 1'b0 ;
  assign n34423 = n4546 | n9969 ;
  assign n34424 = n10480 | n34423 ;
  assign n34425 = n34424 ^ n8572 ^ 1'b0 ;
  assign n34426 = n29150 ^ n18403 ^ 1'b0 ;
  assign n34427 = n34425 & ~n34426 ;
  assign n34428 = n16783 & ~n24537 ;
  assign n34429 = n12167 & ~n14642 ;
  assign n34430 = n34428 & n34429 ;
  assign n34431 = n8372 | n21003 ;
  assign n34432 = n25694 ^ n20026 ^ n3835 ;
  assign n34433 = n11726 ^ n3726 ^ 1'b0 ;
  assign n34434 = ( n15707 & n34159 ) | ( n15707 & ~n34433 ) | ( n34159 & ~n34433 ) ;
  assign n34435 = n15130 ^ n14920 ^ 1'b0 ;
  assign n34436 = n11211 & ~n34435 ;
  assign n34437 = n29988 ^ n4052 ^ 1'b0 ;
  assign n34438 = ~n2302 & n34437 ;
  assign n34439 = n29782 | n30165 ;
  assign n34440 = n34438 | n34439 ;
  assign n34441 = ~x145 & n9610 ;
  assign n34442 = ~x188 & x242 ;
  assign n34443 = n34441 & ~n34442 ;
  assign n34444 = ( n1399 & ~n19582 ) | ( n1399 & n34443 ) | ( ~n19582 & n34443 ) ;
  assign n34445 = n7496 ^ n2758 ^ 1'b0 ;
  assign n34446 = n17188 ^ n15714 ^ n14966 ;
  assign n34447 = n31992 ^ n24345 ^ n1090 ;
  assign n34448 = n7043 & n34447 ;
  assign n34449 = n25028 ^ n9088 ^ 1'b0 ;
  assign n34450 = n20014 & ~n34449 ;
  assign n34451 = n17510 ^ n7617 ^ 1'b0 ;
  assign n34452 = n15263 ^ n7757 ^ 1'b0 ;
  assign n34453 = ( n24740 & ~n26944 ) | ( n24740 & n34452 ) | ( ~n26944 & n34452 ) ;
  assign n34454 = n12525 ^ n10830 ^ 1'b0 ;
  assign n34455 = n9721 | n34454 ;
  assign n34456 = n34455 ^ n16739 ^ n347 ;
  assign n34457 = n11751 ^ n9020 ^ 1'b0 ;
  assign n34459 = n20895 ^ n7113 ^ n2137 ;
  assign n34458 = ~n3904 & n15116 ;
  assign n34460 = n34459 ^ n34458 ^ 1'b0 ;
  assign n34461 = n3339 & ~n15784 ;
  assign n34462 = n26818 & n34461 ;
  assign n34463 = n34462 ^ n10500 ^ 1'b0 ;
  assign n34464 = n11575 ^ n11344 ^ 1'b0 ;
  assign n34465 = n21090 & ~n26201 ;
  assign n34466 = n33889 ^ n8111 ^ 1'b0 ;
  assign n34467 = n34465 & ~n34466 ;
  assign n34468 = n19163 ^ n17140 ^ 1'b0 ;
  assign n34469 = n7263 & ~n34468 ;
  assign n34470 = n34469 ^ n7228 ^ 1'b0 ;
  assign n34471 = n34470 ^ n1638 ^ 1'b0 ;
  assign n34472 = n1751 | n13254 ;
  assign n34473 = n5782 ^ n2236 ^ 1'b0 ;
  assign n34474 = ~n5704 & n34473 ;
  assign n34475 = n34474 ^ n20009 ^ n1579 ;
  assign n34476 = n1424 & n1776 ;
  assign n34477 = n34476 ^ n6889 ^ 1'b0 ;
  assign n34478 = n17928 & n34477 ;
  assign n34479 = ( n26588 & n34475 ) | ( n26588 & ~n34478 ) | ( n34475 & ~n34478 ) ;
  assign n34480 = n24096 ^ n15149 ^ 1'b0 ;
  assign n34481 = n34479 & n34480 ;
  assign n34482 = n34109 | n34481 ;
  assign n34483 = n25824 ^ n13741 ^ 1'b0 ;
  assign n34484 = ( n7066 & n16524 ) | ( n7066 & n21834 ) | ( n16524 & n21834 ) ;
  assign n34485 = n34484 ^ n17086 ^ 1'b0 ;
  assign n34486 = ~n8717 & n27702 ;
  assign n34487 = n12129 & n14321 ;
  assign n34488 = n34487 ^ n7512 ^ 1'b0 ;
  assign n34489 = n34488 ^ n12733 ^ n5844 ;
  assign n34490 = n31062 | n34489 ;
  assign n34491 = n1362 ^ n577 ^ x131 ;
  assign n34492 = n34491 ^ n18757 ^ n3746 ;
  assign n34494 = n10391 & ~n29998 ;
  assign n34495 = n34494 ^ n1510 ^ 1'b0 ;
  assign n34493 = n7617 & ~n9217 ;
  assign n34496 = n34495 ^ n34493 ^ 1'b0 ;
  assign n34497 = ~n25851 & n34496 ;
  assign n34498 = n20466 ^ n13595 ^ 1'b0 ;
  assign n34499 = ~n2531 & n3511 ;
  assign n34500 = n34499 ^ n27861 ^ n23363 ;
  assign n34501 = ~n21671 & n34500 ;
  assign n34502 = ( n7427 & ~n24543 ) | ( n7427 & n26662 ) | ( ~n24543 & n26662 ) ;
  assign n34503 = ~n1503 & n34502 ;
  assign n34504 = n10163 & ~n34503 ;
  assign n34505 = ( n2481 & n21157 ) | ( n2481 & ~n30923 ) | ( n21157 & ~n30923 ) ;
  assign n34506 = n32964 ^ n7101 ^ 1'b0 ;
  assign n34507 = ~n5155 & n32288 ;
  assign n34508 = n34507 ^ n26321 ^ 1'b0 ;
  assign n34509 = n21201 | n34508 ;
  assign n34510 = ~n24166 & n30207 ;
  assign n34511 = n4761 & n34510 ;
  assign n34512 = n4041 ^ x198 ^ x179 ;
  assign n34513 = n7122 | n34512 ;
  assign n34514 = n15524 ^ n6032 ^ 1'b0 ;
  assign n34515 = x149 & ~n15760 ;
  assign n34516 = n5491 & n34515 ;
  assign n34517 = n27523 ^ n16315 ^ 1'b0 ;
  assign n34518 = n16840 | n34517 ;
  assign n34519 = ( x1 & n1129 ) | ( x1 & ~n5072 ) | ( n1129 & ~n5072 ) ;
  assign n34520 = n34519 ^ n5258 ^ 1'b0 ;
  assign n34521 = ~n12396 & n34520 ;
  assign n34522 = ~n6896 & n34521 ;
  assign n34523 = n19402 ^ n2688 ^ 1'b0 ;
  assign n34524 = n12805 & ~n34523 ;
  assign n34525 = ( n2931 & n5830 ) | ( n2931 & ~n14559 ) | ( n5830 & ~n14559 ) ;
  assign n34526 = ( ~n16493 & n34524 ) | ( ~n16493 & n34525 ) | ( n34524 & n34525 ) ;
  assign n34527 = n13607 | n22349 ;
  assign n34528 = n24698 | n34527 ;
  assign n34529 = n30836 ^ n6988 ^ n6629 ;
  assign n34530 = n34528 & n34529 ;
  assign n34531 = n34530 ^ n22442 ^ 1'b0 ;
  assign n34532 = n21487 ^ n6983 ^ 1'b0 ;
  assign n34533 = n18561 ^ n5190 ^ 1'b0 ;
  assign n34534 = n10621 & n34533 ;
  assign n34535 = n26930 ^ x35 ^ 1'b0 ;
  assign n34536 = n28704 | n33002 ;
  assign n34537 = n34536 ^ n24565 ^ 1'b0 ;
  assign n34538 = n20905 ^ n20773 ^ n16640 ;
  assign n34539 = n17562 | n34538 ;
  assign n34540 = n34539 ^ n12032 ^ 1'b0 ;
  assign n34541 = n34540 ^ n29042 ^ n24789 ;
  assign n34542 = n16190 ^ n6558 ^ 1'b0 ;
  assign n34543 = n4448 | n34542 ;
  assign n34544 = n8928 | n14011 ;
  assign n34545 = n34544 ^ n7172 ^ 1'b0 ;
  assign n34546 = n34545 ^ n14170 ^ 1'b0 ;
  assign n34547 = n30459 | n34546 ;
  assign n34548 = n34547 ^ n14912 ^ 1'b0 ;
  assign n34549 = ( n14770 & ~n34543 ) | ( n14770 & n34548 ) | ( ~n34543 & n34548 ) ;
  assign n34550 = n18164 & ~n34549 ;
  assign n34551 = ( n13974 & n26881 ) | ( n13974 & n34550 ) | ( n26881 & n34550 ) ;
  assign n34552 = ( n933 & n4592 ) | ( n933 & n7142 ) | ( n4592 & n7142 ) ;
  assign n34553 = n20139 & ~n34552 ;
  assign n34554 = n34553 ^ n27530 ^ n20276 ;
  assign n34555 = n31482 ^ n5840 ^ n5265 ;
  assign n34556 = n2925 & ~n34555 ;
  assign n34557 = n8688 | n28789 ;
  assign n34558 = n4591 & n9955 ;
  assign n34559 = n12677 ^ n9071 ^ 1'b0 ;
  assign n34560 = n34559 ^ n6892 ^ 1'b0 ;
  assign n34561 = ~n34558 & n34560 ;
  assign n34562 = n21793 ^ n1105 ^ 1'b0 ;
  assign n34563 = n34562 ^ n28305 ^ 1'b0 ;
  assign n34564 = n14741 | n34563 ;
  assign n34565 = n455 | n2152 ;
  assign n34566 = n2422 & ~n34565 ;
  assign n34567 = n34566 ^ n8626 ^ n1429 ;
  assign n34568 = n2873 & ~n3401 ;
  assign n34569 = n21994 & n22703 ;
  assign n34570 = ~n10085 & n15717 ;
  assign n34571 = n3662 & ~n34570 ;
  assign n34572 = n34569 & n34571 ;
  assign n34573 = ( n4020 & n6109 ) | ( n4020 & ~n28668 ) | ( n6109 & ~n28668 ) ;
  assign n34574 = x247 & n6796 ;
  assign n34575 = ~n2529 & n34574 ;
  assign n34576 = n34575 ^ n28608 ^ n2720 ;
  assign n34577 = ~n9460 & n16911 ;
  assign n34578 = n34577 ^ n3073 ^ 1'b0 ;
  assign n34579 = n34578 ^ n29277 ^ 1'b0 ;
  assign n34580 = n11823 | n15278 ;
  assign n34581 = n32804 ^ n1197 ^ 1'b0 ;
  assign n34582 = n9503 & n30037 ;
  assign n34583 = n12575 & n13617 ;
  assign n34584 = n10218 ^ n7994 ^ 1'b0 ;
  assign n34585 = n26365 ^ n8043 ^ n7293 ;
  assign n34586 = n6930 & n25048 ;
  assign n34587 = n8459 & n34586 ;
  assign n34588 = ~n18668 & n18972 ;
  assign n34589 = n34588 ^ n10102 ^ 1'b0 ;
  assign n34590 = n34589 ^ n19194 ^ 1'b0 ;
  assign n34591 = ~n31053 & n34590 ;
  assign n34592 = n33978 ^ n16750 ^ 1'b0 ;
  assign n34593 = n17185 & ~n34592 ;
  assign n34594 = n3631 & ~n6779 ;
  assign n34595 = n9050 & n34594 ;
  assign n34596 = n764 & ~n5451 ;
  assign n34597 = ~n4723 & n9666 ;
  assign n34598 = n5434 & n34597 ;
  assign n34599 = n30832 & n34598 ;
  assign n34600 = ( n29578 & n34596 ) | ( n29578 & ~n34599 ) | ( n34596 & ~n34599 ) ;
  assign n34605 = n14065 ^ n11951 ^ 1'b0 ;
  assign n34606 = n34605 ^ n7044 ^ 1'b0 ;
  assign n34607 = n5975 & n34606 ;
  assign n34601 = n4117 | n19900 ;
  assign n34602 = n34601 ^ n21341 ^ 1'b0 ;
  assign n34603 = n13114 & ~n31769 ;
  assign n34604 = n34602 & n34603 ;
  assign n34608 = n34607 ^ n34604 ^ 1'b0 ;
  assign n34609 = ~n13262 & n28250 ;
  assign n34610 = n17902 & ~n21462 ;
  assign n34612 = ( n4097 & n7575 ) | ( n4097 & ~n13170 ) | ( n7575 & ~n13170 ) ;
  assign n34611 = ~n16555 & n19641 ;
  assign n34613 = n34612 ^ n34611 ^ n14237 ;
  assign n34614 = n34613 ^ n31456 ^ 1'b0 ;
  assign n34618 = n14869 ^ n5054 ^ 1'b0 ;
  assign n34615 = ~n17027 & n29106 ;
  assign n34616 = n27600 & n34615 ;
  assign n34617 = ( ~n18728 & n19759 ) | ( ~n18728 & n34616 ) | ( n19759 & n34616 ) ;
  assign n34619 = n34618 ^ n34617 ^ n1369 ;
  assign n34620 = n34619 ^ n15533 ^ 1'b0 ;
  assign n34621 = x109 & n11141 ;
  assign n34622 = ~n11500 & n34621 ;
  assign n34623 = n23294 ^ n330 ^ 1'b0 ;
  assign n34624 = n34623 ^ n34093 ^ 1'b0 ;
  assign n34625 = ~n1399 & n34624 ;
  assign n34626 = n16702 & n26780 ;
  assign n34627 = n17514 | n33430 ;
  assign n34628 = n1538 & n7500 ;
  assign n34629 = n34628 ^ n304 ^ 1'b0 ;
  assign n34630 = ( n10269 & ~n26910 ) | ( n10269 & n34629 ) | ( ~n26910 & n34629 ) ;
  assign n34631 = n22469 | n25743 ;
  assign n34632 = ( n3952 & n7647 ) | ( n3952 & n8843 ) | ( n7647 & n8843 ) ;
  assign n34633 = ( n21591 & n25725 ) | ( n21591 & ~n34632 ) | ( n25725 & ~n34632 ) ;
  assign n34634 = n21260 ^ n14372 ^ 1'b0 ;
  assign n34635 = n4979 & ~n6835 ;
  assign n34636 = n29399 & n34635 ;
  assign n34637 = n21213 ^ n15115 ^ n8784 ;
  assign n34638 = n26413 & n34637 ;
  assign n34639 = n18046 ^ n2179 ^ 1'b0 ;
  assign n34640 = n34639 ^ n32572 ^ n21106 ;
  assign n34641 = n393 ^ x56 ^ 1'b0 ;
  assign n34642 = n13279 ^ n4564 ^ 1'b0 ;
  assign n34643 = n34642 ^ n16529 ^ 1'b0 ;
  assign n34644 = n34641 & ~n34643 ;
  assign n34645 = n23677 & n34644 ;
  assign n34646 = ~n5373 & n34645 ;
  assign n34647 = ( n3305 & n34640 ) | ( n3305 & ~n34646 ) | ( n34640 & ~n34646 ) ;
  assign n34648 = ~n15279 & n20499 ;
  assign n34649 = n34648 ^ n11380 ^ 1'b0 ;
  assign n34650 = ~n14958 & n34649 ;
  assign n34651 = ( n1041 & ~n30339 ) | ( n1041 & n34650 ) | ( ~n30339 & n34650 ) ;
  assign n34652 = ~n17209 & n33124 ;
  assign n34653 = n34652 ^ n3517 ^ 1'b0 ;
  assign n34654 = ( ~n3049 & n5153 ) | ( ~n3049 & n18715 ) | ( n5153 & n18715 ) ;
  assign n34655 = n1237 & ~n14580 ;
  assign n34656 = n34654 & n34655 ;
  assign n34661 = n4024 & ~n28905 ;
  assign n34662 = ~n5456 & n34661 ;
  assign n34657 = n13968 & ~n17562 ;
  assign n34658 = n476 & ~n1236 ;
  assign n34659 = n34658 ^ n15556 ^ 1'b0 ;
  assign n34660 = n34657 & n34659 ;
  assign n34663 = n34662 ^ n34660 ^ 1'b0 ;
  assign n34664 = n31113 & ~n34663 ;
  assign n34665 = n5052 & n15639 ;
  assign n34666 = ( n1462 & n5291 ) | ( n1462 & ~n34665 ) | ( n5291 & ~n34665 ) ;
  assign n34667 = ( n24575 & ~n31664 ) | ( n24575 & n34666 ) | ( ~n31664 & n34666 ) ;
  assign n34668 = ( n17993 & n33330 ) | ( n17993 & n34667 ) | ( n33330 & n34667 ) ;
  assign n34669 = n29429 ^ n13197 ^ n1276 ;
  assign n34670 = ( n966 & ~n17702 ) | ( n966 & n34375 ) | ( ~n17702 & n34375 ) ;
  assign n34671 = n17230 ^ n2939 ^ n1113 ;
  assign n34672 = ~n8168 & n34671 ;
  assign n34673 = n34672 ^ n17134 ^ n9824 ;
  assign n34674 = n16829 | n19679 ;
  assign n34675 = n8145 & ~n15505 ;
  assign n34676 = n7638 & n34675 ;
  assign n34677 = n34631 ^ n25657 ^ n13505 ;
  assign n34678 = x71 & n2772 ;
  assign n34679 = ( n642 & ~n10909 ) | ( n642 & n34678 ) | ( ~n10909 & n34678 ) ;
  assign n34680 = n10174 | n34679 ;
  assign n34681 = n34680 ^ n11371 ^ 1'b0 ;
  assign n34682 = n18243 | n34681 ;
  assign n34683 = n34682 ^ n27764 ^ n16027 ;
  assign n34684 = n5163 & n22310 ;
  assign n34685 = n18861 ^ n16362 ^ n6016 ;
  assign n34686 = n34685 ^ n20453 ^ n1722 ;
  assign n34687 = ( n9972 & n15186 ) | ( n9972 & ~n16259 ) | ( n15186 & ~n16259 ) ;
  assign n34688 = n16857 | n34687 ;
  assign n34689 = n34688 ^ n5813 ^ 1'b0 ;
  assign n34690 = n23981 ^ n3059 ^ n1040 ;
  assign n34691 = ( x172 & n10351 ) | ( x172 & ~n34690 ) | ( n10351 & ~n34690 ) ;
  assign n34692 = ( ~n1253 & n6563 ) | ( ~n1253 & n9765 ) | ( n6563 & n9765 ) ;
  assign n34693 = ~n29905 & n34692 ;
  assign n34694 = n34693 ^ n8025 ^ 1'b0 ;
  assign n34695 = n10328 ^ n1302 ^ 1'b0 ;
  assign n34696 = ~n3051 & n34695 ;
  assign n34697 = n32266 ^ n904 ^ 1'b0 ;
  assign n34698 = ~n18307 & n19980 ;
  assign n34699 = ( ~x47 & n5030 ) | ( ~x47 & n27527 ) | ( n5030 & n27527 ) ;
  assign n34700 = n5234 & n5969 ;
  assign n34701 = n34700 ^ n22679 ^ 1'b0 ;
  assign n34702 = n4443 & n34701 ;
  assign n34703 = n9230 | n26602 ;
  assign n34704 = ~n2433 & n8260 ;
  assign n34705 = n21057 & n34704 ;
  assign n34706 = ~n7503 & n19689 ;
  assign n34707 = ~n34705 & n34706 ;
  assign n34708 = n25987 ^ x125 ^ 1'b0 ;
  assign n34709 = n13553 & n34708 ;
  assign n34710 = ~n11992 & n34709 ;
  assign n34711 = n17517 ^ n14275 ^ n14125 ;
  assign n34712 = n34711 ^ n28504 ^ 1'b0 ;
  assign n34713 = n10863 ^ n6205 ^ 1'b0 ;
  assign n34714 = n28686 ^ n28087 ^ 1'b0 ;
  assign n34715 = n9138 & n34714 ;
  assign n34716 = n33599 ^ n18394 ^ 1'b0 ;
  assign n34717 = ( n8799 & n14244 ) | ( n8799 & n34716 ) | ( n14244 & n34716 ) ;
  assign n34718 = ( n14481 & n17468 ) | ( n14481 & ~n28718 ) | ( n17468 & ~n28718 ) ;
  assign n34719 = n16165 & n22310 ;
  assign n34720 = n4626 & n34719 ;
  assign n34721 = n34720 ^ n13182 ^ 1'b0 ;
  assign n34722 = n10922 ^ n6638 ^ 1'b0 ;
  assign n34723 = n7051 | n34722 ;
  assign n34724 = n22697 & n34723 ;
  assign n34725 = n29305 ^ n28813 ^ 1'b0 ;
  assign n34726 = n3312 | n28339 ;
  assign n34727 = n10188 | n26660 ;
  assign n34728 = n19871 ^ n17013 ^ 1'b0 ;
  assign n34729 = n5827 | n6357 ;
  assign n34730 = n34729 ^ n507 ^ 1'b0 ;
  assign n34731 = n22497 & ~n34730 ;
  assign n34732 = n34731 ^ n33884 ^ n14692 ;
  assign n34733 = n34732 ^ n26200 ^ n19421 ;
  assign n34734 = n13226 | n21382 ;
  assign n34735 = ~n15630 & n34734 ;
  assign n34736 = n3953 & n34735 ;
  assign n34737 = n34736 ^ n10860 ^ 1'b0 ;
  assign n34738 = n6701 ^ n3045 ^ 1'b0 ;
  assign n34739 = ~n4274 & n34738 ;
  assign n34740 = n9467 | n34739 ;
  assign n34741 = n12642 & n15069 ;
  assign n34743 = n10963 ^ n3408 ^ 1'b0 ;
  assign n34742 = ( n6430 & n8509 ) | ( n6430 & ~n16961 ) | ( n8509 & ~n16961 ) ;
  assign n34744 = n34743 ^ n34742 ^ 1'b0 ;
  assign n34745 = ~n26086 & n34744 ;
  assign n34746 = n1452 & n3157 ;
  assign n34747 = n34746 ^ n15086 ^ 1'b0 ;
  assign n34748 = n34747 ^ n12034 ^ n2818 ;
  assign n34749 = n34748 ^ n15303 ^ 1'b0 ;
  assign n34750 = ~n4162 & n7888 ;
  assign n34751 = n34750 ^ n28276 ^ n28130 ;
  assign n34752 = n20983 & n23400 ;
  assign n34753 = n34751 & n34752 ;
  assign n34754 = n34753 ^ n7528 ^ 1'b0 ;
  assign n34755 = n586 & ~n34754 ;
  assign n34756 = n34755 ^ x243 ^ 1'b0 ;
  assign n34757 = ( ~n7616 & n7864 ) | ( ~n7616 & n8045 ) | ( n7864 & n8045 ) ;
  assign n34758 = ( n900 & ~n34743 ) | ( n900 & n34757 ) | ( ~n34743 & n34757 ) ;
  assign n34759 = x135 & n11050 ;
  assign n34760 = ~n25018 & n34759 ;
  assign n34761 = n30596 ^ n7697 ^ 1'b0 ;
  assign n34762 = n11456 | n34503 ;
  assign n34763 = n34762 ^ n29681 ^ 1'b0 ;
  assign n34764 = n2077 | n17103 ;
  assign n34765 = n3851 | n34764 ;
  assign n34766 = n13360 ^ n2386 ^ 1'b0 ;
  assign n34767 = n23360 & ~n34766 ;
  assign n34768 = n34767 ^ n17926 ^ 1'b0 ;
  assign n34769 = n34768 ^ n20059 ^ 1'b0 ;
  assign n34770 = n28386 ^ n13409 ^ 1'b0 ;
  assign n34771 = ~n9707 & n25726 ;
  assign n34772 = n10058 | n19495 ;
  assign n34773 = n27115 ^ n23013 ^ n5649 ;
  assign n34774 = n4079 & ~n34773 ;
  assign n34775 = n23799 & n34774 ;
  assign n34776 = n4989 ^ n4565 ^ 1'b0 ;
  assign n34777 = n3271 & ~n34776 ;
  assign n34778 = n1231 & n34777 ;
  assign n34779 = n12556 ^ n12059 ^ n3970 ;
  assign n34780 = n12387 ^ n9522 ^ 1'b0 ;
  assign n34781 = ~n1538 & n24966 ;
  assign n34785 = n9545 ^ n6874 ^ 1'b0 ;
  assign n34786 = ~n17199 & n34785 ;
  assign n34782 = n4016 | n22824 ;
  assign n34783 = n34782 ^ n17750 ^ 1'b0 ;
  assign n34784 = n3628 | n34783 ;
  assign n34787 = n34786 ^ n34784 ^ 1'b0 ;
  assign n34788 = n15630 | n31945 ;
  assign n34789 = n34788 ^ n18142 ^ 1'b0 ;
  assign n34791 = n5371 ^ x31 ^ 1'b0 ;
  assign n34790 = x18 & ~n6191 ;
  assign n34792 = n34791 ^ n34790 ^ n13521 ;
  assign n34793 = n4079 & ~n34792 ;
  assign n34794 = n1936 & ~n9263 ;
  assign n34795 = n2942 & ~n9941 ;
  assign n34796 = n34795 ^ n12917 ^ 1'b0 ;
  assign n34797 = ( x83 & n34794 ) | ( x83 & ~n34796 ) | ( n34794 & ~n34796 ) ;
  assign n34798 = n7823 ^ n2943 ^ 1'b0 ;
  assign n34799 = n34798 ^ n19440 ^ n4098 ;
  assign n34800 = n34799 ^ n2277 ^ n587 ;
  assign n34801 = n1939 | n34800 ;
  assign n34802 = n11849 & ~n15279 ;
  assign n34803 = n34802 ^ n26027 ^ 1'b0 ;
  assign n34804 = ( n15461 & n34459 ) | ( n15461 & n34803 ) | ( n34459 & n34803 ) ;
  assign n34805 = n32686 ^ n30254 ^ n23427 ;
  assign n34806 = n9719 ^ n5258 ^ n3531 ;
  assign n34807 = ~n12358 & n34806 ;
  assign n34808 = n18360 ^ n10284 ^ 1'b0 ;
  assign n34809 = n24846 & n28986 ;
  assign n34810 = n34809 ^ n31443 ^ 1'b0 ;
  assign n34811 = n9354 & ~n21717 ;
  assign n34812 = n34811 ^ n6432 ^ 1'b0 ;
  assign n34813 = n3698 & ~n10106 ;
  assign n34814 = n18432 & n34813 ;
  assign n34815 = n34814 ^ n18895 ^ 1'b0 ;
  assign n34816 = n27788 ^ n7975 ^ 1'b0 ;
  assign n34817 = n30926 ^ n5031 ^ 1'b0 ;
  assign n34818 = n6291 ^ n1797 ^ 1'b0 ;
  assign n34819 = ( n6506 & n28625 ) | ( n6506 & ~n34818 ) | ( n28625 & ~n34818 ) ;
  assign n34820 = n30208 ^ n26086 ^ n17571 ;
  assign n34821 = n18628 ^ n7970 ^ 1'b0 ;
  assign n34822 = ~n14069 & n34821 ;
  assign n34823 = n12558 & n22332 ;
  assign n34824 = n8284 & ~n11285 ;
  assign n34825 = ~n6515 & n21465 ;
  assign n34826 = n17716 ^ n13250 ^ n12267 ;
  assign n34827 = n4833 & n23764 ;
  assign n34828 = n9176 & n34827 ;
  assign n34829 = ( x202 & ~n3596 ) | ( x202 & n8471 ) | ( ~n3596 & n8471 ) ;
  assign n34830 = ~n5684 & n5889 ;
  assign n34831 = ~n11058 & n34830 ;
  assign n34832 = n13857 ^ n7856 ^ n7850 ;
  assign n34833 = n34832 ^ n29602 ^ 1'b0 ;
  assign n34834 = n11061 ^ n1241 ^ 1'b0 ;
  assign n34835 = ~n5762 & n34834 ;
  assign n34836 = n34835 ^ n10265 ^ 1'b0 ;
  assign n34837 = n34833 | n34836 ;
  assign n34838 = n34837 ^ n32700 ^ 1'b0 ;
  assign n34839 = n34831 & ~n34838 ;
  assign n34840 = n22418 ^ n12002 ^ n8105 ;
  assign n34841 = ( n8685 & n19428 ) | ( n8685 & n32961 ) | ( n19428 & n32961 ) ;
  assign n34842 = ~n28617 & n34841 ;
  assign n34843 = n12433 & n23562 ;
  assign n34844 = ~n3698 & n34843 ;
  assign n34845 = n31237 & n34844 ;
  assign n34846 = n10619 ^ n4200 ^ 1'b0 ;
  assign n34847 = n28718 ^ n8572 ^ 1'b0 ;
  assign n34848 = ~n29827 & n34847 ;
  assign n34849 = n8867 & ~n20752 ;
  assign n34850 = n1168 | n29894 ;
  assign n34852 = n6667 & n19915 ;
  assign n34853 = ~n407 & n34852 ;
  assign n34851 = n3828 | n27523 ;
  assign n34854 = n34853 ^ n34851 ^ 1'b0 ;
  assign n34855 = n20726 & ~n34854 ;
  assign n34856 = n13017 ^ n10829 ^ n2976 ;
  assign n34857 = n34856 ^ n6626 ^ 1'b0 ;
  assign n34858 = n13363 ^ n6779 ^ 1'b0 ;
  assign n34859 = ~n6398 & n34858 ;
  assign n34860 = n34859 ^ n8916 ^ 1'b0 ;
  assign n34861 = x108 & ~n11152 ;
  assign n34862 = ~n895 & n34861 ;
  assign n34863 = n15135 | n34862 ;
  assign n34864 = n34863 ^ n374 ^ 1'b0 ;
  assign n34865 = ~n1192 & n34864 ;
  assign n34866 = n503 | n15963 ;
  assign n34867 = n34866 ^ n13694 ^ n9076 ;
  assign n34868 = n34867 ^ n18801 ^ n2774 ;
  assign n34869 = n22276 | n34868 ;
  assign n34870 = n12203 & ~n34869 ;
  assign n34871 = n34870 ^ n26953 ^ n9417 ;
  assign n34872 = n4567 | n22908 ;
  assign n34873 = ~n612 & n20323 ;
  assign n34874 = n34873 ^ n17116 ^ 1'b0 ;
  assign n34875 = n18073 ^ n17517 ^ n3726 ;
  assign n34876 = ~n8958 & n34875 ;
  assign n34877 = n34876 ^ n21330 ^ 1'b0 ;
  assign n34878 = n34877 ^ n24168 ^ 1'b0 ;
  assign n34879 = n9445 | n14386 ;
  assign n34880 = n17758 | n34879 ;
  assign n34881 = n28444 ^ n26080 ^ 1'b0 ;
  assign n34882 = ~n7189 & n34881 ;
  assign n34883 = n34882 ^ n6339 ^ 1'b0 ;
  assign n34884 = n1613 & n34883 ;
  assign n34885 = n3107 & n14201 ;
  assign n34886 = ~n25379 & n34885 ;
  assign n34887 = n1888 | n34886 ;
  assign n34888 = n34887 ^ n25434 ^ 1'b0 ;
  assign n34894 = ( n1859 & ~n3016 ) | ( n1859 & n7263 ) | ( ~n3016 & n7263 ) ;
  assign n34895 = n32831 & n34894 ;
  assign n34896 = n34895 ^ n24767 ^ 1'b0 ;
  assign n34889 = n10014 ^ n8554 ^ 1'b0 ;
  assign n34890 = n16342 ^ n5992 ^ n5359 ;
  assign n34891 = n34890 ^ n11469 ^ 1'b0 ;
  assign n34892 = n34891 ^ n957 ^ 1'b0 ;
  assign n34893 = n34889 | n34892 ;
  assign n34897 = n34896 ^ n34893 ^ 1'b0 ;
  assign n34898 = ( n22999 & n28574 ) | ( n22999 & n32568 ) | ( n28574 & n32568 ) ;
  assign n34899 = n17756 ^ n15054 ^ 1'b0 ;
  assign n34900 = x213 & n8084 ;
  assign n34901 = n12812 & n34900 ;
  assign n34902 = n34901 ^ n10644 ^ 1'b0 ;
  assign n34903 = n16031 | n16202 ;
  assign n34904 = n33484 | n34903 ;
  assign n34915 = n12544 & ~n22556 ;
  assign n34916 = ~n19975 & n34915 ;
  assign n34910 = n28969 & ~n34679 ;
  assign n34911 = ( n13822 & n22337 ) | ( n13822 & ~n34910 ) | ( n22337 & ~n34910 ) ;
  assign n34905 = n25444 ^ n4623 ^ 1'b0 ;
  assign n34906 = n7231 & n34905 ;
  assign n34907 = n5297 | n13399 ;
  assign n34908 = n34906 & n34907 ;
  assign n34909 = ~n8702 & n34908 ;
  assign n34912 = n34911 ^ n34909 ^ 1'b0 ;
  assign n34913 = ~n21772 & n34912 ;
  assign n34914 = ~n21553 & n34913 ;
  assign n34917 = n34916 ^ n34914 ^ 1'b0 ;
  assign n34918 = n23239 ^ n11201 ^ 1'b0 ;
  assign n34919 = n23665 ^ n8358 ^ n5031 ;
  assign n34920 = n15293 & n29552 ;
  assign n34921 = ~n3766 & n34920 ;
  assign n34922 = n17049 ^ n11370 ^ n3294 ;
  assign n34923 = n894 | n34922 ;
  assign n34924 = n34923 ^ n5245 ^ 1'b0 ;
  assign n34925 = n25106 ^ n5987 ^ 1'b0 ;
  assign n34926 = n34925 ^ n15357 ^ n14259 ;
  assign n34927 = n15421 | n34926 ;
  assign n34928 = n18158 & n34169 ;
  assign n34929 = n11351 | n13497 ;
  assign n34930 = n25233 & ~n34929 ;
  assign n34931 = ( ~n1584 & n5146 ) | ( ~n1584 & n34930 ) | ( n5146 & n34930 ) ;
  assign n34932 = n2268 & n26759 ;
  assign n34933 = ( n5584 & ~n6008 ) | ( n5584 & n34932 ) | ( ~n6008 & n34932 ) ;
  assign n34934 = n31374 ^ n6444 ^ 1'b0 ;
  assign n34935 = n6695 & n18430 ;
  assign n34936 = n9467 & ~n34935 ;
  assign n34937 = n21552 ^ n13821 ^ n13099 ;
  assign n34938 = ~n28481 & n34937 ;
  assign n34939 = n17938 ^ n10100 ^ 1'b0 ;
  assign n34940 = n6298 & n34939 ;
  assign n34941 = x82 & ~n1105 ;
  assign n34942 = n4039 | n11256 ;
  assign n34943 = n34942 ^ n15807 ^ 1'b0 ;
  assign n34944 = ( ~n5894 & n34941 ) | ( ~n5894 & n34943 ) | ( n34941 & n34943 ) ;
  assign n34945 = ( n5156 & n10539 ) | ( n5156 & n34944 ) | ( n10539 & n34944 ) ;
  assign n34946 = n34945 ^ n22180 ^ 1'b0 ;
  assign n34947 = n4890 & ~n8903 ;
  assign n34948 = n34947 ^ n9731 ^ 1'b0 ;
  assign n34949 = n11032 & ~n34948 ;
  assign n34950 = n34949 ^ n17654 ^ n6738 ;
  assign n34951 = n24796 ^ n2331 ^ 1'b0 ;
  assign n34954 = ~n14208 & n28828 ;
  assign n34955 = n34954 ^ n11532 ^ 1'b0 ;
  assign n34952 = ~n21350 & n31059 ;
  assign n34953 = n34952 ^ n32031 ^ 1'b0 ;
  assign n34956 = n34955 ^ n34953 ^ 1'b0 ;
  assign n34957 = n3589 & ~n7326 ;
  assign n34958 = n25769 ^ n8979 ^ 1'b0 ;
  assign n34959 = ~n16047 & n34958 ;
  assign n34962 = n29968 ^ n1734 ^ 1'b0 ;
  assign n34963 = n3521 | n34962 ;
  assign n34960 = n1874 | n15732 ;
  assign n34961 = n3135 & ~n34960 ;
  assign n34964 = n34963 ^ n34961 ^ 1'b0 ;
  assign n34965 = ( ~n5464 & n7986 ) | ( ~n5464 & n14094 ) | ( n7986 & n14094 ) ;
  assign n34966 = ( ~x209 & n29268 ) | ( ~x209 & n34965 ) | ( n29268 & n34965 ) ;
  assign n34967 = ~n2538 & n9404 ;
  assign n34968 = ~n1951 & n34967 ;
  assign n34969 = n16874 | n34968 ;
  assign n34970 = ( ~n1895 & n3456 ) | ( ~n1895 & n16637 ) | ( n3456 & n16637 ) ;
  assign n34971 = n12980 | n14585 ;
  assign n34972 = n34971 ^ n6015 ^ 1'b0 ;
  assign n34973 = ( n2182 & ~n2491 ) | ( n2182 & n10120 ) | ( ~n2491 & n10120 ) ;
  assign n34974 = n34973 ^ n10380 ^ 1'b0 ;
  assign n34975 = ~x57 & n3190 ;
  assign n34976 = n34975 ^ n30486 ^ n3859 ;
  assign n34977 = ( n7440 & n11989 ) | ( n7440 & n17796 ) | ( n11989 & n17796 ) ;
  assign n34978 = ( n3211 & n5631 ) | ( n3211 & ~n34977 ) | ( n5631 & ~n34977 ) ;
  assign n34979 = n5385 | n34978 ;
  assign n34980 = n34976 & ~n34979 ;
  assign n34981 = n24002 ^ n8295 ^ 1'b0 ;
  assign n34982 = n9645 & n34981 ;
  assign n34983 = n34982 ^ n27130 ^ 1'b0 ;
  assign n34984 = ~n29640 & n34983 ;
  assign n34985 = n30046 | n31666 ;
  assign n34986 = n9092 & ~n12134 ;
  assign n34987 = n4861 & ~n18419 ;
  assign n34988 = n10285 | n25546 ;
  assign n34989 = n10544 & ~n34988 ;
  assign n34990 = n34989 ^ n9807 ^ 1'b0 ;
  assign n34991 = n20180 ^ n10405 ^ 1'b0 ;
  assign n34992 = ( n15026 & n19018 ) | ( n15026 & ~n34991 ) | ( n19018 & ~n34991 ) ;
  assign n34993 = n21414 ^ n19572 ^ 1'b0 ;
  assign n34994 = ( n8957 & n27368 ) | ( n8957 & ~n34993 ) | ( n27368 & ~n34993 ) ;
  assign n34995 = ( ~n279 & n2616 ) | ( ~n279 & n5368 ) | ( n2616 & n5368 ) ;
  assign n34996 = n5175 & ~n34995 ;
  assign n34997 = ~n5632 & n34996 ;
  assign n34998 = n5073 & n9561 ;
  assign n34999 = ~x113 & n34998 ;
  assign n35000 = n14968 ^ n5878 ^ 1'b0 ;
  assign n35001 = n34999 | n35000 ;
  assign n35002 = ~n34997 & n35001 ;
  assign n35003 = n22850 ^ n18755 ^ n18558 ;
  assign n35004 = n35003 ^ x146 ^ 1'b0 ;
  assign n35005 = n24746 ^ n10636 ^ 1'b0 ;
  assign n35006 = n7087 & ~n35005 ;
  assign n35007 = n35006 ^ n3498 ^ 1'b0 ;
  assign n35008 = n32442 ^ n11888 ^ n6077 ;
  assign n35009 = n35008 ^ n34650 ^ n26555 ;
  assign n35012 = n20433 ^ n10211 ^ n7080 ;
  assign n35013 = n35012 ^ n1272 ^ 1'b0 ;
  assign n35014 = n13225 & n35013 ;
  assign n35015 = n35014 ^ n293 ^ 1'b0 ;
  assign n35011 = n16003 | n22801 ;
  assign n35016 = n35015 ^ n35011 ^ 1'b0 ;
  assign n35017 = n35016 ^ n17174 ^ n14839 ;
  assign n35018 = n7035 | n27882 ;
  assign n35019 = n35017 | n35018 ;
  assign n35010 = n15550 & n20207 ;
  assign n35020 = n35019 ^ n35010 ^ 1'b0 ;
  assign n35021 = n8718 & n28198 ;
  assign n35022 = ~n24894 & n35021 ;
  assign n35023 = n26329 ^ n9073 ^ 1'b0 ;
  assign n35024 = n35023 ^ n16695 ^ 1'b0 ;
  assign n35025 = ~n19858 & n35024 ;
  assign n35026 = n35025 ^ n23791 ^ 1'b0 ;
  assign n35027 = ~n4878 & n35026 ;
  assign n35028 = ~n7912 & n35027 ;
  assign n35029 = n14855 & n35028 ;
  assign n35030 = n27904 ^ n633 ^ 1'b0 ;
  assign n35031 = n34961 | n35030 ;
  assign n35032 = n15394 ^ n13132 ^ n8307 ;
  assign n35033 = ( n4378 & n8416 ) | ( n4378 & n28262 ) | ( n8416 & n28262 ) ;
  assign n35034 = n17086 ^ n3113 ^ 1'b0 ;
  assign n35035 = ~n3770 & n35034 ;
  assign n35036 = n17623 ^ n6415 ^ 1'b0 ;
  assign n35037 = n35035 & n35036 ;
  assign n35038 = n14989 & ~n35037 ;
  assign n35039 = n35038 ^ n1843 ^ 1'b0 ;
  assign n35041 = n17907 | n18872 ;
  assign n35040 = ( ~n1603 & n1896 ) | ( ~n1603 & n12610 ) | ( n1896 & n12610 ) ;
  assign n35042 = n35041 ^ n35040 ^ 1'b0 ;
  assign n35043 = n30211 & n35042 ;
  assign n35044 = n11345 ^ n2798 ^ 1'b0 ;
  assign n35045 = x120 | n1554 ;
  assign n35046 = n35045 ^ n4193 ^ x25 ;
  assign n35047 = n1224 & ~n35046 ;
  assign n35048 = n35047 ^ n22120 ^ 1'b0 ;
  assign n35049 = ( n12801 & ~n20298 ) | ( n12801 & n22095 ) | ( ~n20298 & n22095 ) ;
  assign n35050 = n35048 | n35049 ;
  assign n35051 = n1416 & n20399 ;
  assign n35052 = n35051 ^ n18917 ^ n3393 ;
  assign n35053 = n11782 ^ x222 ^ 1'b0 ;
  assign n35054 = n25002 | n35053 ;
  assign n35055 = n35054 ^ n30404 ^ 1'b0 ;
  assign n35056 = ( n5658 & ~n6791 ) | ( n5658 & n16949 ) | ( ~n6791 & n16949 ) ;
  assign n35057 = ( ~n31119 & n32424 ) | ( ~n31119 & n35056 ) | ( n32424 & n35056 ) ;
  assign n35058 = n7716 & ~n12321 ;
  assign n35059 = n35058 ^ n5420 ^ 1'b0 ;
  assign n35060 = ( n7240 & n26458 ) | ( n7240 & ~n35059 ) | ( n26458 & ~n35059 ) ;
  assign n35061 = n25527 ^ n2828 ^ 1'b0 ;
  assign n35062 = n33413 | n35061 ;
  assign n35063 = n9037 | n12887 ;
  assign n35064 = n16482 ^ n13216 ^ 1'b0 ;
  assign n35065 = ~n13915 & n35064 ;
  assign n35066 = n3881 & n35065 ;
  assign n35067 = n35066 ^ n13872 ^ 1'b0 ;
  assign n35068 = n27338 ^ n3286 ^ 1'b0 ;
  assign n35070 = ~n2660 & n5755 ;
  assign n35069 = n9444 | n11574 ;
  assign n35071 = n35070 ^ n35069 ^ n13497 ;
  assign n35076 = ( n10304 & n16653 ) | ( n10304 & ~n27775 ) | ( n16653 & ~n27775 ) ;
  assign n35073 = n17960 ^ n16105 ^ 1'b0 ;
  assign n35074 = n27620 & n35073 ;
  assign n35075 = n1536 & n35074 ;
  assign n35077 = n35076 ^ n35075 ^ 1'b0 ;
  assign n35072 = n16006 & n19079 ;
  assign n35078 = n35077 ^ n35072 ^ 1'b0 ;
  assign n35079 = n13448 & n20569 ;
  assign n35080 = ~n24916 & n35079 ;
  assign n35081 = ~n9606 & n10546 ;
  assign n35082 = ~n13560 & n35081 ;
  assign n35083 = ( n1860 & ~n12279 ) | ( n1860 & n29543 ) | ( ~n12279 & n29543 ) ;
  assign n35084 = n8480 & n35083 ;
  assign n35085 = n5589 & ~n26329 ;
  assign n35086 = n9538 & n35085 ;
  assign n35087 = n12611 ^ n4398 ^ n3654 ;
  assign n35088 = ~n11854 & n35087 ;
  assign n35089 = n8679 & ~n26635 ;
  assign n35090 = ( n11758 & n19236 ) | ( n11758 & n33735 ) | ( n19236 & n33735 ) ;
  assign n35091 = n26773 ^ n14470 ^ 1'b0 ;
  assign n35092 = n20853 | n35091 ;
  assign n35093 = n13102 & ~n35092 ;
  assign n35094 = n34488 & ~n35093 ;
  assign n35095 = n21782 ^ n10398 ^ 1'b0 ;
  assign n35096 = ~n20596 & n35095 ;
  assign n35097 = n10851 & n35096 ;
  assign n35098 = ( n18982 & n26828 ) | ( n18982 & ~n35097 ) | ( n26828 & ~n35097 ) ;
  assign n35099 = n21985 ^ n17381 ^ 1'b0 ;
  assign n35100 = n8294 & n35099 ;
  assign n35101 = n6450 & ~n31669 ;
  assign n35102 = n35101 ^ n1519 ^ 1'b0 ;
  assign n35103 = ( n2769 & n6642 ) | ( n2769 & n15936 ) | ( n6642 & n15936 ) ;
  assign n35104 = n35103 ^ n32633 ^ 1'b0 ;
  assign n35105 = ( n6080 & n9068 ) | ( n6080 & n35104 ) | ( n9068 & n35104 ) ;
  assign n35106 = x25 & n7992 ;
  assign n35107 = n35106 ^ n16536 ^ n4837 ;
  assign n35108 = n33411 ^ n14005 ^ n9104 ;
  assign n35109 = n7707 & n8556 ;
  assign n35110 = n11736 & n19696 ;
  assign n35111 = n23481 & n35110 ;
  assign n35112 = n7758 | n8473 ;
  assign n35113 = n9059 | n35112 ;
  assign n35114 = x109 & x228 ;
  assign n35115 = ~n2783 & n35114 ;
  assign n35116 = n35115 ^ n6540 ^ 1'b0 ;
  assign n35117 = ~n19191 & n35116 ;
  assign n35118 = n35117 ^ n897 ^ 1'b0 ;
  assign n35119 = ~n3774 & n35118 ;
  assign n35120 = ~n35113 & n35119 ;
  assign n35121 = n25379 ^ n17840 ^ 1'b0 ;
  assign n35122 = ( n5376 & n29631 ) | ( n5376 & ~n35121 ) | ( n29631 & ~n35121 ) ;
  assign n35123 = n12036 & ~n26495 ;
  assign n35124 = n2261 ^ n374 ^ 1'b0 ;
  assign n35125 = n35124 ^ n19659 ^ n5874 ;
  assign n35126 = n12680 & ~n15767 ;
  assign n35127 = n35126 ^ n783 ^ 1'b0 ;
  assign n35128 = n12786 | n35127 ;
  assign n35129 = ~n6904 & n7243 ;
  assign n35130 = n5162 & n35129 ;
  assign n35131 = n549 | n35130 ;
  assign n35132 = n35131 ^ n21773 ^ 1'b0 ;
  assign n35133 = ~n9466 & n22161 ;
  assign n35134 = ~n440 & n23972 ;
  assign n35135 = n35134 ^ n9129 ^ 1'b0 ;
  assign n35136 = n21963 & n23245 ;
  assign n35137 = ~n35135 & n35136 ;
  assign n35138 = n12382 ^ n11013 ^ n7325 ;
  assign n35139 = n34988 ^ n2126 ^ 1'b0 ;
  assign n35140 = n35138 & n35139 ;
  assign n35141 = n28727 ^ n15887 ^ 1'b0 ;
  assign n35142 = n13167 & ~n35141 ;
  assign n35143 = ( n19764 & n22323 ) | ( n19764 & ~n35142 ) | ( n22323 & ~n35142 ) ;
  assign n35144 = n28281 ^ n2594 ^ 1'b0 ;
  assign n35145 = n33453 ^ n26610 ^ 1'b0 ;
  assign n35146 = ( ~n27003 & n35144 ) | ( ~n27003 & n35145 ) | ( n35144 & n35145 ) ;
  assign n35147 = n16928 ^ n8418 ^ n8047 ;
  assign n35148 = n2089 | n9699 ;
  assign n35149 = n35148 ^ n2978 ^ 1'b0 ;
  assign n35150 = ~n31796 & n35149 ;
  assign n35151 = ~n14139 & n35150 ;
  assign n35152 = n32767 & ~n35151 ;
  assign n35153 = ~n35147 & n35152 ;
  assign n35154 = n27600 ^ n18114 ^ n2847 ;
  assign n35155 = n3857 & ~n5927 ;
  assign n35156 = ~n35154 & n35155 ;
  assign n35157 = n24126 ^ n20671 ^ n1739 ;
  assign n35158 = n35157 ^ n8764 ^ 1'b0 ;
  assign n35159 = n12167 & n35158 ;
  assign n35160 = n21472 ^ n12350 ^ n994 ;
  assign n35161 = n12359 & ~n35160 ;
  assign n35162 = n30730 & n31099 ;
  assign n35164 = n18663 ^ n8829 ^ n5865 ;
  assign n35163 = n15387 & n16869 ;
  assign n35165 = n35164 ^ n35163 ^ 1'b0 ;
  assign n35166 = n35165 ^ n12010 ^ n6603 ;
  assign n35167 = n35166 ^ n10862 ^ n962 ;
  assign n35168 = ( n21816 & ~n33828 ) | ( n21816 & n35167 ) | ( ~n33828 & n35167 ) ;
  assign n35169 = ~n6710 & n8528 ;
  assign n35170 = ( n1506 & n9894 ) | ( n1506 & ~n35169 ) | ( n9894 & ~n35169 ) ;
  assign n35171 = n35170 ^ n11898 ^ 1'b0 ;
  assign n35172 = n17307 & ~n35171 ;
  assign n35173 = ( n6975 & ~n7099 ) | ( n6975 & n34692 ) | ( ~n7099 & n34692 ) ;
  assign n35174 = ~n18936 & n35173 ;
  assign n35175 = n35174 ^ n14136 ^ 1'b0 ;
  assign n35176 = n35175 ^ n31681 ^ n21003 ;
  assign n35177 = n35176 ^ n17865 ^ 1'b0 ;
  assign n35178 = n1888 | n35177 ;
  assign n35179 = n18913 ^ n1624 ^ 1'b0 ;
  assign n35180 = ( n7522 & n18372 ) | ( n7522 & ~n25376 ) | ( n18372 & ~n25376 ) ;
  assign n35181 = ~n22497 & n35180 ;
  assign n35182 = n35179 & n35181 ;
  assign n35183 = n35182 ^ n853 ^ 1'b0 ;
  assign n35184 = n941 & n7883 ;
  assign n35185 = ~n7883 & n35184 ;
  assign n35186 = n11529 ^ n9356 ^ 1'b0 ;
  assign n35187 = n35185 | n35186 ;
  assign n35188 = n35187 ^ n19721 ^ 1'b0 ;
  assign n35189 = ( ~n3344 & n10358 ) | ( ~n3344 & n35188 ) | ( n10358 & n35188 ) ;
  assign n35190 = n11137 ^ n1919 ^ 1'b0 ;
  assign n35191 = ~n19768 & n35190 ;
  assign n35192 = n35191 ^ n26184 ^ 1'b0 ;
  assign n35193 = n19495 & ~n35192 ;
  assign n35194 = ~n29890 & n31185 ;
  assign n35195 = ~n6878 & n35194 ;
  assign n35196 = ( n11044 & n15720 ) | ( n11044 & ~n27891 ) | ( n15720 & ~n27891 ) ;
  assign n35197 = n35196 ^ n720 ^ 1'b0 ;
  assign n35198 = n30284 & ~n35197 ;
  assign n35201 = n13788 ^ n10465 ^ 1'b0 ;
  assign n35202 = ~n2052 & n35201 ;
  assign n35199 = n2125 & ~n11793 ;
  assign n35200 = n20641 & n35199 ;
  assign n35203 = n35202 ^ n35200 ^ n6339 ;
  assign n35204 = n12321 ^ n4460 ^ 1'b0 ;
  assign n35205 = n11351 ^ n2639 ^ 1'b0 ;
  assign n35206 = n9943 & ~n33636 ;
  assign n35207 = n35205 & n35206 ;
  assign n35208 = n18310 | n35207 ;
  assign n35209 = n35204 | n35208 ;
  assign n35210 = ~n7667 & n22389 ;
  assign n35211 = n23284 & n35210 ;
  assign n35212 = n35211 ^ n14319 ^ 1'b0 ;
  assign n35213 = ( n23132 & ~n35209 ) | ( n23132 & n35212 ) | ( ~n35209 & n35212 ) ;
  assign n35214 = ( n17605 & n29525 ) | ( n17605 & ~n31192 ) | ( n29525 & ~n31192 ) ;
  assign n35215 = n31646 ^ n5867 ^ 1'b0 ;
  assign n35216 = ~n17007 & n35215 ;
  assign n35217 = n35216 ^ n34613 ^ 1'b0 ;
  assign n35218 = n14635 | n29453 ;
  assign n35219 = n5749 & ~n35218 ;
  assign n35220 = n9685 & n35219 ;
  assign n35221 = n6733 | n11315 ;
  assign n35222 = ( n4270 & ~n12531 ) | ( n4270 & n35221 ) | ( ~n12531 & n35221 ) ;
  assign n35223 = n26671 | n35222 ;
  assign n35224 = n27302 | n35223 ;
  assign n35225 = n8315 & ~n26646 ;
  assign n35226 = n35225 ^ n17246 ^ 1'b0 ;
  assign n35227 = n19353 ^ n1361 ^ 1'b0 ;
  assign n35228 = n31320 ^ n22398 ^ 1'b0 ;
  assign n35229 = n12092 ^ n3892 ^ n1253 ;
  assign n35230 = ( n5163 & n10142 ) | ( n5163 & ~n35229 ) | ( n10142 & ~n35229 ) ;
  assign n35231 = n9814 ^ n2095 ^ 1'b0 ;
  assign n35232 = n35230 & ~n35231 ;
  assign n35233 = n7639 ^ n4476 ^ 1'b0 ;
  assign n35234 = n17126 & n35233 ;
  assign n35235 = ( n3937 & n15350 ) | ( n3937 & ~n35234 ) | ( n15350 & ~n35234 ) ;
  assign n35236 = ~n9173 & n31540 ;
  assign n35237 = n23675 ^ n13331 ^ 1'b0 ;
  assign n35238 = ~n2931 & n35237 ;
  assign n35239 = n9382 & ~n18517 ;
  assign n35240 = n35239 ^ n28784 ^ 1'b0 ;
  assign n35241 = n10010 & ~n35240 ;
  assign n35242 = ~n5098 & n16645 ;
  assign n35243 = n14415 ^ n775 ^ 1'b0 ;
  assign n35244 = n12976 | n35243 ;
  assign n35245 = n22747 ^ n15356 ^ 1'b0 ;
  assign n35246 = n4153 & ~n35245 ;
  assign n35247 = n35246 ^ n4257 ^ 1'b0 ;
  assign n35249 = n20576 ^ n11854 ^ 1'b0 ;
  assign n35250 = n3056 & ~n35249 ;
  assign n35248 = ~n6683 & n30641 ;
  assign n35251 = n35250 ^ n35248 ^ 1'b0 ;
  assign n35253 = n2111 & n10844 ;
  assign n35254 = n35253 ^ n9332 ^ 1'b0 ;
  assign n35252 = n29108 ^ n10640 ^ 1'b0 ;
  assign n35255 = n35254 ^ n35252 ^ 1'b0 ;
  assign n35256 = n20297 ^ n11680 ^ 1'b0 ;
  assign n35257 = n12034 | n35256 ;
  assign n35258 = n35255 | n35257 ;
  assign n35259 = n27420 | n31562 ;
  assign n35260 = n22114 & n27106 ;
  assign n35261 = n30956 ^ n9858 ^ 1'b0 ;
  assign n35262 = n35260 & ~n35261 ;
  assign n35263 = n13182 & n34214 ;
  assign n35264 = ~n3060 & n9393 ;
  assign n35265 = n35264 ^ n27021 ^ 1'b0 ;
  assign n35266 = ( n16284 & n35263 ) | ( n16284 & n35265 ) | ( n35263 & n35265 ) ;
  assign n35267 = n35266 ^ n16923 ^ 1'b0 ;
  assign n35268 = ( n3605 & ~n10784 ) | ( n3605 & n21460 ) | ( ~n10784 & n21460 ) ;
  assign n35269 = ~n1655 & n23616 ;
  assign n35270 = n35269 ^ n5659 ^ 1'b0 ;
  assign n35271 = n5519 & n9529 ;
  assign n35272 = ~n35270 & n35271 ;
  assign n35273 = n35272 ^ n3649 ^ n1010 ;
  assign n35274 = n20966 & ~n35273 ;
  assign n35275 = ( n25619 & n26408 ) | ( n25619 & n35274 ) | ( n26408 & n35274 ) ;
  assign n35276 = n21180 ^ n13129 ^ n3940 ;
  assign n35277 = ~n22865 & n35276 ;
  assign n35278 = n2107 & ~n16940 ;
  assign n35279 = n35278 ^ n14045 ^ 1'b0 ;
  assign n35280 = n5185 & n6382 ;
  assign n35281 = n35280 ^ n30066 ^ 1'b0 ;
  assign n35282 = n11097 & n27361 ;
  assign n35283 = ~n35281 & n35282 ;
  assign n35284 = ( n10603 & n14809 ) | ( n10603 & n24327 ) | ( n14809 & n24327 ) ;
  assign n35285 = n5818 & ~n35284 ;
  assign n35286 = n24998 | n33003 ;
  assign n35287 = ( ~n11937 & n27158 ) | ( ~n11937 & n35286 ) | ( n27158 & n35286 ) ;
  assign n35288 = n22496 ^ n20747 ^ 1'b0 ;
  assign n35289 = n35287 | n35288 ;
  assign n35290 = n13260 ^ n3490 ^ 1'b0 ;
  assign n35291 = n35290 ^ n16524 ^ n6088 ;
  assign n35292 = n20595 ^ n20008 ^ n1740 ;
  assign n35293 = n27352 ^ n3416 ^ 1'b0 ;
  assign n35294 = n11441 ^ n8717 ^ 1'b0 ;
  assign n35295 = n35294 ^ n2396 ^ 1'b0 ;
  assign n35296 = n18073 & ~n35295 ;
  assign n35297 = n12926 ^ n6326 ^ 1'b0 ;
  assign n35298 = ~n10539 & n35297 ;
  assign n35299 = n8155 ^ n3688 ^ 1'b0 ;
  assign n35300 = n13395 | n35299 ;
  assign n35301 = n2906 & ~n13800 ;
  assign n35302 = ( ~n35298 & n35300 ) | ( ~n35298 & n35301 ) | ( n35300 & n35301 ) ;
  assign n35303 = ( n9780 & n21463 ) | ( n9780 & n28314 ) | ( n21463 & n28314 ) ;
  assign n35304 = n23659 ^ n22952 ^ n15690 ;
  assign n35305 = ~n5443 & n16759 ;
  assign n35306 = ~n25686 & n35305 ;
  assign n35307 = n24246 ^ n8433 ^ 1'b0 ;
  assign n35308 = n21180 & ~n35307 ;
  assign n35309 = n7811 | n8494 ;
  assign n35310 = n9356 ^ n3980 ^ 1'b0 ;
  assign n35311 = ( n28483 & n35309 ) | ( n28483 & n35310 ) | ( n35309 & n35310 ) ;
  assign n35312 = n35311 ^ n33043 ^ 1'b0 ;
  assign n35313 = n15154 & n35312 ;
  assign n35314 = n2584 | n15438 ;
  assign n35315 = ( ~n8845 & n28235 ) | ( ~n8845 & n35314 ) | ( n28235 & n35314 ) ;
  assign n35316 = n14467 ^ n13806 ^ 1'b0 ;
  assign n35317 = n35316 ^ n26348 ^ n3047 ;
  assign n35318 = n31164 ^ n25917 ^ 1'b0 ;
  assign n35319 = ~n9335 & n35318 ;
  assign n35320 = n35319 ^ n14731 ^ 1'b0 ;
  assign n35321 = n35317 & n35320 ;
  assign n35322 = n26926 ^ n14489 ^ 1'b0 ;
  assign n35323 = n4638 & n27921 ;
  assign n35324 = n19793 ^ n12635 ^ n12010 ;
  assign n35325 = ~n35323 & n35324 ;
  assign n35326 = n13345 & ~n16455 ;
  assign n35327 = n35326 ^ n10758 ^ 1'b0 ;
  assign n35328 = n35327 ^ n6071 ^ 1'b0 ;
  assign n35329 = ~n20072 & n35328 ;
  assign n35330 = n35329 ^ n25436 ^ n2278 ;
  assign n35331 = n35330 ^ n12601 ^ 1'b0 ;
  assign n35332 = ~n34442 & n35331 ;
  assign n35333 = n4072 & n14636 ;
  assign n35334 = n35333 ^ n7661 ^ 1'b0 ;
  assign n35335 = n13505 & n35334 ;
  assign n35336 = n35335 ^ n2399 ^ 1'b0 ;
  assign n35340 = n3327 & n12764 ;
  assign n35341 = ~n997 & n35340 ;
  assign n35342 = n35341 ^ n7497 ^ 1'b0 ;
  assign n35343 = ~n5732 & n35342 ;
  assign n35337 = ( n1925 & n9872 ) | ( n1925 & ~n11022 ) | ( n9872 & ~n11022 ) ;
  assign n35338 = n3182 & ~n35337 ;
  assign n35339 = ~n8222 & n35338 ;
  assign n35344 = n35343 ^ n35339 ^ 1'b0 ;
  assign n35345 = n19897 | n29750 ;
  assign n35346 = n35345 ^ n17496 ^ 1'b0 ;
  assign n35347 = n9277 ^ n6817 ^ 1'b0 ;
  assign n35348 = n3344 & n35347 ;
  assign n35349 = n35348 ^ n4361 ^ 1'b0 ;
  assign n35350 = ( n10372 & ~n28269 ) | ( n10372 & n35349 ) | ( ~n28269 & n35349 ) ;
  assign n35351 = n3826 & ~n7325 ;
  assign n35352 = n17597 & ~n21487 ;
  assign n35353 = n35352 ^ n24269 ^ 1'b0 ;
  assign n35354 = ~n9709 & n22820 ;
  assign n35355 = n35353 & n35354 ;
  assign n35356 = n12037 ^ n4469 ^ 1'b0 ;
  assign n35357 = n2964 | n35356 ;
  assign n35360 = n10762 ^ n10220 ^ n9012 ;
  assign n35358 = ~n3051 & n8198 ;
  assign n35359 = n7132 & n35358 ;
  assign n35361 = n35360 ^ n35359 ^ n13308 ;
  assign n35362 = n5246 & n11475 ;
  assign n35363 = n35362 ^ n26346 ^ 1'b0 ;
  assign n35364 = n13734 ^ n4991 ^ n3854 ;
  assign n35365 = n35115 ^ n21156 ^ n14038 ;
  assign n35366 = n35365 ^ n17700 ^ 1'b0 ;
  assign n35367 = n13877 & n35366 ;
  assign n35368 = x90 | n11187 ;
  assign n35369 = n21067 & ~n35368 ;
  assign n35370 = ( n6530 & n31985 ) | ( n6530 & n35369 ) | ( n31985 & n35369 ) ;
  assign n35371 = ( n616 & ~n9777 ) | ( n616 & n29958 ) | ( ~n9777 & n29958 ) ;
  assign n35372 = n35370 & n35371 ;
  assign n35373 = n35372 ^ n23702 ^ 1'b0 ;
  assign n35374 = n7218 & ~n9743 ;
  assign n35375 = n26496 & n35374 ;
  assign n35376 = ( n24271 & n25125 ) | ( n24271 & ~n35375 ) | ( n25125 & ~n35375 ) ;
  assign n35377 = n35376 ^ n19752 ^ 1'b0 ;
  assign n35378 = ~n9146 & n35377 ;
  assign n35379 = n12642 | n15571 ;
  assign n35380 = n30221 | n35379 ;
  assign n35381 = n31161 ^ n12218 ^ 1'b0 ;
  assign n35382 = n33069 ^ n8819 ^ 1'b0 ;
  assign n35383 = n17317 & ~n35382 ;
  assign n35384 = n4677 & ~n12232 ;
  assign n35385 = n18872 & n35384 ;
  assign n35386 = n11266 ^ n5702 ^ 1'b0 ;
  assign n35387 = n3924 | n35386 ;
  assign n35388 = n22913 ^ n18913 ^ 1'b0 ;
  assign n35389 = ~n7391 & n18770 ;
  assign n35390 = n34862 & n35389 ;
  assign n35391 = n14528 ^ n9860 ^ n8665 ;
  assign n35394 = ~n7320 & n13105 ;
  assign n35395 = n4425 & ~n30369 ;
  assign n35396 = ~n35394 & n35395 ;
  assign n35392 = n22442 ^ n21075 ^ 1'b0 ;
  assign n35393 = ( ~n6068 & n16617 ) | ( ~n6068 & n35392 ) | ( n16617 & n35392 ) ;
  assign n35397 = n35396 ^ n35393 ^ n10606 ;
  assign n35398 = x57 & ~n22483 ;
  assign n35399 = n29999 ^ n8681 ^ 1'b0 ;
  assign n35400 = n10032 ^ n6764 ^ 1'b0 ;
  assign n35401 = n17006 | n35400 ;
  assign n35402 = n26296 ^ n1168 ^ 1'b0 ;
  assign n35403 = n9061 ^ n4129 ^ 1'b0 ;
  assign n35404 = n35403 ^ n9668 ^ n5416 ;
  assign n35405 = ( ~n1871 & n4556 ) | ( ~n1871 & n15198 ) | ( n4556 & n15198 ) ;
  assign n35406 = n5476 & ~n10157 ;
  assign n35407 = n35405 & n35406 ;
  assign n35408 = n19806 ^ n7009 ^ 1'b0 ;
  assign n35411 = n35234 ^ n677 ^ 1'b0 ;
  assign n35409 = n33041 ^ n5337 ^ n3771 ;
  assign n35410 = ~n33541 & n35409 ;
  assign n35412 = n35411 ^ n35410 ^ 1'b0 ;
  assign n35413 = n1553 | n9746 ;
  assign n35414 = n19642 | n33867 ;
  assign n35416 = ~n1859 & n5172 ;
  assign n35415 = n7523 & n24487 ;
  assign n35417 = n35416 ^ n35415 ^ 1'b0 ;
  assign n35418 = ( n7725 & n19851 ) | ( n7725 & n20334 ) | ( n19851 & n20334 ) ;
  assign n35419 = ~n27170 & n35418 ;
  assign n35420 = n15971 & n24400 ;
  assign n35421 = n12147 & ~n31148 ;
  assign n35422 = n35421 ^ n22265 ^ 1'b0 ;
  assign n35423 = n1243 & n9131 ;
  assign n35424 = ~n22598 & n35423 ;
  assign n35425 = n3915 & ~n35424 ;
  assign n35426 = n16140 | n35425 ;
  assign n35427 = n18374 | n35426 ;
  assign n35428 = n35427 ^ n10381 ^ 1'b0 ;
  assign n35429 = n6898 ^ n5384 ^ n5094 ;
  assign n35430 = ( n2103 & n28982 ) | ( n2103 & ~n35429 ) | ( n28982 & ~n35429 ) ;
  assign n35431 = n7780 | n34098 ;
  assign n35432 = n35431 ^ n30434 ^ 1'b0 ;
  assign n35433 = n3203 | n15694 ;
  assign n35434 = n6065 & ~n35433 ;
  assign n35435 = n35434 ^ n8362 ^ 1'b0 ;
  assign n35436 = n27103 & n35435 ;
  assign n35437 = n32744 ^ n9716 ^ 1'b0 ;
  assign n35438 = ~n3628 & n35437 ;
  assign n35439 = n33704 ^ n15936 ^ n14689 ;
  assign n35440 = ( n20576 & ~n26638 ) | ( n20576 & n32433 ) | ( ~n26638 & n32433 ) ;
  assign n35441 = n35440 ^ n16027 ^ n9266 ;
  assign n35443 = ~n3232 & n23468 ;
  assign n35444 = n14722 & n35443 ;
  assign n35442 = ~n3203 & n31787 ;
  assign n35445 = n35444 ^ n35442 ^ 1'b0 ;
  assign n35447 = n29040 ^ n4446 ^ 1'b0 ;
  assign n35446 = n4717 & ~n17674 ;
  assign n35448 = n35447 ^ n35446 ^ 1'b0 ;
  assign n35449 = n27136 ^ n790 ^ 1'b0 ;
  assign n35450 = n5618 | n18635 ;
  assign n35451 = n1880 & ~n35450 ;
  assign n35452 = n34891 & ~n35451 ;
  assign n35453 = n15134 ^ n14243 ^ n4153 ;
  assign n35454 = n35453 ^ n31192 ^ 1'b0 ;
  assign n35455 = n33084 & ~n35454 ;
  assign n35456 = ( n4825 & n14374 ) | ( n4825 & n35455 ) | ( n14374 & n35455 ) ;
  assign n35457 = n21749 & n22293 ;
  assign n35458 = n2481 | n4293 ;
  assign n35459 = n35458 ^ n2546 ^ 1'b0 ;
  assign n35460 = n19670 & ~n35459 ;
  assign n35461 = ~n35457 & n35460 ;
  assign n35462 = ( x100 & n16205 ) | ( x100 & n18728 ) | ( n16205 & n18728 ) ;
  assign n35463 = n11470 | n35462 ;
  assign n35464 = n18650 & ~n22879 ;
  assign n35465 = n35464 ^ n31909 ^ 1'b0 ;
  assign n35466 = n1845 & ~n11448 ;
  assign n35467 = n33756 ^ n1106 ^ 1'b0 ;
  assign n35468 = n10199 | n35467 ;
  assign n35469 = ( ~n1786 & n35466 ) | ( ~n1786 & n35468 ) | ( n35466 & n35468 ) ;
  assign n35470 = n35469 ^ n17874 ^ n16662 ;
  assign n35471 = ( n5112 & n16844 ) | ( n5112 & ~n35470 ) | ( n16844 & ~n35470 ) ;
  assign n35472 = n1879 ^ x207 ^ 1'b0 ;
  assign n35473 = n7182 & ~n35472 ;
  assign n35474 = n35473 ^ n2103 ^ 1'b0 ;
  assign n35475 = n29299 & ~n35474 ;
  assign n35476 = n13127 ^ n2169 ^ 1'b0 ;
  assign n35477 = ~n3523 & n5613 ;
  assign n35478 = n8346 & n35477 ;
  assign n35479 = n35478 ^ n27907 ^ 1'b0 ;
  assign n35480 = n35476 & n35479 ;
  assign n35481 = n7472 & n23509 ;
  assign n35482 = ( n1060 & n16678 ) | ( n1060 & n35481 ) | ( n16678 & n35481 ) ;
  assign n35483 = n10075 & ~n20992 ;
  assign n35484 = n35483 ^ n19101 ^ n12197 ;
  assign n35485 = n1111 & ~n14779 ;
  assign n35486 = n7966 & n35485 ;
  assign n35487 = n17938 | n33608 ;
  assign n35488 = n18861 ^ n1270 ^ 1'b0 ;
  assign n35489 = ( n813 & ~n7564 ) | ( n813 & n26412 ) | ( ~n7564 & n26412 ) ;
  assign n35490 = n20471 ^ n15713 ^ n7386 ;
  assign n35491 = ( n16161 & n35489 ) | ( n16161 & n35490 ) | ( n35489 & n35490 ) ;
  assign n35492 = n35491 ^ n29280 ^ n2605 ;
  assign n35493 = n5608 & ~n12214 ;
  assign n35494 = n35493 ^ n22896 ^ n17669 ;
  assign n35495 = n23541 | n35494 ;
  assign n35497 = n18793 ^ n18552 ^ 1'b0 ;
  assign n35498 = n4934 & n35497 ;
  assign n35499 = ~n17172 & n35498 ;
  assign n35496 = n6253 | n17642 ;
  assign n35500 = n35499 ^ n35496 ^ 1'b0 ;
  assign n35501 = n12535 ^ n11110 ^ 1'b0 ;
  assign n35502 = ~n6069 & n19775 ;
  assign n35503 = n11214 & n35502 ;
  assign n35504 = n35503 ^ n13167 ^ 1'b0 ;
  assign n35505 = n35501 | n35504 ;
  assign n35506 = ( n1247 & ~n8490 ) | ( n1247 & n12378 ) | ( ~n8490 & n12378 ) ;
  assign n35507 = n35506 ^ n26916 ^ n5798 ;
  assign n35508 = n35507 ^ n31945 ^ 1'b0 ;
  assign n35509 = n4812 | n35508 ;
  assign n35510 = n10164 ^ n3576 ^ x162 ;
  assign n35511 = ( n3847 & n5929 ) | ( n3847 & ~n35510 ) | ( n5929 & ~n35510 ) ;
  assign n35516 = n1953 & n9892 ;
  assign n35515 = n1161 | n10099 ;
  assign n35517 = n35516 ^ n35515 ^ n13144 ;
  assign n35512 = n23852 ^ n2293 ^ 1'b0 ;
  assign n35513 = n35512 ^ n16635 ^ 1'b0 ;
  assign n35514 = ( n14587 & ~n16499 ) | ( n14587 & n35513 ) | ( ~n16499 & n35513 ) ;
  assign n35518 = n35517 ^ n35514 ^ n22016 ;
  assign n35519 = ~n10160 & n10683 ;
  assign n35520 = n35519 ^ n18552 ^ 1'b0 ;
  assign n35521 = n12646 | n23468 ;
  assign n35522 = n35521 ^ n9552 ^ 1'b0 ;
  assign n35523 = n35522 ^ n11726 ^ 1'b0 ;
  assign n35524 = n609 | n1289 ;
  assign n35525 = n5824 | n35524 ;
  assign n35526 = n24949 & n35525 ;
  assign n35527 = n13140 & n35526 ;
  assign n35528 = n8076 & n35527 ;
  assign n35529 = ( n4108 & n6213 ) | ( n4108 & n27435 ) | ( n6213 & n27435 ) ;
  assign n35530 = n24394 | n35529 ;
  assign n35531 = n35530 ^ n17619 ^ 1'b0 ;
  assign n35532 = n22415 ^ n18568 ^ n9326 ;
  assign n35533 = n34925 ^ n14226 ^ n5551 ;
  assign n35534 = n10645 | n35533 ;
  assign n35535 = n292 & n18366 ;
  assign n35536 = n22790 ^ n19507 ^ n12670 ;
  assign n35537 = ~n10194 & n35536 ;
  assign n35538 = n21886 & n27099 ;
  assign n35539 = ~n1802 & n35538 ;
  assign n35540 = n27194 ^ n11133 ^ 1'b0 ;
  assign n35541 = n11397 & ~n35540 ;
  assign n35542 = n9048 & n14135 ;
  assign n35543 = n22439 ^ n6436 ^ 1'b0 ;
  assign n35544 = n15796 & ~n35543 ;
  assign n35545 = n35542 & n35544 ;
  assign n35546 = n23244 ^ n16880 ^ 1'b0 ;
  assign n35547 = n19239 ^ n709 ^ 1'b0 ;
  assign n35548 = n718 & ~n35547 ;
  assign n35549 = n23550 ^ n13321 ^ 1'b0 ;
  assign n35550 = ( n12032 & n35548 ) | ( n12032 & n35549 ) | ( n35548 & n35549 ) ;
  assign n35551 = ( n9700 & n14672 ) | ( n9700 & ~n18594 ) | ( n14672 & ~n18594 ) ;
  assign n35552 = n8272 & n9572 ;
  assign n35553 = n20433 ^ n10450 ^ 1'b0 ;
  assign n35554 = n17767 | n35553 ;
  assign n35555 = n7932 | n20115 ;
  assign n35556 = n35555 ^ n6453 ^ 1'b0 ;
  assign n35557 = n35556 ^ n27269 ^ 1'b0 ;
  assign n35558 = ~n282 & n35557 ;
  assign n35559 = n454 & n3211 ;
  assign n35560 = n35559 ^ n1657 ^ 1'b0 ;
  assign n35561 = n10356 & ~n35560 ;
  assign n35562 = n35561 ^ n27523 ^ n24103 ;
  assign n35563 = ~n10234 & n35562 ;
  assign n35564 = ~n35558 & n35563 ;
  assign n35565 = n11823 & ~n21056 ;
  assign n35566 = n32439 ^ n24583 ^ n20878 ;
  assign n35567 = n2746 & n9260 ;
  assign n35568 = n8580 & n10311 ;
  assign n35569 = n35568 ^ n22498 ^ n18435 ;
  assign n35570 = ( n5062 & n5767 ) | ( n5062 & n12035 ) | ( n5767 & n12035 ) ;
  assign n35571 = ~n5126 & n35570 ;
  assign n35572 = ~n25911 & n35571 ;
  assign n35573 = n10434 & ~n10712 ;
  assign n35574 = n35573 ^ n2462 ^ 1'b0 ;
  assign n35575 = ( n3054 & ~n3268 ) | ( n3054 & n7182 ) | ( ~n3268 & n7182 ) ;
  assign n35576 = n31587 & ~n35575 ;
  assign n35577 = n35576 ^ n31698 ^ 1'b0 ;
  assign n35578 = ~n26108 & n35577 ;
  assign n35579 = n5684 | n16837 ;
  assign n35580 = n35579 ^ n20049 ^ 1'b0 ;
  assign n35581 = n35580 ^ n27420 ^ n6723 ;
  assign n35582 = n16531 ^ n8278 ^ 1'b0 ;
  assign n35583 = ( n862 & n2538 ) | ( n862 & n35582 ) | ( n2538 & n35582 ) ;
  assign n35584 = ~n18586 & n22407 ;
  assign n35585 = n26308 ^ n16927 ^ 1'b0 ;
  assign n35586 = n14452 | n35585 ;
  assign n35587 = n8009 & ~n9582 ;
  assign n35588 = ~n1045 & n35587 ;
  assign n35589 = n4039 | n35588 ;
  assign n35590 = n35589 ^ n18026 ^ 1'b0 ;
  assign n35591 = ~n9300 & n23988 ;
  assign n35592 = n35591 ^ n6453 ^ 1'b0 ;
  assign n35594 = n8161 & n9272 ;
  assign n35595 = n16497 & n35594 ;
  assign n35593 = n12908 & ~n34138 ;
  assign n35596 = n35595 ^ n35593 ^ 1'b0 ;
  assign n35597 = ~n8017 & n20138 ;
  assign n35598 = n6428 & n7592 ;
  assign n35599 = n35598 ^ n27561 ^ n4904 ;
  assign n35600 = ( ~n263 & n1054 ) | ( ~n263 & n22554 ) | ( n1054 & n22554 ) ;
  assign n35601 = ( n1596 & n4790 ) | ( n1596 & ~n35600 ) | ( n4790 & ~n35600 ) ;
  assign n35602 = n28737 ^ n21345 ^ n1890 ;
  assign n35603 = n22568 | n31398 ;
  assign n35604 = n25585 & ~n26042 ;
  assign n35605 = n35604 ^ n10571 ^ 1'b0 ;
  assign n35606 = n17633 & ~n35605 ;
  assign n35607 = n5370 & n18224 ;
  assign n35608 = ~n8805 & n35607 ;
  assign n35609 = ~n23785 & n33209 ;
  assign n35610 = n15590 ^ n7893 ^ 1'b0 ;
  assign n35611 = ~n25450 & n35610 ;
  assign n35612 = ~n2850 & n5969 ;
  assign n35613 = n35612 ^ n10662 ^ 1'b0 ;
  assign n35614 = n6910 | n31820 ;
  assign n35615 = n25237 ^ n1388 ^ 1'b0 ;
  assign n35617 = n7504 | n15750 ;
  assign n35616 = n3566 | n7267 ;
  assign n35618 = n35617 ^ n35616 ^ 1'b0 ;
  assign n35619 = n3666 & n4896 ;
  assign n35620 = n35619 ^ n27977 ^ 1'b0 ;
  assign n35621 = n34540 ^ n8634 ^ 1'b0 ;
  assign n35622 = n22866 | n35621 ;
  assign n35623 = n4346 & ~n35622 ;
  assign n35624 = n19501 ^ n18395 ^ 1'b0 ;
  assign n35625 = n35624 ^ n23086 ^ 1'b0 ;
  assign n35626 = n23237 & ~n35625 ;
  assign n35627 = ~n30489 & n35626 ;
  assign n35628 = ~n16682 & n35627 ;
  assign n35629 = n26812 ^ n10372 ^ 1'b0 ;
  assign n35630 = n26590 | n35629 ;
  assign n35631 = n10408 ^ n5538 ^ n455 ;
  assign n35632 = n7553 ^ n266 ^ 1'b0 ;
  assign n35633 = n35632 ^ n32961 ^ n3332 ;
  assign n35634 = n35633 ^ n31303 ^ n4024 ;
  assign n35635 = ( ~n5815 & n31262 ) | ( ~n5815 & n35634 ) | ( n31262 & n35634 ) ;
  assign n35636 = n24374 ^ n619 ^ 1'b0 ;
  assign n35637 = n35636 ^ n18931 ^ n5998 ;
  assign n35638 = n35637 ^ n34164 ^ n2289 ;
  assign n35639 = ~n3943 & n24609 ;
  assign n35640 = ~n7358 & n12799 ;
  assign n35641 = n14993 ^ n3016 ^ 1'b0 ;
  assign n35642 = n5607 & ~n25611 ;
  assign n35643 = n35641 & n35642 ;
  assign n35647 = n2090 & n2645 ;
  assign n35648 = ~n1366 & n35647 ;
  assign n35649 = n3159 ^ n2769 ^ n807 ;
  assign n35650 = n12831 & n35649 ;
  assign n35651 = ( ~n8275 & n35648 ) | ( ~n8275 & n35650 ) | ( n35648 & n35650 ) ;
  assign n35644 = n16171 & n20901 ;
  assign n35645 = ~n19346 & n35644 ;
  assign n35646 = n16422 | n35645 ;
  assign n35652 = n35651 ^ n35646 ^ 1'b0 ;
  assign n35653 = n1388 | n20115 ;
  assign n35654 = n11101 ^ n8481 ^ 1'b0 ;
  assign n35655 = n26021 & n35654 ;
  assign n35656 = ~n25037 & n35655 ;
  assign n35657 = n2580 | n3797 ;
  assign n35658 = n2687 | n35657 ;
  assign n35659 = ( n1247 & n20437 ) | ( n1247 & ~n35658 ) | ( n20437 & ~n35658 ) ;
  assign n35660 = ~n22186 & n23494 ;
  assign n35661 = ( n1657 & n3402 ) | ( n1657 & n8484 ) | ( n3402 & n8484 ) ;
  assign n35662 = ~n4120 & n35661 ;
  assign n35663 = n35662 ^ n25019 ^ 1'b0 ;
  assign n35664 = n978 | n35663 ;
  assign n35665 = ( n21894 & n22590 ) | ( n21894 & ~n28507 ) | ( n22590 & ~n28507 ) ;
  assign n35666 = ~n2313 & n35665 ;
  assign n35669 = ~n1617 & n6866 ;
  assign n35667 = n5206 & n8588 ;
  assign n35668 = n35667 ^ n22917 ^ n12373 ;
  assign n35670 = n35669 ^ n35668 ^ 1'b0 ;
  assign n35671 = n35670 ^ n3429 ^ n2498 ;
  assign n35672 = n1203 & n16869 ;
  assign n35673 = n35672 ^ n34680 ^ 1'b0 ;
  assign n35674 = n2431 & n15015 ;
  assign n35675 = n2323 & n35674 ;
  assign n35676 = ( n12794 & n17033 ) | ( n12794 & ~n24089 ) | ( n17033 & ~n24089 ) ;
  assign n35677 = n917 & ~n35676 ;
  assign n35678 = n4799 | n29693 ;
  assign n35679 = n7029 | n35678 ;
  assign n35680 = n23497 & n32253 ;
  assign n35681 = n13205 & n35680 ;
  assign n35682 = ( n2401 & n27116 ) | ( n2401 & n35681 ) | ( n27116 & n35681 ) ;
  assign n35683 = n3947 | n13533 ;
  assign n35684 = n35683 ^ n27573 ^ n4391 ;
  assign n35685 = n9196 ^ n6759 ^ 1'b0 ;
  assign n35686 = n11353 & ~n35685 ;
  assign n35687 = n28906 ^ n22663 ^ 1'b0 ;
  assign n35688 = n2245 & n16248 ;
  assign n35689 = n19801 & n35688 ;
  assign n35690 = n7987 & ~n35689 ;
  assign n35691 = n12508 ^ n11912 ^ 1'b0 ;
  assign n35692 = ~n35690 & n35691 ;
  assign n35693 = n34297 ^ n16977 ^ 1'b0 ;
  assign n35694 = ~n21656 & n35693 ;
  assign n35695 = n13461 | n16937 ;
  assign n35696 = n35695 ^ n20055 ^ 1'b0 ;
  assign n35697 = n35696 ^ n32398 ^ n19692 ;
  assign n35698 = n33711 ^ n7943 ^ 1'b0 ;
  assign n35699 = n6597 ^ n3093 ^ x253 ;
  assign n35700 = n13012 ^ n5459 ^ n1814 ;
  assign n35701 = n3364 & n7948 ;
  assign n35702 = ( n35699 & ~n35700 ) | ( n35699 & n35701 ) | ( ~n35700 & n35701 ) ;
  assign n35703 = n8120 | n33447 ;
  assign n35704 = n35703 ^ n24347 ^ 1'b0 ;
  assign n35705 = ~n16118 & n28224 ;
  assign n35706 = ~x116 & n35705 ;
  assign n35707 = n8679 | n8883 ;
  assign n35708 = n35707 ^ n7813 ^ 1'b0 ;
  assign n35709 = n24250 & n35708 ;
  assign n35710 = n3614 & n18589 ;
  assign n35711 = ~n35709 & n35710 ;
  assign n35712 = n27774 ^ n2835 ^ 1'b0 ;
  assign n35713 = n19704 ^ n13604 ^ n1076 ;
  assign n35714 = n656 & ~n12673 ;
  assign n35715 = ~n26609 & n35714 ;
  assign n35716 = n2874 | n35715 ;
  assign n35717 = n35713 | n35716 ;
  assign n35718 = n1422 & ~n13862 ;
  assign n35719 = n15802 & n35718 ;
  assign n35720 = n35719 ^ n13475 ^ 1'b0 ;
  assign n35721 = ( n17104 & n17315 ) | ( n17104 & n29257 ) | ( n17315 & n29257 ) ;
  assign n35722 = n1034 ^ x181 ^ 1'b0 ;
  assign n35723 = n5128 ^ n482 ^ 1'b0 ;
  assign n35724 = n5119 & n35723 ;
  assign n35725 = ( x113 & n35722 ) | ( x113 & ~n35724 ) | ( n35722 & ~n35724 ) ;
  assign n35726 = ( ~n17832 & n35721 ) | ( ~n17832 & n35725 ) | ( n35721 & n35725 ) ;
  assign n35727 = n35726 ^ n33287 ^ 1'b0 ;
  assign n35728 = n11046 & n35727 ;
  assign n35729 = n12995 ^ n3585 ^ 1'b0 ;
  assign n35730 = ( n5411 & ~n9751 ) | ( n5411 & n35729 ) | ( ~n9751 & n35729 ) ;
  assign n35731 = n32906 ^ n6436 ^ n3767 ;
  assign n35732 = n33762 ^ n2326 ^ 1'b0 ;
  assign n35733 = n27526 | n35732 ;
  assign n35736 = n6422 | n24949 ;
  assign n35734 = n18452 ^ n16844 ^ 1'b0 ;
  assign n35735 = ~n7959 & n35734 ;
  assign n35737 = n35736 ^ n35735 ^ 1'b0 ;
  assign n35738 = n4118 & ~n29733 ;
  assign n35739 = n19134 ^ n15578 ^ 1'b0 ;
  assign n35740 = n1220 | n20100 ;
  assign n35741 = n17627 & n35008 ;
  assign n35742 = ~n21015 & n26341 ;
  assign n35743 = n35742 ^ n20601 ^ 1'b0 ;
  assign n35744 = n5973 | n6350 ;
  assign n35745 = n35744 ^ n13221 ^ n1636 ;
  assign n35747 = n1325 | n15219 ;
  assign n35746 = ~n13970 & n25042 ;
  assign n35748 = n35747 ^ n35746 ^ n18525 ;
  assign n35749 = n35748 ^ n3634 ^ 1'b0 ;
  assign n35750 = ( n9356 & n15782 ) | ( n9356 & ~n19810 ) | ( n15782 & ~n19810 ) ;
  assign n35751 = ~n2315 & n17862 ;
  assign n35752 = n29351 & n35751 ;
  assign n35753 = n5022 | n12301 ;
  assign n35757 = n13779 ^ n12296 ^ 1'b0 ;
  assign n35755 = n19428 ^ n2349 ^ 1'b0 ;
  assign n35756 = n15347 & ~n35755 ;
  assign n35758 = n35757 ^ n35756 ^ n6944 ;
  assign n35754 = x150 | n5398 ;
  assign n35759 = n35758 ^ n35754 ^ 1'b0 ;
  assign n35760 = n25552 ^ n14725 ^ 1'b0 ;
  assign n35761 = n20742 ^ n16713 ^ n1005 ;
  assign n35762 = n23588 ^ n10334 ^ n6332 ;
  assign n35763 = n8477 ^ n6524 ^ 1'b0 ;
  assign n35764 = n20323 & ~n35763 ;
  assign n35765 = n35764 ^ x155 ^ 1'b0 ;
  assign n35766 = n2877 ^ n2423 ^ 1'b0 ;
  assign n35767 = ( n13358 & ~n16347 ) | ( n13358 & n35766 ) | ( ~n16347 & n35766 ) ;
  assign n35768 = n4469 & ~n35767 ;
  assign n35769 = n16363 ^ n12049 ^ 1'b0 ;
  assign n35770 = n3389 & ~n5548 ;
  assign n35771 = n7895 & n35770 ;
  assign n35772 = n35771 ^ n17326 ^ n14637 ;
  assign n35773 = ( n981 & n35769 ) | ( n981 & n35772 ) | ( n35769 & n35772 ) ;
  assign n35777 = ~n10860 & n12220 ;
  assign n35774 = n32253 ^ n12550 ^ 1'b0 ;
  assign n35775 = n5991 & ~n35774 ;
  assign n35776 = n672 | n35775 ;
  assign n35778 = n35777 ^ n35776 ^ n29150 ;
  assign n35779 = n35778 ^ n25471 ^ n5504 ;
  assign n35780 = n11582 | n22908 ;
  assign n35782 = ( n8143 & n8466 ) | ( n8143 & n10130 ) | ( n8466 & n10130 ) ;
  assign n35781 = n1793 & ~n29972 ;
  assign n35783 = n35782 ^ n35781 ^ 1'b0 ;
  assign n35784 = n33880 & n35783 ;
  assign n35785 = n716 & n26045 ;
  assign n35786 = n35785 ^ n6303 ^ 1'b0 ;
  assign n35787 = n1981 | n6562 ;
  assign n35788 = n15584 ^ x240 ^ 1'b0 ;
  assign n35789 = ( ~n11052 & n12491 ) | ( ~n11052 & n35788 ) | ( n12491 & n35788 ) ;
  assign n35790 = n19926 ^ n3580 ^ 1'b0 ;
  assign n35791 = ( n4302 & ~n14804 ) | ( n4302 & n20144 ) | ( ~n14804 & n20144 ) ;
  assign n35792 = n15033 & n35791 ;
  assign n35793 = n10258 | n21042 ;
  assign n35794 = n23335 ^ n2717 ^ 1'b0 ;
  assign n35795 = n13640 & n35794 ;
  assign n35796 = n10563 ^ n2435 ^ 1'b0 ;
  assign n35797 = n11697 | n30019 ;
  assign n35798 = n35796 & n35797 ;
  assign n35799 = n7946 & ~n18742 ;
  assign n35800 = n12066 & n35799 ;
  assign n35801 = ( n8191 & n16682 ) | ( n8191 & ~n35800 ) | ( n16682 & ~n35800 ) ;
  assign n35802 = ~n2616 & n35801 ;
  assign n35803 = ( n19685 & n29428 ) | ( n19685 & n35802 ) | ( n29428 & n35802 ) ;
  assign n35804 = n21892 ^ n17333 ^ 1'b0 ;
  assign n35805 = ( x13 & n23448 ) | ( x13 & ~n35804 ) | ( n23448 & ~n35804 ) ;
  assign n35806 = n12576 & n32363 ;
  assign n35807 = ( ~n14032 & n21651 ) | ( ~n14032 & n31547 ) | ( n21651 & n31547 ) ;
  assign n35808 = n5624 | n35807 ;
  assign n35809 = n9260 ^ n6074 ^ 1'b0 ;
  assign n35810 = n35808 & ~n35809 ;
  assign n35812 = n35529 ^ n23117 ^ 1'b0 ;
  assign n35813 = n28754 & ~n35812 ;
  assign n35811 = n15969 ^ n14059 ^ 1'b0 ;
  assign n35814 = n35813 ^ n35811 ^ 1'b0 ;
  assign n35815 = n10919 ^ n4611 ^ 1'b0 ;
  assign n35816 = n7858 & n25690 ;
  assign n35817 = n35816 ^ n17532 ^ 1'b0 ;
  assign n35818 = n12768 ^ n9954 ^ 1'b0 ;
  assign n35819 = n3217 | n35818 ;
  assign n35820 = n35819 ^ n447 ^ 1'b0 ;
  assign n35821 = n2178 & n29199 ;
  assign n35822 = n35821 ^ n14698 ^ 1'b0 ;
  assign n35823 = ( n356 & ~n3079 ) | ( n356 & n4516 ) | ( ~n3079 & n4516 ) ;
  assign n35824 = ( n968 & n21048 ) | ( n968 & ~n35823 ) | ( n21048 & ~n35823 ) ;
  assign n35825 = n14816 | n35824 ;
  assign n35826 = n35825 ^ n15562 ^ 1'b0 ;
  assign n35827 = ~n3357 & n12888 ;
  assign n35828 = n35827 ^ n18159 ^ 1'b0 ;
  assign n35829 = n6246 & n9539 ;
  assign n35830 = n11540 & ~n16717 ;
  assign n35831 = n35829 & n35830 ;
  assign n35832 = n35831 ^ n4659 ^ 1'b0 ;
  assign n35833 = n7391 & n35832 ;
  assign n35834 = ( n8155 & ~n22692 ) | ( n8155 & n30722 ) | ( ~n22692 & n30722 ) ;
  assign n35835 = n30133 | n35834 ;
  assign n35836 = n28040 ^ n23099 ^ 1'b0 ;
  assign n35837 = n6783 & ~n23848 ;
  assign n35838 = n32693 & n35837 ;
  assign n35839 = ~n1227 & n31170 ;
  assign n35840 = n35839 ^ n7839 ^ 1'b0 ;
  assign n35841 = n25189 ^ n23007 ^ 1'b0 ;
  assign n35842 = ~n35164 & n35655 ;
  assign n35843 = ( ~n20797 & n35841 ) | ( ~n20797 & n35842 ) | ( n35841 & n35842 ) ;
  assign n35844 = n27188 | n30605 ;
  assign n35845 = n17994 ^ n7549 ^ n2701 ;
  assign n35846 = x28 & n16252 ;
  assign n35847 = n35846 ^ n20158 ^ 1'b0 ;
  assign n35848 = n12702 ^ n5342 ^ 1'b0 ;
  assign n35849 = n1886 | n35848 ;
  assign n35850 = n35847 & ~n35849 ;
  assign n35851 = ~n14344 & n35850 ;
  assign n35852 = ~n2691 & n8303 ;
  assign n35853 = ~n8520 & n35852 ;
  assign n35854 = n35853 ^ n22699 ^ 1'b0 ;
  assign n35855 = n27851 & n35854 ;
  assign n35856 = n35855 ^ n6779 ^ 1'b0 ;
  assign n35859 = n10966 & ~n13142 ;
  assign n35860 = n35859 ^ n11285 ^ 1'b0 ;
  assign n35858 = n7906 | n27852 ;
  assign n35857 = ( n1128 & n11276 ) | ( n1128 & ~n28693 ) | ( n11276 & ~n28693 ) ;
  assign n35861 = n35860 ^ n35858 ^ n35857 ;
  assign n35862 = ( n13391 & n14709 ) | ( n13391 & ~n24916 ) | ( n14709 & ~n24916 ) ;
  assign n35863 = n25975 ^ n13278 ^ 1'b0 ;
  assign n35864 = n8449 ^ n3553 ^ 1'b0 ;
  assign n35865 = n14405 | n35864 ;
  assign n35866 = n35865 ^ n24456 ^ 1'b0 ;
  assign n35867 = n3837 & n35866 ;
  assign n35868 = ~n35863 & n35867 ;
  assign n35869 = ( ~n11863 & n18266 ) | ( ~n11863 & n19873 ) | ( n18266 & n19873 ) ;
  assign n35870 = n31881 ^ n17678 ^ 1'b0 ;
  assign n35871 = n14019 ^ n6523 ^ n4014 ;
  assign n35872 = n2679 & ~n22357 ;
  assign n35873 = ~n35871 & n35872 ;
  assign n35875 = ( n10495 & n13858 ) | ( n10495 & n26966 ) | ( n13858 & n26966 ) ;
  assign n35874 = ~n9221 & n11457 ;
  assign n35876 = n35875 ^ n35874 ^ 1'b0 ;
  assign n35879 = ( ~n6930 & n18420 ) | ( ~n6930 & n20157 ) | ( n18420 & n20157 ) ;
  assign n35877 = n15032 & n19768 ;
  assign n35878 = n34287 & n35877 ;
  assign n35880 = n35879 ^ n35878 ^ 1'b0 ;
  assign n35881 = ~n8713 & n35880 ;
  assign n35882 = n8049 & n10243 ;
  assign n35883 = n35882 ^ n20443 ^ 1'b0 ;
  assign n35884 = n29100 ^ n4991 ^ 1'b0 ;
  assign n35885 = n35883 | n35884 ;
  assign n35886 = n35885 ^ n9666 ^ 1'b0 ;
  assign n35887 = n20767 & n35886 ;
  assign n35888 = n35887 ^ n23978 ^ 1'b0 ;
  assign n35889 = n34468 ^ n33663 ^ 1'b0 ;
  assign n35890 = n10629 & n23741 ;
  assign n35891 = n35890 ^ n10395 ^ 1'b0 ;
  assign n35892 = ( n6053 & n14527 ) | ( n6053 & ~n34922 ) | ( n14527 & ~n34922 ) ;
  assign n35893 = n29624 & ~n35892 ;
  assign n35894 = ( n329 & ~n35767 ) | ( n329 & n35893 ) | ( ~n35767 & n35893 ) ;
  assign n35895 = n35894 ^ n10121 ^ 1'b0 ;
  assign n35896 = n35891 & ~n35895 ;
  assign n35897 = n35896 ^ n27209 ^ 1'b0 ;
  assign n35898 = n12796 ^ x231 ^ 1'b0 ;
  assign n35899 = n12543 | n35898 ;
  assign n35900 = n2401 ^ n738 ^ 1'b0 ;
  assign n35901 = ~n35899 & n35900 ;
  assign n35902 = n35901 ^ n23852 ^ n19640 ;
  assign n35903 = n15532 ^ n7480 ^ n6182 ;
  assign n35904 = n35903 ^ n35494 ^ 1'b0 ;
  assign n35905 = n1450 & ~n18700 ;
  assign n35906 = ~n1886 & n15213 ;
  assign n35907 = ( n34374 & ~n35905 ) | ( n34374 & n35906 ) | ( ~n35905 & n35906 ) ;
  assign n35908 = n1385 | n7798 ;
  assign n35909 = n25762 & ~n35908 ;
  assign n35910 = n11357 | n35909 ;
  assign n35911 = n35910 ^ n19529 ^ 1'b0 ;
  assign n35912 = ~n2735 & n4581 ;
  assign n35913 = n35912 ^ n6015 ^ 1'b0 ;
  assign n35914 = n29109 & n33772 ;
  assign n35915 = ~n9030 & n19435 ;
  assign n35916 = ( n5662 & n35139 ) | ( n5662 & ~n35915 ) | ( n35139 & ~n35915 ) ;
  assign n35918 = n30700 & n34078 ;
  assign n35919 = n35918 ^ n12768 ^ 1'b0 ;
  assign n35917 = ~n12094 & n20680 ;
  assign n35920 = n35919 ^ n35917 ^ n12619 ;
  assign n35921 = ( n10335 & n34161 ) | ( n10335 & ~n35920 ) | ( n34161 & ~n35920 ) ;
  assign n35923 = n21489 ^ n9842 ^ 1'b0 ;
  assign n35924 = ~n34495 & n35923 ;
  assign n35922 = ~n17750 & n21305 ;
  assign n35925 = n35924 ^ n35922 ^ 1'b0 ;
  assign n35926 = ( n1891 & n6848 ) | ( n1891 & n32334 ) | ( n6848 & n32334 ) ;
  assign n35927 = n10642 & ~n14454 ;
  assign n35928 = n2210 ^ x227 ^ 1'b0 ;
  assign n35929 = n35928 ^ n20829 ^ 1'b0 ;
  assign n35930 = n2818 & n19070 ;
  assign n35931 = n35930 ^ n35347 ^ 1'b0 ;
  assign n35932 = n11017 & ~n19491 ;
  assign n35933 = n2840 | n9719 ;
  assign n35934 = n10910 | n20438 ;
  assign n35935 = n35933 | n35934 ;
  assign n35936 = n35935 ^ n14986 ^ 1'b0 ;
  assign n35937 = n35932 & ~n35936 ;
  assign n35939 = n9963 & ~n25877 ;
  assign n35938 = n9398 & ~n23238 ;
  assign n35940 = n35939 ^ n35938 ^ 1'b0 ;
  assign n35941 = n15894 | n20858 ;
  assign n35942 = n25010 | n35941 ;
  assign n35943 = n18960 ^ n2242 ^ 1'b0 ;
  assign n35944 = ~n1906 & n7047 ;
  assign n35945 = n35944 ^ n3740 ^ 1'b0 ;
  assign n35946 = n27270 ^ n14880 ^ 1'b0 ;
  assign n35947 = ~n28148 & n35946 ;
  assign n35948 = ( ~n19734 & n22017 ) | ( ~n19734 & n34391 ) | ( n22017 & n34391 ) ;
  assign n35949 = n7769 & ~n21604 ;
  assign n35950 = n13887 | n23545 ;
  assign n35951 = n35950 ^ n12099 ^ 1'b0 ;
  assign n35952 = ( n13092 & n26550 ) | ( n13092 & n35951 ) | ( n26550 & n35951 ) ;
  assign n35953 = n13006 ^ n1928 ^ 1'b0 ;
  assign n35954 = n35953 ^ n22251 ^ 1'b0 ;
  assign n35955 = n11242 & n35954 ;
  assign n35956 = ( n5752 & n19411 ) | ( n5752 & ~n30988 ) | ( n19411 & ~n30988 ) ;
  assign n35957 = n35956 ^ n3641 ^ 1'b0 ;
  assign n35958 = n29506 & n35957 ;
  assign n35960 = n14796 | n24158 ;
  assign n35961 = n26370 | n35960 ;
  assign n35962 = n35961 ^ n34618 ^ 1'b0 ;
  assign n35959 = ~n10624 & n27225 ;
  assign n35963 = n35962 ^ n35959 ^ n26083 ;
  assign n35965 = n4492 | n31905 ;
  assign n35966 = n15919 & ~n35965 ;
  assign n35967 = n8351 & n35966 ;
  assign n35964 = n27101 ^ n21123 ^ 1'b0 ;
  assign n35968 = n35967 ^ n35964 ^ 1'b0 ;
  assign n35969 = ~n10998 & n19781 ;
  assign n35971 = ~n4034 & n7366 ;
  assign n35972 = n35971 ^ n3771 ^ 1'b0 ;
  assign n35970 = n13593 & n16556 ;
  assign n35973 = n35972 ^ n35970 ^ n533 ;
  assign n35974 = n17039 & ~n35973 ;
  assign n35975 = n4247 | n8213 ;
  assign n35976 = n4247 & ~n35975 ;
  assign n35977 = n7345 & ~n35976 ;
  assign n35978 = n17639 & n35977 ;
  assign n35979 = ~n1463 & n15410 ;
  assign n35980 = n35978 & n35979 ;
  assign n35981 = x249 & ~n35980 ;
  assign n35982 = n31022 ^ n866 ^ 1'b0 ;
  assign n35983 = ~n4635 & n35982 ;
  assign n35984 = n14743 | n17383 ;
  assign n35985 = n6043 & ~n35984 ;
  assign n35988 = n2857 & ~n8157 ;
  assign n35989 = n35988 ^ n6856 ^ 1'b0 ;
  assign n35990 = n35989 ^ n10768 ^ n1476 ;
  assign n35986 = n12207 | n23587 ;
  assign n35987 = n2277 & ~n35986 ;
  assign n35991 = n35990 ^ n35987 ^ n21506 ;
  assign n35992 = n5333 & ~n35991 ;
  assign n35993 = n19674 | n24113 ;
  assign n35994 = n4902 & ~n23422 ;
  assign n35995 = ~n35993 & n35994 ;
  assign n35996 = ( ~n22267 & n23343 ) | ( ~n22267 & n35995 ) | ( n23343 & n35995 ) ;
  assign n35997 = ~n2987 & n35996 ;
  assign n35998 = n1536 & ~n27010 ;
  assign n35999 = n16360 ^ n14586 ^ n12084 ;
  assign n36000 = ~n9764 & n12591 ;
  assign n36001 = n11285 | n36000 ;
  assign n36002 = n30972 ^ x217 ^ 1'b0 ;
  assign n36003 = ~n32012 & n36002 ;
  assign n36004 = n36003 ^ n7060 ^ 1'b0 ;
  assign n36005 = n25415 ^ n11973 ^ n11322 ;
  assign n36006 = n956 | n36005 ;
  assign n36007 = n36006 ^ n1350 ^ 1'b0 ;
  assign n36008 = n36007 ^ n25049 ^ 1'b0 ;
  assign n36009 = ~n36004 & n36008 ;
  assign n36010 = ( n9035 & n15378 ) | ( n9035 & n17736 ) | ( n15378 & n17736 ) ;
  assign n36011 = n11801 ^ n11719 ^ 1'b0 ;
  assign n36012 = n879 & ~n36011 ;
  assign n36013 = ~n32607 & n36012 ;
  assign n36014 = n36013 ^ n3657 ^ 1'b0 ;
  assign n36015 = ( n13749 & ~n14159 ) | ( n13749 & n14170 ) | ( ~n14159 & n14170 ) ;
  assign n36016 = n24367 & n36015 ;
  assign n36017 = n14863 | n34833 ;
  assign n36018 = n4585 & ~n36017 ;
  assign n36019 = x193 & ~n36018 ;
  assign n36020 = n14889 ^ n4001 ^ 1'b0 ;
  assign n36021 = n36019 & n36020 ;
  assign n36022 = n22937 & n36021 ;
  assign n36025 = n18850 ^ n11945 ^ 1'b0 ;
  assign n36023 = n10266 ^ n1496 ^ 1'b0 ;
  assign n36024 = n1387 & n36023 ;
  assign n36026 = n36025 ^ n36024 ^ 1'b0 ;
  assign n36027 = ~n17443 & n24907 ;
  assign n36028 = n284 | n10243 ;
  assign n36029 = ( n18668 & n34174 ) | ( n18668 & n36028 ) | ( n34174 & n36028 ) ;
  assign n36030 = n16044 ^ n3883 ^ 1'b0 ;
  assign n36031 = ~n9604 & n36030 ;
  assign n36032 = n36031 ^ n1378 ^ 1'b0 ;
  assign n36033 = n14791 | n36032 ;
  assign n36034 = n11133 | n36033 ;
  assign n36035 = n34308 | n36034 ;
  assign n36036 = n17899 ^ n5593 ^ 1'b0 ;
  assign n36037 = n2244 & ~n36036 ;
  assign n36038 = n36037 ^ n29782 ^ 1'b0 ;
  assign n36039 = n36035 & ~n36038 ;
  assign n36040 = ~n5848 & n16882 ;
  assign n36041 = n36040 ^ n26232 ^ 1'b0 ;
  assign n36042 = ~n21951 & n36041 ;
  assign n36043 = ~n36039 & n36042 ;
  assign n36044 = n8589 ^ n2586 ^ 1'b0 ;
  assign n36045 = ~n6537 & n6557 ;
  assign n36046 = n36045 ^ n29196 ^ 1'b0 ;
  assign n36047 = ( n5185 & ~n6724 ) | ( n5185 & n16559 ) | ( ~n6724 & n16559 ) ;
  assign n36048 = n36047 ^ n15273 ^ 1'b0 ;
  assign n36049 = n6373 & n36048 ;
  assign n36050 = n887 & n16899 ;
  assign n36051 = ~n27701 & n30427 ;
  assign n36052 = n36051 ^ n25579 ^ 1'b0 ;
  assign n36053 = n36052 ^ x10 ^ 1'b0 ;
  assign n36054 = n15217 & n24599 ;
  assign n36055 = n5153 ^ n338 ^ 1'b0 ;
  assign n36057 = n30928 ^ n11128 ^ 1'b0 ;
  assign n36058 = ~n5128 & n36057 ;
  assign n36056 = ~n5081 & n29922 ;
  assign n36059 = n36058 ^ n36056 ^ n17674 ;
  assign n36060 = n32617 ^ n24035 ^ n844 ;
  assign n36061 = n13063 | n13546 ;
  assign n36062 = n36061 ^ n31922 ^ n11884 ;
  assign n36063 = ( n2385 & n5141 ) | ( n2385 & n36062 ) | ( n5141 & n36062 ) ;
  assign n36064 = n15059 ^ n3862 ^ 1'b0 ;
  assign n36065 = n20450 & ~n36064 ;
  assign n36066 = ( ~n911 & n2256 ) | ( ~n911 & n9626 ) | ( n2256 & n9626 ) ;
  assign n36067 = n36066 ^ n9644 ^ 1'b0 ;
  assign n36068 = n26657 | n36067 ;
  assign n36069 = n18120 ^ n2212 ^ n1082 ;
  assign n36070 = n27797 & ~n36069 ;
  assign n36071 = n1875 & n36070 ;
  assign n36072 = ~n24513 & n36071 ;
  assign n36073 = n18276 ^ n14880 ^ 1'b0 ;
  assign n36074 = n2385 | n35588 ;
  assign n36075 = n36074 ^ n1671 ^ 1'b0 ;
  assign n36076 = n11215 & ~n26009 ;
  assign n36077 = n6262 & ~n36076 ;
  assign n36078 = n36077 ^ n12764 ^ 1'b0 ;
  assign n36079 = ( n5658 & ~n19123 ) | ( n5658 & n22160 ) | ( ~n19123 & n22160 ) ;
  assign n36080 = n36079 ^ n23494 ^ n3047 ;
  assign n36081 = n18817 ^ n13116 ^ n9333 ;
  assign n36082 = n28462 ^ n5263 ^ 1'b0 ;
  assign n36083 = n22951 | n36082 ;
  assign n36084 = n23745 ^ n16649 ^ 1'b0 ;
  assign n36085 = n8362 | n34639 ;
  assign n36086 = n10272 & ~n36085 ;
  assign n36089 = n5522 ^ n3466 ^ 1'b0 ;
  assign n36087 = ( n12306 & ~n17822 ) | ( n12306 & n29963 ) | ( ~n17822 & n29963 ) ;
  assign n36088 = n36087 ^ n33738 ^ n15283 ;
  assign n36090 = n36089 ^ n36088 ^ n4612 ;
  assign n36092 = n10785 & ~n25710 ;
  assign n36093 = n476 & n36092 ;
  assign n36091 = n18858 & ~n27005 ;
  assign n36094 = n36093 ^ n36091 ^ n9316 ;
  assign n36095 = n10539 | n15807 ;
  assign n36096 = n4804 & n12145 ;
  assign n36097 = n36096 ^ n21508 ^ 1'b0 ;
  assign n36098 = n33484 & n36097 ;
  assign n36099 = n396 | n14168 ;
  assign n36100 = n36099 ^ x184 ^ 1'b0 ;
  assign n36101 = ~n11242 & n20506 ;
  assign n36102 = n28129 ^ n20453 ^ 1'b0 ;
  assign n36103 = n36101 & ~n36102 ;
  assign n36104 = n26287 & ~n36103 ;
  assign n36105 = ~n13731 & n18120 ;
  assign n36106 = ~n33373 & n36105 ;
  assign n36107 = n9682 ^ n9562 ^ 1'b0 ;
  assign n36108 = n18861 ^ n3960 ^ 1'b0 ;
  assign n36109 = n33145 ^ n16642 ^ n4237 ;
  assign n36110 = n9165 | n27345 ;
  assign n36111 = ~n20119 & n24160 ;
  assign n36112 = n36111 ^ n10691 ^ 1'b0 ;
  assign n36114 = n725 | n14002 ;
  assign n36115 = ~n10860 & n35516 ;
  assign n36116 = n36115 ^ n15991 ^ 1'b0 ;
  assign n36117 = ( n11437 & n36114 ) | ( n11437 & ~n36116 ) | ( n36114 & ~n36116 ) ;
  assign n36113 = n1385 | n1989 ;
  assign n36118 = n36117 ^ n36113 ^ 1'b0 ;
  assign n36119 = n12886 ^ n7119 ^ 1'b0 ;
  assign n36120 = n6514 | n36119 ;
  assign n36121 = n36120 ^ n1746 ^ 1'b0 ;
  assign n36122 = ~n9858 & n27775 ;
  assign n36123 = ( n7554 & n12305 ) | ( n7554 & ~n36122 ) | ( n12305 & ~n36122 ) ;
  assign n36124 = n18483 & n25421 ;
  assign n36125 = n36124 ^ n35113 ^ 1'b0 ;
  assign n36126 = ( n23438 & n31897 ) | ( n23438 & n36125 ) | ( n31897 & n36125 ) ;
  assign n36127 = n1388 & ~n8284 ;
  assign n36128 = n36127 ^ n10847 ^ n8121 ;
  assign n36129 = n11510 & ~n36128 ;
  assign n36130 = n36126 & n36129 ;
  assign n36131 = ( ~n11446 & n17965 ) | ( ~n11446 & n36130 ) | ( n17965 & n36130 ) ;
  assign n36132 = ~n5408 & n20336 ;
  assign n36133 = n10355 & n36132 ;
  assign n36134 = n31664 | n32639 ;
  assign n36135 = n22251 & ~n36134 ;
  assign n36136 = n1154 & ~n36135 ;
  assign n36137 = n36136 ^ n16073 ^ 1'b0 ;
  assign n36138 = n18656 ^ n16363 ^ n4423 ;
  assign n36139 = n457 & n24213 ;
  assign n36140 = ~n10932 & n36139 ;
  assign n36141 = ( n15575 & ~n24037 ) | ( n15575 & n36140 ) | ( ~n24037 & n36140 ) ;
  assign n36142 = n8438 & ~n11105 ;
  assign n36143 = ( ~n24024 & n36141 ) | ( ~n24024 & n36142 ) | ( n36141 & n36142 ) ;
  assign n36144 = n34308 & n36143 ;
  assign n36145 = ~n6124 & n20238 ;
  assign n36146 = ~n451 & n36145 ;
  assign n36147 = ~n30412 & n35448 ;
  assign n36148 = ~n19278 & n36147 ;
  assign n36149 = n19461 ^ n18666 ^ 1'b0 ;
  assign n36150 = n9117 | n24432 ;
  assign n36151 = n36150 ^ n12698 ^ 1'b0 ;
  assign n36153 = ( ~n20076 & n22469 ) | ( ~n20076 & n24445 ) | ( n22469 & n24445 ) ;
  assign n36152 = n5752 & ~n17146 ;
  assign n36154 = n36153 ^ n36152 ^ 1'b0 ;
  assign n36155 = n36154 ^ n32651 ^ 1'b0 ;
  assign n36156 = ~n36151 & n36155 ;
  assign n36157 = n3138 | n25110 ;
  assign n36158 = n36157 ^ n8488 ^ 1'b0 ;
  assign n36159 = n6157 | n25592 ;
  assign n36160 = n616 & n36159 ;
  assign n36161 = n36158 & n36160 ;
  assign n36162 = ~n15597 & n24098 ;
  assign n36163 = n36162 ^ n19115 ^ 1'b0 ;
  assign n36164 = n5347 & n21188 ;
  assign n36165 = n36164 ^ n32182 ^ 1'b0 ;
  assign n36166 = n26949 | n36165 ;
  assign n36168 = ( ~n13012 & n35205 ) | ( ~n13012 & n35892 ) | ( n35205 & n35892 ) ;
  assign n36169 = n11883 & n36168 ;
  assign n36170 = n36169 ^ n20404 ^ 1'b0 ;
  assign n36167 = n9142 & n12831 ;
  assign n36171 = n36170 ^ n36167 ^ 1'b0 ;
  assign n36172 = n17796 ^ x81 ^ 1'b0 ;
  assign n36173 = ~n14684 & n36172 ;
  assign n36174 = n1107 & ~n22847 ;
  assign n36175 = ~n13618 & n36174 ;
  assign n36176 = n14226 & ~n36175 ;
  assign n36177 = n18476 & ~n23452 ;
  assign n36178 = n11223 & ~n11377 ;
  assign n36179 = n28125 ^ n9360 ^ 1'b0 ;
  assign n36180 = n36178 | n36179 ;
  assign n36181 = n3322 & ~n15206 ;
  assign n36182 = n36181 ^ n22453 ^ 1'b0 ;
  assign n36183 = n24259 ^ n8391 ^ n5386 ;
  assign n36184 = ~n36182 & n36183 ;
  assign n36185 = ~n2178 & n29501 ;
  assign n36186 = n36185 ^ n15438 ^ 1'b0 ;
  assign n36187 = n18383 ^ n12841 ^ 1'b0 ;
  assign n36188 = ( ~n7240 & n27380 ) | ( ~n7240 & n36187 ) | ( n27380 & n36187 ) ;
  assign n36189 = n2993 ^ n2885 ^ 1'b0 ;
  assign n36190 = ( n1979 & n11451 ) | ( n1979 & ~n36189 ) | ( n11451 & ~n36189 ) ;
  assign n36191 = n36190 ^ n21105 ^ 1'b0 ;
  assign n36192 = n36188 & n36191 ;
  assign n36193 = ( n28020 & n36186 ) | ( n28020 & n36192 ) | ( n36186 & n36192 ) ;
  assign n36195 = n1308 & ~n22546 ;
  assign n36196 = n6904 & n36195 ;
  assign n36194 = n5377 & n17212 ;
  assign n36197 = n36196 ^ n36194 ^ n11837 ;
  assign n36198 = n8128 ^ n1116 ^ 1'b0 ;
  assign n36199 = n15579 | n36198 ;
  assign n36200 = n34479 ^ n28040 ^ 1'b0 ;
  assign n36201 = ~n36199 & n36200 ;
  assign n36202 = n2082 | n5987 ;
  assign n36203 = x125 | n36202 ;
  assign n36204 = n18631 ^ n10986 ^ 1'b0 ;
  assign n36205 = n36203 & n36204 ;
  assign n36206 = n1367 | n11666 ;
  assign n36207 = n36206 ^ n11159 ^ 1'b0 ;
  assign n36208 = n16969 & ~n18496 ;
  assign n36209 = n36208 ^ n34791 ^ 1'b0 ;
  assign n36210 = n15944 ^ n15730 ^ 1'b0 ;
  assign n36211 = ( n6201 & ~n8026 ) | ( n6201 & n27515 ) | ( ~n8026 & n27515 ) ;
  assign n36212 = n27226 & n36211 ;
  assign n36213 = n12579 ^ n11149 ^ 1'b0 ;
  assign n36214 = ~n3291 & n36213 ;
  assign n36215 = ~n17239 & n36214 ;
  assign n36216 = n36215 ^ n7848 ^ 1'b0 ;
  assign n36217 = ( ~x105 & n19413 ) | ( ~x105 & n32441 ) | ( n19413 & n32441 ) ;
  assign n36218 = n27594 ^ n18365 ^ n13041 ;
  assign n36219 = n36218 ^ n15526 ^ n9139 ;
  assign n36220 = n3095 & ~n23106 ;
  assign n36221 = n36220 ^ n22478 ^ n264 ;
  assign n36225 = n19529 ^ n5739 ^ n4197 ;
  assign n36222 = n5066 & ~n15136 ;
  assign n36223 = ~n24429 & n36222 ;
  assign n36224 = n3597 & ~n36223 ;
  assign n36226 = n36225 ^ n36224 ^ 1'b0 ;
  assign n36228 = n12359 ^ n9850 ^ n1650 ;
  assign n36227 = ( n6037 & n6351 ) | ( n6037 & ~n12391 ) | ( n6351 & ~n12391 ) ;
  assign n36229 = n36228 ^ n36227 ^ n10416 ;
  assign n36231 = n12953 ^ n4870 ^ n445 ;
  assign n36230 = n3368 | n14300 ;
  assign n36232 = n36231 ^ n36230 ^ 1'b0 ;
  assign n36233 = n36232 ^ n30987 ^ n810 ;
  assign n36234 = n29037 ^ n27166 ^ n12197 ;
  assign n36235 = n15517 & ~n36234 ;
  assign n36236 = n36235 ^ n14754 ^ 1'b0 ;
  assign n36237 = n30530 & n36236 ;
  assign n36238 = n18204 & n36237 ;
  assign n36239 = n3172 & n17821 ;
  assign n36240 = n10214 ^ n5183 ^ 1'b0 ;
  assign n36241 = n6919 & n36240 ;
  assign n36242 = n30092 ^ n3299 ^ n3072 ;
  assign n36243 = ( n13050 & ~n13164 ) | ( n13050 & n16570 ) | ( ~n13164 & n16570 ) ;
  assign n36244 = n36242 | n36243 ;
  assign n36245 = n1784 & n20501 ;
  assign n36246 = n36245 ^ n4561 ^ 1'b0 ;
  assign n36247 = n36246 ^ n30109 ^ n2682 ;
  assign n36248 = ~n18948 & n19431 ;
  assign n36249 = ~n25372 & n36248 ;
  assign n36250 = n36249 ^ n35019 ^ 1'b0 ;
  assign n36251 = ~n36247 & n36250 ;
  assign n36252 = n6865 ^ n6106 ^ 1'b0 ;
  assign n36253 = ~n16470 & n36252 ;
  assign n36254 = n26756 ^ n16168 ^ 1'b0 ;
  assign n36255 = n13521 | n36254 ;
  assign n36261 = n2445 & n14161 ;
  assign n36256 = n13148 ^ n1325 ^ 1'b0 ;
  assign n36257 = n3669 & ~n36256 ;
  assign n36258 = n36257 ^ n3552 ^ 1'b0 ;
  assign n36259 = ~n4449 & n36258 ;
  assign n36260 = n36259 ^ n22782 ^ n6664 ;
  assign n36262 = n36261 ^ n36260 ^ 1'b0 ;
  assign n36263 = ~n15115 & n36262 ;
  assign n36266 = n26162 ^ n9866 ^ 1'b0 ;
  assign n36267 = ~n8965 & n36266 ;
  assign n36264 = n9185 & ~n17353 ;
  assign n36265 = ( n29325 & ~n29983 ) | ( n29325 & n36264 ) | ( ~n29983 & n36264 ) ;
  assign n36268 = n36267 ^ n36265 ^ n2643 ;
  assign n36269 = ~n23098 & n29642 ;
  assign n36270 = n424 | n25627 ;
  assign n36271 = n13119 ^ n11840 ^ n8116 ;
  assign n36272 = n36271 ^ n2680 ^ 1'b0 ;
  assign n36273 = n30013 & n36272 ;
  assign n36274 = n4807 | n11707 ;
  assign n36275 = n36274 ^ n4612 ^ 1'b0 ;
  assign n36276 = n20779 ^ n13554 ^ n450 ;
  assign n36277 = ~n3651 & n27899 ;
  assign n36278 = n36277 ^ n33903 ^ 1'b0 ;
  assign n36279 = n20143 | n30322 ;
  assign n36280 = n23616 & ~n36279 ;
  assign n36281 = ~n19754 & n36280 ;
  assign n36282 = n7315 & ~n9776 ;
  assign n36283 = ~n25338 & n36282 ;
  assign n36284 = ( n9634 & n13860 ) | ( n9634 & n36283 ) | ( n13860 & n36283 ) ;
  assign n36285 = n18800 & ~n36284 ;
  assign n36286 = n36281 & n36285 ;
  assign n36287 = ~n2387 & n3000 ;
  assign n36288 = n23631 ^ n8341 ^ 1'b0 ;
  assign n36289 = n23505 & n36288 ;
  assign n36290 = ~n8538 & n36289 ;
  assign n36291 = n36290 ^ n14801 ^ 1'b0 ;
  assign n36292 = n36291 ^ n35079 ^ n2051 ;
  assign n36293 = n28441 ^ n13444 ^ n12522 ;
  assign n36294 = n23351 | n36293 ;
  assign n36295 = n36294 ^ n6310 ^ 1'b0 ;
  assign n36296 = n24093 ^ n20861 ^ 1'b0 ;
  assign n36297 = ~n5842 & n36296 ;
  assign n36298 = ~n10503 & n13066 ;
  assign n36299 = n8507 ^ n7304 ^ 1'b0 ;
  assign n36300 = ~n15671 & n36299 ;
  assign n36301 = n5171 | n36300 ;
  assign n36302 = n19520 ^ n10547 ^ 1'b0 ;
  assign n36303 = ~n14728 & n27702 ;
  assign n36304 = n15516 & n36303 ;
  assign n36305 = n6846 & ~n36304 ;
  assign n36306 = n6875 & n13251 ;
  assign n36307 = n36306 ^ n1334 ^ 1'b0 ;
  assign n36308 = n11330 & ~n22658 ;
  assign n36309 = ~n23039 & n36308 ;
  assign n36310 = n16796 | n34965 ;
  assign n36311 = ~n15712 & n22186 ;
  assign n36312 = n2452 & n36311 ;
  assign n36313 = n13137 ^ n10496 ^ 1'b0 ;
  assign n36314 = n36312 | n36313 ;
  assign n36315 = ~n17436 & n36314 ;
  assign n36316 = n3750 & ~n10142 ;
  assign n36317 = n36315 & n36316 ;
  assign n36318 = ( x22 & n5341 ) | ( x22 & ~n29327 ) | ( n5341 & ~n29327 ) ;
  assign n36319 = n21128 & n36318 ;
  assign n36320 = n36317 & n36319 ;
  assign n36321 = ~n5509 & n20075 ;
  assign n36322 = n36320 & n36321 ;
  assign n36323 = ( ~n10663 & n17076 ) | ( ~n10663 & n36164 ) | ( n17076 & n36164 ) ;
  assign n36324 = n3063 | n16086 ;
  assign n36325 = n36323 & ~n36324 ;
  assign n36326 = n36325 ^ n5223 ^ 1'b0 ;
  assign n36330 = x56 & ~n22184 ;
  assign n36331 = n36330 ^ n7382 ^ 1'b0 ;
  assign n36327 = n35157 ^ n3662 ^ n1258 ;
  assign n36328 = n6962 ^ n2782 ^ n1403 ;
  assign n36329 = n36327 | n36328 ;
  assign n36332 = n36331 ^ n36329 ^ n34512 ;
  assign n36333 = ( n2441 & n10558 ) | ( n2441 & ~n18646 ) | ( n10558 & ~n18646 ) ;
  assign n36334 = n27422 ^ n10910 ^ n6352 ;
  assign n36335 = n6040 | n22481 ;
  assign n36336 = n20647 | n36335 ;
  assign n36337 = n36336 ^ n31723 ^ 1'b0 ;
  assign n36338 = n7212 & n29025 ;
  assign n36340 = n20688 ^ n1561 ^ 1'b0 ;
  assign n36339 = ~n3636 & n4563 ;
  assign n36341 = n36340 ^ n36339 ^ n16898 ;
  assign n36342 = n14691 & n36341 ;
  assign n36343 = n30988 ^ n27895 ^ 1'b0 ;
  assign n36344 = ~n35558 & n36343 ;
  assign n36345 = n35310 ^ n7189 ^ 1'b0 ;
  assign n36346 = ( n13665 & ~n31759 ) | ( n13665 & n36345 ) | ( ~n31759 & n36345 ) ;
  assign n36347 = n28396 & ~n31053 ;
  assign n36348 = ~n6326 & n36347 ;
  assign n36349 = ( ~n1492 & n23625 ) | ( ~n1492 & n36348 ) | ( n23625 & n36348 ) ;
  assign n36351 = n25531 ^ n11152 ^ 1'b0 ;
  assign n36352 = n708 | n36351 ;
  assign n36353 = ( n5894 & n8025 ) | ( n5894 & ~n14084 ) | ( n8025 & ~n14084 ) ;
  assign n36354 = n36352 | n36353 ;
  assign n36350 = n659 & ~n4424 ;
  assign n36355 = n36354 ^ n36350 ^ 1'b0 ;
  assign n36356 = n2843 & ~n5095 ;
  assign n36357 = n36356 ^ n18092 ^ 1'b0 ;
  assign n36358 = n16687 & n29201 ;
  assign n36359 = n36358 ^ n21637 ^ 1'b0 ;
  assign n36360 = n16270 ^ n629 ^ 1'b0 ;
  assign n36361 = n19968 ^ n3969 ^ 1'b0 ;
  assign n36362 = n36361 ^ n26298 ^ n8683 ;
  assign n36363 = ( n8442 & n9149 ) | ( n8442 & ~n36362 ) | ( n9149 & ~n36362 ) ;
  assign n36364 = n34976 ^ n3967 ^ 1'b0 ;
  assign n36365 = n34341 ^ n15291 ^ 1'b0 ;
  assign n36366 = n25471 ^ n9338 ^ 1'b0 ;
  assign n36367 = n13152 ^ n8381 ^ 1'b0 ;
  assign n36368 = n6866 & n36367 ;
  assign n36369 = n36368 ^ n8940 ^ 1'b0 ;
  assign n36370 = ~n1378 & n23619 ;
  assign n36371 = ~n18465 & n36370 ;
  assign n36372 = n19698 | n36371 ;
  assign n36373 = n28191 & ~n36372 ;
  assign n36374 = ~n9707 & n13277 ;
  assign n36375 = n16929 ^ n16429 ^ 1'b0 ;
  assign n36376 = n36374 & n36375 ;
  assign n36377 = ( ~n4893 & n7010 ) | ( ~n4893 & n13930 ) | ( n7010 & n13930 ) ;
  assign n36380 = n14506 ^ n13981 ^ n10429 ;
  assign n36381 = ( n6781 & ~n23254 ) | ( n6781 & n36380 ) | ( ~n23254 & n36380 ) ;
  assign n36378 = n5752 | n11910 ;
  assign n36379 = n17553 | n36378 ;
  assign n36382 = n36381 ^ n36379 ^ n20546 ;
  assign n36383 = n10016 ^ n5349 ^ 1'b0 ;
  assign n36384 = ~n5325 & n23470 ;
  assign n36385 = n36384 ^ n33309 ^ 1'b0 ;
  assign n36386 = n36385 ^ n29837 ^ n623 ;
  assign n36387 = ( n15938 & ~n36383 ) | ( n15938 & n36386 ) | ( ~n36383 & n36386 ) ;
  assign n36388 = n1800 & n23400 ;
  assign n36389 = n18646 | n36388 ;
  assign n36390 = n36389 ^ n36089 ^ 1'b0 ;
  assign n36391 = n19558 ^ n14677 ^ 1'b0 ;
  assign n36392 = n15675 | n36391 ;
  assign n36393 = n8185 & ~n9024 ;
  assign n36394 = n32854 & ~n36393 ;
  assign n36395 = n4637 | n36394 ;
  assign n36396 = n36395 ^ n23620 ^ 1'b0 ;
  assign n36399 = n11480 ^ n6206 ^ 1'b0 ;
  assign n36400 = n36399 ^ n5044 ^ 1'b0 ;
  assign n36401 = n2171 | n28379 ;
  assign n36402 = n36400 & ~n36401 ;
  assign n36397 = n13521 | n34453 ;
  assign n36398 = n29266 & ~n36397 ;
  assign n36403 = n36402 ^ n36398 ^ n33897 ;
  assign n36406 = n4840 | n25710 ;
  assign n36404 = n1183 & n11682 ;
  assign n36405 = n36404 ^ n10888 ^ 1'b0 ;
  assign n36407 = n36406 ^ n36405 ^ 1'b0 ;
  assign n36408 = n34692 ^ n17963 ^ 1'b0 ;
  assign n36409 = n31170 & ~n36408 ;
  assign n36410 = n6896 ^ n4083 ^ 1'b0 ;
  assign n36411 = ~n2050 & n36410 ;
  assign n36412 = n11103 & n22554 ;
  assign n36413 = ~n36411 & n36412 ;
  assign n36414 = n36413 ^ n30419 ^ n5211 ;
  assign n36415 = n20998 | n36414 ;
  assign n36416 = n8124 | n36415 ;
  assign n36417 = n19977 ^ n1487 ^ 1'b0 ;
  assign n36418 = n29820 & n36417 ;
  assign n36419 = n30276 ^ n8144 ^ 1'b0 ;
  assign n36420 = n17304 | n33092 ;
  assign n36421 = n14489 ^ n8989 ^ 1'b0 ;
  assign n36422 = ( ~n2092 & n36420 ) | ( ~n2092 & n36421 ) | ( n36420 & n36421 ) ;
  assign n36423 = n19755 | n24982 ;
  assign n36424 = n36423 ^ n1050 ^ 1'b0 ;
  assign n36425 = n36424 ^ n4431 ^ n3905 ;
  assign n36426 = n20994 ^ n8668 ^ 1'b0 ;
  assign n36427 = n7799 & ~n12666 ;
  assign n36429 = ~n8430 & n29399 ;
  assign n36428 = n7388 | n12672 ;
  assign n36430 = n36429 ^ n36428 ^ 1'b0 ;
  assign n36431 = n5883 & ~n13884 ;
  assign n36432 = n36431 ^ n6788 ^ n2418 ;
  assign n36434 = n6154 & n6972 ;
  assign n36435 = n36434 ^ n24583 ^ 1'b0 ;
  assign n36433 = n3471 & n30630 ;
  assign n36436 = n36435 ^ n36433 ^ 1'b0 ;
  assign n36437 = n36436 ^ n28395 ^ n17585 ;
  assign n36438 = n23608 ^ n3622 ^ 1'b0 ;
  assign n36439 = n36438 ^ n17589 ^ n8929 ;
  assign n36440 = n3912 | n25552 ;
  assign n36441 = n36440 ^ n5712 ^ 1'b0 ;
  assign n36442 = n21327 ^ n20572 ^ 1'b0 ;
  assign n36443 = ~n3689 & n36442 ;
  assign n36444 = n36441 & n36443 ;
  assign n36447 = x104 & ~n11392 ;
  assign n36448 = n36447 ^ n15967 ^ 1'b0 ;
  assign n36449 = n36448 ^ n3307 ^ n282 ;
  assign n36445 = n33064 ^ x111 ^ 1'b0 ;
  assign n36446 = n5815 | n36445 ;
  assign n36450 = n36449 ^ n36446 ^ n2906 ;
  assign n36451 = n4767 & ~n11870 ;
  assign n36452 = n36451 ^ n23106 ^ n16967 ;
  assign n36453 = n2670 & n14533 ;
  assign n36454 = ~n20163 & n27540 ;
  assign n36455 = n13004 & n27256 ;
  assign n36456 = ~n24310 & n35293 ;
  assign n36457 = n5638 | n6424 ;
  assign n36458 = n36457 ^ n2113 ^ 1'b0 ;
  assign n36459 = ( n8079 & ~n22590 ) | ( n8079 & n36458 ) | ( ~n22590 & n36458 ) ;
  assign n36460 = n36459 ^ n11578 ^ 1'b0 ;
  assign n36461 = n23105 ^ n3461 ^ n1239 ;
  assign n36462 = ( n6765 & ~n28481 ) | ( n6765 & n36461 ) | ( ~n28481 & n36461 ) ;
  assign n36466 = n20022 ^ n12140 ^ n2130 ;
  assign n36463 = ( n7384 & n21153 ) | ( n7384 & n29408 ) | ( n21153 & n29408 ) ;
  assign n36464 = n2466 | n4061 ;
  assign n36465 = n36463 | n36464 ;
  assign n36467 = n36466 ^ n36465 ^ n29875 ;
  assign n36468 = n20354 ^ n5858 ^ n2406 ;
  assign n36469 = n12771 | n36468 ;
  assign n36470 = ( n11389 & ~n19849 ) | ( n11389 & n24573 ) | ( ~n19849 & n24573 ) ;
  assign n36471 = n8909 ^ n8697 ^ 1'b0 ;
  assign n36472 = ~n8622 & n36471 ;
  assign n36473 = n13146 & n36472 ;
  assign n36474 = ~n17572 & n36473 ;
  assign n36475 = n25183 | n36474 ;
  assign n36476 = n36475 ^ n34489 ^ 1'b0 ;
  assign n36477 = ( n5139 & n27099 ) | ( n5139 & ~n28681 ) | ( n27099 & ~n28681 ) ;
  assign n36478 = n36477 ^ n21711 ^ n6622 ;
  assign n36479 = n7361 & n36478 ;
  assign n36480 = n17817 ^ n11408 ^ 1'b0 ;
  assign n36481 = n9193 | n27530 ;
  assign n36482 = n1301 | n21592 ;
  assign n36483 = x93 & n11511 ;
  assign n36484 = n36483 ^ n13605 ^ 1'b0 ;
  assign n36485 = n11875 | n36484 ;
  assign n36486 = n36485 ^ n26509 ^ 1'b0 ;
  assign n36487 = ~n4579 & n18465 ;
  assign n36488 = n36487 ^ n3316 ^ 1'b0 ;
  assign n36489 = n36488 ^ n24079 ^ n4558 ;
  assign n36490 = n12939 & ~n17727 ;
  assign n36491 = n2821 & n36490 ;
  assign n36492 = n36491 ^ n20874 ^ n20323 ;
  assign n36493 = n27363 ^ n4468 ^ 1'b0 ;
  assign n36494 = ~n18256 & n27487 ;
  assign n36495 = ~n6929 & n36494 ;
  assign n36496 = ~n1350 & n2145 ;
  assign n36497 = n2379 & n36496 ;
  assign n36498 = n10401 | n24959 ;
  assign n36499 = ~n36497 & n36498 ;
  assign n36500 = n7848 & n36499 ;
  assign n36501 = ~n6839 & n7096 ;
  assign n36502 = n36501 ^ n15291 ^ 1'b0 ;
  assign n36503 = n2833 & ~n36502 ;
  assign n36504 = n24338 ^ n2830 ^ 1'b0 ;
  assign n36505 = n13488 | n36504 ;
  assign n36506 = n14749 ^ n8962 ^ 1'b0 ;
  assign n36507 = ~n26569 & n36506 ;
  assign n36508 = n34521 ^ n24782 ^ n8116 ;
  assign n36509 = ( n19342 & n36507 ) | ( n19342 & ~n36508 ) | ( n36507 & ~n36508 ) ;
  assign n36510 = n15652 ^ n5723 ^ 1'b0 ;
  assign n36511 = n2551 & n6143 ;
  assign n36512 = n513 & n36511 ;
  assign n36513 = n36512 ^ n28924 ^ n6894 ;
  assign n36514 = n1496 & ~n9045 ;
  assign n36515 = n16688 & ~n23012 ;
  assign n36516 = n36515 ^ n3707 ^ 1'b0 ;
  assign n36517 = n16869 ^ n9641 ^ n2012 ;
  assign n36518 = n3255 & ~n5003 ;
  assign n36519 = n13444 ^ n9037 ^ n3248 ;
  assign n36520 = n33938 & ~n36519 ;
  assign n36521 = n2323 | n6357 ;
  assign n36522 = n36521 ^ n15810 ^ 1'b0 ;
  assign n36523 = n5725 | n36522 ;
  assign n36524 = n36523 ^ n28293 ^ 1'b0 ;
  assign n36525 = n13990 & ~n36524 ;
  assign n36526 = n16408 & ~n25193 ;
  assign n36527 = ~x121 & n36526 ;
  assign n36528 = n11791 ^ n7923 ^ 1'b0 ;
  assign n36529 = n15734 & ~n36528 ;
  assign n36530 = ~n4799 & n11590 ;
  assign n36531 = ~n2585 & n36530 ;
  assign n36532 = n36531 ^ n17545 ^ n1387 ;
  assign n36533 = n14131 & n36532 ;
  assign n36534 = ~n20852 & n36533 ;
  assign n36535 = ( n15913 & ~n27980 ) | ( n15913 & n36534 ) | ( ~n27980 & n36534 ) ;
  assign n36536 = n18818 & n23096 ;
  assign n36537 = ( n14275 & n36331 ) | ( n14275 & ~n36536 ) | ( n36331 & ~n36536 ) ;
  assign n36538 = n3664 | n28728 ;
  assign n36539 = n36538 ^ n11546 ^ 1'b0 ;
  assign n36540 = n13693 & n36539 ;
  assign n36541 = n15648 ^ n4910 ^ 1'b0 ;
  assign n36542 = ( ~x158 & n4695 ) | ( ~x158 & n8437 ) | ( n4695 & n8437 ) ;
  assign n36543 = ( ~n15836 & n19157 ) | ( ~n15836 & n36542 ) | ( n19157 & n36542 ) ;
  assign n36544 = n8757 & ~n36543 ;
  assign n36545 = n36541 & n36544 ;
  assign n36546 = n490 | n20875 ;
  assign n36547 = n36546 ^ n675 ^ 1'b0 ;
  assign n36548 = ( n24371 & n29660 ) | ( n24371 & ~n36547 ) | ( n29660 & ~n36547 ) ;
  assign n36549 = n31953 ^ n27479 ^ n5601 ;
  assign n36550 = n12499 & n25866 ;
  assign n36551 = n6370 ^ n4781 ^ 1'b0 ;
  assign n36552 = n8368 & ~n36551 ;
  assign n36553 = n36552 ^ n26724 ^ n8673 ;
  assign n36554 = ~n36550 & n36553 ;
  assign n36555 = n29956 ^ n10608 ^ n5846 ;
  assign n36556 = ( n4645 & n10245 ) | ( n4645 & n14575 ) | ( n10245 & n14575 ) ;
  assign n36557 = n18075 | n36556 ;
  assign n36558 = n36557 ^ n15325 ^ n1862 ;
  assign n36559 = n9864 & ~n12392 ;
  assign n36560 = n21255 & n36559 ;
  assign n36561 = n36560 ^ n12207 ^ n1638 ;
  assign n36562 = ( n18840 & n24234 ) | ( n18840 & ~n32433 ) | ( n24234 & ~n32433 ) ;
  assign n36563 = n19254 | n23180 ;
  assign n36564 = ( n16130 & n36562 ) | ( n16130 & n36563 ) | ( n36562 & n36563 ) ;
  assign n36565 = n17390 ^ n16701 ^ 1'b0 ;
  assign n36566 = ~n15175 & n36565 ;
  assign n36567 = n5842 | n36566 ;
  assign n36568 = n7016 & n13360 ;
  assign n36569 = ( n15368 & n15820 ) | ( n15368 & n22469 ) | ( n15820 & n22469 ) ;
  assign n36570 = n36569 ^ n1759 ^ n1276 ;
  assign n36571 = ( ~n16058 & n23184 ) | ( ~n16058 & n26408 ) | ( n23184 & n26408 ) ;
  assign n36572 = ( n10457 & n13162 ) | ( n10457 & ~n29723 ) | ( n13162 & ~n29723 ) ;
  assign n36573 = n36572 ^ n31188 ^ n16172 ;
  assign n36574 = ~n31547 & n32158 ;
  assign n36575 = n1354 & n36574 ;
  assign n36576 = n36575 ^ n8774 ^ 1'b0 ;
  assign n36578 = ( n2878 & n5400 ) | ( n2878 & ~n6913 ) | ( n5400 & ~n6913 ) ;
  assign n36579 = n2517 & n36578 ;
  assign n36580 = n36579 ^ n3570 ^ 1'b0 ;
  assign n36577 = n17292 ^ n14919 ^ n11338 ;
  assign n36581 = n36580 ^ n36577 ^ 1'b0 ;
  assign n36582 = n9250 | n36581 ;
  assign n36583 = n36279 ^ n7086 ^ 1'b0 ;
  assign n36584 = ~n15013 & n22602 ;
  assign n36585 = ~n3810 & n32022 ;
  assign n36586 = ~n10059 & n36585 ;
  assign n36587 = ~n36585 & n36586 ;
  assign n36588 = n775 | n36587 ;
  assign n36589 = n775 & ~n36588 ;
  assign n36590 = n36589 ^ n24849 ^ 1'b0 ;
  assign n36591 = n14550 & ~n36590 ;
  assign n36592 = n36591 ^ n20720 ^ 1'b0 ;
  assign n36593 = n27579 ^ n15737 ^ 1'b0 ;
  assign n36594 = ( n13691 & n36592 ) | ( n13691 & ~n36593 ) | ( n36592 & ~n36593 ) ;
  assign n36595 = n8467 | n30754 ;
  assign n36596 = n36595 ^ n12230 ^ 1'b0 ;
  assign n36597 = ~n18953 & n36596 ;
  assign n36598 = n33024 & n36597 ;
  assign n36599 = ( n2806 & ~n20300 ) | ( n2806 & n36598 ) | ( ~n20300 & n36598 ) ;
  assign n36600 = n13227 ^ n2207 ^ 1'b0 ;
  assign n36601 = ( n7078 & ~n28614 ) | ( n7078 & n32806 ) | ( ~n28614 & n32806 ) ;
  assign n36602 = n25807 & n28214 ;
  assign n36603 = n30045 ^ n3950 ^ 1'b0 ;
  assign n36604 = ( n341 & n5362 ) | ( n341 & ~n7257 ) | ( n5362 & ~n7257 ) ;
  assign n36605 = n36604 ^ n14641 ^ n10465 ;
  assign n36606 = n36232 ^ n17920 ^ n9215 ;
  assign n36607 = n9551 & ~n36606 ;
  assign n36608 = ~n4390 & n14040 ;
  assign n36609 = n36608 ^ n12041 ^ 1'b0 ;
  assign n36610 = n21372 ^ n16592 ^ 1'b0 ;
  assign n36611 = n3771 & ~n36610 ;
  assign n36612 = n13959 ^ n6459 ^ n4101 ;
  assign n36613 = n3494 & n3736 ;
  assign n36614 = ( n6066 & n22575 ) | ( n6066 & ~n36613 ) | ( n22575 & ~n36613 ) ;
  assign n36615 = n36612 | n36614 ;
  assign n36616 = n5755 | n36615 ;
  assign n36617 = n36616 ^ n10162 ^ 1'b0 ;
  assign n36618 = n8054 & n9224 ;
  assign n36619 = n36618 ^ n4481 ^ 1'b0 ;
  assign n36620 = n36619 ^ n14395 ^ n3523 ;
  assign n36621 = n3496 & n13516 ;
  assign n36622 = n36621 ^ n16749 ^ 1'b0 ;
  assign n36623 = n36622 ^ n21859 ^ n3725 ;
  assign n36624 = n36623 ^ n22168 ^ n2841 ;
  assign n36625 = ~n7721 & n19600 ;
  assign n36626 = ~n15307 & n36625 ;
  assign n36627 = n36626 ^ n12219 ^ 1'b0 ;
  assign n36628 = ~n5302 & n36627 ;
  assign n36629 = n4754 | n36628 ;
  assign n36630 = n2123 & n23154 ;
  assign n36631 = ~n12981 & n19806 ;
  assign n36632 = n29428 & n36631 ;
  assign n36633 = n11611 & ~n14926 ;
  assign n36634 = n36633 ^ n13078 ^ 1'b0 ;
  assign n36635 = ( n13664 & ~n16977 ) | ( n13664 & n25190 ) | ( ~n16977 & n25190 ) ;
  assign n36636 = ~n9411 & n36635 ;
  assign n36638 = n26724 ^ n5458 ^ 1'b0 ;
  assign n36637 = n6609 ^ n3708 ^ 1'b0 ;
  assign n36639 = n36638 ^ n36637 ^ 1'b0 ;
  assign n36640 = n36639 ^ n14395 ^ 1'b0 ;
  assign n36644 = n15135 | n21004 ;
  assign n36641 = ( ~n3370 & n7761 ) | ( ~n3370 & n19424 ) | ( n7761 & n19424 ) ;
  assign n36642 = n36641 ^ n16600 ^ n9253 ;
  assign n36643 = n3472 & ~n36642 ;
  assign n36645 = n36644 ^ n36643 ^ n4479 ;
  assign n36646 = ( ~n642 & n5334 ) | ( ~n642 & n21459 ) | ( n5334 & n21459 ) ;
  assign n36647 = n21563 & n36646 ;
  assign n36648 = n30165 ^ n1870 ^ 1'b0 ;
  assign n36649 = n5965 | n36648 ;
  assign n36650 = n36647 | n36649 ;
  assign n36651 = n28294 ^ n18452 ^ 1'b0 ;
  assign n36652 = n15710 | n36651 ;
  assign n36653 = n22365 ^ n2227 ^ n1585 ;
  assign n36654 = n17361 ^ n5391 ^ 1'b0 ;
  assign n36655 = ~n7883 & n23333 ;
  assign n36656 = ( n14960 & n23944 ) | ( n14960 & ~n36655 ) | ( n23944 & ~n36655 ) ;
  assign n36657 = n7637 ^ n4696 ^ n2901 ;
  assign n36658 = n7899 | n36657 ;
  assign n36659 = n8834 | n36658 ;
  assign n36660 = n4654 | n18850 ;
  assign n36661 = n36659 | n36660 ;
  assign n36662 = n16488 | n19661 ;
  assign n36663 = n5183 | n36662 ;
  assign n36664 = n3417 & n33617 ;
  assign n36665 = n36664 ^ n31939 ^ 1'b0 ;
  assign n36666 = n21805 ^ n18917 ^ n801 ;
  assign n36667 = n23468 & ~n36666 ;
  assign n36668 = n24769 ^ n17191 ^ 1'b0 ;
  assign n36669 = ~n11410 & n36668 ;
  assign n36670 = ( n5448 & ~n13535 ) | ( n5448 & n27575 ) | ( ~n13535 & n27575 ) ;
  assign n36671 = ~n2045 & n18766 ;
  assign n36672 = ~n2845 & n22796 ;
  assign n36673 = ~n16710 & n36672 ;
  assign n36674 = n36673 ^ n36143 ^ n25674 ;
  assign n36675 = ( n5609 & ~n11698 ) | ( n5609 & n27015 ) | ( ~n11698 & n27015 ) ;
  assign n36676 = n9292 & ~n11976 ;
  assign n36677 = ~n36675 & n36676 ;
  assign n36678 = n36677 ^ n3878 ^ 1'b0 ;
  assign n36679 = n8329 ^ n6065 ^ 1'b0 ;
  assign n36680 = n20115 ^ n9880 ^ 1'b0 ;
  assign n36681 = n36679 & n36680 ;
  assign n36682 = n16701 | n18151 ;
  assign n36683 = n32194 ^ n560 ^ 1'b0 ;
  assign n36684 = ~n36682 & n36683 ;
  assign n36688 = n733 | n11917 ;
  assign n36689 = n36688 ^ n4147 ^ 1'b0 ;
  assign n36685 = n4948 & ~n5527 ;
  assign n36686 = ~n5324 & n36685 ;
  assign n36687 = n36686 ^ n8319 ^ n4616 ;
  assign n36690 = n36689 ^ n36687 ^ n7277 ;
  assign n36691 = ( ~n4836 & n6720 ) | ( ~n4836 & n19402 ) | ( n6720 & n19402 ) ;
  assign n36692 = n396 & ~n36691 ;
  assign n36693 = n20357 | n33493 ;
  assign n36694 = n17683 | n36693 ;
  assign n36695 = n36694 ^ n8060 ^ 1'b0 ;
  assign n36696 = n21908 ^ n2422 ^ n471 ;
  assign n36697 = n5593 & ~n20381 ;
  assign n36698 = n36696 & n36697 ;
  assign n36699 = ~n6596 & n19066 ;
  assign n36700 = n36699 ^ n7983 ^ 1'b0 ;
  assign n36701 = n17987 ^ n11985 ^ 1'b0 ;
  assign n36702 = n20895 ^ n19510 ^ n16516 ;
  assign n36703 = n11548 ^ n3716 ^ 1'b0 ;
  assign n36704 = n27727 ^ n23207 ^ 1'b0 ;
  assign n36705 = n23398 ^ n10060 ^ n8996 ;
  assign n36706 = n16642 & n32227 ;
  assign n36707 = ~n21460 & n36706 ;
  assign n36710 = n14422 ^ n3617 ^ 1'b0 ;
  assign n36708 = n20870 ^ n18142 ^ n11283 ;
  assign n36709 = n27537 & n36708 ;
  assign n36711 = n36710 ^ n36709 ^ n4852 ;
  assign n36712 = n13411 | n36711 ;
  assign n36713 = n3234 & ~n6624 ;
  assign n36714 = n36713 ^ n20566 ^ 1'b0 ;
  assign n36715 = ( n2677 & n6627 ) | ( n2677 & n36714 ) | ( n6627 & n36714 ) ;
  assign n36716 = ( ~n6944 & n32781 ) | ( ~n6944 & n36715 ) | ( n32781 & n36715 ) ;
  assign n36717 = ( n6643 & ~n12412 ) | ( n6643 & n19245 ) | ( ~n12412 & n19245 ) ;
  assign n36718 = n10230 & n22262 ;
  assign n36719 = n13488 ^ n12263 ^ n9714 ;
  assign n36720 = n2274 & ~n36719 ;
  assign n36721 = n4191 & ~n15954 ;
  assign n36722 = n35746 & ~n36721 ;
  assign n36723 = ~x198 & n36722 ;
  assign n36724 = n22308 | n36723 ;
  assign n36725 = n36724 ^ n29853 ^ 1'b0 ;
  assign n36726 = n36725 ^ n22264 ^ n14967 ;
  assign n36728 = n15519 ^ n5406 ^ 1'b0 ;
  assign n36729 = n36728 ^ n17256 ^ n12102 ;
  assign n36727 = n4501 | n18326 ;
  assign n36730 = n36729 ^ n36727 ^ 1'b0 ;
  assign n36731 = n6477 ^ n2570 ^ 1'b0 ;
  assign n36732 = n13984 & n36731 ;
  assign n36733 = ~n3862 & n9347 ;
  assign n36734 = n36733 ^ n2192 ^ 1'b0 ;
  assign n36736 = n7677 | n17064 ;
  assign n36737 = n26480 & n36736 ;
  assign n36735 = n7420 | n28699 ;
  assign n36738 = n36737 ^ n36735 ^ 1'b0 ;
  assign n36739 = ~n5643 & n36738 ;
  assign n36740 = n5355 & n36739 ;
  assign n36741 = n2310 & n11172 ;
  assign n36742 = n36740 & n36741 ;
  assign n36743 = n34293 ^ n17027 ^ 1'b0 ;
  assign n36744 = n9574 & ~n14048 ;
  assign n36745 = n17731 | n36744 ;
  assign n36748 = n7248 ^ n5797 ^ 1'b0 ;
  assign n36746 = n11121 | n25534 ;
  assign n36747 = n36746 ^ n24358 ^ 1'b0 ;
  assign n36749 = n36748 ^ n36747 ^ n31741 ;
  assign n36750 = ( ~n13865 & n28887 ) | ( ~n13865 & n34101 ) | ( n28887 & n34101 ) ;
  assign n36751 = n2443 | n7723 ;
  assign n36752 = n36751 ^ n1174 ^ 1'b0 ;
  assign n36753 = n36267 & n36752 ;
  assign n36754 = n7979 ^ n5863 ^ 1'b0 ;
  assign n36755 = n30218 & n36754 ;
  assign n36756 = n24375 & n25416 ;
  assign n36757 = ~n3410 & n36756 ;
  assign n36758 = n34174 ^ n18421 ^ 1'b0 ;
  assign n36759 = n2595 & n36758 ;
  assign n36760 = n2173 & n36759 ;
  assign n36761 = ~n3919 & n36760 ;
  assign n36762 = n17401 ^ n8213 ^ n4876 ;
  assign n36763 = n36762 ^ n36300 ^ 1'b0 ;
  assign n36764 = n9844 & ~n18589 ;
  assign n36765 = n23961 ^ n8475 ^ 1'b0 ;
  assign n36766 = n11317 & ~n36765 ;
  assign n36767 = ( ~n18481 & n36764 ) | ( ~n18481 & n36766 ) | ( n36764 & n36766 ) ;
  assign n36768 = n31723 ^ n1154 ^ 1'b0 ;
  assign n36769 = n1424 & ~n3023 ;
  assign n36770 = n36769 ^ n12285 ^ 1'b0 ;
  assign n36771 = n13290 & ~n14772 ;
  assign n36772 = n26125 ^ n2217 ^ 1'b0 ;
  assign n36773 = ~n35462 & n36772 ;
  assign n36774 = n2962 & n36773 ;
  assign n36775 = n36771 & n36774 ;
  assign n36776 = n27066 ^ n4904 ^ 1'b0 ;
  assign n36777 = n1677 ^ n1397 ^ 1'b0 ;
  assign n36778 = n3444 & ~n36777 ;
  assign n36779 = n3833 & ~n36778 ;
  assign n36780 = n36779 ^ n4072 ^ 1'b0 ;
  assign n36781 = n17618 ^ n13604 ^ 1'b0 ;
  assign n36782 = n2554 & n10376 ;
  assign n36783 = n36782 ^ n7051 ^ 1'b0 ;
  assign n36784 = n36781 | n36783 ;
  assign n36785 = ~n20742 & n27458 ;
  assign n36786 = ( n21201 & n28558 ) | ( n21201 & n36785 ) | ( n28558 & n36785 ) ;
  assign n36787 = n15184 ^ n2775 ^ 1'b0 ;
  assign n36788 = n36786 & ~n36787 ;
  assign n36789 = n8246 ^ n4433 ^ 1'b0 ;
  assign n36790 = n701 & n36789 ;
  assign n36791 = ( ~n3881 & n23417 ) | ( ~n3881 & n36790 ) | ( n23417 & n36790 ) ;
  assign n36792 = n3256 ^ n3050 ^ n826 ;
  assign n36795 = n10834 ^ n1515 ^ x182 ;
  assign n36796 = ~n13715 & n36795 ;
  assign n36793 = n14714 ^ n7591 ^ n3681 ;
  assign n36794 = n27643 | n36793 ;
  assign n36797 = n36796 ^ n36794 ^ n28967 ;
  assign n36798 = ~n10713 & n29180 ;
  assign n36799 = ~n24846 & n36798 ;
  assign n36800 = n36799 ^ n21998 ^ 1'b0 ;
  assign n36801 = ~n7257 & n32386 ;
  assign n36802 = n36470 ^ n2240 ^ 1'b0 ;
  assign n36803 = ~n36801 & n36802 ;
  assign n36805 = n11285 ^ n11149 ^ n3404 ;
  assign n36804 = ~n8412 & n12611 ;
  assign n36806 = n36805 ^ n36804 ^ 1'b0 ;
  assign n36807 = n13675 ^ n7794 ^ n1863 ;
  assign n36808 = ~n14279 & n17412 ;
  assign n36809 = ~n26354 & n36808 ;
  assign n36813 = n14669 ^ n288 ^ 1'b0 ;
  assign n36814 = n6183 & ~n36813 ;
  assign n36810 = n30800 ^ n26518 ^ 1'b0 ;
  assign n36811 = n932 & ~n36810 ;
  assign n36812 = n16568 & n36811 ;
  assign n36815 = n36814 ^ n36812 ^ 1'b0 ;
  assign n36816 = ( n21283 & ~n36809 ) | ( n21283 & n36815 ) | ( ~n36809 & n36815 ) ;
  assign n36817 = n2573 & ~n33727 ;
  assign n36818 = n36817 ^ n7632 ^ 1'b0 ;
  assign n36819 = n5111 | n36818 ;
  assign n36820 = n36819 ^ n11457 ^ 1'b0 ;
  assign n36821 = n36820 ^ n27372 ^ n2543 ;
  assign n36822 = n26097 ^ n5805 ^ 1'b0 ;
  assign n36823 = n36822 ^ n13949 ^ 1'b0 ;
  assign n36824 = n6415 | n27215 ;
  assign n36825 = n17140 ^ n2024 ^ 1'b0 ;
  assign n36826 = n36824 & ~n36825 ;
  assign n36827 = n14185 | n36826 ;
  assign n36828 = ~n2140 & n9103 ;
  assign n36829 = n17015 & n36828 ;
  assign n36830 = n16600 ^ n7457 ^ 1'b0 ;
  assign n36831 = n16429 & n36830 ;
  assign n36832 = ~n432 & n12202 ;
  assign n36833 = ~n3510 & n29867 ;
  assign n36834 = n36833 ^ n5398 ^ 1'b0 ;
  assign n36835 = ~n12420 & n14057 ;
  assign n36836 = ~n36834 & n36835 ;
  assign n36837 = ( n6310 & n36832 ) | ( n6310 & ~n36836 ) | ( n36832 & ~n36836 ) ;
  assign n36838 = n21769 & n36837 ;
  assign n36839 = n36838 ^ n21337 ^ 1'b0 ;
  assign n36840 = n24698 ^ n22560 ^ n820 ;
  assign n36841 = n36840 ^ n21951 ^ 1'b0 ;
  assign n36845 = n14923 ^ n9153 ^ 1'b0 ;
  assign n36844 = ( n4006 & n14704 ) | ( n4006 & n24314 ) | ( n14704 & n24314 ) ;
  assign n36846 = n36845 ^ n36844 ^ 1'b0 ;
  assign n36842 = n15715 ^ n15272 ^ 1'b0 ;
  assign n36843 = n11403 & n36842 ;
  assign n36847 = n36846 ^ n36843 ^ n1881 ;
  assign n36848 = n10100 & ~n19541 ;
  assign n36849 = ( n7957 & ~n16908 ) | ( n7957 & n36848 ) | ( ~n16908 & n36848 ) ;
  assign n36850 = n36849 ^ n28082 ^ n19993 ;
  assign n36851 = ( ~n15472 & n23265 ) | ( ~n15472 & n24577 ) | ( n23265 & n24577 ) ;
  assign n36852 = n14259 ^ n9527 ^ 1'b0 ;
  assign n36853 = ~n5736 & n36852 ;
  assign n36854 = ( ~n6606 & n36851 ) | ( ~n6606 & n36853 ) | ( n36851 & n36853 ) ;
  assign n36855 = n26317 ^ n10188 ^ 1'b0 ;
  assign n36856 = n14224 & ~n36855 ;
  assign n36857 = ~n4832 & n36856 ;
  assign n36858 = n18466 & n36857 ;
  assign n36859 = n21249 ^ n20226 ^ 1'b0 ;
  assign n36860 = ~n23674 & n36859 ;
  assign n36861 = n22527 & ~n24518 ;
  assign n36863 = ( n4692 & ~n5852 ) | ( n4692 & n30195 ) | ( ~n5852 & n30195 ) ;
  assign n36862 = ~n2205 & n4598 ;
  assign n36864 = n36863 ^ n36862 ^ 1'b0 ;
  assign n36865 = n11351 ^ n4707 ^ n3410 ;
  assign n36866 = n14201 & n36865 ;
  assign n36867 = n36866 ^ n32349 ^ 1'b0 ;
  assign n36868 = n36864 & n36867 ;
  assign n36869 = n3344 & ~n18302 ;
  assign n36870 = n36869 ^ n1343 ^ 1'b0 ;
  assign n36871 = n8492 | n36870 ;
  assign n36872 = n1770 | n36871 ;
  assign n36873 = n21304 | n36872 ;
  assign n36874 = n14364 ^ n14324 ^ 1'b0 ;
  assign n36875 = n12214 ^ n5863 ^ n4069 ;
  assign n36876 = n5043 & ~n9858 ;
  assign n36877 = n36876 ^ n17769 ^ 1'b0 ;
  assign n36878 = n10272 & n36877 ;
  assign n36879 = n36878 ^ n27024 ^ n13583 ;
  assign n36880 = n20167 | n34953 ;
  assign n36881 = n17381 & ~n32467 ;
  assign n36882 = n36881 ^ n31825 ^ 1'b0 ;
  assign n36883 = n13481 & n26760 ;
  assign n36884 = n36883 ^ n6901 ^ 1'b0 ;
  assign n36885 = ( n8757 & n9158 ) | ( n8757 & ~n36884 ) | ( n9158 & ~n36884 ) ;
  assign n36886 = n35800 ^ n30182 ^ n3498 ;
  assign n36887 = n34153 ^ n29000 ^ 1'b0 ;
  assign n36888 = ~n10106 & n36887 ;
  assign n36889 = n11148 ^ n5629 ^ 1'b0 ;
  assign n36890 = n36889 ^ n28070 ^ n8000 ;
  assign n36891 = n36890 ^ n14044 ^ n2865 ;
  assign n36892 = n18818 & ~n36891 ;
  assign n36893 = ~n36888 & n36892 ;
  assign n36894 = x211 & n5333 ;
  assign n36895 = ~n10172 & n36894 ;
  assign n36896 = n9277 | n36895 ;
  assign n36897 = n5448 & ~n36896 ;
  assign n36898 = n36897 ^ n25256 ^ 1'b0 ;
  assign n36899 = n31495 | n36898 ;
  assign n36900 = n3768 & ~n7246 ;
  assign n36901 = ~n34610 & n36900 ;
  assign n36902 = n21701 ^ n10663 ^ n7624 ;
  assign n36903 = n36902 ^ n25151 ^ n6221 ;
  assign n36904 = ( ~n4720 & n8548 ) | ( ~n4720 & n21180 ) | ( n8548 & n21180 ) ;
  assign n36905 = ( ~n2901 & n18626 ) | ( ~n2901 & n27359 ) | ( n18626 & n27359 ) ;
  assign n36906 = n36905 ^ n22928 ^ n15003 ;
  assign n36907 = n34844 ^ n25434 ^ n12981 ;
  assign n36908 = n15525 & n35173 ;
  assign n36909 = n33732 ^ n25591 ^ 1'b0 ;
  assign n36910 = n36908 & ~n36909 ;
  assign n36911 = n2831 & n10287 ;
  assign n36912 = n36911 ^ n6878 ^ 1'b0 ;
  assign n36913 = n5114 | n18390 ;
  assign n36914 = n34508 ^ n3690 ^ n1962 ;
  assign n36915 = n5090 | n6222 ;
  assign n36916 = n18594 | n25810 ;
  assign n36917 = n3199 | n36916 ;
  assign n36918 = n27999 ^ n25316 ^ 1'b0 ;
  assign n36919 = n18240 ^ n829 ^ 1'b0 ;
  assign n36920 = n21981 & ~n36919 ;
  assign n36921 = n36920 ^ n28639 ^ n1032 ;
  assign n36922 = ( x113 & ~n610 ) | ( x113 & n35473 ) | ( ~n610 & n35473 ) ;
  assign n36923 = n36922 ^ n24879 ^ n1604 ;
  assign n36924 = n18939 | n25404 ;
  assign n36925 = n36923 & ~n36924 ;
  assign n36926 = ~n14049 & n26137 ;
  assign n36927 = ~n36925 & n36926 ;
  assign n36928 = n6100 | n7362 ;
  assign n36929 = n36928 ^ n17108 ^ 1'b0 ;
  assign n36930 = n36929 ^ n31083 ^ 1'b0 ;
  assign n36931 = n18541 & ~n35899 ;
  assign n36932 = n10375 & n36931 ;
  assign n36933 = n36932 ^ n32366 ^ 1'b0 ;
  assign n36934 = n13158 ^ n8905 ^ 1'b0 ;
  assign n36935 = ( ~n20023 & n29905 ) | ( ~n20023 & n36934 ) | ( n29905 & n36934 ) ;
  assign n36936 = n6752 ^ n2859 ^ 1'b0 ;
  assign n36937 = n8769 | n28836 ;
  assign n36938 = n4600 | n33088 ;
  assign n36939 = n36938 ^ n23862 ^ 1'b0 ;
  assign n36940 = ~n24196 & n32350 ;
  assign n36941 = n36940 ^ n7837 ^ 1'b0 ;
  assign n36942 = n6634 & ~n15586 ;
  assign n36943 = n36941 & n36942 ;
  assign n36944 = n5014 ^ n1788 ^ 1'b0 ;
  assign n36945 = n30001 | n36944 ;
  assign n36946 = n17999 | n19157 ;
  assign n36947 = n2634 & n36946 ;
  assign n36948 = n20097 ^ n19713 ^ n6682 ;
  assign n36949 = n22410 ^ n8622 ^ 1'b0 ;
  assign n36950 = n2150 & n36949 ;
  assign n36951 = n18824 | n36950 ;
  assign n36952 = n17727 | n23617 ;
  assign n36953 = n10974 & ~n36952 ;
  assign n36954 = n36951 | n36953 ;
  assign n36955 = ( ~n5865 & n10212 ) | ( ~n5865 & n10405 ) | ( n10212 & n10405 ) ;
  assign n36956 = n13346 | n36955 ;
  assign n36957 = n18586 & ~n36956 ;
  assign n36958 = n3719 & n36957 ;
  assign n36960 = ( x56 & n8715 ) | ( x56 & n19889 ) | ( n8715 & n19889 ) ;
  assign n36959 = n4310 & ~n35520 ;
  assign n36961 = n36960 ^ n36959 ^ 1'b0 ;
  assign n36962 = ~n11019 & n16694 ;
  assign n36963 = ~n16827 & n36962 ;
  assign n36964 = n6875 ^ n5628 ^ n4190 ;
  assign n36965 = n1452 & n2321 ;
  assign n36966 = ~n36964 & n36965 ;
  assign n36967 = n11388 & ~n36966 ;
  assign n36968 = n36963 & n36967 ;
  assign n36969 = n756 | n8187 ;
  assign n36970 = n15724 & ~n36969 ;
  assign n36971 = n36970 ^ n8312 ^ n6828 ;
  assign n36972 = n6399 & n36971 ;
  assign n36973 = n8920 ^ n5777 ^ 1'b0 ;
  assign n36974 = ( ~n9897 & n25356 ) | ( ~n9897 & n36973 ) | ( n25356 & n36973 ) ;
  assign n36975 = n36974 ^ n35145 ^ n21929 ;
  assign n36976 = n22908 ^ n9732 ^ 1'b0 ;
  assign n36977 = ~n31729 & n36976 ;
  assign n36980 = n9945 ^ n4411 ^ 1'b0 ;
  assign n36981 = n1407 & n36980 ;
  assign n36982 = n12467 | n33779 ;
  assign n36983 = n36981 | n36982 ;
  assign n36979 = ( n9696 & ~n25776 ) | ( n9696 & n31201 ) | ( ~n25776 & n31201 ) ;
  assign n36984 = n36983 ^ n36979 ^ n7008 ;
  assign n36978 = n16519 & ~n34854 ;
  assign n36985 = n36984 ^ n36978 ^ 1'b0 ;
  assign n36989 = ( n2006 & n3793 ) | ( n2006 & n5042 ) | ( n3793 & n5042 ) ;
  assign n36987 = n24745 ^ n8940 ^ n818 ;
  assign n36986 = n15022 | n29373 ;
  assign n36988 = n36987 ^ n36986 ^ 1'b0 ;
  assign n36990 = n36989 ^ n36988 ^ n4034 ;
  assign n36991 = n23683 ^ n5199 ^ 1'b0 ;
  assign n36992 = n32753 ^ n32355 ^ n21822 ;
  assign n36993 = n36371 & ~n36992 ;
  assign n36997 = n21343 ^ n661 ^ 1'b0 ;
  assign n36998 = n20568 & n36997 ;
  assign n36994 = n3738 & ~n4164 ;
  assign n36995 = n36994 ^ n15334 ^ 1'b0 ;
  assign n36996 = n36995 ^ n18586 ^ 1'b0 ;
  assign n36999 = n36998 ^ n36996 ^ n3016 ;
  assign n37000 = ~n9740 & n18425 ;
  assign n37001 = n7622 ^ n2925 ^ 1'b0 ;
  assign n37002 = n37000 & ~n37001 ;
  assign n37003 = n33722 ^ n27356 ^ n18486 ;
  assign n37004 = n37003 ^ n21592 ^ 1'b0 ;
  assign n37005 = n2133 & ~n24454 ;
  assign n37006 = n25946 ^ n12419 ^ 1'b0 ;
  assign n37007 = n22907 & n37006 ;
  assign n37008 = ~n402 & n37007 ;
  assign n37009 = n9144 & ~n25016 ;
  assign n37010 = n16340 & ~n37009 ;
  assign n37011 = n7067 & n7485 ;
  assign n37012 = ( n2222 & n24530 ) | ( n2222 & n37011 ) | ( n24530 & n37011 ) ;
  assign n37013 = n25433 & n37012 ;
  assign n37014 = n20008 ^ n7209 ^ 1'b0 ;
  assign n37015 = ~n9608 & n37014 ;
  assign n37016 = ~n1966 & n18231 ;
  assign n37017 = n18057 | n37016 ;
  assign n37018 = n37015 | n37017 ;
  assign n37019 = n20357 & n24224 ;
  assign n37020 = n37019 ^ n23111 ^ 1'b0 ;
  assign n37021 = n21346 ^ n11965 ^ 1'b0 ;
  assign n37022 = n18675 ^ n4123 ^ 1'b0 ;
  assign n37023 = n20139 ^ n14605 ^ 1'b0 ;
  assign n37024 = ( n2769 & ~n37022 ) | ( n2769 & n37023 ) | ( ~n37022 & n37023 ) ;
  assign n37025 = n35302 ^ n9937 ^ n4298 ;
  assign n37030 = n10889 | n26638 ;
  assign n37031 = x10 | n37030 ;
  assign n37026 = n17493 & ~n22058 ;
  assign n37027 = ~n22413 & n37026 ;
  assign n37028 = n31732 | n37027 ;
  assign n37029 = n37028 ^ n29074 ^ 1'b0 ;
  assign n37032 = n37031 ^ n37029 ^ n12439 ;
  assign n37033 = n10281 ^ n9219 ^ 1'b0 ;
  assign n37034 = n11317 & n37033 ;
  assign n37035 = ~n11135 & n37034 ;
  assign n37041 = n12904 ^ n10045 ^ 1'b0 ;
  assign n37042 = n37041 ^ n19826 ^ 1'b0 ;
  assign n37036 = n663 | n3602 ;
  assign n37037 = n37036 ^ n3747 ^ 1'b0 ;
  assign n37038 = n23556 ^ n21346 ^ 1'b0 ;
  assign n37039 = ( ~n4397 & n37037 ) | ( ~n4397 & n37038 ) | ( n37037 & n37038 ) ;
  assign n37040 = n12959 & n37039 ;
  assign n37043 = n37042 ^ n37040 ^ 1'b0 ;
  assign n37044 = ~n8149 & n17126 ;
  assign n37045 = n37044 ^ n3816 ^ 1'b0 ;
  assign n37046 = x85 & ~n9803 ;
  assign n37047 = n37046 ^ n22961 ^ 1'b0 ;
  assign n37048 = n15134 ^ n857 ^ 1'b0 ;
  assign n37049 = n11841 ^ n10135 ^ 1'b0 ;
  assign n37050 = n37048 & ~n37049 ;
  assign n37051 = n11061 | n27725 ;
  assign n37052 = ( n26779 & n32257 ) | ( n26779 & n37051 ) | ( n32257 & n37051 ) ;
  assign n37053 = ( n1959 & n2068 ) | ( n1959 & ~n11775 ) | ( n2068 & ~n11775 ) ;
  assign n37054 = n671 & ~n13839 ;
  assign n37055 = n13839 & n37054 ;
  assign n37056 = ( n26017 & n37053 ) | ( n26017 & n37055 ) | ( n37053 & n37055 ) ;
  assign n37057 = n22262 ^ x63 ^ 1'b0 ;
  assign n37058 = n4203 & n32792 ;
  assign n37059 = ~n6732 & n37058 ;
  assign n37060 = n26944 & ~n37059 ;
  assign n37061 = n31638 & n37060 ;
  assign n37062 = n13174 ^ n6893 ^ 1'b0 ;
  assign n37063 = n37061 | n37062 ;
  assign n37064 = n854 & n18887 ;
  assign n37065 = n34747 ^ n18248 ^ n11141 ;
  assign n37066 = ~n9850 & n37065 ;
  assign n37067 = n19696 ^ n6395 ^ 1'b0 ;
  assign n37068 = n37067 ^ n2978 ^ 1'b0 ;
  assign n37069 = n10927 & n37068 ;
  assign n37075 = n24697 ^ x85 ^ 1'b0 ;
  assign n37070 = n23049 ^ n15394 ^ 1'b0 ;
  assign n37071 = n36271 | n37070 ;
  assign n37072 = n34337 ^ n27194 ^ 1'b0 ;
  assign n37073 = n32735 & ~n37072 ;
  assign n37074 = n37071 & n37073 ;
  assign n37076 = n37075 ^ n37074 ^ n7179 ;
  assign n37077 = n15601 ^ n14698 ^ 1'b0 ;
  assign n37078 = n37077 ^ n27362 ^ n14846 ;
  assign n37079 = n20691 ^ n8610 ^ 1'b0 ;
  assign n37080 = n1284 & n10031 ;
  assign n37081 = n37080 ^ n7111 ^ 1'b0 ;
  assign n37082 = n23947 & ~n37081 ;
  assign n37083 = ~n12077 & n37082 ;
  assign n37084 = n6205 | n23653 ;
  assign n37085 = n263 | n37084 ;
  assign n37086 = n13789 | n19765 ;
  assign n37087 = n37085 | n37086 ;
  assign n37088 = ~n2118 & n22912 ;
  assign n37089 = n21214 ^ n20713 ^ 1'b0 ;
  assign n37090 = n37089 ^ n19135 ^ n5793 ;
  assign n37091 = ( n3335 & ~n5211 ) | ( n3335 & n37090 ) | ( ~n5211 & n37090 ) ;
  assign n37092 = n24897 ^ n23703 ^ n19070 ;
  assign n37093 = n2663 & ~n10011 ;
  assign n37094 = n37093 ^ n4283 ^ 1'b0 ;
  assign n37095 = ( n5773 & n7395 ) | ( n5773 & n37094 ) | ( n7395 & n37094 ) ;
  assign n37096 = ~n12826 & n34459 ;
  assign n37097 = ~n11838 & n37096 ;
  assign n37098 = n14821 & n34540 ;
  assign n37099 = n37098 ^ n3452 ^ 1'b0 ;
  assign n37101 = n13785 ^ n12272 ^ 1'b0 ;
  assign n37100 = n12284 | n21999 ;
  assign n37102 = n37101 ^ n37100 ^ 1'b0 ;
  assign n37103 = n23335 ^ n4164 ^ 1'b0 ;
  assign n37104 = n37102 | n37103 ;
  assign n37105 = n9709 & ~n23844 ;
  assign n37106 = n16721 & ~n32904 ;
  assign n37107 = n37106 ^ n25867 ^ 1'b0 ;
  assign n37108 = n37107 ^ n20122 ^ 1'b0 ;
  assign n37109 = n7707 & n37108 ;
  assign n37110 = n37109 ^ n7317 ^ 1'b0 ;
  assign n37111 = n3941 & ~n37110 ;
  assign n37112 = n10546 & n29229 ;
  assign n37113 = n10822 & n37112 ;
  assign n37114 = n18308 ^ n832 ^ 1'b0 ;
  assign n37115 = ~n17898 & n37114 ;
  assign n37119 = n19542 ^ n2124 ^ 1'b0 ;
  assign n37120 = n10232 | n37119 ;
  assign n37116 = n3139 | n7974 ;
  assign n37117 = n10266 | n37116 ;
  assign n37118 = ~n18468 & n37117 ;
  assign n37121 = n37120 ^ n37118 ^ 1'b0 ;
  assign n37122 = n37121 ^ n33594 ^ n17875 ;
  assign n37123 = ( n4014 & n17756 ) | ( n4014 & n37122 ) | ( n17756 & n37122 ) ;
  assign n37124 = ( ~n37113 & n37115 ) | ( ~n37113 & n37123 ) | ( n37115 & n37123 ) ;
  assign n37125 = n33740 ^ n19634 ^ n9349 ;
  assign n37126 = n11733 & n16136 ;
  assign n37127 = n37126 ^ n33189 ^ 1'b0 ;
  assign n37129 = n29386 ^ n6015 ^ 1'b0 ;
  assign n37130 = n17903 & n37129 ;
  assign n37128 = n7798 & ~n19212 ;
  assign n37131 = n37130 ^ n37128 ^ 1'b0 ;
  assign n37132 = n514 | n12458 ;
  assign n37133 = ( ~n15487 & n22478 ) | ( ~n15487 & n37132 ) | ( n22478 & n37132 ) ;
  assign n37134 = n4746 & ~n37133 ;
  assign n37135 = ~n7586 & n17678 ;
  assign n37136 = n10611 ^ n5397 ^ 1'b0 ;
  assign n37137 = n710 & n27086 ;
  assign n37138 = n37137 ^ n4668 ^ 1'b0 ;
  assign n37139 = n17674 ^ n11511 ^ 1'b0 ;
  assign n37140 = n11761 & ~n37139 ;
  assign n37141 = n37140 ^ n6522 ^ 1'b0 ;
  assign n37142 = n37138 & ~n37141 ;
  assign n37143 = n18557 & n21453 ;
  assign n37144 = n16144 | n29766 ;
  assign n37145 = n37144 ^ n14698 ^ 1'b0 ;
  assign n37147 = n36225 ^ n10547 ^ 1'b0 ;
  assign n37148 = n15550 & n37147 ;
  assign n37146 = n9257 & n17976 ;
  assign n37149 = n37148 ^ n37146 ^ n24753 ;
  assign n37150 = ( n2769 & ~n23893 ) | ( n2769 & n30304 ) | ( ~n23893 & n30304 ) ;
  assign n37151 = n9415 | n12662 ;
  assign n37152 = n37151 ^ n3715 ^ 1'b0 ;
  assign n37153 = n22048 | n37152 ;
  assign n37154 = n37153 ^ x70 ^ 1'b0 ;
  assign n37155 = n37154 ^ n7676 ^ 1'b0 ;
  assign n37156 = n37155 ^ n640 ^ 1'b0 ;
  assign n37157 = n8646 ^ n3666 ^ 1'b0 ;
  assign n37158 = ~n14932 & n37157 ;
  assign n37159 = n14576 | n29717 ;
  assign n37160 = n1104 & n1605 ;
  assign n37161 = ~n1104 & n37160 ;
  assign n37162 = n9411 ^ n4898 ^ 1'b0 ;
  assign n37163 = n37161 | n37162 ;
  assign n37164 = n13320 | n37163 ;
  assign n37165 = ~n8328 & n11178 ;
  assign n37166 = n23584 ^ n11325 ^ 1'b0 ;
  assign n37167 = n37166 ^ n28860 ^ 1'b0 ;
  assign n37168 = n37165 & n37167 ;
  assign n37169 = n35118 ^ n29424 ^ 1'b0 ;
  assign n37170 = ~n10172 & n11140 ;
  assign n37171 = n15121 | n37170 ;
  assign n37172 = n3052 & ~n3739 ;
  assign n37173 = n9443 & n31733 ;
  assign n37174 = n37173 ^ n33224 ^ 1'b0 ;
  assign n37175 = n13559 | n37174 ;
  assign n37176 = ( n3938 & ~n8573 ) | ( n3938 & n11751 ) | ( ~n8573 & n11751 ) ;
  assign n37177 = n37176 ^ n7992 ^ 1'b0 ;
  assign n37178 = n17901 | n37177 ;
  assign n37179 = n37178 ^ n12587 ^ 1'b0 ;
  assign n37180 = n29636 ^ n15870 ^ 1'b0 ;
  assign n37181 = n37179 & ~n37180 ;
  assign n37182 = n9522 & n19480 ;
  assign n37183 = ( n18476 & ~n25529 ) | ( n18476 & n37182 ) | ( ~n25529 & n37182 ) ;
  assign n37184 = n24437 ^ n4361 ^ n837 ;
  assign n37185 = n8539 ^ n3604 ^ 1'b0 ;
  assign n37186 = ~n7805 & n37185 ;
  assign n37187 = n37186 ^ n8923 ^ 1'b0 ;
  assign n37188 = ~n13763 & n32503 ;
  assign n37189 = n23677 ^ n17847 ^ 1'b0 ;
  assign n37190 = n27897 ^ n5601 ^ 1'b0 ;
  assign n37191 = n36349 | n37190 ;
  assign n37192 = n11361 ^ n3546 ^ 1'b0 ;
  assign n37193 = n7291 & ~n11686 ;
  assign n37194 = n37193 ^ n17071 ^ 1'b0 ;
  assign n37195 = n1201 & ~n7598 ;
  assign n37196 = ~n1201 & n37195 ;
  assign n37197 = n14104 | n37196 ;
  assign n37198 = n26900 | n37197 ;
  assign n37199 = n7102 & n8143 ;
  assign n37200 = n27248 & n37199 ;
  assign n37201 = ~n17144 & n28113 ;
  assign n37202 = n37201 ^ n574 ^ 1'b0 ;
  assign n37203 = ( n9255 & n10243 ) | ( n9255 & ~n25618 ) | ( n10243 & ~n25618 ) ;
  assign n37204 = n36952 ^ n27349 ^ 1'b0 ;
  assign n37205 = ~n28407 & n36528 ;
  assign n37206 = ~n30691 & n37205 ;
  assign n37207 = n4045 & ~n6770 ;
  assign n37211 = ~n28542 & n30075 ;
  assign n37212 = n36491 | n37211 ;
  assign n37209 = ( n1174 & ~n2362 ) | ( n1174 & n12123 ) | ( ~n2362 & n12123 ) ;
  assign n37208 = n18201 & ~n25100 ;
  assign n37210 = n37209 ^ n37208 ^ 1'b0 ;
  assign n37213 = n37212 ^ n37210 ^ 1'b0 ;
  assign n37214 = n37207 & ~n37213 ;
  assign n37215 = n26561 ^ n7711 ^ 1'b0 ;
  assign n37216 = n14077 ^ n12807 ^ 1'b0 ;
  assign n37217 = n1635 & ~n16482 ;
  assign n37218 = n12828 & ~n37217 ;
  assign n37219 = ~n37216 & n37218 ;
  assign n37220 = n23649 ^ n1336 ^ 1'b0 ;
  assign n37221 = n30433 ^ n17271 ^ 1'b0 ;
  assign n37222 = n37220 & ~n37221 ;
  assign n37223 = n26777 ^ n13975 ^ 1'b0 ;
  assign n37224 = n9897 & ~n9955 ;
  assign n37225 = n6756 & n37224 ;
  assign n37226 = n37225 ^ n32497 ^ n5153 ;
  assign n37227 = n12841 | n17924 ;
  assign n37228 = n19242 ^ n3014 ^ 1'b0 ;
  assign n37229 = n14063 | n21904 ;
  assign n37230 = n37229 ^ n12214 ^ 1'b0 ;
  assign n37234 = n10579 ^ n5662 ^ 1'b0 ;
  assign n37235 = n37234 ^ n10755 ^ 1'b0 ;
  assign n37236 = x123 & n37235 ;
  assign n37237 = n37236 ^ n13659 ^ 1'b0 ;
  assign n37231 = n10368 ^ n9302 ^ n2821 ;
  assign n37232 = n10507 & ~n37231 ;
  assign n37233 = n37232 ^ n5940 ^ 1'b0 ;
  assign n37238 = n37237 ^ n37233 ^ 1'b0 ;
  assign n37239 = n36394 | n37238 ;
  assign n37240 = ~n11318 & n13409 ;
  assign n37241 = ~n3299 & n12298 ;
  assign n37242 = ( ~n6854 & n33543 ) | ( ~n6854 & n37241 ) | ( n33543 & n37241 ) ;
  assign n37243 = n1820 | n6821 ;
  assign n37244 = n1941 & n2305 ;
  assign n37245 = n37244 ^ n3641 ^ 1'b0 ;
  assign n37246 = ( ~n34488 & n37243 ) | ( ~n34488 & n37245 ) | ( n37243 & n37245 ) ;
  assign n37247 = ~n574 & n37246 ;
  assign n37254 = n2758 ^ n2588 ^ 1'b0 ;
  assign n37255 = n6613 & n37254 ;
  assign n37256 = n13756 & n37255 ;
  assign n37248 = n15818 ^ n8411 ^ 1'b0 ;
  assign n37249 = n37248 ^ n26622 ^ n2294 ;
  assign n37250 = n17234 ^ n1578 ^ 1'b0 ;
  assign n37251 = n32959 & n37250 ;
  assign n37252 = n37249 & n37251 ;
  assign n37253 = n11122 | n37252 ;
  assign n37257 = n37256 ^ n37253 ^ 1'b0 ;
  assign n37258 = n15831 & ~n21366 ;
  assign n37259 = n37258 ^ n33813 ^ 1'b0 ;
  assign n37260 = n3271 & ~n18208 ;
  assign n37261 = n4215 & n37260 ;
  assign n37262 = n729 & n3471 ;
  assign n37263 = n6854 ^ n5872 ^ 1'b0 ;
  assign n37264 = n9659 & n37263 ;
  assign n37265 = n37264 ^ n22697 ^ 1'b0 ;
  assign n37266 = ( n9776 & n31138 ) | ( n9776 & ~n34119 ) | ( n31138 & ~n34119 ) ;
  assign n37267 = n15881 ^ n3595 ^ n614 ;
  assign n37268 = n37267 ^ n11008 ^ 1'b0 ;
  assign n37269 = n8478 & ~n37268 ;
  assign n37270 = ( n1376 & n13499 ) | ( n1376 & n16174 ) | ( n13499 & n16174 ) ;
  assign n37271 = n32833 & n37270 ;
  assign n37272 = n9276 | n28272 ;
  assign n37273 = n37271 | n37272 ;
  assign n37274 = n29839 ^ n14686 ^ 1'b0 ;
  assign n37275 = n10474 & n37274 ;
  assign n37276 = n37275 ^ n24101 ^ n13114 ;
  assign n37277 = n1972 | n23565 ;
  assign n37278 = n29224 & ~n37277 ;
  assign n37279 = n20938 ^ n16958 ^ 1'b0 ;
  assign n37280 = ~n5257 & n37279 ;
  assign n37281 = n6341 ^ n5399 ^ 1'b0 ;
  assign n37286 = n10483 ^ n621 ^ 1'b0 ;
  assign n37287 = n37286 ^ n2539 ^ 1'b0 ;
  assign n37284 = n19706 ^ n5860 ^ n5344 ;
  assign n37285 = n37284 ^ n9736 ^ n8572 ;
  assign n37282 = n4296 & n7404 ;
  assign n37283 = n37282 ^ n22929 ^ 1'b0 ;
  assign n37288 = n37287 ^ n37285 ^ n37283 ;
  assign n37289 = n24432 | n24555 ;
  assign n37290 = ( ~n2016 & n36956 ) | ( ~n2016 & n37289 ) | ( n36956 & n37289 ) ;
  assign n37291 = ( n5114 & n17799 ) | ( n5114 & ~n20238 ) | ( n17799 & ~n20238 ) ;
  assign n37292 = n37290 | n37291 ;
  assign n37293 = n32954 | n37050 ;
  assign n37294 = n7273 & ~n12529 ;
  assign n37295 = ~n18854 & n37294 ;
  assign n37296 = n35534 & n37295 ;
  assign n37297 = n1907 & ~n6697 ;
  assign n37298 = ~n4405 & n37297 ;
  assign n37299 = n7218 & ~n15933 ;
  assign n37300 = n37299 ^ n36686 ^ 1'b0 ;
  assign n37301 = ~n9785 & n37300 ;
  assign n37302 = n37301 ^ n16249 ^ 1'b0 ;
  assign n37303 = n25135 ^ n19769 ^ 1'b0 ;
  assign n37304 = n22372 & n37303 ;
  assign n37305 = n6306 & n8713 ;
  assign n37306 = n37305 ^ n32787 ^ n16087 ;
  assign n37307 = n37306 ^ n27116 ^ 1'b0 ;
  assign n37310 = n26811 ^ n9765 ^ 1'b0 ;
  assign n37311 = ( n8182 & n10409 ) | ( n8182 & ~n37310 ) | ( n10409 & ~n37310 ) ;
  assign n37312 = n37311 ^ n19681 ^ 1'b0 ;
  assign n37308 = n1454 & n8363 ;
  assign n37309 = n37308 ^ n4931 ^ 1'b0 ;
  assign n37313 = n37312 ^ n37309 ^ n16883 ;
  assign n37314 = n6786 | n12703 ;
  assign n37315 = n31034 ^ n4013 ^ 1'b0 ;
  assign n37316 = n29135 & n30074 ;
  assign n37317 = ~n30749 & n37316 ;
  assign n37320 = n24790 | n25020 ;
  assign n37321 = n37320 ^ n1066 ^ 1'b0 ;
  assign n37318 = n8749 ^ n1963 ^ 1'b0 ;
  assign n37319 = n15832 | n37318 ;
  assign n37322 = n37321 ^ n37319 ^ 1'b0 ;
  assign n37325 = n519 & n15517 ;
  assign n37323 = n7880 | n33240 ;
  assign n37324 = n37323 ^ n13579 ^ 1'b0 ;
  assign n37326 = n37325 ^ n37324 ^ 1'b0 ;
  assign n37328 = ( n5294 & n15392 ) | ( n5294 & n28658 ) | ( n15392 & n28658 ) ;
  assign n37327 = ( x238 & n12622 ) | ( x238 & ~n13000 ) | ( n12622 & ~n13000 ) ;
  assign n37329 = n37328 ^ n37327 ^ n27273 ;
  assign n37330 = ~n17293 & n35212 ;
  assign n37331 = n27034 ^ n4434 ^ 1'b0 ;
  assign n37332 = n11968 | n37331 ;
  assign n37333 = n37332 ^ n13380 ^ 1'b0 ;
  assign n37334 = ~n4592 & n37333 ;
  assign n37335 = n14387 ^ n9176 ^ 1'b0 ;
  assign n37342 = n16006 & ~n20115 ;
  assign n37336 = n31047 ^ n18856 ^ 1'b0 ;
  assign n37337 = n8872 | n37336 ;
  assign n37338 = n13295 & ~n22404 ;
  assign n37339 = ~n21790 & n37338 ;
  assign n37340 = n5624 | n37339 ;
  assign n37341 = ( n16106 & n37337 ) | ( n16106 & n37340 ) | ( n37337 & n37340 ) ;
  assign n37343 = n37342 ^ n37341 ^ n2867 ;
  assign n37344 = n10526 ^ n1294 ^ 1'b0 ;
  assign n37345 = n36342 ^ n29715 ^ n20879 ;
  assign n37346 = ~n615 & n24792 ;
  assign n37347 = n37346 ^ n9586 ^ 1'b0 ;
  assign n37348 = ~n976 & n37347 ;
  assign n37349 = ( n14476 & n20718 ) | ( n14476 & ~n37348 ) | ( n20718 & ~n37348 ) ;
  assign n37350 = n13923 ^ n10412 ^ 1'b0 ;
  assign n37351 = n10228 ^ n1543 ^ 1'b0 ;
  assign n37352 = ( ~n552 & n26809 ) | ( ~n552 & n31135 ) | ( n26809 & n31135 ) ;
  assign n37353 = ~n37351 & n37352 ;
  assign n37354 = ~n18903 & n20597 ;
  assign n37355 = n8155 | n31749 ;
  assign n37356 = n11393 ^ n7452 ^ n3654 ;
  assign n37357 = ~n604 & n37356 ;
  assign n37358 = ~n34841 & n37357 ;
  assign n37359 = n7324 | n24608 ;
  assign n37360 = n28563 & ~n37359 ;
  assign n37361 = n24580 & ~n37360 ;
  assign n37362 = n25065 ^ n19709 ^ 1'b0 ;
  assign n37363 = n21594 ^ n290 ^ 1'b0 ;
  assign n37364 = n8143 & ~n37363 ;
  assign n37365 = ~n21654 & n26515 ;
  assign n37366 = n37365 ^ n27115 ^ 1'b0 ;
  assign n37367 = ~n15609 & n37366 ;
  assign n37368 = n37367 ^ n2547 ^ 1'b0 ;
  assign n37369 = ~n4662 & n23107 ;
  assign n37370 = ~n16919 & n37369 ;
  assign n37371 = n37370 ^ n327 ^ 1'b0 ;
  assign n37372 = n17292 | n37371 ;
  assign n37373 = n18931 & n20631 ;
  assign n37374 = n3641 & n37373 ;
  assign n37375 = ( n5476 & n10516 ) | ( n5476 & n37374 ) | ( n10516 & n37374 ) ;
  assign n37376 = n34159 ^ n18780 ^ n7876 ;
  assign n37377 = n28944 ^ n26365 ^ n18798 ;
  assign n37378 = ~n4943 & n13475 ;
  assign n37379 = ~n7466 & n37378 ;
  assign n37380 = n10432 ^ n7835 ^ 1'b0 ;
  assign n37381 = n18924 & ~n37380 ;
  assign n37382 = n30203 ^ n4836 ^ n1304 ;
  assign n37383 = n37381 & ~n37382 ;
  assign n37384 = n10135 | n17892 ;
  assign n37385 = n37384 ^ x104 ^ 1'b0 ;
  assign n37386 = n14938 ^ n968 ^ 1'b0 ;
  assign n37387 = n24114 | n37386 ;
  assign n37388 = n2094 & ~n8739 ;
  assign n37389 = n37388 ^ n8387 ^ 1'b0 ;
  assign n37390 = ( n23074 & n31611 ) | ( n23074 & ~n37389 ) | ( n31611 & ~n37389 ) ;
  assign n37391 = n37390 ^ n7299 ^ n5099 ;
  assign n37392 = n37391 ^ n15383 ^ 1'b0 ;
  assign n37393 = n4751 & n37392 ;
  assign n37394 = ( ~n21699 & n37387 ) | ( ~n21699 & n37393 ) | ( n37387 & n37393 ) ;
  assign n37395 = ( ~n9656 & n13569 ) | ( ~n9656 & n18418 ) | ( n13569 & n18418 ) ;
  assign n37396 = n36845 ^ n1460 ^ 1'b0 ;
  assign n37397 = n23792 ^ n9296 ^ n6098 ;
  assign n37398 = n375 & n37397 ;
  assign n37399 = n3630 & n37398 ;
  assign n37400 = n37399 ^ n3873 ^ 1'b0 ;
  assign n37401 = n9849 & n28230 ;
  assign n37402 = ~n25127 & n37401 ;
  assign n37403 = ( n13478 & n13494 ) | ( n13478 & ~n29694 ) | ( n13494 & ~n29694 ) ;
  assign n37404 = n37403 ^ n24322 ^ n6917 ;
  assign n37405 = n22798 ^ n11167 ^ 1'b0 ;
  assign n37406 = ~n18573 & n37405 ;
  assign n37407 = n37404 | n37406 ;
  assign n37408 = n35570 ^ n26944 ^ n20655 ;
  assign n37409 = x175 & n6030 ;
  assign n37410 = n14185 & n37409 ;
  assign n37411 = ~n11432 & n37410 ;
  assign n37412 = ( n6982 & n25359 ) | ( n6982 & ~n37411 ) | ( n25359 & ~n37411 ) ;
  assign n37413 = n2383 & ~n22172 ;
  assign n37414 = ~n9492 & n37413 ;
  assign n37415 = ( ~n11037 & n11426 ) | ( ~n11037 & n37414 ) | ( n11426 & n37414 ) ;
  assign n37416 = n36981 ^ n15060 ^ n9174 ;
  assign n37417 = n7830 & n20849 ;
  assign n37418 = n1727 & n37417 ;
  assign n37419 = ~n3408 & n15747 ;
  assign n37420 = n20929 ^ n2461 ^ 1'b0 ;
  assign n37421 = n37419 & n37420 ;
  assign n37422 = n8926 & n11020 ;
  assign n37423 = ~n9628 & n22146 ;
  assign n37424 = ~n1543 & n37423 ;
  assign n37425 = n37424 ^ n10696 ^ 1'b0 ;
  assign n37427 = n11728 ^ n5341 ^ 1'b0 ;
  assign n37426 = x24 & ~n12454 ;
  assign n37428 = n37427 ^ n37426 ^ 1'b0 ;
  assign n37429 = n28523 | n37428 ;
  assign n37430 = n27810 & ~n37429 ;
  assign n37431 = n2056 & ~n25169 ;
  assign n37432 = n37431 ^ n18721 ^ n9732 ;
  assign n37433 = x20 & ~n37432 ;
  assign n37434 = ~n36125 & n37433 ;
  assign n37435 = ~n7794 & n20040 ;
  assign n37436 = n37435 ^ n25164 ^ 1'b0 ;
  assign n37437 = n7798 | n37436 ;
  assign n37438 = n9927 ^ n1590 ^ n850 ;
  assign n37439 = n11273 | n37438 ;
  assign n37440 = ~n7465 & n37439 ;
  assign n37441 = n18745 & n37440 ;
  assign n37442 = n16126 & ~n34732 ;
  assign n37445 = ~n4216 & n7712 ;
  assign n37446 = ~n7712 & n37445 ;
  assign n37447 = n4426 & n6326 ;
  assign n37448 = ~n6326 & n37447 ;
  assign n37449 = n4097 & ~n37448 ;
  assign n37450 = n37448 & n37449 ;
  assign n37451 = n9533 | n19270 ;
  assign n37452 = n37451 ^ n11381 ^ 1'b0 ;
  assign n37453 = ( n37446 & ~n37450 ) | ( n37446 & n37452 ) | ( ~n37450 & n37452 ) ;
  assign n37443 = n10632 ^ n766 ^ 1'b0 ;
  assign n37444 = n37443 ^ n28312 ^ n2921 ;
  assign n37454 = n37453 ^ n37444 ^ n24819 ;
  assign n37456 = n5682 | n8243 ;
  assign n37457 = n37456 ^ n16370 ^ 1'b0 ;
  assign n37455 = n6613 & ~n27575 ;
  assign n37458 = n37457 ^ n37455 ^ 1'b0 ;
  assign n37459 = n13830 ^ n6236 ^ 1'b0 ;
  assign n37460 = ~n6628 & n37459 ;
  assign n37461 = n37460 ^ n545 ^ 1'b0 ;
  assign n37462 = n21978 ^ n8755 ^ 1'b0 ;
  assign n37463 = ~n18984 & n37462 ;
  assign n37464 = n14679 & n37463 ;
  assign n37465 = n1635 | n5412 ;
  assign n37466 = n1709 | n37465 ;
  assign n37467 = n37466 ^ n23096 ^ n931 ;
  assign n37468 = n21661 ^ n10543 ^ 1'b0 ;
  assign n37469 = ~n28217 & n37468 ;
  assign n37470 = ~n7026 & n15073 ;
  assign n37471 = ~n37469 & n37470 ;
  assign n37472 = ( n703 & n6804 ) | ( n703 & ~n37471 ) | ( n6804 & ~n37471 ) ;
  assign n37473 = n8341 & ~n8375 ;
  assign n37474 = n14715 & n37473 ;
  assign n37475 = ( ~n5679 & n37472 ) | ( ~n5679 & n37474 ) | ( n37472 & n37474 ) ;
  assign n37476 = ~n678 & n2125 ;
  assign n37477 = n37476 ^ n23199 ^ n17806 ;
  assign n37478 = n13680 ^ n12174 ^ 1'b0 ;
  assign n37479 = n2178 ^ n1886 ^ 1'b0 ;
  assign n37480 = n16969 & n22661 ;
  assign n37481 = n1955 & n37480 ;
  assign n37482 = n10921 ^ n1390 ^ 1'b0 ;
  assign n37483 = n37255 & n37482 ;
  assign n37484 = n14246 & n37483 ;
  assign n37485 = n16032 ^ n7549 ^ 1'b0 ;
  assign n37486 = n17115 & ~n18443 ;
  assign n37487 = n3774 & n37486 ;
  assign n37488 = ( n5854 & ~n23506 ) | ( n5854 & n37487 ) | ( ~n23506 & n37487 ) ;
  assign n37489 = n29817 ^ n9153 ^ 1'b0 ;
  assign n37490 = n19421 | n37489 ;
  assign n37491 = n30571 ^ n5470 ^ 1'b0 ;
  assign n37492 = n16732 & ~n34724 ;
  assign n37493 = n37492 ^ n22883 ^ 1'b0 ;
  assign n37494 = ( n37490 & ~n37491 ) | ( n37490 & n37493 ) | ( ~n37491 & n37493 ) ;
  assign n37495 = ( ~n986 & n7906 ) | ( ~n986 & n13375 ) | ( n7906 & n13375 ) ;
  assign n37496 = n28925 | n37495 ;
  assign n37497 = n37496 ^ n25380 ^ 1'b0 ;
  assign n37498 = ~n29916 & n37497 ;
  assign n37499 = n11976 ^ n8228 ^ 1'b0 ;
  assign n37500 = ~n12784 & n37499 ;
  assign n37501 = n17046 ^ n9381 ^ 1'b0 ;
  assign n37502 = n37500 & n37501 ;
  assign n37503 = n16362 & n23561 ;
  assign n37504 = n37503 ^ n12696 ^ 1'b0 ;
  assign n37505 = n24904 | n37504 ;
  assign n37506 = ~n16500 & n37505 ;
  assign n37507 = ~n37502 & n37506 ;
  assign n37508 = n17422 & n34479 ;
  assign n37509 = n37508 ^ n951 ^ 1'b0 ;
  assign n37511 = n7303 & n11240 ;
  assign n37510 = n15031 & n22560 ;
  assign n37512 = n37511 ^ n37510 ^ 1'b0 ;
  assign n37513 = n17507 ^ n10632 ^ 1'b0 ;
  assign n37514 = n8442 & n37513 ;
  assign n37515 = n26133 & n37514 ;
  assign n37516 = n35076 ^ n8049 ^ 1'b0 ;
  assign n37517 = n14324 & n37516 ;
  assign n37518 = ( n6030 & n24248 ) | ( n6030 & ~n37517 ) | ( n24248 & ~n37517 ) ;
  assign n37519 = ( n24811 & n37515 ) | ( n24811 & ~n37518 ) | ( n37515 & ~n37518 ) ;
  assign n37520 = n11418 ^ n9762 ^ n3767 ;
  assign n37521 = ~n26984 & n37520 ;
  assign n37522 = n9542 ^ x66 ^ 1'b0 ;
  assign n37523 = n4953 ^ n2275 ^ 1'b0 ;
  assign n37524 = n16765 & n37523 ;
  assign n37525 = ~n37522 & n37524 ;
  assign n37526 = n18291 & n37525 ;
  assign n37527 = n31972 ^ n24232 ^ 1'b0 ;
  assign n37528 = n1653 | n3210 ;
  assign n37529 = ( ~n26027 & n32757 ) | ( ~n26027 & n37528 ) | ( n32757 & n37528 ) ;
  assign n37530 = n37529 ^ n11449 ^ 1'b0 ;
  assign n37531 = n24114 | n37530 ;
  assign n37537 = ~n23481 & n24666 ;
  assign n37533 = n4966 | n25231 ;
  assign n37534 = n37533 ^ n7996 ^ 1'b0 ;
  assign n37535 = n37534 ^ n5355 ^ 1'b0 ;
  assign n37536 = n9709 | n37535 ;
  assign n37532 = n4153 & n9393 ;
  assign n37538 = n37537 ^ n37536 ^ n37532 ;
  assign n37539 = n23355 ^ n20174 ^ n9426 ;
  assign n37540 = n37539 ^ n7284 ^ 1'b0 ;
  assign n37542 = n2970 & n24949 ;
  assign n37543 = ~n11072 & n37542 ;
  assign n37541 = n6062 ^ n1944 ^ 1'b0 ;
  assign n37544 = n37543 ^ n37541 ^ 1'b0 ;
  assign n37545 = n26019 ^ n20556 ^ 1'b0 ;
  assign n37546 = ( n15901 & n25424 ) | ( n15901 & n33734 ) | ( n25424 & n33734 ) ;
  assign n37547 = n8834 ^ n2575 ^ 1'b0 ;
  assign n37548 = ~n468 & n3614 ;
  assign n37549 = n6921 & n37548 ;
  assign n37550 = n37549 ^ n32332 ^ 1'b0 ;
  assign n37551 = n16139 & ~n37550 ;
  assign n37552 = n5298 ^ n2005 ^ 1'b0 ;
  assign n37553 = n28789 | n37552 ;
  assign n37554 = n536 & ~n37553 ;
  assign n37555 = n37554 ^ n11664 ^ 1'b0 ;
  assign n37556 = n27136 | n37555 ;
  assign n37557 = n19761 | n37556 ;
  assign n37558 = n19300 ^ x251 ^ 1'b0 ;
  assign n37559 = ( n1024 & n12528 ) | ( n1024 & n34890 ) | ( n12528 & n34890 ) ;
  assign n37560 = n12575 & n23310 ;
  assign n37561 = n37560 ^ n21949 ^ 1'b0 ;
  assign n37562 = n37561 ^ n15123 ^ n6337 ;
  assign n37563 = ( ~n18487 & n37559 ) | ( ~n18487 & n37562 ) | ( n37559 & n37562 ) ;
  assign n37564 = n29078 ^ n26623 ^ 1'b0 ;
  assign n37565 = n9219 & ~n37564 ;
  assign n37566 = n37565 ^ n34298 ^ 1'b0 ;
  assign n37567 = n6697 | n13321 ;
  assign n37568 = n37567 ^ n26298 ^ n18304 ;
  assign n37569 = n37568 ^ n26969 ^ n13664 ;
  assign n37570 = ( n5672 & n24609 ) | ( n5672 & n37541 ) | ( n24609 & n37541 ) ;
  assign n37571 = ~n1427 & n19204 ;
  assign n37572 = n6260 ^ n5518 ^ 1'b0 ;
  assign n37573 = n3099 & n37572 ;
  assign n37574 = n27921 ^ n1285 ^ n994 ;
  assign n37575 = ( n13662 & n15347 ) | ( n13662 & ~n32767 ) | ( n15347 & ~n32767 ) ;
  assign n37576 = n1074 & ~n2895 ;
  assign n37577 = n37576 ^ n7715 ^ 1'b0 ;
  assign n37578 = n8370 | n29795 ;
  assign n37579 = n37577 & ~n37578 ;
  assign n37580 = n2917 ^ n2677 ^ 1'b0 ;
  assign n37581 = ~n14422 & n37580 ;
  assign n37582 = n13886 & ~n24159 ;
  assign n37583 = n5929 | n23467 ;
  assign n37584 = n25597 ^ n18174 ^ 1'b0 ;
  assign n37585 = ( n11913 & n32758 ) | ( n11913 & ~n37584 ) | ( n32758 & ~n37584 ) ;
  assign n37586 = n20888 ^ n18362 ^ 1'b0 ;
  assign n37587 = n37586 ^ n7034 ^ n5188 ;
  assign n37588 = n37587 ^ n37429 ^ 1'b0 ;
  assign n37589 = n29168 ^ n23264 ^ 1'b0 ;
  assign n37590 = ( ~n312 & n1489 ) | ( ~n312 & n37589 ) | ( n1489 & n37589 ) ;
  assign n37591 = n10113 | n37590 ;
  assign n37592 = n32732 ^ n24347 ^ 1'b0 ;
  assign n37593 = ~n10711 & n37592 ;
  assign n37594 = n31552 & n37593 ;
  assign n37595 = n37594 ^ n7740 ^ 1'b0 ;
  assign n37597 = n9627 | n17381 ;
  assign n37596 = ~n9092 & n11172 ;
  assign n37598 = n37597 ^ n37596 ^ 1'b0 ;
  assign n37599 = n20414 | n30278 ;
  assign n37600 = n36089 ^ n9078 ^ n2138 ;
  assign n37601 = n9075 | n37600 ;
  assign n37602 = n37601 ^ n27449 ^ 1'b0 ;
  assign n37603 = n16825 ^ n7189 ^ 1'b0 ;
  assign n37604 = n1388 & ~n9002 ;
  assign n37605 = ( n24241 & n37603 ) | ( n24241 & n37604 ) | ( n37603 & n37604 ) ;
  assign n37610 = ( ~n1082 & n12541 ) | ( ~n1082 & n32658 ) | ( n12541 & n32658 ) ;
  assign n37606 = n18395 ^ n10581 ^ 1'b0 ;
  assign n37607 = n8537 | n37606 ;
  assign n37608 = n20157 ^ n19118 ^ 1'b0 ;
  assign n37609 = ( ~n6602 & n37607 ) | ( ~n6602 & n37608 ) | ( n37607 & n37608 ) ;
  assign n37611 = n37610 ^ n37609 ^ n25003 ;
  assign n37612 = n20235 & n21259 ;
  assign n37613 = n13706 & n37612 ;
  assign n37614 = n20747 ^ n5869 ^ 1'b0 ;
  assign n37615 = ~n37613 & n37614 ;
  assign n37616 = ~n24651 & n26605 ;
  assign n37617 = ~n4280 & n37616 ;
  assign n37618 = n33559 | n34935 ;
  assign n37619 = n13930 ^ n12477 ^ 1'b0 ;
  assign n37620 = n23807 | n37619 ;
  assign n37621 = n37620 ^ n16041 ^ 1'b0 ;
  assign n37622 = n31486 ^ n986 ^ 1'b0 ;
  assign n37628 = n25294 ^ n24651 ^ n5094 ;
  assign n37629 = n5118 & ~n37628 ;
  assign n37630 = ~n12450 & n37629 ;
  assign n37625 = n5377 ^ n516 ^ 1'b0 ;
  assign n37626 = ~n6392 & n37625 ;
  assign n37623 = ( n3607 & n10854 ) | ( n3607 & ~n36870 ) | ( n10854 & ~n36870 ) ;
  assign n37624 = ( ~n2005 & n22320 ) | ( ~n2005 & n37623 ) | ( n22320 & n37623 ) ;
  assign n37627 = n37626 ^ n37624 ^ 1'b0 ;
  assign n37631 = n37630 ^ n37627 ^ n17795 ;
  assign n37632 = ~n6335 & n7232 ;
  assign n37633 = n37632 ^ n30748 ^ n22147 ;
  assign n37634 = n34500 ^ n3341 ^ 1'b0 ;
  assign n37635 = n14829 & ~n28991 ;
  assign n37636 = n9924 & n34319 ;
  assign n37637 = n37636 ^ n28693 ^ 1'b0 ;
  assign n37638 = ~n8119 & n15820 ;
  assign n37639 = n4863 & n37638 ;
  assign n37640 = n37639 ^ n18061 ^ n12292 ;
  assign n37641 = n17626 & n30743 ;
  assign n37642 = n29029 & n37641 ;
  assign n37643 = ( n17599 & n37640 ) | ( n17599 & n37642 ) | ( n37640 & n37642 ) ;
  assign n37644 = n37620 ^ n29788 ^ n25084 ;
  assign n37645 = n7087 & ~n9062 ;
  assign n37646 = ~n27333 & n37645 ;
  assign n37647 = ( ~n11358 & n18143 ) | ( ~n11358 & n37646 ) | ( n18143 & n37646 ) ;
  assign n37649 = n12331 ^ n6431 ^ n1598 ;
  assign n37648 = n13109 & ~n17773 ;
  assign n37650 = n37649 ^ n37648 ^ 1'b0 ;
  assign n37651 = n13716 ^ n3166 ^ 1'b0 ;
  assign n37652 = x24 | n37651 ;
  assign n37653 = ~n14135 & n31071 ;
  assign n37654 = ~n37652 & n37653 ;
  assign n37655 = n22835 ^ n18405 ^ 1'b0 ;
  assign n37656 = n24587 ^ n17078 ^ 1'b0 ;
  assign n37657 = n22949 & n37656 ;
  assign n37658 = n37657 ^ n11229 ^ 1'b0 ;
  assign n37659 = n6869 | n29123 ;
  assign n37660 = n3361 & ~n15586 ;
  assign n37661 = n13869 & ~n26179 ;
  assign n37662 = ~n37660 & n37661 ;
  assign n37663 = n3705 ^ n2601 ^ 1'b0 ;
  assign n37664 = ~n20659 & n37663 ;
  assign n37665 = n8942 & n18589 ;
  assign n37666 = n11596 & n37665 ;
  assign n37667 = n828 & ~n37666 ;
  assign n37668 = ~n16827 & n37667 ;
  assign n37669 = n27601 | n37668 ;
  assign n37670 = n21192 ^ n8250 ^ 1'b0 ;
  assign n37671 = ( ~n2160 & n14170 ) | ( ~n2160 & n35932 ) | ( n14170 & n35932 ) ;
  assign n37672 = n9736 & n27099 ;
  assign n37673 = ~n15311 & n37672 ;
  assign n37674 = n7932 & ~n37673 ;
  assign n37675 = n14259 | n27602 ;
  assign n37676 = n37675 ^ n25901 ^ 1'b0 ;
  assign n37677 = ~n9219 & n15590 ;
  assign n37678 = n1066 & n37677 ;
  assign n37679 = ~n1693 & n17742 ;
  assign n37680 = n7847 & n37679 ;
  assign n37681 = n37680 ^ n15206 ^ 1'b0 ;
  assign n37682 = n22165 ^ n17078 ^ 1'b0 ;
  assign n37683 = ~n25579 & n37682 ;
  assign n37684 = n33614 ^ n10805 ^ 1'b0 ;
  assign n37685 = n6105 & n37684 ;
  assign n37686 = ( ~n20168 & n28556 ) | ( ~n20168 & n37685 ) | ( n28556 & n37685 ) ;
  assign n37687 = n32215 ^ n6093 ^ 1'b0 ;
  assign n37688 = n13708 ^ n12594 ^ n4407 ;
  assign n37689 = n22099 ^ n10208 ^ 1'b0 ;
  assign n37690 = ~n37688 & n37689 ;
  assign n37691 = n24633 | n25838 ;
  assign n37692 = n16761 & n18656 ;
  assign n37693 = n37692 ^ n22381 ^ 1'b0 ;
  assign n37694 = ~n14992 & n37693 ;
  assign n37695 = n37694 ^ n11044 ^ 1'b0 ;
  assign n37696 = n37695 ^ n26872 ^ n11371 ;
  assign n37697 = ( n7739 & n18687 ) | ( n7739 & ~n19261 ) | ( n18687 & ~n19261 ) ;
  assign n37698 = ~n9707 & n17277 ;
  assign n37699 = ~n4987 & n37698 ;
  assign n37700 = n11491 & ~n37699 ;
  assign n37701 = ~n9038 & n37700 ;
  assign n37702 = n37701 ^ n12284 ^ n10932 ;
  assign n37703 = ~n1289 & n2606 ;
  assign n37704 = n32923 ^ n475 ^ 1'b0 ;
  assign n37705 = x182 & n37704 ;
  assign n37706 = n24389 ^ x47 ^ 1'b0 ;
  assign n37707 = ~n7080 & n37706 ;
  assign n37708 = n24776 ^ n19156 ^ 1'b0 ;
  assign n37709 = n7388 | n12079 ;
  assign n37710 = n5793 & n6147 ;
  assign n37711 = n11324 & n25770 ;
  assign n37712 = n10805 & ~n24068 ;
  assign n37713 = n33771 | n37712 ;
  assign n37714 = n1234 | n1525 ;
  assign n37715 = ( ~n17013 & n24154 ) | ( ~n17013 & n37714 ) | ( n24154 & n37714 ) ;
  assign n37721 = n4963 & ~n22289 ;
  assign n37722 = n37721 ^ n20810 ^ 1'b0 ;
  assign n37716 = n22929 ^ n18864 ^ 1'b0 ;
  assign n37717 = ( n3255 & n22736 ) | ( n3255 & n24241 ) | ( n22736 & n24241 ) ;
  assign n37718 = n37717 ^ n26934 ^ n8207 ;
  assign n37719 = n37718 ^ n22837 ^ 1'b0 ;
  assign n37720 = n37716 & n37719 ;
  assign n37723 = n37722 ^ n37720 ^ 1'b0 ;
  assign n37724 = n12587 ^ n4817 ^ 1'b0 ;
  assign n37725 = n17174 ^ n12823 ^ 1'b0 ;
  assign n37726 = n17412 ^ n5428 ^ 1'b0 ;
  assign n37727 = n2740 & ~n20316 ;
  assign n37728 = n21879 | n37727 ;
  assign n37729 = n37728 ^ n25534 ^ 1'b0 ;
  assign n37730 = n37729 ^ n20257 ^ 1'b0 ;
  assign n37731 = n37726 | n37730 ;
  assign n37732 = ~n3638 & n27058 ;
  assign n37733 = n31349 & n37732 ;
  assign n37734 = ( ~n8429 & n14953 ) | ( ~n8429 & n25986 ) | ( n14953 & n25986 ) ;
  assign n37735 = n5215 & n37734 ;
  assign n37736 = n21525 ^ n14100 ^ 1'b0 ;
  assign n37737 = n10498 ^ n5069 ^ 1'b0 ;
  assign n37738 = n4398 & ~n37737 ;
  assign n37739 = n31388 ^ n8364 ^ 1'b0 ;
  assign n37740 = ~n15843 & n37739 ;
  assign n37741 = n37740 ^ n6056 ^ 1'b0 ;
  assign n37742 = n26513 ^ n5404 ^ 1'b0 ;
  assign n37743 = n37485 & ~n37742 ;
  assign n37748 = ( n22897 & n35543 ) | ( n22897 & n36897 ) | ( n35543 & n36897 ) ;
  assign n37749 = n1486 & ~n37748 ;
  assign n37750 = ~n11841 & n37749 ;
  assign n37751 = n37750 ^ n6253 ^ 1'b0 ;
  assign n37744 = ~n7245 & n30427 ;
  assign n37745 = n27372 ^ n356 ^ 1'b0 ;
  assign n37746 = n37744 & n37745 ;
  assign n37747 = ~n25314 & n37746 ;
  assign n37752 = n37751 ^ n37747 ^ 1'b0 ;
  assign n37753 = n9010 & n30820 ;
  assign n37754 = n37753 ^ n19772 ^ 1'b0 ;
  assign n37755 = n19479 & ~n21941 ;
  assign n37756 = n24086 ^ n13689 ^ n13255 ;
  assign n37758 = n21160 | n29584 ;
  assign n37757 = n4485 ^ n3512 ^ 1'b0 ;
  assign n37759 = n37758 ^ n37757 ^ n8446 ;
  assign n37760 = ( ~n1257 & n8473 ) | ( ~n1257 & n19936 ) | ( n8473 & n19936 ) ;
  assign n37761 = n12270 & ~n20219 ;
  assign n37762 = n37761 ^ n30405 ^ n16641 ;
  assign n37763 = n37762 ^ n13949 ^ 1'b0 ;
  assign n37764 = n7099 & ~n37763 ;
  assign n37765 = n3980 | n37764 ;
  assign n37766 = ~n11472 & n15237 ;
  assign n37767 = n8748 & n37766 ;
  assign n37768 = n37767 ^ n12051 ^ 1'b0 ;
  assign n37769 = n25974 | n37768 ;
  assign n37770 = n7857 ^ n4973 ^ 1'b0 ;
  assign n37771 = n7437 | n37770 ;
  assign n37772 = n24953 ^ n9492 ^ n4934 ;
  assign n37773 = ( n21774 & n30318 ) | ( n21774 & ~n37772 ) | ( n30318 & ~n37772 ) ;
  assign n37774 = ( n3483 & n5060 ) | ( n3483 & ~n5623 ) | ( n5060 & ~n5623 ) ;
  assign n37775 = n26129 ^ n471 ^ 1'b0 ;
  assign n37776 = ~n25640 & n37775 ;
  assign n37777 = n37776 ^ n24843 ^ n11432 ;
  assign n37778 = ~n11380 & n19573 ;
  assign n37779 = ~n23956 & n37778 ;
  assign n37780 = n33053 ^ n10621 ^ 1'b0 ;
  assign n37781 = ~n464 & n37780 ;
  assign n37782 = n29748 ^ n15826 ^ n1596 ;
  assign n37783 = n37782 ^ n2262 ^ 1'b0 ;
  assign n37784 = n37781 | n37783 ;
  assign n37785 = n9540 ^ n1447 ^ 1'b0 ;
  assign n37786 = ~n2822 & n37785 ;
  assign n37787 = n24846 ^ n24536 ^ 1'b0 ;
  assign n37788 = ~n1890 & n37787 ;
  assign n37790 = ~n6569 & n7814 ;
  assign n37789 = x115 & n9443 ;
  assign n37791 = n37790 ^ n37789 ^ 1'b0 ;
  assign n37792 = n4844 & n37170 ;
  assign n37794 = n15800 ^ n12898 ^ n3404 ;
  assign n37793 = n37553 ^ n4980 ^ 1'b0 ;
  assign n37795 = n37794 ^ n37793 ^ n8110 ;
  assign n37796 = ( n3376 & n14104 ) | ( n3376 & n37795 ) | ( n14104 & n37795 ) ;
  assign n37797 = ~n18181 & n36550 ;
  assign n37798 = ~n37796 & n37797 ;
  assign n37799 = n37798 ^ n31364 ^ n12183 ;
  assign n37800 = n14999 | n18813 ;
  assign n37801 = n37800 ^ n18654 ^ 1'b0 ;
  assign n37802 = n37801 ^ n22527 ^ n17504 ;
  assign n37803 = n30387 ^ n24429 ^ 1'b0 ;
  assign n37804 = n28539 ^ n1023 ^ 1'b0 ;
  assign n37807 = ~n5956 & n16186 ;
  assign n37805 = ( n24375 & n32753 ) | ( n24375 & n33742 ) | ( n32753 & n33742 ) ;
  assign n37806 = n4147 | n37805 ;
  assign n37808 = n37807 ^ n37806 ^ 1'b0 ;
  assign n37809 = n18364 ^ n12896 ^ n1298 ;
  assign n37810 = n15429 & n37809 ;
  assign n37811 = n37810 ^ n24190 ^ 1'b0 ;
  assign n37812 = n32723 & n37811 ;
  assign n37813 = n20045 ^ n3182 ^ 1'b0 ;
  assign n37821 = n33444 ^ n7391 ^ 1'b0 ;
  assign n37814 = n28602 ^ n1731 ^ 1'b0 ;
  assign n37815 = n2595 & ~n37814 ;
  assign n37816 = n33325 ^ n31948 ^ n24184 ;
  assign n37817 = n37816 ^ n3800 ^ 1'b0 ;
  assign n37818 = n37815 & n37817 ;
  assign n37819 = ~n10092 & n29321 ;
  assign n37820 = ~n37818 & n37819 ;
  assign n37822 = n37821 ^ n37820 ^ n17121 ;
  assign n37825 = n37534 ^ n8922 ^ n4533 ;
  assign n37823 = ~n1687 & n30838 ;
  assign n37824 = n37823 ^ n3813 ^ 1'b0 ;
  assign n37826 = n37825 ^ n37824 ^ 1'b0 ;
  assign n37827 = ~n729 & n6656 ;
  assign n37828 = ~n3691 & n37827 ;
  assign n37829 = ( n9772 & n13704 ) | ( n9772 & ~n28702 ) | ( n13704 & ~n28702 ) ;
  assign n37830 = n37828 | n37829 ;
  assign n37831 = n31881 ^ n4006 ^ 1'b0 ;
  assign n37832 = n37830 | n37831 ;
  assign n37833 = n17214 | n17674 ;
  assign n37834 = n35939 | n37833 ;
  assign n37835 = n10801 ^ n7284 ^ 1'b0 ;
  assign n37837 = n21277 ^ n11582 ^ n6496 ;
  assign n37836 = n15632 & ~n17153 ;
  assign n37838 = n37837 ^ n37836 ^ n24390 ;
  assign n37839 = n27435 | n32572 ;
  assign n37840 = n37839 ^ n16287 ^ 1'b0 ;
  assign n37841 = ( n9363 & ~n14553 ) | ( n9363 & n37840 ) | ( ~n14553 & n37840 ) ;
  assign n37843 = n11328 ^ n5725 ^ 1'b0 ;
  assign n37842 = n7002 & n15798 ;
  assign n37844 = n37843 ^ n37842 ^ 1'b0 ;
  assign n37845 = n4553 ^ n4214 ^ 1'b0 ;
  assign n37846 = n29518 & n37845 ;
  assign n37847 = ~n11052 & n25221 ;
  assign n37848 = ~n18972 & n37847 ;
  assign n37849 = ( ~n8690 & n13072 ) | ( ~n8690 & n31583 ) | ( n13072 & n31583 ) ;
  assign n37850 = n36140 ^ n1701 ^ n968 ;
  assign n37851 = n37850 ^ n29002 ^ n24546 ;
  assign n37852 = n6913 ^ n2005 ^ n1276 ;
  assign n37853 = n37852 ^ n20473 ^ 1'b0 ;
  assign n37854 = n26540 & ~n37853 ;
  assign n37855 = n14914 ^ n9088 ^ 1'b0 ;
  assign n37856 = ~n30143 & n37855 ;
  assign n37857 = ~n28036 & n37856 ;
  assign n37858 = ~n29307 & n37857 ;
  assign n37859 = n1478 | n27749 ;
  assign n37860 = n1979 & ~n13542 ;
  assign n37861 = n37860 ^ n18941 ^ 1'b0 ;
  assign n37862 = ( n24502 & n25383 ) | ( n24502 & ~n37861 ) | ( n25383 & ~n37861 ) ;
  assign n37863 = ~n19135 & n37862 ;
  assign n37864 = n18915 ^ n798 ^ 1'b0 ;
  assign n37865 = ( n10495 & ~n19823 ) | ( n10495 & n37864 ) | ( ~n19823 & n37864 ) ;
  assign n37866 = n21140 ^ n17833 ^ 1'b0 ;
  assign n37870 = n3590 ^ n943 ^ 1'b0 ;
  assign n37867 = n29241 ^ n24312 ^ 1'b0 ;
  assign n37868 = n14960 & ~n37867 ;
  assign n37869 = n37868 ^ n5134 ^ n3723 ;
  assign n37871 = n37870 ^ n37869 ^ n32009 ;
  assign n37875 = n1978 | n4719 ;
  assign n37876 = n22629 & ~n37875 ;
  assign n37873 = ~n8697 & n18073 ;
  assign n37874 = ~x153 & n37873 ;
  assign n37872 = n14318 | n23173 ;
  assign n37877 = n37876 ^ n37874 ^ n37872 ;
  assign n37878 = ~x250 & n6400 ;
  assign n37879 = n37878 ^ n29898 ^ 1'b0 ;
  assign n37884 = n16155 ^ n3919 ^ 1'b0 ;
  assign n37885 = n22822 | n37884 ;
  assign n37880 = n8729 & ~n18853 ;
  assign n37881 = n7252 & n37880 ;
  assign n37882 = ~n16471 & n27465 ;
  assign n37883 = ~n37881 & n37882 ;
  assign n37886 = n37885 ^ n37883 ^ 1'b0 ;
  assign n37887 = n3604 | n34199 ;
  assign n37888 = n22380 ^ n11448 ^ 1'b0 ;
  assign n37889 = n11729 & ~n37888 ;
  assign n37890 = n37889 ^ n9874 ^ 1'b0 ;
  assign n37891 = x137 & ~n27519 ;
  assign n37892 = ( ~n15646 & n21637 ) | ( ~n15646 & n37891 ) | ( n21637 & n37891 ) ;
  assign n37893 = n10426 ^ x139 ^ 1'b0 ;
  assign n37894 = ( ~n6246 & n13979 ) | ( ~n6246 & n37893 ) | ( n13979 & n37893 ) ;
  assign n37895 = ~x120 & n27622 ;
  assign n37896 = ~n15778 & n37895 ;
  assign n37897 = ( n19943 & ~n33408 ) | ( n19943 & n37896 ) | ( ~n33408 & n37896 ) ;
  assign n37898 = n7378 | n7496 ;
  assign n37899 = n36837 ^ n23123 ^ 1'b0 ;
  assign n37900 = n26306 ^ x37 ^ 1'b0 ;
  assign n37901 = n8593 | n37900 ;
  assign n37902 = n4979 | n37901 ;
  assign n37903 = ~n5484 & n11592 ;
  assign n37904 = n4435 & ~n37903 ;
  assign n37905 = n37904 ^ n12575 ^ n9197 ;
  assign n37906 = ~n31675 & n37905 ;
  assign n37907 = ~n2092 & n20315 ;
  assign n37908 = n37907 ^ n550 ^ 1'b0 ;
  assign n37909 = n3605 | n15933 ;
  assign n37910 = n7282 & ~n37909 ;
  assign n37911 = ( n32407 & ~n37908 ) | ( n32407 & n37910 ) | ( ~n37908 & n37910 ) ;
  assign n37912 = n20442 & ~n21984 ;
  assign n37913 = n23808 ^ n9901 ^ n1416 ;
  assign n37914 = ( ~n3984 & n25164 ) | ( ~n3984 & n37913 ) | ( n25164 & n37913 ) ;
  assign n37915 = n5646 & ~n30387 ;
  assign n37916 = ~n34136 & n37915 ;
  assign n37917 = ( n37912 & ~n37914 ) | ( n37912 & n37916 ) | ( ~n37914 & n37916 ) ;
  assign n37918 = n9831 & n32320 ;
  assign n37919 = n738 & n15621 ;
  assign n37920 = n37919 ^ n12417 ^ n11634 ;
  assign n37921 = n22190 | n37920 ;
  assign n37922 = n4434 & n26372 ;
  assign n37923 = n37921 & n37922 ;
  assign n37924 = n36999 ^ n8300 ^ 1'b0 ;
  assign n37929 = ~n5964 & n22990 ;
  assign n37927 = ~x82 & n5239 ;
  assign n37925 = ~n539 & n15590 ;
  assign n37926 = n8060 & n37925 ;
  assign n37928 = n37927 ^ n37926 ^ n31587 ;
  assign n37930 = n37929 ^ n37928 ^ 1'b0 ;
  assign n37931 = n11318 ^ n9803 ^ x9 ;
  assign n37932 = n37931 ^ n30310 ^ n3151 ;
  assign n37933 = n13320 & ~n37932 ;
  assign n37934 = n3740 | n37933 ;
  assign n37935 = n31418 ^ n7976 ^ n1176 ;
  assign n37936 = n18425 & ~n37935 ;
  assign n37937 = n37936 ^ n27310 ^ 1'b0 ;
  assign n37938 = n11804 & n33069 ;
  assign n37939 = n4063 & n37938 ;
  assign n37940 = n18592 | n29040 ;
  assign n37941 = n12664 ^ n12298 ^ n7745 ;
  assign n37942 = n27366 ^ n25394 ^ n24126 ;
  assign n37943 = ~n4361 & n8895 ;
  assign n37944 = n37942 & n37943 ;
  assign n37945 = n37944 ^ n15517 ^ 1'b0 ;
  assign n37946 = n36782 ^ n9376 ^ 1'b0 ;
  assign n37947 = ~n11747 & n37946 ;
  assign n37948 = n6982 | n16100 ;
  assign n37949 = n14151 | n37948 ;
  assign n37950 = n20990 ^ n6326 ^ 1'b0 ;
  assign n37951 = n6866 & ~n37950 ;
  assign n37952 = n12046 ^ n5270 ^ x160 ;
  assign n37953 = n37952 ^ n13774 ^ 1'b0 ;
  assign n37954 = n9341 ^ n5889 ^ 1'b0 ;
  assign n37955 = n1661 | n21286 ;
  assign n37956 = ( ~n15791 & n17727 ) | ( ~n15791 & n34136 ) | ( n17727 & n34136 ) ;
  assign n37957 = n37639 | n37956 ;
  assign n37958 = n37955 & ~n37957 ;
  assign n37959 = n7881 ^ n6568 ^ 1'b0 ;
  assign n37960 = n37959 ^ n20292 ^ n5097 ;
  assign n37961 = n37960 ^ n14423 ^ 1'b0 ;
  assign n37962 = n25739 & n37961 ;
  assign n37963 = n20250 ^ n13050 ^ n10629 ;
  assign n37964 = n37963 ^ n19785 ^ 1'b0 ;
  assign n37965 = n15031 & ~n37964 ;
  assign n37966 = n17579 ^ n9885 ^ 1'b0 ;
  assign n37967 = n24504 ^ n13414 ^ 1'b0 ;
  assign n37970 = n10092 ^ n4343 ^ 1'b0 ;
  assign n37971 = n17277 & n37970 ;
  assign n37969 = n21850 ^ n5433 ^ 1'b0 ;
  assign n37968 = n11714 ^ n2691 ^ n337 ;
  assign n37972 = n37971 ^ n37969 ^ n37968 ;
  assign n37973 = n12291 ^ n9889 ^ 1'b0 ;
  assign n37974 = n9244 ^ n4417 ^ 1'b0 ;
  assign n37975 = ( n3182 & ~n13494 ) | ( n3182 & n37974 ) | ( ~n13494 & n37974 ) ;
  assign n37976 = n37975 ^ n22297 ^ 1'b0 ;
  assign n37977 = n37973 | n37976 ;
  assign n37978 = n7466 & ~n37977 ;
  assign n37979 = n37978 ^ n654 ^ 1'b0 ;
  assign n37980 = ~n20208 & n28075 ;
  assign n37981 = n21926 | n35444 ;
  assign n37982 = n20714 | n37981 ;
  assign n37983 = n27238 ^ n23468 ^ n3674 ;
  assign n37984 = ~n18814 & n21168 ;
  assign n37985 = n37983 & n37984 ;
  assign n37986 = n37985 ^ n10168 ^ 1'b0 ;
  assign n37987 = ~n17562 & n37986 ;
  assign n37988 = n36061 ^ n6613 ^ 1'b0 ;
  assign n37989 = n37988 ^ n13678 ^ 1'b0 ;
  assign n37990 = ( n10121 & ~n11572 ) | ( n10121 & n32254 ) | ( ~n11572 & n32254 ) ;
  assign n37991 = n15023 & n32422 ;
  assign n37992 = n37991 ^ n8447 ^ 1'b0 ;
  assign n37996 = n11084 | n25063 ;
  assign n37997 = n15039 | n37996 ;
  assign n37998 = n23000 & n37997 ;
  assign n37999 = n19985 & n37998 ;
  assign n38000 = ( n16017 & n23774 ) | ( n16017 & ~n37999 ) | ( n23774 & ~n37999 ) ;
  assign n37993 = n9044 & ~n11066 ;
  assign n37994 = n37993 ^ n27169 ^ 1'b0 ;
  assign n37995 = ~n29956 & n37994 ;
  assign n38001 = n38000 ^ n37995 ^ 1'b0 ;
  assign n38002 = n31842 ^ n23185 ^ 1'b0 ;
  assign n38003 = n10670 | n14634 ;
  assign n38004 = n38003 ^ n11852 ^ n10566 ;
  assign n38005 = n24981 ^ n18604 ^ n13581 ;
  assign n38006 = n20538 ^ n18734 ^ 1'b0 ;
  assign n38007 = n7864 & n38006 ;
  assign n38008 = n38007 ^ n34836 ^ n5973 ;
  assign n38009 = n15706 | n32476 ;
  assign n38010 = n22856 ^ n16528 ^ 1'b0 ;
  assign n38011 = ~n38009 & n38010 ;
  assign n38012 = n10024 & n38011 ;
  assign n38013 = ( ~n13061 & n36709 ) | ( ~n13061 & n38012 ) | ( n36709 & n38012 ) ;
  assign n38014 = n6647 ^ n6184 ^ 1'b0 ;
  assign n38015 = n3073 ^ n2731 ^ 1'b0 ;
  assign n38016 = n38014 & ~n38015 ;
  assign n38017 = n30968 ^ n18161 ^ 1'b0 ;
  assign n38018 = n13698 & ~n17450 ;
  assign n38020 = n23153 ^ n20703 ^ 1'b0 ;
  assign n38019 = n25424 & ~n27089 ;
  assign n38021 = n38020 ^ n38019 ^ 1'b0 ;
  assign n38022 = n11058 & ~n33296 ;
  assign n38023 = ~n11072 & n38022 ;
  assign n38024 = n38023 ^ n14363 ^ 1'b0 ;
  assign n38025 = n8999 ^ n8603 ^ 1'b0 ;
  assign n38026 = n29849 ^ n13881 ^ 1'b0 ;
  assign n38027 = n36309 ^ n5424 ^ 1'b0 ;
  assign n38028 = n38026 & n38027 ;
  assign n38029 = ( n1733 & n9062 ) | ( n1733 & ~n16746 ) | ( n9062 & ~n16746 ) ;
  assign n38030 = n13319 ^ n4386 ^ 1'b0 ;
  assign n38031 = ~n38029 & n38030 ;
  assign n38032 = n38031 ^ n1671 ^ x225 ;
  assign n38033 = n9538 | n38032 ;
  assign n38034 = n10250 ^ n4836 ^ 1'b0 ;
  assign n38035 = n38033 & ~n38034 ;
  assign n38036 = ~n955 & n26495 ;
  assign n38037 = ~n21231 & n38036 ;
  assign n38038 = n38037 ^ n5976 ^ 1'b0 ;
  assign n38039 = n6907 & ~n38038 ;
  assign n38040 = n37660 ^ n21426 ^ 1'b0 ;
  assign n38041 = n16081 & n21275 ;
  assign n38042 = n38041 ^ n8357 ^ 1'b0 ;
  assign n38043 = n38042 ^ n4326 ^ 1'b0 ;
  assign n38044 = n18405 | n38043 ;
  assign n38045 = ~n11148 & n36563 ;
  assign n38049 = n2647 | n11803 ;
  assign n38050 = n6720 & ~n38049 ;
  assign n38047 = n29534 ^ n24815 ^ n16874 ;
  assign n38048 = n6351 & ~n38047 ;
  assign n38051 = n38050 ^ n38048 ^ 1'b0 ;
  assign n38046 = n2891 & ~n27287 ;
  assign n38052 = n38051 ^ n38046 ^ 1'b0 ;
  assign n38053 = ( n7111 & n9264 ) | ( n7111 & n26641 ) | ( n9264 & n26641 ) ;
  assign n38054 = n36917 ^ n20802 ^ 1'b0 ;
  assign n38055 = n29125 & n30529 ;
  assign n38056 = n21622 ^ n13368 ^ 1'b0 ;
  assign n38057 = ( ~n3678 & n17953 ) | ( ~n3678 & n24168 ) | ( n17953 & n24168 ) ;
  assign n38058 = n38056 & ~n38057 ;
  assign n38059 = n15855 & n38058 ;
  assign n38060 = n21062 | n35390 ;
  assign n38061 = n11243 | n38060 ;
  assign n38062 = n24216 & ~n27106 ;
  assign n38063 = n21579 ^ n10595 ^ 1'b0 ;
  assign n38064 = n18711 & ~n38063 ;
  assign n38065 = ( n273 & ~n17148 ) | ( n273 & n38064 ) | ( ~n17148 & n38064 ) ;
  assign n38066 = ~n7665 & n14489 ;
  assign n38067 = n38066 ^ n3557 ^ 1'b0 ;
  assign n38068 = n38067 ^ n35513 ^ n33428 ;
  assign n38069 = ( n14050 & ~n15931 ) | ( n14050 & n35747 ) | ( ~n15931 & n35747 ) ;
  assign n38070 = n8732 ^ n2766 ^ 1'b0 ;
  assign n38071 = n21291 & n35860 ;
  assign n38072 = ~n38070 & n38071 ;
  assign n38073 = n27797 ^ n25953 ^ 1'b0 ;
  assign n38074 = n5472 | n38073 ;
  assign n38075 = ~n15252 & n24784 ;
  assign n38076 = n38075 ^ n6482 ^ 1'b0 ;
  assign n38077 = n18109 ^ n4318 ^ 1'b0 ;
  assign n38078 = n24953 & ~n38077 ;
  assign n38079 = ( n27221 & n33003 ) | ( n27221 & n38078 ) | ( n33003 & n38078 ) ;
  assign n38080 = n18209 ^ n511 ^ 1'b0 ;
  assign n38081 = ( n11186 & ~n25688 ) | ( n11186 & n38080 ) | ( ~n25688 & n38080 ) ;
  assign n38082 = n31320 ^ n30464 ^ 1'b0 ;
  assign n38083 = n31359 | n38082 ;
  assign n38084 = n38081 & ~n38083 ;
  assign n38085 = n13952 ^ n4829 ^ 1'b0 ;
  assign n38086 = n14866 & n38085 ;
  assign n38087 = n5752 ^ n1452 ^ 1'b0 ;
  assign n38088 = ~n15549 & n38087 ;
  assign n38089 = n38088 ^ n11630 ^ n1083 ;
  assign n38090 = n6770 & ~n38089 ;
  assign n38091 = ~n6945 & n38090 ;
  assign n38092 = n7094 & ~n20647 ;
  assign n38093 = n38092 ^ n4155 ^ 1'b0 ;
  assign n38094 = n15106 & n38093 ;
  assign n38095 = n27221 & n38094 ;
  assign n38096 = n35427 ^ n26165 ^ n10659 ;
  assign n38097 = ~n16757 & n38096 ;
  assign n38098 = n38097 ^ n36623 ^ 1'b0 ;
  assign n38099 = n10837 ^ n4477 ^ 1'b0 ;
  assign n38100 = n32786 & n38099 ;
  assign n38101 = n30662 & n38100 ;
  assign n38102 = n6094 & ~n24372 ;
  assign n38103 = n38101 & n38102 ;
  assign n38104 = n23123 & ~n24674 ;
  assign n38105 = n38104 ^ n4957 ^ 1'b0 ;
  assign n38109 = ~n12792 & n37469 ;
  assign n38110 = n38109 ^ n6125 ^ 1'b0 ;
  assign n38107 = ( n3475 & ~n6532 ) | ( n3475 & n9986 ) | ( ~n6532 & n9986 ) ;
  assign n38108 = ( ~n6752 & n12225 ) | ( ~n6752 & n38107 ) | ( n12225 & n38107 ) ;
  assign n38106 = n19916 ^ n1106 ^ 1'b0 ;
  assign n38111 = n38110 ^ n38108 ^ n38106 ;
  assign n38112 = n5371 ^ n3926 ^ 1'b0 ;
  assign n38113 = n26025 & ~n38112 ;
  assign n38114 = n21624 ^ n13866 ^ 1'b0 ;
  assign n38115 = ~n2649 & n38114 ;
  assign n38116 = n38115 ^ n4482 ^ 1'b0 ;
  assign n38117 = ~n8634 & n16095 ;
  assign n38118 = n38117 ^ n14578 ^ 1'b0 ;
  assign n38119 = n12547 | n38118 ;
  assign n38120 = ( n5394 & ~n16404 ) | ( n5394 & n20024 ) | ( ~n16404 & n20024 ) ;
  assign n38121 = n38120 ^ n5239 ^ 1'b0 ;
  assign n38122 = ~n10609 & n38121 ;
  assign n38123 = ( n35716 & n38119 ) | ( n35716 & n38122 ) | ( n38119 & n38122 ) ;
  assign n38124 = n9857 ^ n2039 ^ 1'b0 ;
  assign n38125 = n37444 & n38124 ;
  assign n38126 = ~n3030 & n38125 ;
  assign n38127 = n5885 & ~n12513 ;
  assign n38128 = n38127 ^ n10982 ^ 1'b0 ;
  assign n38129 = n13274 | n38128 ;
  assign n38130 = n24888 ^ n11242 ^ 1'b0 ;
  assign n38131 = ~n11437 & n38130 ;
  assign n38132 = n38131 ^ n13377 ^ n6699 ;
  assign n38134 = ( n4390 & ~n6018 ) | ( n4390 & n8647 ) | ( ~n6018 & n8647 ) ;
  assign n38133 = ( n4317 & ~n6113 ) | ( n4317 & n8751 ) | ( ~n6113 & n8751 ) ;
  assign n38135 = n38134 ^ n38133 ^ n2491 ;
  assign n38136 = n15954 & ~n23043 ;
  assign n38137 = n38135 & n38136 ;
  assign n38138 = n11068 ^ n4553 ^ 1'b0 ;
  assign n38139 = n3899 & n38138 ;
  assign n38140 = n36736 & n38139 ;
  assign n38141 = n38140 ^ n22961 ^ n10735 ;
  assign n38146 = n8319 & ~n29748 ;
  assign n38147 = ~n9125 & n38146 ;
  assign n38142 = n18657 & ~n24003 ;
  assign n38143 = n38142 ^ n26071 ^ 1'b0 ;
  assign n38144 = n18126 & ~n38143 ;
  assign n38145 = ~n1711 & n38144 ;
  assign n38148 = n38147 ^ n38145 ^ 1'b0 ;
  assign n38150 = ( n10064 & n17627 ) | ( n10064 & ~n27705 ) | ( n17627 & ~n27705 ) ;
  assign n38149 = n24630 ^ n2580 ^ 1'b0 ;
  assign n38151 = n38150 ^ n38149 ^ 1'b0 ;
  assign n38152 = ~n29956 & n38151 ;
  assign n38153 = n14381 ^ n10053 ^ 1'b0 ;
  assign n38154 = n3792 | n38153 ;
  assign n38155 = n22163 ^ n14660 ^ 1'b0 ;
  assign n38156 = ~n14600 & n18120 ;
  assign n38157 = n38156 ^ n13170 ^ 1'b0 ;
  assign n38158 = ( n1018 & n1671 ) | ( n1018 & n38157 ) | ( n1671 & n38157 ) ;
  assign n38159 = n19752 & ~n24883 ;
  assign n38160 = n7562 & n38159 ;
  assign n38161 = n33186 ^ n20678 ^ n1533 ;
  assign n38162 = n38161 ^ n9236 ^ 1'b0 ;
  assign n38163 = ~n5377 & n10629 ;
  assign n38165 = n12528 & n37398 ;
  assign n38164 = n6706 & n14136 ;
  assign n38166 = n38165 ^ n38164 ^ 1'b0 ;
  assign n38167 = n11443 | n20075 ;
  assign n38168 = n38031 ^ n21763 ^ 1'b0 ;
  assign n38169 = n7961 | n19607 ;
  assign n38170 = n38169 ^ n6152 ^ 1'b0 ;
  assign n38171 = n26023 ^ n3040 ^ 1'b0 ;
  assign n38172 = ~n7035 & n38171 ;
  assign n38173 = n9468 & ~n24169 ;
  assign n38174 = n1194 & ~n16073 ;
  assign n38175 = n6569 & n38174 ;
  assign n38176 = n17099 | n38175 ;
  assign n38177 = n18577 & ~n38176 ;
  assign n38178 = n22164 & ~n38177 ;
  assign n38179 = ~n29109 & n38178 ;
  assign n38180 = n3751 | n38179 ;
  assign n38181 = n38173 & ~n38180 ;
  assign n38182 = n16144 ^ n13620 ^ n5034 ;
  assign n38183 = ( n5269 & n16109 ) | ( n5269 & n18833 ) | ( n16109 & n18833 ) ;
  assign n38184 = ( n25874 & n38182 ) | ( n25874 & n38183 ) | ( n38182 & n38183 ) ;
  assign n38185 = ~n24667 & n34618 ;
  assign n38186 = n5809 & n6090 ;
  assign n38187 = n28243 & n38186 ;
  assign n38188 = n38187 ^ n28910 ^ n18696 ;
  assign n38189 = n21863 ^ n2135 ^ 1'b0 ;
  assign n38190 = ~n38188 & n38189 ;
  assign n38191 = n29241 ^ n9392 ^ 1'b0 ;
  assign n38192 = n25106 & ~n38191 ;
  assign n38193 = n3776 & n38192 ;
  assign n38194 = ~n38190 & n38193 ;
  assign n38195 = ~n19598 & n28647 ;
  assign n38196 = n35404 & ~n38195 ;
  assign n38197 = n38196 ^ n13402 ^ 1'b0 ;
  assign n38198 = n35367 ^ n30115 ^ 1'b0 ;
  assign n38199 = n31059 ^ n21345 ^ 1'b0 ;
  assign n38200 = n38198 & n38199 ;
  assign n38201 = n37879 ^ n3958 ^ 1'b0 ;
  assign n38202 = ~n8157 & n38201 ;
  assign n38203 = n29064 ^ n17047 ^ 1'b0 ;
  assign n38204 = x31 & n15151 ;
  assign n38205 = n38204 ^ n17621 ^ 1'b0 ;
  assign n38207 = n12315 ^ n9422 ^ n7035 ;
  assign n38206 = n567 & n11210 ;
  assign n38208 = n38207 ^ n38206 ^ n29844 ;
  assign n38209 = n20751 ^ n843 ^ 1'b0 ;
  assign n38210 = ~n30856 & n38209 ;
  assign n38211 = n14690 ^ n9879 ^ n3394 ;
  assign n38212 = n24872 & ~n38211 ;
  assign n38213 = n38212 ^ n4590 ^ 1'b0 ;
  assign n38216 = ( ~n5586 & n7216 ) | ( ~n5586 & n8732 ) | ( n7216 & n8732 ) ;
  assign n38214 = n25328 ^ n10179 ^ 1'b0 ;
  assign n38215 = ~n32569 & n38214 ;
  assign n38217 = n38216 ^ n38215 ^ 1'b0 ;
  assign n38218 = n23616 ^ n7525 ^ 1'b0 ;
  assign n38219 = n18001 & ~n38218 ;
  assign n38220 = n27932 & n36729 ;
  assign n38221 = n24425 & n38220 ;
  assign n38222 = n13142 | n15936 ;
  assign n38223 = n6498 & ~n38222 ;
  assign n38224 = n15382 | n21375 ;
  assign n38225 = ~n8312 & n35164 ;
  assign n38226 = n1409 | n17047 ;
  assign n38227 = n15714 | n38226 ;
  assign n38228 = n32781 ^ n32364 ^ x20 ;
  assign n38229 = n35139 ^ n30929 ^ 1'b0 ;
  assign n38233 = n30561 | n32308 ;
  assign n38230 = n10562 & n28602 ;
  assign n38231 = n15050 & ~n38230 ;
  assign n38232 = n38231 ^ n8733 ^ 1'b0 ;
  assign n38234 = n38233 ^ n38232 ^ n12666 ;
  assign n38235 = n38234 ^ n25455 ^ n25046 ;
  assign n38236 = n16121 ^ n7244 ^ 1'b0 ;
  assign n38237 = n7639 | n38236 ;
  assign n38238 = n38237 ^ n34850 ^ n29440 ;
  assign n38239 = n1832 | n4472 ;
  assign n38240 = n11555 & ~n38239 ;
  assign n38241 = n38240 ^ n37974 ^ 1'b0 ;
  assign n38242 = n7801 ^ n3910 ^ 1'b0 ;
  assign n38243 = n35157 & n38242 ;
  assign n38244 = ~n14762 & n33404 ;
  assign n38245 = ~n38243 & n38244 ;
  assign n38247 = ( n2103 & n2225 ) | ( n2103 & n23274 ) | ( n2225 & n23274 ) ;
  assign n38246 = ~n10817 & n21245 ;
  assign n38248 = n38247 ^ n38246 ^ 1'b0 ;
  assign n38249 = n8251 ^ n423 ^ 1'b0 ;
  assign n38250 = n38249 ^ n8975 ^ n6799 ;
  assign n38251 = n6776 & n22725 ;
  assign n38252 = n8075 ^ n5044 ^ 1'b0 ;
  assign n38253 = n27058 & n38252 ;
  assign n38254 = n19977 & n38253 ;
  assign n38255 = ( n7801 & n17517 ) | ( n7801 & n38254 ) | ( n17517 & n38254 ) ;
  assign n38256 = n3766 | n18821 ;
  assign n38257 = n13762 & n38256 ;
  assign n38258 = n18409 & n38257 ;
  assign n38259 = n18726 ^ n11777 ^ 1'b0 ;
  assign n38260 = n38259 ^ n9944 ^ 1'b0 ;
  assign n38261 = n4575 & n6062 ;
  assign n38262 = n10839 & n38261 ;
  assign n38263 = n38262 ^ n17035 ^ 1'b0 ;
  assign n38264 = n11966 | n15065 ;
  assign n38265 = n38263 & n38264 ;
  assign n38266 = ~n36477 & n38265 ;
  assign n38267 = ( n593 & ~n17290 ) | ( n593 & n22469 ) | ( ~n17290 & n22469 ) ;
  assign n38270 = n13152 ^ n1602 ^ 1'b0 ;
  assign n38268 = n11007 ^ n6172 ^ 1'b0 ;
  assign n38269 = n22052 & ~n38268 ;
  assign n38271 = n38270 ^ n38269 ^ n13660 ;
  assign n38272 = ( x219 & ~n2363 ) | ( x219 & n15746 ) | ( ~n2363 & n15746 ) ;
  assign n38273 = n38272 ^ n20718 ^ 1'b0 ;
  assign n38274 = n2708 | n4673 ;
  assign n38275 = n14440 | n38274 ;
  assign n38276 = n1304 & n7715 ;
  assign n38277 = n22207 ^ n18949 ^ n7677 ;
  assign n38278 = n12131 | n38277 ;
  assign n38279 = n38278 ^ n30348 ^ 1'b0 ;
  assign n38280 = ( n38275 & n38276 ) | ( n38275 & n38279 ) | ( n38276 & n38279 ) ;
  assign n38281 = ( n1142 & ~n9861 ) | ( n1142 & n36474 ) | ( ~n9861 & n36474 ) ;
  assign n38282 = n17144 ^ n11296 ^ n10579 ;
  assign n38283 = x226 & n5430 ;
  assign n38284 = n2958 & n3418 ;
  assign n38285 = n16644 & n38284 ;
  assign n38286 = n23439 ^ n13816 ^ 1'b0 ;
  assign n38287 = n38285 | n38286 ;
  assign n38288 = ( ~n7553 & n22957 ) | ( ~n7553 & n34211 ) | ( n22957 & n34211 ) ;
  assign n38289 = n28668 ^ n675 ^ 1'b0 ;
  assign n38290 = n38288 & n38289 ;
  assign n38291 = ( n7466 & ~n16739 ) | ( n7466 & n32599 ) | ( ~n16739 & n32599 ) ;
  assign n38292 = n14878 & ~n38291 ;
  assign n38293 = ~n32227 & n38292 ;
  assign n38294 = n7004 ^ n1327 ^ 1'b0 ;
  assign n38295 = n3864 & n38294 ;
  assign n38296 = n38293 | n38295 ;
  assign n38297 = ( ~n12736 & n22462 ) | ( ~n12736 & n24195 ) | ( n22462 & n24195 ) ;
  assign n38298 = n34447 ^ n1775 ^ n711 ;
  assign n38299 = ( n28312 & n34368 ) | ( n28312 & ~n38298 ) | ( n34368 & ~n38298 ) ;
  assign n38300 = n6576 & n38134 ;
  assign n38301 = n10509 | n21252 ;
  assign n38302 = n4916 & ~n38301 ;
  assign n38303 = n38302 ^ n23112 ^ 1'b0 ;
  assign n38304 = n38300 | n38303 ;
  assign n38305 = n38304 ^ n29836 ^ 1'b0 ;
  assign n38306 = n21003 & ~n38305 ;
  assign n38307 = n16290 & ~n35907 ;
  assign n38308 = n38307 ^ n20630 ^ 1'b0 ;
  assign n38309 = n6048 ^ x183 ^ 1'b0 ;
  assign n38310 = n11898 & n38309 ;
  assign n38311 = ~n8286 & n38310 ;
  assign n38312 = n25913 & ~n38311 ;
  assign n38313 = n8732 ^ n2744 ^ 1'b0 ;
  assign n38314 = ~n2396 & n3547 ;
  assign n38315 = ~n10826 & n38314 ;
  assign n38316 = ~n38313 & n38315 ;
  assign n38317 = n38312 & ~n38316 ;
  assign n38318 = n38317 ^ n32095 ^ 1'b0 ;
  assign n38319 = n28622 ^ n4032 ^ 1'b0 ;
  assign n38320 = n11984 ^ n4963 ^ 1'b0 ;
  assign n38321 = n36824 ^ n24070 ^ n15785 ;
  assign n38325 = ~n5564 & n6074 ;
  assign n38326 = n38325 ^ n26621 ^ 1'b0 ;
  assign n38327 = ~n3535 & n38326 ;
  assign n38323 = ( n11474 & ~n16096 ) | ( n11474 & n37138 ) | ( ~n16096 & n37138 ) ;
  assign n38324 = n38323 ^ n12498 ^ n8587 ;
  assign n38322 = n18825 & n20613 ;
  assign n38328 = n38327 ^ n38324 ^ n38322 ;
  assign n38330 = ~n16423 & n26265 ;
  assign n38329 = n4294 & n33053 ;
  assign n38331 = n38330 ^ n38329 ^ 1'b0 ;
  assign n38332 = n36422 ^ n18418 ^ 1'b0 ;
  assign n38333 = n14131 & ~n38332 ;
  assign n38334 = n1045 | n14333 ;
  assign n38335 = n19261 | n38334 ;
  assign n38336 = n38335 ^ n15859 ^ 1'b0 ;
  assign n38337 = n9263 | n38336 ;
  assign n38338 = n7220 | n13956 ;
  assign n38339 = n38338 ^ n28214 ^ 1'b0 ;
  assign n38340 = n14811 & n38339 ;
  assign n38341 = n10353 ^ n6021 ^ 1'b0 ;
  assign n38342 = n5012 | n38341 ;
  assign n38343 = ( n8633 & n23469 ) | ( n8633 & n27679 ) | ( n23469 & n27679 ) ;
  assign n38344 = n14172 ^ n2735 ^ 1'b0 ;
  assign n38345 = ~n38343 & n38344 ;
  assign n38346 = n8446 & n19724 ;
  assign n38347 = ~n6411 & n34806 ;
  assign n38348 = n21450 & n38347 ;
  assign n38349 = n38348 ^ n22861 ^ n12264 ;
  assign n38353 = n14497 ^ n6921 ^ 1'b0 ;
  assign n38354 = n15668 | n38353 ;
  assign n38350 = ( n4462 & n5087 ) | ( n4462 & ~n14606 ) | ( n5087 & ~n14606 ) ;
  assign n38351 = ~n27861 & n38350 ;
  assign n38352 = ~n27702 & n38351 ;
  assign n38355 = n38354 ^ n38352 ^ n37744 ;
  assign n38356 = n4881 & ~n13395 ;
  assign n38357 = n5454 & n38356 ;
  assign n38358 = ( n1830 & n8737 ) | ( n1830 & n12746 ) | ( n8737 & n12746 ) ;
  assign n38359 = ~n7069 & n38358 ;
  assign n38360 = ~n21382 & n38359 ;
  assign n38361 = n5675 & ~n38360 ;
  assign n38362 = n38361 ^ n3019 ^ 1'b0 ;
  assign n38363 = n23047 ^ n20199 ^ 1'b0 ;
  assign n38364 = n6082 | n38363 ;
  assign n38365 = n8368 & n25153 ;
  assign n38366 = ~n6856 & n38365 ;
  assign n38367 = n38366 ^ n10824 ^ n8927 ;
  assign n38368 = n19680 & ~n32257 ;
  assign n38369 = ( n3198 & n36381 ) | ( n3198 & ~n38368 ) | ( n36381 & ~n38368 ) ;
  assign n38370 = n21980 ^ n15022 ^ n14266 ;
  assign n38371 = n34973 ^ n29625 ^ n14393 ;
  assign n38372 = n38371 ^ n25582 ^ n735 ;
  assign n38373 = ~n20404 & n32133 ;
  assign n38374 = n3307 | n15203 ;
  assign n38375 = n38374 ^ n25876 ^ 1'b0 ;
  assign n38376 = n3207 & n29025 ;
  assign n38377 = ~n7320 & n38376 ;
  assign n38378 = ( n8952 & n24490 ) | ( n8952 & ~n38377 ) | ( n24490 & ~n38377 ) ;
  assign n38379 = ~n21573 & n38378 ;
  assign n38380 = ~n38375 & n38379 ;
  assign n38381 = n14742 & ~n38380 ;
  assign n38382 = n16095 ^ n3610 ^ n2257 ;
  assign n38383 = n38382 ^ n10391 ^ 1'b0 ;
  assign n38384 = ~n3636 & n38383 ;
  assign n38385 = n14138 | n15654 ;
  assign n38386 = n38385 ^ n20379 ^ 1'b0 ;
  assign n38387 = n4496 & n11920 ;
  assign n38388 = n38387 ^ n29747 ^ 1'b0 ;
  assign n38389 = ( ~n38384 & n38386 ) | ( ~n38384 & n38388 ) | ( n38386 & n38388 ) ;
  assign n38390 = ~n1908 & n7254 ;
  assign n38391 = n17589 & n38390 ;
  assign n38392 = n38391 ^ n16017 ^ 1'b0 ;
  assign n38393 = n24250 ^ n13625 ^ n4520 ;
  assign n38394 = x219 & n38393 ;
  assign n38395 = n3739 & ~n12255 ;
  assign n38396 = ~n2733 & n38395 ;
  assign n38397 = n17806 | n19679 ;
  assign n38398 = n38397 ^ n6204 ^ 1'b0 ;
  assign n38399 = ~n20785 & n38398 ;
  assign n38400 = ( ~n6458 & n7282 ) | ( ~n6458 & n8843 ) | ( n7282 & n8843 ) ;
  assign n38401 = n29173 & n38400 ;
  assign n38402 = n16059 ^ n3688 ^ 1'b0 ;
  assign n38403 = n21070 & ~n38402 ;
  assign n38404 = n37639 ^ n25583 ^ 1'b0 ;
  assign n38405 = n12701 | n38404 ;
  assign n38406 = n23455 ^ n3046 ^ 1'b0 ;
  assign n38407 = n12550 ^ n4363 ^ 1'b0 ;
  assign n38408 = n1022 | n38407 ;
  assign n38409 = n38406 & ~n38408 ;
  assign n38410 = n38409 ^ n28857 ^ n28187 ;
  assign n38411 = n15739 ^ n4565 ^ 1'b0 ;
  assign n38412 = n38411 ^ n1115 ^ 1'b0 ;
  assign n38419 = ~n12474 & n20813 ;
  assign n38420 = n28753 & ~n38419 ;
  assign n38421 = n38420 ^ n15590 ^ 1'b0 ;
  assign n38413 = ~n3702 & n12289 ;
  assign n38414 = n2734 & n7210 ;
  assign n38415 = ~n17394 & n38414 ;
  assign n38416 = n25984 | n38415 ;
  assign n38417 = n38413 & ~n38416 ;
  assign n38418 = n5259 & ~n38417 ;
  assign n38422 = n38421 ^ n38418 ^ 1'b0 ;
  assign n38423 = n37379 & n38422 ;
  assign n38424 = n38423 ^ n10465 ^ 1'b0 ;
  assign n38425 = ~n23342 & n31161 ;
  assign n38426 = n14596 ^ n9614 ^ 1'b0 ;
  assign n38427 = n630 | n34311 ;
  assign n38428 = n31961 ^ n9002 ^ 1'b0 ;
  assign n38429 = ( n2071 & ~n6658 ) | ( n2071 & n24394 ) | ( ~n6658 & n24394 ) ;
  assign n38430 = n12473 | n27636 ;
  assign n38431 = n7917 & ~n12587 ;
  assign n38432 = n15421 ^ n9812 ^ 1'b0 ;
  assign n38433 = n20897 & n38432 ;
  assign n38434 = n11159 ^ n5263 ^ 1'b0 ;
  assign n38435 = n848 | n38434 ;
  assign n38436 = n27832 ^ n7189 ^ 1'b0 ;
  assign n38437 = ~n38435 & n38436 ;
  assign n38438 = n2672 & ~n6127 ;
  assign n38439 = n38438 ^ n10428 ^ 1'b0 ;
  assign n38440 = ~n13409 & n38439 ;
  assign n38441 = ( x62 & n19284 ) | ( x62 & n38440 ) | ( n19284 & n38440 ) ;
  assign n38442 = n1562 | n18960 ;
  assign n38443 = n7915 & n38442 ;
  assign n38444 = n32477 & n38443 ;
  assign n38445 = n38441 & ~n38444 ;
  assign n38446 = n27923 & n38445 ;
  assign n38447 = n3106 | n37639 ;
  assign n38448 = n27058 | n38447 ;
  assign n38449 = ( n3268 & ~n6775 ) | ( n3268 & n24291 ) | ( ~n6775 & n24291 ) ;
  assign n38450 = n4700 | n21131 ;
  assign n38451 = n38450 ^ n22438 ^ n805 ;
  assign n38452 = n3891 & ~n17592 ;
  assign n38453 = ~n26503 & n38452 ;
  assign n38454 = n1145 & n38453 ;
  assign n38455 = ( n6127 & n7982 ) | ( n6127 & n36846 ) | ( n7982 & n36846 ) ;
  assign n38456 = n38455 ^ n22628 ^ n16926 ;
  assign n38457 = n38456 ^ n38273 ^ 1'b0 ;
  assign n38458 = ( n6034 & n9709 ) | ( n6034 & n10599 ) | ( n9709 & n10599 ) ;
  assign n38459 = n675 & n4816 ;
  assign n38460 = ~n344 & n38459 ;
  assign n38461 = ( ~n1000 & n30282 ) | ( ~n1000 & n38460 ) | ( n30282 & n38460 ) ;
  assign n38462 = n16032 & n35992 ;
  assign n38463 = ~n6201 & n31463 ;
  assign n38464 = ( n26799 & n30361 ) | ( n26799 & n38463 ) | ( n30361 & n38463 ) ;
  assign n38465 = ~n2682 & n5121 ;
  assign n38466 = n35420 ^ n3067 ^ 1'b0 ;
  assign n38467 = ( n6938 & n7168 ) | ( n6938 & ~n23825 ) | ( n7168 & ~n23825 ) ;
  assign n38468 = n2883 | n20168 ;
  assign n38469 = ( n34238 & n34357 ) | ( n34238 & ~n38468 ) | ( n34357 & ~n38468 ) ;
  assign n38470 = n29501 ^ n9109 ^ 1'b0 ;
  assign n38471 = n7380 & ~n18915 ;
  assign n38472 = ( n4736 & n30278 ) | ( n4736 & n38471 ) | ( n30278 & n38471 ) ;
  assign n38476 = n25937 ^ n21648 ^ 1'b0 ;
  assign n38473 = n20621 ^ n2299 ^ 1'b0 ;
  assign n38474 = ~n19993 & n38473 ;
  assign n38475 = n38474 ^ n8276 ^ n5370 ;
  assign n38477 = n38476 ^ n38475 ^ 1'b0 ;
  assign n38478 = n38472 & ~n38477 ;
  assign n38479 = ~n7723 & n22821 ;
  assign n38480 = n14688 ^ n7855 ^ 1'b0 ;
  assign n38481 = n10516 & n38480 ;
  assign n38482 = n20641 ^ n11072 ^ 1'b0 ;
  assign n38483 = n2628 | n38482 ;
  assign n38484 = n9987 ^ n7057 ^ 1'b0 ;
  assign n38485 = ~n38483 & n38484 ;
  assign n38486 = n26806 ^ n4515 ^ 1'b0 ;
  assign n38487 = n38485 & ~n38486 ;
  assign n38488 = n9004 & n38487 ;
  assign n38489 = n38488 ^ n3470 ^ 1'b0 ;
  assign n38490 = n5944 ^ n4379 ^ n3986 ;
  assign n38491 = n38490 ^ n2356 ^ 1'b0 ;
  assign n38492 = n19872 & ~n38491 ;
  assign n38493 = n5291 | n6791 ;
  assign n38494 = n15060 ^ n5397 ^ 1'b0 ;
  assign n38495 = n12853 & n38494 ;
  assign n38496 = n19453 & n38495 ;
  assign n38497 = ( n38492 & n38493 ) | ( n38492 & ~n38496 ) | ( n38493 & ~n38496 ) ;
  assign n38498 = n24558 ^ n13041 ^ 1'b0 ;
  assign n38499 = n38498 ^ n16592 ^ n5439 ;
  assign n38500 = n10401 | n38499 ;
  assign n38501 = n25793 ^ n18860 ^ 1'b0 ;
  assign n38502 = ~n16548 & n30044 ;
  assign n38503 = n34377 ^ n2259 ^ 1'b0 ;
  assign n38504 = n20924 & ~n38503 ;
  assign n38505 = ( n24667 & n27138 ) | ( n24667 & n35855 ) | ( n27138 & n35855 ) ;
  assign n38506 = n356 & n7471 ;
  assign n38507 = n38506 ^ n33663 ^ 1'b0 ;
  assign n38509 = n7556 & ~n19801 ;
  assign n38510 = n38509 ^ n31806 ^ 1'b0 ;
  assign n38508 = n23774 ^ n23274 ^ 1'b0 ;
  assign n38511 = n38510 ^ n38508 ^ n20186 ;
  assign n38512 = n10014 ^ n2372 ^ 1'b0 ;
  assign n38513 = n2822 & n38512 ;
  assign n38514 = n37325 ^ n2328 ^ 1'b0 ;
  assign n38515 = n2906 | n38514 ;
  assign n38516 = ~n14127 & n29851 ;
  assign n38517 = n38515 & n38516 ;
  assign n38518 = n5362 | n33720 ;
  assign n38519 = n36260 ^ n7904 ^ 1'b0 ;
  assign n38520 = n16543 & n34401 ;
  assign n38521 = n2500 & ~n9071 ;
  assign n38522 = n38521 ^ n18639 ^ 1'b0 ;
  assign n38524 = n25742 ^ n18797 ^ n9777 ;
  assign n38523 = n5255 ^ n4477 ^ 1'b0 ;
  assign n38525 = n38524 ^ n38523 ^ n8956 ;
  assign n38526 = ( n19013 & ~n20168 ) | ( n19013 & n23936 ) | ( ~n20168 & n23936 ) ;
  assign n38527 = ~n2790 & n12094 ;
  assign n38528 = n10437 & ~n35126 ;
  assign n38529 = n4041 & n38528 ;
  assign n38530 = n9280 & n34488 ;
  assign n38531 = n4369 & n38530 ;
  assign n38532 = n16429 & n17533 ;
  assign n38533 = n38531 & n38532 ;
  assign n38534 = n16019 & n25033 ;
  assign n38535 = n8389 | n38534 ;
  assign n38536 = n38533 & ~n38535 ;
  assign n38537 = n32682 ^ n20382 ^ n15738 ;
  assign n38538 = ( ~n12362 & n25853 ) | ( ~n12362 & n36143 ) | ( n25853 & n36143 ) ;
  assign n38539 = n29949 & ~n30282 ;
  assign n38540 = n38539 ^ n30650 ^ n16878 ;
  assign n38541 = n7958 & ~n23967 ;
  assign n38542 = n38541 ^ n425 ^ 1'b0 ;
  assign n38543 = n38542 ^ n22631 ^ 1'b0 ;
  assign n38544 = n12691 & n38543 ;
  assign n38545 = n38544 ^ n6547 ^ 1'b0 ;
  assign n38546 = n38545 ^ n8067 ^ 1'b0 ;
  assign n38547 = ( n9206 & n16390 ) | ( n9206 & ~n35622 ) | ( n16390 & ~n35622 ) ;
  assign n38548 = n38546 & n38547 ;
  assign n38549 = n21326 ^ n16261 ^ 1'b0 ;
  assign n38550 = n11536 & ~n38549 ;
  assign n38551 = n38550 ^ n33670 ^ 1'b0 ;
  assign n38552 = n11447 & ~n12011 ;
  assign n38553 = n30899 ^ n15902 ^ 1'b0 ;
  assign n38554 = n9237 ^ n2463 ^ 1'b0 ;
  assign n38555 = ( n10789 & n14637 ) | ( n10789 & n38554 ) | ( n14637 & n38554 ) ;
  assign n38556 = n26462 & ~n38555 ;
  assign n38557 = n38556 ^ n13879 ^ 1'b0 ;
  assign n38558 = n15971 & ~n38557 ;
  assign n38559 = ~x103 & n38558 ;
  assign n38560 = n38559 ^ n31463 ^ n14466 ;
  assign n38561 = n18853 ^ n5223 ^ 1'b0 ;
  assign n38562 = ( ~n1465 & n5277 ) | ( ~n1465 & n38561 ) | ( n5277 & n38561 ) ;
  assign n38563 = n36574 ^ n7499 ^ n4244 ;
  assign n38564 = ( n14912 & n32063 ) | ( n14912 & ~n38563 ) | ( n32063 & ~n38563 ) ;
  assign n38565 = n22438 & n34891 ;
  assign n38566 = n2228 | n10931 ;
  assign n38567 = n38565 | n38566 ;
  assign n38569 = n8303 ^ n5746 ^ 1'b0 ;
  assign n38568 = ~n10355 & n20992 ;
  assign n38570 = n38569 ^ n38568 ^ 1'b0 ;
  assign n38571 = n29615 ^ n25411 ^ 1'b0 ;
  assign n38572 = n18123 & n38571 ;
  assign n38573 = n1751 & n19878 ;
  assign n38574 = n2221 & n10154 ;
  assign n38575 = ~n1666 & n38574 ;
  assign n38576 = n38575 ^ n15290 ^ n5698 ;
  assign n38577 = ( n14898 & n18617 ) | ( n14898 & n22946 ) | ( n18617 & n22946 ) ;
  assign n38578 = n38577 ^ n2272 ^ 1'b0 ;
  assign n38581 = n23669 & n27530 ;
  assign n38579 = ~n7394 & n18887 ;
  assign n38580 = ~n3197 & n38579 ;
  assign n38582 = n38581 ^ n38580 ^ 1'b0 ;
  assign n38583 = n13397 & ~n20958 ;
  assign n38584 = ~n5163 & n38583 ;
  assign n38585 = ~n4448 & n8531 ;
  assign n38586 = n27776 & ~n38585 ;
  assign n38587 = n16885 ^ n10794 ^ 1'b0 ;
  assign n38588 = n14304 & ~n38587 ;
  assign n38589 = n34551 ^ n25306 ^ 1'b0 ;
  assign n38590 = n2717 & ~n38589 ;
  assign n38591 = n10764 | n30467 ;
  assign n38592 = n21470 & n38591 ;
  assign n38593 = n38592 ^ n35370 ^ 1'b0 ;
  assign n38594 = ~n22935 & n26916 ;
  assign n38597 = n10457 ^ n5973 ^ 1'b0 ;
  assign n38595 = ( n8463 & ~n17136 ) | ( n8463 & n28979 ) | ( ~n17136 & n28979 ) ;
  assign n38596 = n10794 | n38595 ;
  assign n38598 = n38597 ^ n38596 ^ 1'b0 ;
  assign n38599 = n5424 | n7976 ;
  assign n38600 = ~n20319 & n38599 ;
  assign n38601 = n38600 ^ n30160 ^ n24037 ;
  assign n38602 = n1827 ^ n877 ^ 1'b0 ;
  assign n38603 = ~n11710 & n38602 ;
  assign n38604 = ~n4063 & n38603 ;
  assign n38605 = n22482 ^ n5215 ^ 1'b0 ;
  assign n38606 = ~n3851 & n25220 ;
  assign n38607 = ( n25850 & ~n33414 ) | ( n25850 & n38606 ) | ( ~n33414 & n38606 ) ;
  assign n38608 = n13736 & ~n38607 ;
  assign n38609 = n7177 & n36411 ;
  assign n38610 = n2465 & n38609 ;
  assign n38611 = n38610 ^ n22784 ^ 1'b0 ;
  assign n38612 = n38611 ^ n13167 ^ n8644 ;
  assign n38614 = n24370 | n28459 ;
  assign n38615 = n38614 ^ n16469 ^ 1'b0 ;
  assign n38613 = n30367 ^ n5108 ^ 1'b0 ;
  assign n38616 = n38615 ^ n38613 ^ n9015 ;
  assign n38617 = ( n4338 & n5233 ) | ( n4338 & ~n12858 ) | ( n5233 & ~n12858 ) ;
  assign n38618 = n38617 ^ n5481 ^ 1'b0 ;
  assign n38619 = n2909 & n23092 ;
  assign n38620 = n38619 ^ n12526 ^ 1'b0 ;
  assign n38621 = n493 & n13130 ;
  assign n38622 = n24499 & ~n38621 ;
  assign n38623 = n38622 ^ n22595 ^ 1'b0 ;
  assign n38624 = n29810 ^ n15738 ^ 1'b0 ;
  assign n38625 = n38624 ^ n2119 ^ 1'b0 ;
  assign n38626 = n13201 & ~n22150 ;
  assign n38627 = n4097 & n16599 ;
  assign n38628 = n38627 ^ n945 ^ 1'b0 ;
  assign n38629 = n6980 & ~n38628 ;
  assign n38630 = ~n27769 & n37888 ;
  assign n38631 = n17903 & n27620 ;
  assign n38632 = n879 | n17642 ;
  assign n38633 = n3935 & ~n5405 ;
  assign n38634 = ( ~n2705 & n3190 ) | ( ~n2705 & n38633 ) | ( n3190 & n38633 ) ;
  assign n38635 = ~n30702 & n38634 ;
  assign n38636 = n38635 ^ n13461 ^ 1'b0 ;
  assign n38637 = n36572 ^ n23398 ^ n1133 ;
  assign n38638 = ~n2381 & n23665 ;
  assign n38639 = ~n955 & n2957 ;
  assign n38640 = ~n38638 & n38639 ;
  assign n38641 = n21523 | n38640 ;
  assign n38642 = n12064 & n22352 ;
  assign n38643 = ~n23223 & n25770 ;
  assign n38644 = n11328 & ~n20438 ;
  assign n38645 = n25171 & n38644 ;
  assign n38646 = n21045 & n38645 ;
  assign n38647 = n38646 ^ n9003 ^ 1'b0 ;
  assign n38649 = n17620 ^ n1927 ^ 1'b0 ;
  assign n38648 = n38211 ^ n9936 ^ n754 ;
  assign n38650 = n38649 ^ n38648 ^ n2754 ;
  assign n38651 = n8038 & ~n29553 ;
  assign n38652 = n14004 ^ n9245 ^ 1'b0 ;
  assign n38653 = n10321 & ~n38652 ;
  assign n38654 = n9228 & n22785 ;
  assign n38655 = n7513 & ~n10485 ;
  assign n38656 = ~n26591 & n38655 ;
  assign n38657 = n17621 ^ n13968 ^ 1'b0 ;
  assign n38658 = n12676 ^ n11463 ^ n4827 ;
  assign n38659 = n35478 ^ n7976 ^ 1'b0 ;
  assign n38660 = n10464 & ~n13731 ;
  assign n38661 = n8981 & n12194 ;
  assign n38662 = n5294 | n25528 ;
  assign n38663 = n15800 & ~n38662 ;
  assign n38664 = n12273 & ~n38663 ;
  assign n38665 = ~n38661 & n38664 ;
  assign n38666 = n3567 | n11567 ;
  assign n38667 = n38666 ^ n9591 ^ 1'b0 ;
  assign n38668 = n12303 ^ n6473 ^ 1'b0 ;
  assign n38669 = n38667 & ~n38668 ;
  assign n38670 = n12648 ^ n7637 ^ 1'b0 ;
  assign n38671 = n19753 ^ n7569 ^ 1'b0 ;
  assign n38672 = ~n38670 & n38671 ;
  assign n38673 = n1103 | n9952 ;
  assign n38674 = n38673 ^ n30611 ^ 1'b0 ;
  assign n38675 = n38672 & ~n38674 ;
  assign n38676 = n3469 ^ n2075 ^ 1'b0 ;
  assign n38677 = n38676 ^ n34093 ^ 1'b0 ;
  assign n38678 = n23732 ^ n3203 ^ 1'b0 ;
  assign n38679 = n5672 & ~n13976 ;
  assign n38680 = ~n4469 & n38679 ;
  assign n38681 = x26 | n38680 ;
  assign n38682 = n1154 & ~n7789 ;
  assign n38683 = n38682 ^ n19419 ^ 1'b0 ;
  assign n38684 = ( ~n7137 & n32863 ) | ( ~n7137 & n38683 ) | ( n32863 & n38683 ) ;
  assign n38685 = ( ~n9341 & n11982 ) | ( ~n9341 & n38684 ) | ( n11982 & n38684 ) ;
  assign n38686 = n11584 ^ n10928 ^ n5649 ;
  assign n38687 = n31334 ^ n4614 ^ n2660 ;
  assign n38688 = n18606 ^ n12129 ^ 1'b0 ;
  assign n38689 = n20952 | n38688 ;
  assign n38690 = n12374 ^ n8193 ^ 1'b0 ;
  assign n38691 = n8551 & n38690 ;
  assign n38693 = n1669 | n5999 ;
  assign n38692 = ~n1870 & n18600 ;
  assign n38694 = n38693 ^ n38692 ^ 1'b0 ;
  assign n38695 = n3885 ^ n2240 ^ 1'b0 ;
  assign n38696 = ~n10573 & n38695 ;
  assign n38697 = n5322 & n38696 ;
  assign n38698 = n38697 ^ n17532 ^ 1'b0 ;
  assign n38699 = n10726 & ~n14118 ;
  assign n38700 = ~n14687 & n38699 ;
  assign n38701 = n21549 & n38700 ;
  assign n38702 = ( n12157 & ~n16643 ) | ( n12157 & n38701 ) | ( ~n16643 & n38701 ) ;
  assign n38703 = n11080 ^ n1999 ^ 1'b0 ;
  assign n38704 = n19292 & ~n22209 ;
  assign n38705 = n38704 ^ n30636 ^ 1'b0 ;
  assign n38706 = ( n21866 & n38703 ) | ( n21866 & n38705 ) | ( n38703 & n38705 ) ;
  assign n38707 = n34241 ^ n9709 ^ 1'b0 ;
  assign n38708 = n21566 & n38707 ;
  assign n38709 = ( n7622 & ~n30669 ) | ( n7622 & n38708 ) | ( ~n30669 & n38708 ) ;
  assign n38710 = n38709 ^ n11364 ^ 1'b0 ;
  assign n38711 = n15619 & ~n29896 ;
  assign n38712 = n30078 & n38711 ;
  assign n38713 = ( n2972 & ~n13280 ) | ( n2972 & n38712 ) | ( ~n13280 & n38712 ) ;
  assign n38714 = n28646 & n38713 ;
  assign n38715 = n12999 ^ x206 ^ 1'b0 ;
  assign n38716 = n9316 ^ n3767 ^ 1'b0 ;
  assign n38717 = n38716 ^ n37521 ^ 1'b0 ;
  assign n38718 = n11620 & n27447 ;
  assign n38719 = n38718 ^ n6848 ^ 1'b0 ;
  assign n38720 = n1040 & n9343 ;
  assign n38721 = n2841 & n38720 ;
  assign n38722 = ( ~n6756 & n11551 ) | ( ~n6756 & n19558 ) | ( n11551 & n19558 ) ;
  assign n38723 = n38722 ^ n3633 ^ 1'b0 ;
  assign n38724 = n38721 | n38723 ;
  assign n38725 = n38724 ^ n18256 ^ 1'b0 ;
  assign n38726 = ~n25960 & n38725 ;
  assign n38727 = n3859 | n28602 ;
  assign n38728 = n20196 | n38727 ;
  assign n38729 = ( n7135 & n24792 ) | ( n7135 & n38728 ) | ( n24792 & n38728 ) ;
  assign n38730 = n14804 | n22108 ;
  assign n38731 = n15432 & ~n38730 ;
  assign n38732 = n38731 ^ n11917 ^ n7905 ;
  assign n38733 = ( ~n9699 & n9933 ) | ( ~n9699 & n38732 ) | ( n9933 & n38732 ) ;
  assign n38734 = ( n29603 & ~n36376 ) | ( n29603 & n38733 ) | ( ~n36376 & n38733 ) ;
  assign n38735 = n23156 & n35154 ;
  assign n38736 = n13191 | n25451 ;
  assign n38737 = ~n18032 & n33054 ;
  assign n38738 = n38737 ^ n11597 ^ 1'b0 ;
  assign n38739 = n33779 ^ n18913 ^ 1'b0 ;
  assign n38740 = ~n18208 & n38739 ;
  assign n38742 = n38029 ^ n16524 ^ n3651 ;
  assign n38741 = n5872 & n7548 ;
  assign n38743 = n38742 ^ n38741 ^ n1653 ;
  assign n38744 = n6209 ^ n2570 ^ 1'b0 ;
  assign n38745 = n13493 & ~n38744 ;
  assign n38746 = ~n28067 & n38745 ;
  assign n38747 = n37289 ^ n10168 ^ 1'b0 ;
  assign n38748 = n4361 | n38747 ;
  assign n38749 = ( n3532 & n8179 ) | ( n3532 & ~n38748 ) | ( n8179 & ~n38748 ) ;
  assign n38750 = n38749 ^ n2261 ^ 1'b0 ;
  assign n38751 = ~n25057 & n30472 ;
  assign n38752 = n24606 ^ n7535 ^ 1'b0 ;
  assign n38753 = ( n4495 & n23294 ) | ( n4495 & ~n38752 ) | ( n23294 & ~n38752 ) ;
  assign n38754 = n38753 ^ n9520 ^ 1'b0 ;
  assign n38755 = n26818 | n38754 ;
  assign n38756 = n38755 ^ n6656 ^ 1'b0 ;
  assign n38757 = n326 | n38756 ;
  assign n38758 = n38069 ^ n35522 ^ 1'b0 ;
  assign n38759 = n35807 ^ n24397 ^ 1'b0 ;
  assign n38761 = n4797 & n32930 ;
  assign n38762 = n38761 ^ n12589 ^ 1'b0 ;
  assign n38760 = n9467 & n16681 ;
  assign n38763 = n38762 ^ n38760 ^ 1'b0 ;
  assign n38764 = n38763 ^ n27990 ^ n20157 ;
  assign n38765 = ( ~n6989 & n25302 ) | ( ~n6989 & n38764 ) | ( n25302 & n38764 ) ;
  assign n38768 = n574 | n3473 ;
  assign n38769 = n38768 ^ n11274 ^ 1'b0 ;
  assign n38770 = ~n23057 & n38769 ;
  assign n38771 = n38770 ^ n27427 ^ n6015 ;
  assign n38766 = n6805 & ~n33837 ;
  assign n38767 = ( n980 & ~n10597 ) | ( n980 & n38766 ) | ( ~n10597 & n38766 ) ;
  assign n38772 = n38771 ^ n38767 ^ n4723 ;
  assign n38773 = n22785 ^ n11471 ^ n1576 ;
  assign n38775 = n12863 ^ n10900 ^ 1'b0 ;
  assign n38776 = n1849 & n38775 ;
  assign n38774 = ~n549 & n10281 ;
  assign n38777 = n38776 ^ n38774 ^ 1'b0 ;
  assign n38778 = n38777 ^ n7546 ^ 1'b0 ;
  assign n38779 = n38773 & n38778 ;
  assign n38780 = ~n24057 & n37623 ;
  assign n38781 = n6565 | n13789 ;
  assign n38782 = n38780 & ~n38781 ;
  assign n38783 = ( n1291 & n3589 ) | ( n1291 & n8426 ) | ( n3589 & n8426 ) ;
  assign n38784 = n38783 ^ n13449 ^ 1'b0 ;
  assign n38785 = ~n28248 & n38784 ;
  assign n38786 = n26071 ^ x36 ^ 1'b0 ;
  assign n38787 = n38786 ^ n11981 ^ n1671 ;
  assign n38789 = n5713 & ~n20291 ;
  assign n38790 = n38789 ^ n32397 ^ 1'b0 ;
  assign n38791 = n24577 | n38790 ;
  assign n38788 = n17579 ^ n15313 ^ 1'b0 ;
  assign n38792 = n38791 ^ n38788 ^ n33753 ;
  assign n38793 = ( n1995 & ~n6506 ) | ( n1995 & n15876 ) | ( ~n6506 & n15876 ) ;
  assign n38794 = n4807 | n21833 ;
  assign n38795 = n12939 & n38794 ;
  assign n38796 = n25798 | n35559 ;
  assign n38797 = n19917 | n32619 ;
  assign n38798 = n38796 & ~n38797 ;
  assign n38799 = n17683 | n18465 ;
  assign n38800 = n36816 ^ n9189 ^ 1'b0 ;
  assign n38801 = ~n17259 & n38800 ;
  assign n38802 = n29491 ^ n11366 ^ n8116 ;
  assign n38803 = n38802 ^ n33984 ^ 1'b0 ;
  assign n38804 = ( n13700 & n18503 ) | ( n13700 & ~n38803 ) | ( n18503 & ~n38803 ) ;
  assign n38805 = ( n4832 & ~n10461 ) | ( n4832 & n25223 ) | ( ~n10461 & n25223 ) ;
  assign n38806 = n2527 & n27573 ;
  assign n38807 = ( n31937 & ~n38805 ) | ( n31937 & n38806 ) | ( ~n38805 & n38806 ) ;
  assign n38808 = n8317 & n29518 ;
  assign n38809 = ~n17394 & n38808 ;
  assign n38810 = ( n1618 & n15132 ) | ( n1618 & n38809 ) | ( n15132 & n38809 ) ;
  assign n38811 = n20603 ^ n9917 ^ n2966 ;
  assign n38812 = n38811 ^ n1176 ^ 1'b0 ;
  assign n38813 = n24778 & n38812 ;
  assign n38814 = ( ~n34949 & n38810 ) | ( ~n34949 & n38813 ) | ( n38810 & n38813 ) ;
  assign n38815 = n3150 & n17626 ;
  assign n38816 = n38815 ^ x197 ^ 1'b0 ;
  assign n38817 = n38816 ^ n33207 ^ 1'b0 ;
  assign n38818 = n31831 & n38817 ;
  assign n38819 = n14104 ^ n13146 ^ 1'b0 ;
  assign n38820 = n14043 | n38819 ;
  assign n38821 = n21221 | n38820 ;
  assign n38822 = n7968 & ~n29206 ;
  assign n38823 = n18144 | n18627 ;
  assign n38824 = n38823 ^ n14037 ^ 1'b0 ;
  assign n38825 = n10168 & n35701 ;
  assign n38826 = ( n27695 & ~n38824 ) | ( n27695 & n38825 ) | ( ~n38824 & n38825 ) ;
  assign n38827 = n19230 ^ n5577 ^ 1'b0 ;
  assign n38828 = n36376 ^ n34484 ^ n4050 ;
  assign n38829 = ~n13050 & n20180 ;
  assign n38830 = n21526 & ~n38371 ;
  assign n38833 = n11563 & n25677 ;
  assign n38834 = n12415 & n38833 ;
  assign n38831 = ~n12663 & n34907 ;
  assign n38832 = n23617 & n38831 ;
  assign n38835 = n38834 ^ n38832 ^ 1'b0 ;
  assign n38836 = n20545 ^ n2431 ^ 1'b0 ;
  assign n38837 = n7416 & ~n22831 ;
  assign n38838 = n6129 & n38837 ;
  assign n38839 = n15540 | n18037 ;
  assign n38840 = n2592 ^ n2329 ^ 1'b0 ;
  assign n38841 = n29267 ^ n10082 ^ 1'b0 ;
  assign n38842 = ~n38840 & n38841 ;
  assign n38843 = n14916 ^ n13839 ^ 1'b0 ;
  assign n38844 = n10092 ^ n5752 ^ 1'b0 ;
  assign n38847 = n22930 ^ n21303 ^ 1'b0 ;
  assign n38848 = ( n6117 & n10873 ) | ( n6117 & n38847 ) | ( n10873 & n38847 ) ;
  assign n38845 = n14137 ^ n8969 ^ 1'b0 ;
  assign n38846 = n6411 | n38845 ;
  assign n38849 = n38848 ^ n38846 ^ n3672 ;
  assign n38850 = ~n4771 & n10942 ;
  assign n38851 = n16945 | n38850 ;
  assign n38852 = n38851 ^ n15831 ^ 1'b0 ;
  assign n38853 = n26030 ^ n17483 ^ 1'b0 ;
  assign n38855 = ~n8962 & n10922 ;
  assign n38854 = n10454 | n15951 ;
  assign n38856 = n38855 ^ n38854 ^ 1'b0 ;
  assign n38857 = n37666 ^ n14988 ^ 1'b0 ;
  assign n38858 = n18687 ^ n6879 ^ 1'b0 ;
  assign n38859 = n27007 | n38858 ;
  assign n38860 = n36101 ^ n26599 ^ n11871 ;
  assign n38861 = n13757 & n26811 ;
  assign n38862 = n38861 ^ n22381 ^ 1'b0 ;
  assign n38863 = n7190 & n7345 ;
  assign n38864 = ~n9186 & n38863 ;
  assign n38865 = ~n33663 & n38864 ;
  assign n38866 = ~n922 & n9610 ;
  assign n38867 = n28190 ^ n3483 ^ n2228 ;
  assign n38868 = n15477 & ~n38867 ;
  assign n38869 = n38866 & n38868 ;
  assign n38870 = n18025 ^ n8692 ^ 1'b0 ;
  assign n38871 = n35541 & n38870 ;
  assign n38872 = n18866 | n23476 ;
  assign n38873 = n3674 | n38872 ;
  assign n38874 = n4329 | n9507 ;
  assign n38875 = n32097 & ~n38874 ;
  assign n38876 = n21677 | n38875 ;
  assign n38877 = ( n7613 & n11530 ) | ( n7613 & ~n17516 ) | ( n11530 & ~n17516 ) ;
  assign n38878 = n18380 & ~n38877 ;
  assign n38879 = ~n3547 & n38878 ;
  assign n38880 = n18402 ^ n9273 ^ 1'b0 ;
  assign n38881 = n9399 & n38880 ;
  assign n38882 = ( n38876 & ~n38879 ) | ( n38876 & n38881 ) | ( ~n38879 & n38881 ) ;
  assign n38883 = n15180 ^ n6051 ^ 1'b0 ;
  assign n38884 = n16103 ^ n7680 ^ 1'b0 ;
  assign n38885 = n38884 ^ n37600 ^ n31723 ;
  assign n38886 = n6356 & n10602 ;
  assign n38887 = ~n2943 & n4950 ;
  assign n38888 = ~n38886 & n38887 ;
  assign n38889 = n6913 & n20096 ;
  assign n38890 = n38888 & n38889 ;
  assign n38891 = n4457 & ~n17674 ;
  assign n38892 = n38891 ^ n1090 ^ 1'b0 ;
  assign n38893 = n20726 ^ n260 ^ 1'b0 ;
  assign n38894 = n10470 & n38893 ;
  assign n38895 = n38894 ^ n33543 ^ n29681 ;
  assign n38896 = n9827 ^ n3071 ^ 1'b0 ;
  assign n38899 = n11097 & n24476 ;
  assign n38897 = ~n12196 & n35154 ;
  assign n38898 = ~n13538 & n38897 ;
  assign n38900 = n38899 ^ n38898 ^ n9266 ;
  assign n38901 = n11446 & ~n13402 ;
  assign n38902 = n38901 ^ n9574 ^ 1'b0 ;
  assign n38904 = n7335 & ~n20693 ;
  assign n38903 = n10279 ^ n308 ^ x90 ;
  assign n38905 = n38904 ^ n38903 ^ n17497 ;
  assign n38906 = ~n8894 & n23012 ;
  assign n38907 = n6118 ^ n898 ^ 1'b0 ;
  assign n38908 = n38907 ^ n4604 ^ n1958 ;
  assign n38909 = n38906 | n38908 ;
  assign n38910 = n13040 ^ n6410 ^ 1'b0 ;
  assign n38911 = n25127 & ~n38910 ;
  assign n38912 = n38911 ^ n4373 ^ 1'b0 ;
  assign n38913 = ( n2841 & n38909 ) | ( n2841 & ~n38912 ) | ( n38909 & ~n38912 ) ;
  assign n38914 = n2606 & n22149 ;
  assign n38915 = ~n9764 & n38914 ;
  assign n38916 = n38915 ^ n35746 ^ 1'b0 ;
  assign n38917 = n23909 ^ n12723 ^ n3409 ;
  assign n38918 = n38917 ^ n30627 ^ 1'b0 ;
  assign n38919 = n18631 | n38918 ;
  assign n38920 = n27747 ^ n10431 ^ 1'b0 ;
  assign n38928 = n29763 ^ n8429 ^ 1'b0 ;
  assign n38921 = ~n733 & n3019 ;
  assign n38922 = n38921 ^ n35823 ^ 1'b0 ;
  assign n38923 = ~n706 & n3837 ;
  assign n38924 = n38923 ^ n8920 ^ 1'b0 ;
  assign n38925 = n38924 ^ n32654 ^ 1'b0 ;
  assign n38926 = n292 & n38925 ;
  assign n38927 = ( n3180 & n38922 ) | ( n3180 & n38926 ) | ( n38922 & n38926 ) ;
  assign n38929 = n38928 ^ n38927 ^ 1'b0 ;
  assign n38930 = n37562 ^ n33228 ^ 1'b0 ;
  assign n38931 = ~n24817 & n35782 ;
  assign n38932 = n38931 ^ n14365 ^ 1'b0 ;
  assign n38933 = ~n15853 & n38932 ;
  assign n38934 = n25781 ^ n20844 ^ 1'b0 ;
  assign n38935 = n8255 & n38934 ;
  assign n38936 = n9018 & ~n38935 ;
  assign n38937 = n2133 & ~n21759 ;
  assign n38938 = ~n28693 & n38937 ;
  assign n38939 = n28143 ^ n22824 ^ n694 ;
  assign n38944 = ( n2336 & ~n2940 ) | ( n2336 & n19138 ) | ( ~n2940 & n19138 ) ;
  assign n38942 = n2820 & ~n12621 ;
  assign n38943 = n38942 ^ n15334 ^ 1'b0 ;
  assign n38940 = ( n15949 & ~n23703 ) | ( n15949 & n32233 ) | ( ~n23703 & n32233 ) ;
  assign n38941 = ( n15710 & n34836 ) | ( n15710 & n38940 ) | ( n34836 & n38940 ) ;
  assign n38945 = n38944 ^ n38943 ^ n38941 ;
  assign n38946 = n6344 & n35056 ;
  assign n38947 = ~n20050 & n26126 ;
  assign n38948 = n24666 ^ n717 ^ 1'b0 ;
  assign n38949 = ( n8828 & n11684 ) | ( n8828 & n35807 ) | ( n11684 & n35807 ) ;
  assign n38950 = n10710 & ~n38949 ;
  assign n38951 = n23324 ^ n7252 ^ 1'b0 ;
  assign n38952 = n2516 & ~n24750 ;
  assign n38953 = ~n5659 & n38952 ;
  assign n38954 = n38953 ^ n31093 ^ 1'b0 ;
  assign n38958 = n7195 & ~n27270 ;
  assign n38956 = n649 | n17740 ;
  assign n38957 = n38956 ^ n30037 ^ 1'b0 ;
  assign n38955 = n31939 ^ n11973 ^ 1'b0 ;
  assign n38959 = n38958 ^ n38957 ^ n38955 ;
  assign n38960 = ( n4090 & ~n28902 ) | ( n4090 & n36484 ) | ( ~n28902 & n36484 ) ;
  assign n38961 = n23973 ^ n23117 ^ n19004 ;
  assign n38963 = ~n12072 & n28719 ;
  assign n38962 = n12338 & n24746 ;
  assign n38964 = n38963 ^ n38962 ^ 1'b0 ;
  assign n38965 = n16038 & ~n18646 ;
  assign n38966 = ~n8484 & n33224 ;
  assign n38967 = ~n38965 & n38966 ;
  assign n38968 = ( n31389 & n38964 ) | ( n31389 & ~n38967 ) | ( n38964 & ~n38967 ) ;
  assign n38969 = n35772 ^ n3492 ^ 1'b0 ;
  assign n38970 = n34906 & n37478 ;
  assign n38971 = n3020 & ~n29985 ;
  assign n38972 = n22497 & n38971 ;
  assign n38973 = ~n9969 & n28199 ;
  assign n38974 = n38973 ^ n854 ^ 1'b0 ;
  assign n38975 = ~n1451 & n7457 ;
  assign n38976 = n22201 & ~n38975 ;
  assign n38977 = n38976 ^ n987 ^ 1'b0 ;
  assign n38978 = ( n10961 & n12174 ) | ( n10961 & ~n26887 ) | ( n12174 & ~n26887 ) ;
  assign n38979 = n38978 ^ n5707 ^ 1'b0 ;
  assign n38980 = ~n38977 & n38979 ;
  assign n38981 = ~n5155 & n38980 ;
  assign n38982 = n38974 & n38981 ;
  assign n38984 = n21856 ^ n8798 ^ 1'b0 ;
  assign n38983 = n11401 & ~n38762 ;
  assign n38985 = n38984 ^ n38983 ^ 1'b0 ;
  assign n38986 = ~n6221 & n38985 ;
  assign n38987 = n1576 | n16828 ;
  assign n38988 = n16795 & ~n38987 ;
  assign n38989 = n15714 & ~n17300 ;
  assign n38990 = n37257 | n38099 ;
  assign n38991 = n15208 ^ n14000 ^ x198 ;
  assign n38993 = ~n7032 & n29763 ;
  assign n38994 = n2794 & n38993 ;
  assign n38992 = n31953 & ~n33311 ;
  assign n38995 = n38994 ^ n38992 ^ 1'b0 ;
  assign n38996 = ~n7897 & n13630 ;
  assign n38997 = n38996 ^ n37912 ^ n19144 ;
  assign n38998 = ~n13382 & n26448 ;
  assign n38999 = n38997 & n38998 ;
  assign n39000 = n3496 & ~n4547 ;
  assign n39001 = ~n4948 & n39000 ;
  assign n39002 = n3538 & n10805 ;
  assign n39003 = ( n7790 & n39001 ) | ( n7790 & ~n39002 ) | ( n39001 & ~n39002 ) ;
  assign n39004 = n39003 ^ n13587 ^ 1'b0 ;
  assign n39005 = n28386 ^ n8629 ^ 1'b0 ;
  assign n39006 = n39004 | n39005 ;
  assign n39007 = n7840 & n20369 ;
  assign n39008 = n23688 & n39007 ;
  assign n39009 = ( n1939 & n5377 ) | ( n1939 & ~n39008 ) | ( n5377 & ~n39008 ) ;
  assign n39010 = n13766 ^ n7760 ^ 1'b0 ;
  assign n39011 = n10602 & ~n39010 ;
  assign n39012 = n39011 ^ n17279 ^ 1'b0 ;
  assign n39013 = n21995 ^ n6494 ^ 1'b0 ;
  assign n39014 = ( n3932 & ~n23822 ) | ( n3932 & n39013 ) | ( ~n23822 & n39013 ) ;
  assign n39015 = n39014 ^ n37575 ^ 1'b0 ;
  assign n39016 = n29846 ^ n9008 ^ 1'b0 ;
  assign n39017 = ~n5837 & n30550 ;
  assign n39018 = n39016 & n39017 ;
  assign n39019 = ~n5073 & n34859 ;
  assign n39020 = ( n5565 & n10192 ) | ( n5565 & n24174 ) | ( n10192 & n24174 ) ;
  assign n39021 = n39020 ^ n10064 ^ 1'b0 ;
  assign n39022 = n9308 | n12284 ;
  assign n39023 = n39021 | n39022 ;
  assign n39024 = n24430 ^ n16191 ^ n7886 ;
  assign n39025 = n39023 & n39024 ;
  assign n39026 = ( n1141 & n3475 ) | ( n1141 & ~n25700 ) | ( n3475 & ~n25700 ) ;
  assign n39027 = n33428 ^ n12296 ^ 1'b0 ;
  assign n39028 = ~n32571 & n34604 ;
  assign n39029 = ~n1103 & n12671 ;
  assign n39030 = n33653 ^ n31044 ^ 1'b0 ;
  assign n39033 = x172 & n9608 ;
  assign n39031 = n9721 ^ n4282 ^ 1'b0 ;
  assign n39032 = ~n11064 & n39031 ;
  assign n39034 = n39033 ^ n39032 ^ n14527 ;
  assign n39035 = n13591 | n36547 ;
  assign n39036 = n21724 ^ n986 ^ 1'b0 ;
  assign n39037 = n39036 ^ n3865 ^ 1'b0 ;
  assign n39038 = n13106 | n39037 ;
  assign n39039 = n4932 ^ n4561 ^ 1'b0 ;
  assign n39040 = n39039 ^ n1674 ^ 1'b0 ;
  assign n39041 = ~n4190 & n39040 ;
  assign n39042 = ~n3715 & n39041 ;
  assign n39043 = n39042 ^ n22703 ^ 1'b0 ;
  assign n39044 = ~n6066 & n16311 ;
  assign n39045 = n19524 & n39044 ;
  assign n39046 = n39045 ^ n14621 ^ 1'b0 ;
  assign n39047 = n8343 & n39046 ;
  assign n39048 = ~n4255 & n7978 ;
  assign n39049 = n3997 & n39048 ;
  assign n39050 = n39049 ^ n4153 ^ 1'b0 ;
  assign n39051 = n39050 ^ n5588 ^ 1'b0 ;
  assign n39052 = ~n14235 & n39051 ;
  assign n39053 = n11959 & n31631 ;
  assign n39054 = n39053 ^ n29990 ^ 1'b0 ;
  assign n39055 = n18586 ^ n16926 ^ 1'b0 ;
  assign n39056 = n7257 | n39055 ;
  assign n39057 = n39056 ^ n2642 ^ 1'b0 ;
  assign n39058 = ~n5204 & n27217 ;
  assign n39059 = n7444 & n39058 ;
  assign n39060 = n22969 & ~n39059 ;
  assign n39061 = n17422 ^ n3353 ^ 1'b0 ;
  assign n39062 = ~n30454 & n39061 ;
  assign n39063 = n1190 & ~n33757 ;
  assign n39064 = n39063 ^ n22907 ^ n13050 ;
  assign n39065 = n39062 & n39064 ;
  assign n39066 = ( ~n18694 & n39060 ) | ( ~n18694 & n39065 ) | ( n39060 & n39065 ) ;
  assign n39067 = ~n24089 & n25605 ;
  assign n39068 = n2879 ^ n2294 ^ 1'b0 ;
  assign n39069 = n31764 & ~n39068 ;
  assign n39070 = n39069 ^ n13804 ^ 1'b0 ;
  assign n39071 = ~n3905 & n29987 ;
  assign n39072 = n2256 | n7532 ;
  assign n39073 = n39072 ^ n2162 ^ 1'b0 ;
  assign n39074 = n21379 & ~n34379 ;
  assign n39075 = n39074 ^ n29916 ^ 1'b0 ;
  assign n39076 = ( n10076 & n24430 ) | ( n10076 & n39075 ) | ( n24430 & n39075 ) ;
  assign n39077 = ( n2056 & n21669 ) | ( n2056 & n27847 ) | ( n21669 & n27847 ) ;
  assign n39078 = n39077 ^ n38882 ^ 1'b0 ;
  assign n39079 = n37532 ^ n36291 ^ n2033 ;
  assign n39080 = n10450 ^ n5593 ^ 1'b0 ;
  assign n39081 = n14481 | n39080 ;
  assign n39082 = n1401 | n39081 ;
  assign n39083 = n39082 ^ n7729 ^ 1'b0 ;
  assign n39084 = n31989 ^ n26893 ^ n20925 ;
  assign n39085 = n21611 & ~n28825 ;
  assign n39086 = ~n3989 & n5722 ;
  assign n39087 = ~n10683 & n39086 ;
  assign n39088 = n4350 & ~n11202 ;
  assign n39089 = n39087 & n39088 ;
  assign n39090 = n39089 ^ n21842 ^ n8883 ;
  assign n39091 = n24356 ^ n14938 ^ 1'b0 ;
  assign n39092 = ~n8189 & n32367 ;
  assign n39093 = n39092 ^ n1318 ^ 1'b0 ;
  assign n39094 = n6132 & ~n26340 ;
  assign n39095 = n39094 ^ n2068 ^ 1'b0 ;
  assign n39096 = n12459 | n39095 ;
  assign n39097 = n30542 ^ n23604 ^ 1'b0 ;
  assign n39098 = n39096 & n39097 ;
  assign n39099 = n15687 | n16687 ;
  assign n39104 = n15826 ^ n7571 ^ 1'b0 ;
  assign n39103 = ~n12539 & n25595 ;
  assign n39105 = n39104 ^ n39103 ^ 1'b0 ;
  assign n39100 = n11566 | n37411 ;
  assign n39101 = n39100 ^ n24142 ^ 1'b0 ;
  assign n39102 = n39101 ^ n13881 ^ 1'b0 ;
  assign n39106 = n39105 ^ n39102 ^ 1'b0 ;
  assign n39111 = n18238 ^ n2672 ^ 1'b0 ;
  assign n39107 = n34605 ^ n22673 ^ 1'b0 ;
  assign n39108 = ~n6474 & n39107 ;
  assign n39109 = n31497 | n39108 ;
  assign n39110 = n8914 & n39109 ;
  assign n39112 = n39111 ^ n39110 ^ 1'b0 ;
  assign n39113 = n7108 & ~n37462 ;
  assign n39114 = n32679 ^ n6769 ^ n5595 ;
  assign n39115 = ~n15373 & n39114 ;
  assign n39116 = x127 & n6403 ;
  assign n39117 = ( n2403 & n3161 ) | ( n2403 & n31756 ) | ( n3161 & n31756 ) ;
  assign n39118 = n39117 ^ n37201 ^ 1'b0 ;
  assign n39119 = n9736 & ~n22425 ;
  assign n39120 = n39119 ^ n18476 ^ n16136 ;
  assign n39121 = n6793 | n24606 ;
  assign n39122 = n39121 ^ n15999 ^ 1'b0 ;
  assign n39123 = ~n7879 & n39122 ;
  assign n39124 = n18389 & ~n39123 ;
  assign n39125 = ( n4153 & ~n20911 ) | ( n4153 & n39124 ) | ( ~n20911 & n39124 ) ;
  assign n39126 = ~n16872 & n25220 ;
  assign n39127 = ~n13354 & n39126 ;
  assign n39128 = n39127 ^ n5146 ^ 1'b0 ;
  assign n39130 = n4797 | n4955 ;
  assign n39129 = n23370 & ~n32994 ;
  assign n39131 = n39130 ^ n39129 ^ 1'b0 ;
  assign n39132 = ( n33163 & ~n39128 ) | ( n33163 & n39131 ) | ( ~n39128 & n39131 ) ;
  assign n39133 = n14539 | n36463 ;
  assign n39134 = n1521 ^ n375 ^ 1'b0 ;
  assign n39135 = n20217 & ~n21857 ;
  assign n39136 = ~n39134 & n39135 ;
  assign n39137 = n34465 ^ n17108 ^ 1'b0 ;
  assign n39138 = n39136 | n39137 ;
  assign n39139 = n33541 ^ n27842 ^ n27225 ;
  assign n39140 = ~n2802 & n39139 ;
  assign n39141 = n30508 ^ n14897 ^ 1'b0 ;
  assign n39142 = n9853 & n16408 ;
  assign n39143 = ~n14121 & n39142 ;
  assign n39144 = n13850 ^ n5055 ^ 1'b0 ;
  assign n39145 = n16661 & ~n17223 ;
  assign n39146 = n39144 | n39145 ;
  assign n39147 = n3746 & n22161 ;
  assign n39148 = n9698 ^ n7097 ^ 1'b0 ;
  assign n39149 = ( n1260 & n2250 ) | ( n1260 & n26252 ) | ( n2250 & n26252 ) ;
  assign n39150 = n32914 | n39149 ;
  assign n39151 = ( ~n6992 & n14304 ) | ( ~n6992 & n26633 ) | ( n14304 & n26633 ) ;
  assign n39152 = n2844 & ~n2911 ;
  assign n39153 = n9705 & n39152 ;
  assign n39154 = ~n39152 & n39153 ;
  assign n39155 = n39154 ^ n9457 ^ n7512 ;
  assign n39156 = ~n1711 & n25135 ;
  assign n39157 = n535 & n39156 ;
  assign n39158 = n11684 | n13340 ;
  assign n39159 = n15588 | n39158 ;
  assign n39160 = ( ~x209 & n7265 ) | ( ~x209 & n7696 ) | ( n7265 & n7696 ) ;
  assign n39162 = n28044 ^ n19630 ^ 1'b0 ;
  assign n39161 = n14137 & n31852 ;
  assign n39163 = n39162 ^ n39161 ^ n26484 ;
  assign n39164 = n34616 ^ n28970 ^ x218 ;
  assign n39165 = ( n11285 & n18980 ) | ( n11285 & n39164 ) | ( n18980 & n39164 ) ;
  assign n39166 = n31345 ^ n11766 ^ 1'b0 ;
  assign n39167 = ~n28969 & n37588 ;
  assign n39168 = n39166 & n39167 ;
  assign n39169 = n28602 ^ n5042 ^ n2998 ;
  assign n39170 = ~n12391 & n39169 ;
  assign n39171 = ~n10288 & n39170 ;
  assign n39172 = n36286 ^ n34879 ^ 1'b0 ;
  assign n39173 = n13137 & n21551 ;
  assign n39174 = ~n17961 & n39173 ;
  assign n39175 = n5713 ^ n4473 ^ 1'b0 ;
  assign n39177 = n8733 & ~n22061 ;
  assign n39178 = n12495 & n39177 ;
  assign n39176 = n1650 & n2401 ;
  assign n39179 = n39178 ^ n39176 ^ 1'b0 ;
  assign n39180 = n16431 ^ n14063 ^ n8201 ;
  assign n39181 = ( x8 & ~n28881 ) | ( x8 & n39180 ) | ( ~n28881 & n39180 ) ;
  assign n39182 = n2119 & ~n4754 ;
  assign n39183 = ~x209 & n39182 ;
  assign n39184 = ( ~n6686 & n10474 ) | ( ~n6686 & n39183 ) | ( n10474 & n39183 ) ;
  assign n39187 = n35396 & n35886 ;
  assign n39185 = n33418 ^ n24740 ^ 1'b0 ;
  assign n39186 = ~n27707 & n39185 ;
  assign n39188 = n39187 ^ n39186 ^ 1'b0 ;
  assign n39189 = n11463 & ~n23197 ;
  assign n39190 = ~n9073 & n25302 ;
  assign n39191 = ~n35284 & n39190 ;
  assign n39192 = n6054 | n39191 ;
  assign n39193 = n19161 ^ n7466 ^ 1'b0 ;
  assign n39194 = n12412 & ~n39193 ;
  assign n39195 = n3698 & ~n4546 ;
  assign n39196 = n39195 ^ n6342 ^ 1'b0 ;
  assign n39197 = n5009 ^ x233 ^ 1'b0 ;
  assign n39198 = n5037 & n39197 ;
  assign n39199 = n39198 ^ n12657 ^ 1'b0 ;
  assign n39200 = ~n23394 & n39199 ;
  assign n39201 = n39200 ^ n837 ^ 1'b0 ;
  assign n39202 = n39196 | n39201 ;
  assign n39203 = n39194 | n39202 ;
  assign n39207 = ( n4957 & ~n11450 ) | ( n4957 & n13341 ) | ( ~n11450 & n13341 ) ;
  assign n39208 = n39207 ^ n6921 ^ 1'b0 ;
  assign n39204 = n29787 ^ n3854 ^ n1061 ;
  assign n39205 = n375 & n24060 ;
  assign n39206 = ~n39204 & n39205 ;
  assign n39209 = n39208 ^ n39206 ^ n8447 ;
  assign n39210 = n29518 ^ n22287 ^ n17866 ;
  assign n39211 = n10687 ^ n7011 ^ 1'b0 ;
  assign n39212 = n39211 ^ n26115 ^ 1'b0 ;
  assign n39213 = n13618 ^ n1387 ^ 1'b0 ;
  assign n39214 = ~n6789 & n24713 ;
  assign n39215 = n16858 & ~n29335 ;
  assign n39216 = n39215 ^ n26513 ^ 1'b0 ;
  assign n39217 = ~n10009 & n16454 ;
  assign n39218 = n39217 ^ n6320 ^ 1'b0 ;
  assign n39219 = n11174 ^ n9525 ^ 1'b0 ;
  assign n39220 = n38517 | n39219 ;
  assign n39221 = ~n13201 & n23777 ;
  assign n39222 = n8843 & n39221 ;
  assign n39223 = n39222 ^ n1064 ^ 1'b0 ;
  assign n39224 = n39223 ^ n18706 ^ 1'b0 ;
  assign n39225 = n27246 ^ n5146 ^ n1392 ;
  assign n39226 = n39225 ^ n35290 ^ 1'b0 ;
  assign n39227 = n39226 ^ n10959 ^ 1'b0 ;
  assign n39228 = ( n13879 & n39224 ) | ( n13879 & ~n39227 ) | ( n39224 & ~n39227 ) ;
  assign n39229 = ~n32629 & n39228 ;
  assign n39230 = ~n9757 & n39229 ;
  assign n39231 = ~n21793 & n32626 ;
  assign n39232 = n16466 ^ n6969 ^ 1'b0 ;
  assign n39234 = n10195 ^ n6725 ^ 1'b0 ;
  assign n39235 = ~n16031 & n39234 ;
  assign n39236 = n8590 & n39235 ;
  assign n39233 = ~n13429 & n28897 ;
  assign n39237 = n39236 ^ n39233 ^ 1'b0 ;
  assign n39239 = n9922 | n36421 ;
  assign n39238 = x140 & ~n7440 ;
  assign n39240 = n39239 ^ n39238 ^ 1'b0 ;
  assign n39241 = n39240 ^ n26908 ^ 1'b0 ;
  assign n39242 = n35173 & n39241 ;
  assign n39243 = ( ~n17411 & n28825 ) | ( ~n17411 & n38684 ) | ( n28825 & n38684 ) ;
  assign n39247 = n10124 ^ n7517 ^ n4049 ;
  assign n39248 = n3146 & ~n39247 ;
  assign n39249 = n39248 ^ n13407 ^ 1'b0 ;
  assign n39244 = n7439 | n12792 ;
  assign n39245 = n39244 ^ n5963 ^ 1'b0 ;
  assign n39246 = ( ~n3212 & n11457 ) | ( ~n3212 & n39245 ) | ( n11457 & n39245 ) ;
  assign n39250 = n39249 ^ n39246 ^ n29905 ;
  assign n39251 = ( ~n10757 & n11759 ) | ( ~n10757 & n30454 ) | ( n11759 & n30454 ) ;
  assign n39252 = n33643 ^ n33227 ^ 1'b0 ;
  assign n39253 = n39251 | n39252 ;
  assign n39254 = n3335 | n39253 ;
  assign n39255 = n11445 & ~n39254 ;
  assign n39256 = n8384 & ~n39255 ;
  assign n39257 = n39256 ^ n8531 ^ 1'b0 ;
  assign n39258 = n8551 ^ n5670 ^ n5077 ;
  assign n39259 = n7030 & ~n39258 ;
  assign n39260 = n3370 ^ x198 ^ 1'b0 ;
  assign n39261 = n20640 & ~n39260 ;
  assign n39262 = ~n1378 & n39261 ;
  assign n39263 = ~n33263 & n39262 ;
  assign n39265 = n30130 ^ n13762 ^ 1'b0 ;
  assign n39266 = n11173 & ~n39265 ;
  assign n39264 = ( x57 & n2201 ) | ( x57 & ~n14641 ) | ( n2201 & ~n14641 ) ;
  assign n39267 = n39266 ^ n39264 ^ n18334 ;
  assign n39271 = ~n992 & n11187 ;
  assign n39272 = n39271 ^ n6773 ^ 1'b0 ;
  assign n39273 = n34757 & n39272 ;
  assign n39274 = n17614 & ~n39273 ;
  assign n39275 = ~n18425 & n39274 ;
  assign n39268 = ~n774 & n3722 ;
  assign n39269 = n15838 | n39268 ;
  assign n39270 = n39269 ^ n2724 ^ 1'b0 ;
  assign n39276 = n39275 ^ n39270 ^ n29101 ;
  assign n39277 = n9000 ^ n1176 ^ 1'b0 ;
  assign n39278 = n21360 & ~n39277 ;
  assign n39279 = n21126 ^ n9872 ^ 1'b0 ;
  assign n39280 = ( ~n8165 & n11946 ) | ( ~n8165 & n39279 ) | ( n11946 & n39279 ) ;
  assign n39281 = n34922 ^ n27991 ^ n10061 ;
  assign n39282 = n7240 ^ n5573 ^ 1'b0 ;
  assign n39283 = ~n2847 & n39282 ;
  assign n39284 = ~n39281 & n39283 ;
  assign n39285 = n39284 ^ n28305 ^ 1'b0 ;
  assign n39286 = n20755 ^ n1701 ^ 1'b0 ;
  assign n39287 = n20461 | n39286 ;
  assign n39288 = n18297 ^ n12700 ^ 1'b0 ;
  assign n39289 = n604 | n39288 ;
  assign n39290 = n1542 & n10816 ;
  assign n39291 = n26599 ^ n16637 ^ n16034 ;
  assign n39292 = n39291 ^ n24934 ^ 1'b0 ;
  assign n39293 = n39290 | n39292 ;
  assign n39294 = n3294 & n11104 ;
  assign n39295 = ~n39293 & n39294 ;
  assign n39296 = n2452 & n25120 ;
  assign n39297 = n23914 ^ n10028 ^ n3476 ;
  assign n39298 = n17063 | n25215 ;
  assign n39299 = n39297 & ~n39298 ;
  assign n39300 = n39299 ^ n20553 ^ 1'b0 ;
  assign n39301 = n8329 & ~n39300 ;
  assign n39302 = n35885 ^ n35493 ^ n20936 ;
  assign n39303 = n12901 & ~n16593 ;
  assign n39304 = n39303 ^ n38904 ^ n24083 ;
  assign n39305 = n11303 ^ n818 ^ 1'b0 ;
  assign n39306 = ~n7745 & n39305 ;
  assign n39307 = ( n18365 & ~n22872 ) | ( n18365 & n39306 ) | ( ~n22872 & n39306 ) ;
  assign n39308 = ( n8481 & n10654 ) | ( n8481 & ~n23201 ) | ( n10654 & ~n23201 ) ;
  assign n39309 = n17541 ^ n9206 ^ n1043 ;
  assign n39310 = n39309 ^ n19812 ^ 1'b0 ;
  assign n39311 = ~n12260 & n39310 ;
  assign n39312 = ~n39308 & n39311 ;
  assign n39315 = ( n860 & n1584 ) | ( n860 & ~n34552 ) | ( n1584 & ~n34552 ) ;
  assign n39313 = n9814 & n28094 ;
  assign n39314 = n29559 | n39313 ;
  assign n39316 = n39315 ^ n39314 ^ 1'b0 ;
  assign n39317 = n9224 & n14328 ;
  assign n39318 = n14053 & n39317 ;
  assign n39319 = n19900 ^ n16142 ^ 1'b0 ;
  assign n39320 = n13937 | n32552 ;
  assign n39321 = x150 | n39320 ;
  assign n39322 = n39321 ^ n34241 ^ n21303 ;
  assign n39323 = n39322 ^ n17984 ^ 1'b0 ;
  assign n39325 = n16974 ^ n9444 ^ 1'b0 ;
  assign n39326 = n12607 | n39325 ;
  assign n39324 = n7979 & n36411 ;
  assign n39327 = n39326 ^ n39324 ^ 1'b0 ;
  assign n39328 = n3693 & n6958 ;
  assign n39329 = n9522 & n39328 ;
  assign n39330 = n13284 | n39329 ;
  assign n39331 = n2643 & ~n4330 ;
  assign n39332 = n39331 ^ n12485 ^ 1'b0 ;
  assign n39333 = ( ~n2921 & n19874 ) | ( ~n2921 & n36140 ) | ( n19874 & n36140 ) ;
  assign n39334 = ( x141 & ~n27068 ) | ( x141 & n39333 ) | ( ~n27068 & n39333 ) ;
  assign n39335 = ( n4752 & n28912 ) | ( n4752 & ~n39334 ) | ( n28912 & ~n39334 ) ;
  assign n39336 = n9124 ^ n6183 ^ 1'b0 ;
  assign n39337 = n39336 ^ n5322 ^ n4989 ;
  assign n39338 = ~n5415 & n17626 ;
  assign n39339 = n20098 & n39338 ;
  assign n39340 = ( ~n13082 & n35008 ) | ( ~n13082 & n39339 ) | ( n35008 & n39339 ) ;
  assign n39341 = ( n36744 & n39337 ) | ( n36744 & n39340 ) | ( n39337 & n39340 ) ;
  assign n39342 = n29843 & n33271 ;
  assign n39343 = n39342 ^ n21773 ^ 1'b0 ;
  assign n39344 = n16757 ^ n13878 ^ n5978 ;
  assign n39345 = ~n14482 & n39344 ;
  assign n39346 = n39345 ^ n11450 ^ 1'b0 ;
  assign n39347 = n32957 ^ n2302 ^ 1'b0 ;
  assign n39348 = ( n14632 & ~n17091 ) | ( n14632 & n23064 ) | ( ~n17091 & n23064 ) ;
  assign n39349 = n39348 ^ n9630 ^ 1'b0 ;
  assign n39350 = n38012 | n39349 ;
  assign n39351 = n27761 ^ n17387 ^ 1'b0 ;
  assign n39354 = n26130 ^ n509 ^ 1'b0 ;
  assign n39353 = n10449 ^ x30 ^ 1'b0 ;
  assign n39352 = n24986 ^ n1778 ^ 1'b0 ;
  assign n39355 = n39354 ^ n39353 ^ n39352 ;
  assign n39356 = n25851 & ~n39355 ;
  assign n39358 = ~n2433 & n19828 ;
  assign n39359 = n23807 & n39358 ;
  assign n39357 = n34330 ^ n26867 ^ n1791 ;
  assign n39360 = n39359 ^ n39357 ^ n29048 ;
  assign n39361 = n23784 ^ n15110 ^ 1'b0 ;
  assign n39362 = ~n25214 & n38195 ;
  assign n39363 = n8552 & n20403 ;
  assign n39364 = n39363 ^ n14958 ^ 1'b0 ;
  assign n39365 = n30071 & ~n39364 ;
  assign n39366 = n17475 & n39365 ;
  assign n39367 = ~n22118 & n39366 ;
  assign n39368 = n6797 ^ n1343 ^ 1'b0 ;
  assign n39369 = n39368 ^ n6271 ^ n5197 ;
  assign n39370 = n20367 & ~n39369 ;
  assign n39371 = n39370 ^ n7957 ^ 1'b0 ;
  assign n39372 = ~n22219 & n34003 ;
  assign n39373 = n39372 ^ n39353 ^ 1'b0 ;
  assign n39374 = n12863 & ~n39373 ;
  assign n39375 = n36327 ^ n33271 ^ 1'b0 ;
  assign n39376 = n26233 ^ n25494 ^ 1'b0 ;
  assign n39377 = n27251 | n39376 ;
  assign n39378 = n8624 & ~n38316 ;
  assign n39379 = n19216 & n39378 ;
  assign n39380 = ~n17068 & n32149 ;
  assign n39382 = n16993 | n17050 ;
  assign n39381 = n17324 | n26916 ;
  assign n39383 = n39382 ^ n39381 ^ 1'b0 ;
  assign n39384 = n16997 ^ n2734 ^ 1'b0 ;
  assign n39385 = ~n25850 & n39384 ;
  assign n39386 = ~n26587 & n39385 ;
  assign n39387 = ( ~n9467 & n14397 ) | ( ~n9467 & n31778 ) | ( n14397 & n31778 ) ;
  assign n39388 = n18163 | n30427 ;
  assign n39389 = n29248 ^ n5936 ^ 1'b0 ;
  assign n39390 = n39388 & ~n39389 ;
  assign n39391 = n10510 & ~n24753 ;
  assign n39392 = n39391 ^ n12423 ^ 1'b0 ;
  assign n39393 = x71 & ~n31089 ;
  assign n39394 = n39393 ^ n24615 ^ 1'b0 ;
  assign n39395 = n25117 & ~n39394 ;
  assign n39396 = n10279 | n21676 ;
  assign n39397 = ~n18139 & n38275 ;
  assign n39398 = n39397 ^ n9520 ^ 1'b0 ;
  assign n39399 = n1067 & ~n39398 ;
  assign n39400 = n15530 & ~n39399 ;
  assign n39401 = n16725 & n39400 ;
  assign n39402 = n31087 ^ n16997 ^ 1'b0 ;
  assign n39403 = n7976 & ~n39402 ;
  assign n39404 = n24860 ^ n932 ^ 1'b0 ;
  assign n39405 = n22771 & ~n36748 ;
  assign n39406 = ~x132 & n39405 ;
  assign n39407 = ( n1258 & ~n21404 ) | ( n1258 & n39406 ) | ( ~n21404 & n39406 ) ;
  assign n39408 = n25327 ^ n25106 ^ n14781 ;
  assign n39409 = n22923 ^ n17570 ^ 1'b0 ;
  assign n39410 = n38735 ^ n4034 ^ 1'b0 ;
  assign n39411 = n31101 | n39410 ;
  assign n39412 = n37500 ^ n7944 ^ 1'b0 ;
  assign n39413 = x52 & n39412 ;
  assign n39414 = ~n9949 & n14953 ;
  assign n39415 = n12903 & n39414 ;
  assign n39416 = n39415 ^ n20278 ^ 1'b0 ;
  assign n39417 = n12350 ^ n8806 ^ 1'b0 ;
  assign n39418 = ~n6782 & n39417 ;
  assign n39419 = ~n27885 & n39418 ;
  assign n39420 = ( n1450 & n6413 ) | ( n1450 & n13112 ) | ( n6413 & n13112 ) ;
  assign n39421 = n39420 ^ n1835 ^ 1'b0 ;
  assign n39422 = n4120 ^ n424 ^ 1'b0 ;
  assign n39423 = n11007 ^ n5984 ^ 1'b0 ;
  assign n39424 = n16992 | n39423 ;
  assign n39425 = n39422 & n39424 ;
  assign n39426 = n27933 ^ n5316 ^ 1'b0 ;
  assign n39427 = n39426 ^ n11112 ^ n10446 ;
  assign n39428 = n5844 & ~n7517 ;
  assign n39429 = n27094 & n39428 ;
  assign n39430 = n39429 ^ n3605 ^ 1'b0 ;
  assign n39431 = n10403 & ~n39430 ;
  assign n39432 = n8449 | n12416 ;
  assign n39433 = n39432 ^ n684 ^ 1'b0 ;
  assign n39434 = n37089 | n39433 ;
  assign n39435 = n37256 ^ n19875 ^ 1'b0 ;
  assign n39436 = n2005 & n14275 ;
  assign n39437 = n14465 & n39436 ;
  assign n39438 = n27958 ^ n9881 ^ 1'b0 ;
  assign n39439 = n32895 ^ n31687 ^ n9853 ;
  assign n39440 = n39439 ^ n23092 ^ n11844 ;
  assign n39441 = ~n1388 & n32679 ;
  assign n39442 = ( n11657 & n17737 ) | ( n11657 & ~n22676 ) | ( n17737 & ~n22676 ) ;
  assign n39443 = n13354 ^ n1118 ^ n384 ;
  assign n39444 = n17194 | n39443 ;
  assign n39445 = n39444 ^ n22099 ^ 1'b0 ;
  assign n39446 = n5481 | n26666 ;
  assign n39447 = ~n4734 & n10899 ;
  assign n39448 = ~n27666 & n39447 ;
  assign n39449 = ~n20595 & n35548 ;
  assign n39450 = n13925 & n39449 ;
  assign n39451 = n35175 ^ n28292 ^ n953 ;
  assign n39452 = n20900 ^ n13359 ^ 1'b0 ;
  assign n39453 = ~n13700 & n30956 ;
  assign n39454 = ~n27550 & n39453 ;
  assign n39455 = n39452 & n39454 ;
  assign n39456 = ( n13877 & n28331 ) | ( n13877 & n39455 ) | ( n28331 & n39455 ) ;
  assign n39457 = n11805 & n18597 ;
  assign n39458 = n39457 ^ n24232 ^ 1'b0 ;
  assign n39459 = ~n13310 & n39458 ;
  assign n39460 = n39459 ^ n8150 ^ 1'b0 ;
  assign n39461 = n2308 & ~n39460 ;
  assign n39462 = n39461 ^ n1781 ^ 1'b0 ;
  assign n39463 = n11063 & ~n11854 ;
  assign n39464 = ~n7486 & n39463 ;
  assign n39465 = n28437 ^ n7934 ^ 1'b0 ;
  assign n39466 = ~n17877 & n24263 ;
  assign n39467 = ~n39465 & n39466 ;
  assign n39468 = n30742 ^ n28559 ^ n26996 ;
  assign n39469 = ( x109 & n12674 ) | ( x109 & ~n25057 ) | ( n12674 & ~n25057 ) ;
  assign n39470 = ~n4221 & n32469 ;
  assign n39471 = ( n8167 & n11022 ) | ( n8167 & n13365 ) | ( n11022 & n13365 ) ;
  assign n39472 = ~n5798 & n13172 ;
  assign n39473 = n39472 ^ n9685 ^ 1'b0 ;
  assign n39474 = n33599 & ~n39473 ;
  assign n39475 = n37748 ^ n14424 ^ n9273 ;
  assign n39476 = n12080 ^ n6770 ^ 1'b0 ;
  assign n39477 = n29168 ^ n11165 ^ n4690 ;
  assign n39478 = n39477 ^ n33942 ^ n33380 ;
  assign n39479 = n317 & n3130 ;
  assign n39480 = n18025 ^ n1224 ^ 1'b0 ;
  assign n39481 = n39479 | n39480 ;
  assign n39482 = x226 & n35947 ;
  assign n39483 = ~n20724 & n39482 ;
  assign n39484 = n10971 | n28730 ;
  assign n39488 = ~n27297 & n28312 ;
  assign n39485 = n474 & ~n35972 ;
  assign n39486 = n9773 & n39485 ;
  assign n39487 = n35198 & ~n39486 ;
  assign n39489 = n39488 ^ n39487 ^ 1'b0 ;
  assign n39490 = n5165 | n32691 ;
  assign n39491 = n39490 ^ n9757 ^ 1'b0 ;
  assign n39492 = n38875 & ~n39491 ;
  assign n39495 = ( n13129 & ~n17825 ) | ( n13129 & n23239 ) | ( ~n17825 & n23239 ) ;
  assign n39493 = ~n6892 & n24476 ;
  assign n39494 = n39493 ^ n22154 ^ 1'b0 ;
  assign n39496 = n39495 ^ n39494 ^ n316 ;
  assign n39497 = ( n8207 & ~n13833 ) | ( n8207 & n17841 ) | ( ~n13833 & n17841 ) ;
  assign n39498 = n33967 ^ n2722 ^ 1'b0 ;
  assign n39499 = n12227 ^ n1576 ^ 1'b0 ;
  assign n39500 = n8286 | n39499 ;
  assign n39501 = n26796 | n39500 ;
  assign n39502 = n6109 & ~n25372 ;
  assign n39503 = n3983 & n39502 ;
  assign n39504 = n29723 ^ n19295 ^ n10627 ;
  assign n39505 = n39504 ^ n21685 ^ n1243 ;
  assign n39506 = n2565 & ~n19364 ;
  assign n39507 = n39506 ^ n21381 ^ n20665 ;
  assign n39508 = n26871 | n33211 ;
  assign n39513 = ~n341 & n5102 ;
  assign n39509 = n668 & ~n10755 ;
  assign n39510 = n1269 & n5062 ;
  assign n39511 = n39509 & n39510 ;
  assign n39512 = n5225 & ~n39511 ;
  assign n39514 = n39513 ^ n39512 ^ n36883 ;
  assign n39515 = n23128 ^ n7693 ^ n4286 ;
  assign n39516 = n23039 & n39515 ;
  assign n39517 = ~n16702 & n19640 ;
  assign n39518 = n39517 ^ n6552 ^ 1'b0 ;
  assign n39519 = n10660 & n39518 ;
  assign n39520 = n14379 | n15203 ;
  assign n39521 = n39520 ^ n8112 ^ 1'b0 ;
  assign n39522 = n39521 ^ n25078 ^ 1'b0 ;
  assign n39523 = n21272 & ~n39522 ;
  assign n39524 = n35212 & n39523 ;
  assign n39525 = n39524 ^ n14490 ^ 1'b0 ;
  assign n39531 = x60 & ~n17832 ;
  assign n39526 = n9855 | n24437 ;
  assign n39527 = n6660 & n39526 ;
  assign n39528 = ~n29239 & n39527 ;
  assign n39529 = n33050 ^ n8277 ^ 1'b0 ;
  assign n39530 = n39528 | n39529 ;
  assign n39532 = n39531 ^ n39530 ^ n8829 ;
  assign n39533 = n4070 ^ n994 ^ 1'b0 ;
  assign n39534 = n14236 ^ x248 ^ 1'b0 ;
  assign n39535 = n1197 & ~n39534 ;
  assign n39536 = n27136 ^ n9385 ^ 1'b0 ;
  assign n39537 = ~n30082 & n39536 ;
  assign n39538 = n11389 & n24658 ;
  assign n39539 = n7472 | n21266 ;
  assign n39540 = n39538 & ~n39539 ;
  assign n39541 = n14527 ^ x73 ^ 1'b0 ;
  assign n39542 = n19467 | n39541 ;
  assign n39543 = n36785 & ~n39542 ;
  assign n39544 = n39543 ^ n7639 ^ 1'b0 ;
  assign n39545 = ( n10863 & n14014 ) | ( n10863 & ~n39095 ) | ( n14014 & ~n39095 ) ;
  assign n39546 = n29835 ^ n20230 ^ 1'b0 ;
  assign n39547 = n3847 & n39546 ;
  assign n39548 = n25999 ^ n18335 ^ 1'b0 ;
  assign n39549 = n39547 & n39548 ;
  assign n39550 = n26730 ^ n22680 ^ n7754 ;
  assign n39551 = n34479 ^ n1399 ^ 1'b0 ;
  assign n39552 = n39550 | n39551 ;
  assign n39553 = n36037 ^ n17836 ^ 1'b0 ;
  assign n39554 = n11320 | n39553 ;
  assign n39555 = n7895 ^ n5929 ^ 1'b0 ;
  assign n39556 = n25060 ^ n13099 ^ 1'b0 ;
  assign n39557 = n25138 & ~n39556 ;
  assign n39558 = n29819 ^ n23559 ^ n11525 ;
  assign n39559 = n26556 & n39558 ;
  assign n39560 = n13543 & n31938 ;
  assign n39561 = n13463 & n34082 ;
  assign n39562 = n11480 | n21585 ;
  assign n39563 = n39561 | n39562 ;
  assign n39564 = n39563 ^ n2701 ^ 1'b0 ;
  assign n39565 = n16005 & ~n39564 ;
  assign n39566 = n20261 ^ n17438 ^ 1'b0 ;
  assign n39567 = n30620 | n39566 ;
  assign n39568 = n34582 & ~n39567 ;
  assign n39569 = ~n10909 & n39568 ;
  assign n39572 = n5078 & ~n13329 ;
  assign n39573 = n2677 & n39572 ;
  assign n39570 = n4089 | n5076 ;
  assign n39571 = n11545 | n39570 ;
  assign n39574 = n39573 ^ n39571 ^ 1'b0 ;
  assign n39575 = n30982 | n39574 ;
  assign n39576 = ( n2240 & n5311 ) | ( n2240 & ~n14636 ) | ( n5311 & ~n14636 ) ;
  assign n39577 = n10272 & n23236 ;
  assign n39578 = n39577 ^ n35885 ^ 1'b0 ;
  assign n39579 = n39576 & ~n39578 ;
  assign n39580 = n36832 & n39579 ;
  assign n39581 = n18861 ^ n9927 ^ 1'b0 ;
  assign n39582 = ( n16321 & ~n35265 ) | ( n16321 & n39581 ) | ( ~n35265 & n39581 ) ;
  assign n39583 = n7616 & ~n30826 ;
  assign n39584 = n39583 ^ n31193 ^ n26889 ;
  assign n39585 = n19013 & ~n33555 ;
  assign n39586 = n5710 | n10020 ;
  assign n39587 = ~n14578 & n39586 ;
  assign n39588 = n23823 ^ n6306 ^ 1'b0 ;
  assign n39589 = n17134 | n39588 ;
  assign n39590 = ( n2774 & n13170 ) | ( n2774 & ~n29196 ) | ( n13170 & ~n29196 ) ;
  assign n39591 = n29929 ^ n8821 ^ 1'b0 ;
  assign n39592 = n14490 | n18291 ;
  assign n39593 = n33552 & ~n39592 ;
  assign n39594 = n39593 ^ n785 ^ 1'b0 ;
  assign n39595 = n4340 ^ n920 ^ 1'b0 ;
  assign n39596 = n6681 & ~n15391 ;
  assign n39597 = n8157 & n39596 ;
  assign n39598 = n10639 & ~n39597 ;
  assign n39599 = n31615 & n39598 ;
  assign n39600 = n39595 & n39599 ;
  assign n39601 = n4374 | n39600 ;
  assign n39602 = n39601 ^ n25349 ^ 1'b0 ;
  assign n39603 = n17550 & n31701 ;
  assign n39604 = n39603 ^ n34287 ^ 1'b0 ;
  assign n39605 = n39604 ^ n38377 ^ n2601 ;
  assign n39606 = n38080 ^ n14850 ^ n4084 ;
  assign n39607 = n2443 | n2931 ;
  assign n39608 = n22179 | n39607 ;
  assign n39609 = n39608 ^ n10170 ^ n2233 ;
  assign n39610 = n1250 | n7543 ;
  assign n39611 = n39609 & ~n39610 ;
  assign n39612 = n12155 | n13824 ;
  assign n39613 = n20458 & ~n39612 ;
  assign n39614 = n39613 ^ n38724 ^ 1'b0 ;
  assign n39615 = n24875 ^ n2877 ^ 1'b0 ;
  assign n39616 = n39615 ^ n5195 ^ 1'b0 ;
  assign n39617 = n7308 & ~n11448 ;
  assign n39618 = n7109 ^ n4431 ^ 1'b0 ;
  assign n39619 = ~n7334 & n39618 ;
  assign n39620 = n30384 ^ n22490 ^ 1'b0 ;
  assign n39621 = n39619 & ~n39620 ;
  assign n39622 = n15859 | n39621 ;
  assign n39623 = n1820 & ~n29211 ;
  assign n39624 = ~n11268 & n21058 ;
  assign n39625 = n39624 ^ n19323 ^ 1'b0 ;
  assign n39626 = n22990 ^ x114 ^ 1'b0 ;
  assign n39627 = n10638 & n14539 ;
  assign n39628 = n39627 ^ n11671 ^ n11634 ;
  assign n39629 = n496 | n8894 ;
  assign n39630 = n39629 ^ n12634 ^ 1'b0 ;
  assign n39631 = n39628 & ~n39630 ;
  assign n39632 = n8608 & ~n9350 ;
  assign n39633 = ( ~n12546 & n19524 ) | ( ~n12546 & n39632 ) | ( n19524 & n39632 ) ;
  assign n39634 = n715 & n27810 ;
  assign n39635 = n39634 ^ n38861 ^ 1'b0 ;
  assign n39639 = n7273 | n8228 ;
  assign n39640 = ~n15282 & n39639 ;
  assign n39641 = n39640 ^ n13346 ^ 1'b0 ;
  assign n39642 = n39641 ^ n14479 ^ n2823 ;
  assign n39638 = n21144 ^ n16187 ^ n11295 ;
  assign n39636 = n18463 & ~n26682 ;
  assign n39637 = ~n9799 & n39636 ;
  assign n39643 = n39642 ^ n39638 ^ n39637 ;
  assign n39644 = n17922 ^ n17607 ^ n3054 ;
  assign n39645 = n4255 & n32679 ;
  assign n39646 = ~n29710 & n39645 ;
  assign n39647 = n20174 ^ n11845 ^ 1'b0 ;
  assign n39648 = n32149 ^ n22595 ^ n16673 ;
  assign n39649 = n6611 | n39648 ;
  assign n39650 = n39649 ^ n28924 ^ n23551 ;
  assign n39651 = n15886 & n17061 ;
  assign n39652 = n39651 ^ n36236 ^ 1'b0 ;
  assign n39653 = n30605 & ~n39652 ;
  assign n39654 = ( ~n5884 & n27810 ) | ( ~n5884 & n39653 ) | ( n27810 & n39653 ) ;
  assign n39655 = n15938 ^ n5726 ^ 1'b0 ;
  assign n39656 = n12629 & ~n16759 ;
  assign n39657 = n20299 & ~n21033 ;
  assign n39658 = n39657 ^ n22256 ^ 1'b0 ;
  assign n39659 = n32605 ^ n27602 ^ n11389 ;
  assign n39660 = n39659 ^ n18717 ^ n11163 ;
  assign n39661 = n8737 | n25151 ;
  assign n39662 = ~n14033 & n26083 ;
  assign n39663 = n39662 ^ n2557 ^ 1'b0 ;
  assign n39665 = ~n14144 & n20644 ;
  assign n39666 = n8796 | n39665 ;
  assign n39667 = n39666 ^ n2523 ^ 1'b0 ;
  assign n39664 = n22322 ^ n12188 ^ n4258 ;
  assign n39668 = n39667 ^ n39664 ^ n3705 ;
  assign n39669 = n27548 ^ n450 ^ 1'b0 ;
  assign n39670 = ~n39668 & n39669 ;
  assign n39671 = n31105 ^ n27713 ^ 1'b0 ;
  assign n39672 = n17738 & ~n39671 ;
  assign n39673 = n7586 ^ n423 ^ 1'b0 ;
  assign n39674 = ~n26975 & n39673 ;
  assign n39675 = n26930 & n39674 ;
  assign n39676 = n7368 ^ n1593 ^ 1'b0 ;
  assign n39677 = ~n39675 & n39676 ;
  assign n39678 = n36981 ^ n19913 ^ 1'b0 ;
  assign n39679 = ~n16202 & n25490 ;
  assign n39680 = n1176 | n5732 ;
  assign n39681 = n39679 | n39680 ;
  assign n39682 = ( ~n5819 & n6788 ) | ( ~n5819 & n39681 ) | ( n6788 & n39681 ) ;
  assign n39683 = n7342 & n13109 ;
  assign n39684 = n27612 & n39683 ;
  assign n39685 = n39684 ^ n10959 ^ n3613 ;
  assign n39688 = n2819 | n38542 ;
  assign n39689 = n39688 ^ n7302 ^ 1'b0 ;
  assign n39690 = n15958 ^ n1806 ^ 1'b0 ;
  assign n39691 = ~n5460 & n39690 ;
  assign n39692 = ~n39689 & n39691 ;
  assign n39693 = n12799 | n27812 ;
  assign n39694 = n39692 & ~n39693 ;
  assign n39686 = n9187 | n18017 ;
  assign n39687 = n30348 & ~n39686 ;
  assign n39695 = n39694 ^ n39687 ^ 1'b0 ;
  assign n39696 = ~n11595 & n12460 ;
  assign n39697 = n6842 | n39696 ;
  assign n39698 = n19338 & ~n39697 ;
  assign n39699 = n19784 ^ n8700 ^ 1'b0 ;
  assign n39700 = n13374 ^ x49 ^ 1'b0 ;
  assign n39701 = n29487 ^ n19608 ^ 1'b0 ;
  assign n39702 = ~n16408 & n31475 ;
  assign n39703 = n34317 & ~n39702 ;
  assign n39704 = n15820 & ~n32157 ;
  assign n39705 = n14088 & ~n15722 ;
  assign n39706 = n39705 ^ n10380 ^ 1'b0 ;
  assign n39707 = n1021 | n24844 ;
  assign n39708 = n39707 ^ n9901 ^ 1'b0 ;
  assign n39709 = n14897 ^ n1379 ^ 1'b0 ;
  assign n39710 = n39709 ^ n37491 ^ 1'b0 ;
  assign n39711 = n9996 | n39710 ;
  assign n39712 = ( n8582 & n10088 ) | ( n8582 & ~n20278 ) | ( n10088 & ~n20278 ) ;
  assign n39713 = ~n15963 & n39712 ;
  assign n39714 = n29550 ^ n26518 ^ n7464 ;
  assign n39719 = n10135 & n17738 ;
  assign n39720 = n16673 ^ n15959 ^ 1'b0 ;
  assign n39721 = ~n39719 & n39720 ;
  assign n39715 = ~n5470 & n15157 ;
  assign n39716 = n12943 & n39715 ;
  assign n39717 = n12239 & ~n39716 ;
  assign n39718 = n39717 ^ n1161 ^ 1'b0 ;
  assign n39722 = n39721 ^ n39718 ^ n38042 ;
  assign n39723 = n35457 ^ n8839 ^ 1'b0 ;
  assign n39724 = x7 & ~n1827 ;
  assign n39725 = n14465 & n39724 ;
  assign n39726 = ~n24488 & n26945 ;
  assign n39727 = ~n15840 & n39726 ;
  assign n39728 = ( ~n31618 & n39725 ) | ( ~n31618 & n39727 ) | ( n39725 & n39727 ) ;
  assign n39729 = n12721 & ~n21270 ;
  assign n39730 = n835 | n19380 ;
  assign n39731 = n5954 ^ n4651 ^ 1'b0 ;
  assign n39732 = n500 & n39731 ;
  assign n39733 = n34864 ^ n7750 ^ 1'b0 ;
  assign n39734 = n1387 & ~n39733 ;
  assign n39735 = ~n39732 & n39734 ;
  assign n39736 = n1173 | n39735 ;
  assign n39737 = n29949 & ~n32831 ;
  assign n39738 = ( n13535 & ~n38634 ) | ( n13535 & n39737 ) | ( ~n38634 & n39737 ) ;
  assign n39739 = ( n17491 & n32049 ) | ( n17491 & ~n39738 ) | ( n32049 & ~n39738 ) ;
  assign n39740 = n17108 ^ n14128 ^ n3991 ;
  assign n39741 = n9532 & n32831 ;
  assign n39742 = n15118 & n39261 ;
  assign n39743 = n39742 ^ n16532 ^ 1'b0 ;
  assign n39744 = n39743 ^ n1899 ^ 1'b0 ;
  assign n39745 = n17773 ^ n16233 ^ n6094 ;
  assign n39746 = n12848 & n38275 ;
  assign n39747 = ~n39745 & n39746 ;
  assign n39748 = ( ~n28998 & n39744 ) | ( ~n28998 & n39747 ) | ( n39744 & n39747 ) ;
  assign n39749 = n2846 | n11277 ;
  assign n39752 = ( ~x132 & n5535 ) | ( ~x132 & n14138 ) | ( n5535 & n14138 ) ;
  assign n39750 = n5444 & n9844 ;
  assign n39751 = ~x188 & n39750 ;
  assign n39753 = n39752 ^ n39751 ^ 1'b0 ;
  assign n39754 = n7212 & n39753 ;
  assign n39755 = n13515 & n39754 ;
  assign n39756 = n32322 ^ n16847 ^ 1'b0 ;
  assign n39757 = n10568 & ~n39756 ;
  assign n39758 = n1096 | n3977 ;
  assign n39759 = n39758 ^ n19673 ^ 1'b0 ;
  assign n39760 = ~n14103 & n39759 ;
  assign n39761 = n39760 ^ n29241 ^ 1'b0 ;
  assign n39762 = x95 & ~n28982 ;
  assign n39763 = ~n39761 & n39762 ;
  assign n39765 = n1705 & n20852 ;
  assign n39766 = n12331 & n39765 ;
  assign n39764 = n26643 ^ n6453 ^ 1'b0 ;
  assign n39767 = n39766 ^ n39764 ^ n26244 ;
  assign n39768 = n6769 & n14654 ;
  assign n39769 = n39768 ^ n26602 ^ 1'b0 ;
  assign n39770 = n39769 ^ n17414 ^ 1'b0 ;
  assign n39771 = n39770 ^ x83 ^ 1'b0 ;
  assign n39772 = n5950 & n24899 ;
  assign n39773 = n13106 & n39772 ;
  assign n39774 = n2261 | n16722 ;
  assign n39775 = n39774 ^ n5213 ^ 1'b0 ;
  assign n39776 = n13698 ^ n12906 ^ n2466 ;
  assign n39777 = n28896 ^ n26186 ^ 1'b0 ;
  assign n39778 = n374 & n39777 ;
  assign n39779 = n39778 ^ n3087 ^ 1'b0 ;
  assign n39780 = n39776 & n39779 ;
  assign n39781 = n11410 ^ n9017 ^ n3015 ;
  assign n39782 = n39781 ^ n22916 ^ 1'b0 ;
  assign n39783 = n7965 & n39782 ;
  assign n39784 = n38670 ^ n4045 ^ 1'b0 ;
  assign n39785 = ~n32976 & n39784 ;
  assign n39786 = n3943 | n28627 ;
  assign n39787 = n21042 ^ n16689 ^ n3793 ;
  assign n39788 = n3564 & ~n39787 ;
  assign n39789 = n8088 | n17300 ;
  assign n39790 = ~n18184 & n39789 ;
  assign n39791 = n16852 ^ n13881 ^ 1'b0 ;
  assign n39792 = n24678 ^ n13664 ^ 1'b0 ;
  assign n39793 = n2088 & ~n15756 ;
  assign n39794 = n39792 & n39793 ;
  assign n39795 = n24037 ^ n8175 ^ n2859 ;
  assign n39796 = n23890 & ~n39795 ;
  assign n39797 = n39796 ^ n5017 ^ 1'b0 ;
  assign n39798 = ~n10095 & n34524 ;
  assign n39799 = n39798 ^ n7943 ^ 1'b0 ;
  assign n39800 = n39799 ^ n6722 ^ 1'b0 ;
  assign n39801 = n37009 | n39800 ;
  assign n39802 = n19390 ^ n8345 ^ n5662 ;
  assign n39803 = n13680 | n39802 ;
  assign n39804 = n9624 & ~n39803 ;
  assign n39805 = ~n7189 & n9349 ;
  assign n39806 = n39804 & n39805 ;
  assign n39807 = n22413 ^ n10938 ^ 1'b0 ;
  assign n39808 = n26284 & ~n39807 ;
  assign n39809 = n11758 ^ n8597 ^ 1'b0 ;
  assign n39810 = n29695 & n39809 ;
  assign n39811 = n39810 ^ n25164 ^ n24359 ;
  assign n39812 = n39127 ^ n8415 ^ n3423 ;
  assign n39813 = n39812 ^ n14849 ^ n11739 ;
  assign n39814 = n1956 & ~n5553 ;
  assign n39815 = n25834 ^ n6512 ^ 1'b0 ;
  assign n39816 = ~n3475 & n12057 ;
  assign n39817 = ~n1244 & n7689 ;
  assign n39818 = ~n4457 & n39817 ;
  assign n39819 = ( n6093 & ~n38262 ) | ( n6093 & n39818 ) | ( ~n38262 & n39818 ) ;
  assign n39820 = n12353 ^ n8110 ^ 1'b0 ;
  assign n39821 = ( ~n10201 & n28875 ) | ( ~n10201 & n39820 ) | ( n28875 & n39820 ) ;
  assign n39822 = n24089 | n37396 ;
  assign n39823 = ~n14466 & n25457 ;
  assign n39824 = n39823 ^ n22479 ^ 1'b0 ;
  assign n39825 = n39824 ^ n6295 ^ n5071 ;
  assign n39826 = n21773 | n26269 ;
  assign n39827 = ( n16599 & n17928 ) | ( n16599 & n39826 ) | ( n17928 & n39826 ) ;
  assign n39828 = n18761 & n39827 ;
  assign n39829 = ~n39825 & n39828 ;
  assign n39830 = ~n24584 & n28560 ;
  assign n39831 = ~n9402 & n39830 ;
  assign n39832 = ~n9404 & n26550 ;
  assign n39833 = ( n8168 & n35281 ) | ( n8168 & ~n39832 ) | ( n35281 & ~n39832 ) ;
  assign n39834 = n39833 ^ n29540 ^ n22684 ;
  assign n39835 = n27154 ^ n12680 ^ 1'b0 ;
  assign n39836 = ~n11805 & n39835 ;
  assign n39837 = n39836 ^ n38770 ^ 1'b0 ;
  assign n39838 = n39837 ^ n18182 ^ 1'b0 ;
  assign n39839 = n3344 & n32525 ;
  assign n39840 = n9079 & n39839 ;
  assign n39841 = n9576 | n32814 ;
  assign n39842 = n39841 ^ n24473 ^ 1'b0 ;
  assign n39843 = ~n39840 & n39842 ;
  assign n39844 = ~n16911 & n39843 ;
  assign n39847 = n801 & ~n9454 ;
  assign n39848 = ~n801 & n39847 ;
  assign n39845 = n3436 | n19604 ;
  assign n39846 = n5358 | n39845 ;
  assign n39849 = n39848 ^ n39846 ^ 1'b0 ;
  assign n39850 = n25123 & ~n39849 ;
  assign n39851 = n12483 & n39850 ;
  assign n39852 = ~n33926 & n39851 ;
  assign n39853 = ~n4447 & n8659 ;
  assign n39854 = n39853 ^ x143 ^ 1'b0 ;
  assign n39855 = n21788 ^ n11070 ^ 1'b0 ;
  assign n39856 = n4955 & ~n39855 ;
  assign n39857 = n37074 ^ n11035 ^ 1'b0 ;
  assign n39858 = n24545 ^ n18752 ^ n12893 ;
  assign n39859 = n39858 ^ n26437 ^ n9255 ;
  assign n39860 = n3568 & n13660 ;
  assign n39861 = n39860 ^ n7004 ^ 1'b0 ;
  assign n39862 = n9187 ^ n4014 ^ x197 ;
  assign n39863 = n39862 ^ n15927 ^ 1'b0 ;
  assign n39864 = n3327 & ~n39863 ;
  assign n39865 = n39861 & n39864 ;
  assign n39866 = ~n8337 & n39865 ;
  assign n39867 = ( ~n6487 & n39859 ) | ( ~n6487 & n39866 ) | ( n39859 & n39866 ) ;
  assign n39868 = ~n4683 & n8294 ;
  assign n39869 = n22244 ^ n3605 ^ 1'b0 ;
  assign n39870 = n39868 & n39869 ;
  assign n39871 = n19005 & n25930 ;
  assign n39872 = n39871 ^ n31136 ^ 1'b0 ;
  assign n39873 = n15776 ^ n6232 ^ 1'b0 ;
  assign n39874 = n38944 & n39873 ;
  assign n39875 = ~n22638 & n39874 ;
  assign n39876 = n3282 & n39875 ;
  assign n39877 = ~n20546 & n36128 ;
  assign n39878 = n9996 ^ n4683 ^ 1'b0 ;
  assign n39879 = n15371 ^ x37 ^ 1'b0 ;
  assign n39880 = n29963 & n39879 ;
  assign n39881 = n25464 ^ n21897 ^ n13398 ;
  assign n39882 = ( n9770 & n39880 ) | ( n9770 & n39881 ) | ( n39880 & n39881 ) ;
  assign n39883 = ( n4817 & ~n8114 ) | ( n4817 & n9326 ) | ( ~n8114 & n9326 ) ;
  assign n39884 = ~n19309 & n30670 ;
  assign n39885 = ~n39883 & n39884 ;
  assign n39886 = n23402 ^ n7943 ^ 1'b0 ;
  assign n39887 = n731 & n39886 ;
  assign n39888 = n13600 | n25277 ;
  assign n39889 = n39888 ^ n32254 ^ 1'b0 ;
  assign n39890 = n28862 ^ n9341 ^ 1'b0 ;
  assign n39891 = n25020 ^ n22969 ^ 1'b0 ;
  assign n39892 = n29490 & n39891 ;
  assign n39893 = ( n9237 & ~n19197 ) | ( n9237 & n25052 ) | ( ~n19197 & n25052 ) ;
  assign n39894 = n4142 & ~n24949 ;
  assign n39895 = n4882 | n25300 ;
  assign n39896 = n39895 ^ n14785 ^ 1'b0 ;
  assign n39897 = ( ~n5030 & n11009 ) | ( ~n5030 & n39896 ) | ( n11009 & n39896 ) ;
  assign n39898 = ~n13942 & n18189 ;
  assign n39899 = n39898 ^ n24129 ^ 1'b0 ;
  assign n39900 = n4224 | n30079 ;
  assign n39901 = x37 | n39900 ;
  assign n39902 = n39526 & n39901 ;
  assign n39903 = n39902 ^ n11902 ^ 1'b0 ;
  assign n39904 = n19346 ^ n7122 ^ 1'b0 ;
  assign n39905 = n39903 | n39904 ;
  assign n39906 = n9887 & n39905 ;
  assign n39908 = ~n13382 & n23351 ;
  assign n39907 = ~n1624 & n14839 ;
  assign n39909 = n39908 ^ n39907 ^ 1'b0 ;
  assign n39910 = n38864 ^ n22469 ^ n18895 ;
  assign n39911 = ( n8223 & n25968 ) | ( n8223 & n39910 ) | ( n25968 & n39910 ) ;
  assign n39912 = ( ~n4061 & n4163 ) | ( ~n4061 & n8681 ) | ( n4163 & n8681 ) ;
  assign n39913 = n39912 ^ n22795 ^ n8013 ;
  assign n39914 = n6497 | n16327 ;
  assign n39915 = n12907 & ~n39914 ;
  assign n39917 = ~n14785 & n26099 ;
  assign n39918 = n2338 & n39917 ;
  assign n39919 = n22523 ^ n7040 ^ 1'b0 ;
  assign n39920 = n39918 | n39919 ;
  assign n39916 = n2566 & n20352 ;
  assign n39921 = n39920 ^ n39916 ^ 1'b0 ;
  assign n39923 = ~n14683 & n24350 ;
  assign n39924 = n8837 & n39923 ;
  assign n39925 = ~n26994 & n39924 ;
  assign n39922 = n4411 & n28461 ;
  assign n39926 = n39925 ^ n39922 ^ 1'b0 ;
  assign n39927 = n9949 & ~n11344 ;
  assign n39928 = ~n12998 & n16600 ;
  assign n39929 = ~n13175 & n39928 ;
  assign n39930 = n10848 | n39929 ;
  assign n39931 = ~n3401 & n20566 ;
  assign n39932 = n25714 ^ n16663 ^ n13221 ;
  assign n39933 = n27324 ^ n21822 ^ n7957 ;
  assign n39936 = n29839 ^ n22617 ^ 1'b0 ;
  assign n39934 = n9521 & n20771 ;
  assign n39935 = ~n18818 & n39934 ;
  assign n39937 = n39936 ^ n39935 ^ 1'b0 ;
  assign n39938 = ~n24573 & n35403 ;
  assign n39939 = ~n2580 & n39938 ;
  assign n39940 = n39939 ^ n7084 ^ 1'b0 ;
  assign n39941 = n38729 & n39940 ;
  assign n39942 = n39941 ^ n36970 ^ 1'b0 ;
  assign n39943 = n28391 & n37908 ;
  assign n39944 = n39943 ^ n34893 ^ 1'b0 ;
  assign n39945 = n12091 | n29929 ;
  assign n39946 = n34272 | n39945 ;
  assign n39947 = n2379 | n22432 ;
  assign n39948 = n20120 ^ n5868 ^ n4280 ;
  assign n39949 = n9522 ^ n4174 ^ 1'b0 ;
  assign n39950 = x74 & n39949 ;
  assign n39951 = n39264 ^ n10798 ^ n1514 ;
  assign n39952 = n7792 | n28051 ;
  assign n39953 = n39951 & ~n39952 ;
  assign n39954 = n4439 & ~n4927 ;
  assign n39955 = n39954 ^ n2019 ^ 1'b0 ;
  assign n39956 = n7152 & ~n39955 ;
  assign n39957 = n14203 ^ n9740 ^ n5110 ;
  assign n39958 = n13330 ^ n8895 ^ n3619 ;
  assign n39959 = n39958 ^ n22470 ^ 1'b0 ;
  assign n39960 = n39959 ^ n37693 ^ n14822 ;
  assign n39961 = n27810 ^ n13148 ^ 1'b0 ;
  assign n39962 = n12519 & ~n13012 ;
  assign n39963 = n22835 ^ n7606 ^ 1'b0 ;
  assign n39964 = n39963 ^ n39180 ^ n262 ;
  assign n39965 = ( ~x252 & n10767 ) | ( ~x252 & n24613 ) | ( n10767 & n24613 ) ;
  assign n39966 = n39965 ^ n4591 ^ 1'b0 ;
  assign n39967 = n16847 & ~n30237 ;
  assign n39968 = n35731 ^ n11928 ^ 1'b0 ;
  assign n39969 = n10939 & n17490 ;
  assign n39970 = n39969 ^ n23263 ^ 1'b0 ;
  assign n39971 = n14030 & ~n29603 ;
  assign n39972 = n39971 ^ n36047 ^ n35014 ;
  assign n39973 = ~n20154 & n32874 ;
  assign n39974 = n39973 ^ n7734 ^ n2068 ;
  assign n39975 = n39974 ^ n27581 ^ 1'b0 ;
  assign n39976 = ( n1805 & n4685 ) | ( n1805 & ~n15568 ) | ( n4685 & ~n15568 ) ;
  assign n39977 = n35444 ^ n22713 ^ n6045 ;
  assign n39978 = n15772 ^ n1529 ^ 1'b0 ;
  assign n39979 = n26769 & ~n38915 ;
  assign n39980 = n39979 ^ n1248 ^ 1'b0 ;
  assign n39981 = n15228 | n25994 ;
  assign n39982 = n39981 ^ n35396 ^ 1'b0 ;
  assign n39983 = n33653 ^ x94 ^ 1'b0 ;
  assign n39984 = n39983 ^ n33779 ^ n16532 ;
  assign n39985 = ~n13158 & n39984 ;
  assign n39986 = n31120 ^ n9332 ^ n7371 ;
  assign n39987 = n36128 ^ n19592 ^ n16106 ;
  assign n39988 = n14440 ^ n4153 ^ 1'b0 ;
  assign n39989 = n11063 & n39988 ;
  assign n39990 = ~n3097 & n39989 ;
  assign n39991 = n39990 ^ n1080 ^ 1'b0 ;
  assign n39992 = n39991 ^ n11100 ^ n5432 ;
  assign n39993 = n39992 ^ n12046 ^ 1'b0 ;
  assign n39994 = n2282 & ~n19653 ;
  assign n39995 = n31170 ^ n3255 ^ 1'b0 ;
  assign n39996 = ~n14790 & n29707 ;
  assign n39997 = ( ~n4270 & n6889 ) | ( ~n4270 & n20215 ) | ( n6889 & n20215 ) ;
  assign n39998 = ( n2626 & n2851 ) | ( n2626 & n6328 ) | ( n2851 & n6328 ) ;
  assign n39999 = ( ~n6732 & n29834 ) | ( ~n6732 & n39998 ) | ( n29834 & n39998 ) ;
  assign n40000 = n31947 ^ n21966 ^ n4318 ;
  assign n40001 = n40000 ^ n11523 ^ 1'b0 ;
  assign n40002 = n39605 ^ n1071 ^ 1'b0 ;
  assign n40003 = n12594 | n20846 ;
  assign n40004 = n8855 ^ n741 ^ 1'b0 ;
  assign n40005 = ~n9282 & n14840 ;
  assign n40006 = ~n31024 & n40005 ;
  assign n40007 = n39068 ^ n2151 ^ 1'b0 ;
  assign n40008 = n8956 & n15351 ;
  assign n40009 = n40008 ^ n3254 ^ 1'b0 ;
  assign n40010 = n40009 ^ n19628 ^ 1'b0 ;
  assign n40011 = n27031 ^ n24615 ^ 1'b0 ;
  assign n40012 = n8376 & ~n11449 ;
  assign n40013 = n40012 ^ n33984 ^ 1'b0 ;
  assign n40014 = ~n3312 & n40013 ;
  assign n40015 = n3190 & n8063 ;
  assign n40016 = n40015 ^ n7895 ^ 1'b0 ;
  assign n40017 = n16812 & n40016 ;
  assign n40018 = ~n40014 & n40017 ;
  assign n40019 = n8671 ^ n3934 ^ 1'b0 ;
  assign n40020 = n40019 ^ n22062 ^ n5170 ;
  assign n40021 = n369 | n28223 ;
  assign n40022 = n1272 ^ n973 ^ 1'b0 ;
  assign n40023 = ~n10109 & n40022 ;
  assign n40024 = ~n31780 & n40023 ;
  assign n40025 = ~n35648 & n40024 ;
  assign n40026 = n33957 & n38996 ;
  assign n40027 = n6395 ^ n5291 ^ n533 ;
  assign n40028 = n34057 | n40027 ;
  assign n40029 = n38830 ^ n3274 ^ 1'b0 ;
  assign n40030 = n38233 ^ n14241 ^ 1'b0 ;
  assign n40031 = n16294 & n40030 ;
  assign n40032 = n1093 & ~n6794 ;
  assign n40033 = n40032 ^ n26849 ^ 1'b0 ;
  assign n40034 = ( n6929 & n15184 ) | ( n6929 & ~n28049 ) | ( n15184 & ~n28049 ) ;
  assign n40035 = n28248 & n40034 ;
  assign n40036 = ( n23211 & n28314 ) | ( n23211 & ~n40035 ) | ( n28314 & ~n40035 ) ;
  assign n40037 = n12384 ^ n12231 ^ n11035 ;
  assign n40038 = n31433 ^ n12786 ^ n2919 ;
  assign n40042 = n11072 & ~n18433 ;
  assign n40043 = ~n6361 & n40042 ;
  assign n40039 = n1511 & n10258 ;
  assign n40040 = n40039 ^ x244 ^ 1'b0 ;
  assign n40041 = ~n5090 & n40040 ;
  assign n40044 = n40043 ^ n40041 ^ 1'b0 ;
  assign n40045 = n39281 ^ n8519 ^ 1'b0 ;
  assign n40046 = n26861 & ~n40045 ;
  assign n40047 = ~n40044 & n40046 ;
  assign n40048 = ~n2111 & n23539 ;
  assign n40049 = n7336 & ~n29947 ;
  assign n40050 = n14629 ^ n550 ^ 1'b0 ;
  assign n40051 = n3935 & n40050 ;
  assign n40052 = ~n9413 & n40051 ;
  assign n40053 = n1321 & n40052 ;
  assign n40054 = n36738 & ~n40053 ;
  assign n40055 = ( n273 & ~n20806 ) | ( n273 & n25448 ) | ( ~n20806 & n25448 ) ;
  assign n40056 = n14505 & n25518 ;
  assign n40057 = ( n8017 & n27007 ) | ( n8017 & ~n27861 ) | ( n27007 & ~n27861 ) ;
  assign n40058 = n15825 & ~n24333 ;
  assign n40059 = ~n23606 & n40058 ;
  assign n40060 = ~n3600 & n8206 ;
  assign n40061 = n40060 ^ n34692 ^ 1'b0 ;
  assign n40062 = ( n3044 & n25011 ) | ( n3044 & ~n27058 ) | ( n25011 & ~n27058 ) ;
  assign n40063 = n33835 ^ n23115 ^ 1'b0 ;
  assign n40064 = n40062 & ~n40063 ;
  assign n40066 = n20323 ^ n335 ^ 1'b0 ;
  assign n40067 = ( n5881 & ~n8891 ) | ( n5881 & n40066 ) | ( ~n8891 & n40066 ) ;
  assign n40065 = n4893 | n5784 ;
  assign n40068 = n40067 ^ n40065 ^ 1'b0 ;
  assign n40069 = ( ~n15198 & n16982 ) | ( ~n15198 & n22425 ) | ( n16982 & n22425 ) ;
  assign n40070 = n5050 & n9892 ;
  assign n40071 = ~n40069 & n40070 ;
  assign n40072 = n40071 ^ n20649 ^ n13479 ;
  assign n40073 = n3532 | n11520 ;
  assign n40074 = n40073 ^ n5322 ^ 1'b0 ;
  assign n40075 = n40074 ^ n39704 ^ 1'b0 ;
  assign n40076 = ( ~n3255 & n4094 ) | ( ~n3255 & n9824 ) | ( n4094 & n9824 ) ;
  assign n40077 = ( n3349 & n13863 ) | ( n3349 & ~n40076 ) | ( n13863 & ~n40076 ) ;
  assign n40078 = ~n5843 & n10436 ;
  assign n40079 = n5952 | n30765 ;
  assign n40080 = n40079 ^ n9631 ^ 1'b0 ;
  assign n40081 = n1058 & n4209 ;
  assign n40082 = n40081 ^ n10925 ^ 1'b0 ;
  assign n40083 = n40082 ^ n1827 ^ 1'b0 ;
  assign n40084 = ~n40080 & n40083 ;
  assign n40085 = n40084 ^ n10058 ^ 1'b0 ;
  assign n40089 = ~n12107 & n28280 ;
  assign n40090 = ~n10173 & n40089 ;
  assign n40086 = n26441 ^ n18392 ^ 1'b0 ;
  assign n40087 = ~n26340 & n40086 ;
  assign n40088 = n5812 & ~n40087 ;
  assign n40091 = n40090 ^ n40088 ^ n22131 ;
  assign n40092 = n29544 ^ n19408 ^ 1'b0 ;
  assign n40093 = n29898 ^ n22289 ^ n4692 ;
  assign n40094 = n30323 ^ n27580 ^ 1'b0 ;
  assign n40095 = n8367 & n11053 ;
  assign n40096 = n40095 ^ n19264 ^ 1'b0 ;
  assign n40097 = n14606 ^ n12296 ^ n2443 ;
  assign n40098 = n40097 ^ n10327 ^ n5195 ;
  assign n40099 = n16937 & ~n20742 ;
  assign n40100 = n7653 ^ n6526 ^ 1'b0 ;
  assign n40101 = ( ~n6316 & n40099 ) | ( ~n6316 & n40100 ) | ( n40099 & n40100 ) ;
  assign n40102 = n17835 & n40009 ;
  assign n40103 = n40102 ^ n21230 ^ 1'b0 ;
  assign n40104 = n40103 ^ n31205 ^ n3826 ;
  assign n40106 = n27041 ^ n16095 ^ n7952 ;
  assign n40105 = ~n4670 & n20505 ;
  assign n40107 = n40106 ^ n40105 ^ n11200 ;
  assign n40108 = n40107 ^ n33757 ^ 1'b0 ;
  assign n40109 = n18758 | n40108 ;
  assign n40110 = n358 & ~n4282 ;
  assign n40111 = n10025 ^ n8944 ^ 1'b0 ;
  assign n40112 = n31504 ^ n23142 ^ 1'b0 ;
  assign n40113 = ~n40111 & n40112 ;
  assign n40114 = ~n15198 & n30431 ;
  assign n40115 = n40114 ^ n38777 ^ 1'b0 ;
  assign n40116 = ~n5306 & n10132 ;
  assign n40117 = n40116 ^ n17076 ^ 1'b0 ;
  assign n40118 = ( ~n8978 & n15825 ) | ( ~n8978 & n22701 ) | ( n15825 & n22701 ) ;
  assign n40119 = n40118 ^ n27906 ^ n6251 ;
  assign n40125 = n1004 | n3872 ;
  assign n40126 = n1004 & ~n40125 ;
  assign n40127 = n2827 & ~n40126 ;
  assign n40128 = n40126 & n40127 ;
  assign n40120 = n2275 | n32875 ;
  assign n40121 = n32875 & ~n40120 ;
  assign n40122 = ( n604 & n1129 ) | ( n604 & ~n1806 ) | ( n1129 & ~n1806 ) ;
  assign n40123 = n40121 & n40122 ;
  assign n40124 = n15989 | n40123 ;
  assign n40129 = n40128 ^ n40124 ^ 1'b0 ;
  assign n40130 = n40129 ^ n39348 ^ n36992 ;
  assign n40132 = n857 | n1204 ;
  assign n40133 = n40132 ^ x43 ^ 1'b0 ;
  assign n40134 = ( n7097 & ~n12353 ) | ( n7097 & n40133 ) | ( ~n12353 & n40133 ) ;
  assign n40131 = ( n915 & n16334 ) | ( n915 & ~n37639 ) | ( n16334 & ~n37639 ) ;
  assign n40135 = n40134 ^ n40131 ^ n7081 ;
  assign n40136 = ~n4290 & n15532 ;
  assign n40137 = n33295 ^ n8300 ^ 1'b0 ;
  assign n40138 = n40137 ^ n9445 ^ 1'b0 ;
  assign n40139 = n40136 & ~n40138 ;
  assign n40140 = ~n4597 & n6903 ;
  assign n40141 = ~n14811 & n40140 ;
  assign n40142 = n40141 ^ n18435 ^ n9843 ;
  assign n40143 = n17721 | n40142 ;
  assign n40144 = n16809 | n40143 ;
  assign n40146 = ~n9606 & n14157 ;
  assign n40147 = n40146 ^ n10735 ^ 1'b0 ;
  assign n40145 = ~n11912 & n33357 ;
  assign n40148 = n40147 ^ n40145 ^ 1'b0 ;
  assign n40149 = n17592 | n40148 ;
  assign n40150 = n40149 ^ n31481 ^ 1'b0 ;
  assign n40151 = n16613 ^ n1187 ^ 1'b0 ;
  assign n40152 = n40151 ^ n39096 ^ n7454 ;
  assign n40153 = n37584 ^ n874 ^ 1'b0 ;
  assign n40154 = n31789 ^ n13407 ^ 1'b0 ;
  assign n40155 = n14593 ^ n9358 ^ n3759 ;
  assign n40156 = n6289 & ~n23012 ;
  assign n40157 = n40155 & n40156 ;
  assign n40158 = n3544 | n16937 ;
  assign n40159 = ( n40154 & ~n40157 ) | ( n40154 & n40158 ) | ( ~n40157 & n40158 ) ;
  assign n40160 = n36385 ^ n6254 ^ 1'b0 ;
  assign n40161 = n10002 & n40160 ;
  assign n40162 = n20584 ^ n2200 ^ 1'b0 ;
  assign n40163 = n27490 ^ n2429 ^ 1'b0 ;
  assign n40164 = n5199 & n6933 ;
  assign n40165 = ( n19356 & n21640 ) | ( n19356 & n40164 ) | ( n21640 & n40164 ) ;
  assign n40166 = n40165 ^ n38913 ^ 1'b0 ;
  assign n40167 = n16334 & ~n40166 ;
  assign n40168 = n27774 ^ n11811 ^ 1'b0 ;
  assign n40169 = ( n19642 & n22665 ) | ( n19642 & n25824 ) | ( n22665 & n25824 ) ;
  assign n40170 = n18661 ^ n2929 ^ 1'b0 ;
  assign n40171 = n16642 ^ n3634 ^ 1'b0 ;
  assign n40172 = ( n20301 & ~n25839 ) | ( n20301 & n40171 ) | ( ~n25839 & n40171 ) ;
  assign n40173 = n20530 ^ n15913 ^ 1'b0 ;
  assign n40174 = n40173 ^ n22852 ^ 1'b0 ;
  assign n40175 = ~n604 & n40174 ;
  assign n40176 = n28815 ^ n24347 ^ 1'b0 ;
  assign n40177 = n35905 & ~n40176 ;
  assign n40178 = n4906 & n40177 ;
  assign n40179 = n12901 & ~n22691 ;
  assign n40180 = n40179 ^ n17536 ^ 1'b0 ;
  assign n40182 = n317 | n38554 ;
  assign n40183 = n40182 ^ n9156 ^ 1'b0 ;
  assign n40184 = n10650 & n40183 ;
  assign n40181 = n16668 | n30487 ;
  assign n40185 = n40184 ^ n40181 ^ 1'b0 ;
  assign n40186 = n1474 & ~n17990 ;
  assign n40187 = n40186 ^ n11118 ^ 1'b0 ;
  assign n40188 = n6829 & n18525 ;
  assign n40189 = n20720 & n40188 ;
  assign n40190 = x157 & n40189 ;
  assign n40191 = n30214 ^ n29896 ^ 1'b0 ;
  assign n40192 = n40191 ^ n32412 ^ n371 ;
  assign n40194 = n32885 ^ n8015 ^ 1'b0 ;
  assign n40193 = ~n10741 & n17358 ;
  assign n40195 = n40194 ^ n40193 ^ 1'b0 ;
  assign n40196 = n21804 ^ n901 ^ 1'b0 ;
  assign n40197 = n11587 | n40196 ;
  assign n40198 = n40197 ^ n14370 ^ 1'b0 ;
  assign n40199 = n263 & ~n8654 ;
  assign n40200 = n40199 ^ x46 ^ 1'b0 ;
  assign n40201 = ~n740 & n2119 ;
  assign n40202 = n15577 | n19854 ;
  assign n40203 = n6093 & ~n28634 ;
  assign n40204 = n40203 ^ n33594 ^ 1'b0 ;
  assign n40205 = ( ~n5526 & n28219 ) | ( ~n5526 & n40204 ) | ( n28219 & n40204 ) ;
  assign n40206 = ( n6138 & ~n7639 ) | ( n6138 & n16666 ) | ( ~n7639 & n16666 ) ;
  assign n40207 = ~n3146 & n33627 ;
  assign n40208 = n31838 ^ n23844 ^ 1'b0 ;
  assign n40209 = n24265 | n40208 ;
  assign n40210 = n17042 | n37891 ;
  assign n40211 = n2915 | n40210 ;
  assign n40212 = ( n314 & n888 ) | ( n314 & ~n11181 ) | ( n888 & ~n11181 ) ;
  assign n40213 = ( n792 & n29715 ) | ( n792 & n40212 ) | ( n29715 & n40212 ) ;
  assign n40214 = n10994 & ~n32304 ;
  assign n40215 = n40214 ^ n9740 ^ 1'b0 ;
  assign n40216 = n40215 ^ n39609 ^ n29136 ;
  assign n40217 = n19303 ^ n12077 ^ 1'b0 ;
  assign n40218 = n1663 | n6716 ;
  assign n40221 = n17926 ^ n10170 ^ n5985 ;
  assign n40222 = n40221 ^ n19342 ^ 1'b0 ;
  assign n40219 = n6545 & n11781 ;
  assign n40220 = n6243 | n40219 ;
  assign n40223 = n40222 ^ n40220 ^ 1'b0 ;
  assign n40224 = n40223 ^ n20648 ^ n11483 ;
  assign n40225 = n19542 & n31315 ;
  assign n40226 = n40224 & n40225 ;
  assign n40227 = n5391 & n25098 ;
  assign n40228 = ( n3762 & ~n24839 ) | ( n3762 & n27687 ) | ( ~n24839 & n27687 ) ;
  assign n40229 = n3506 | n10376 ;
  assign n40230 = n40229 ^ n35877 ^ n11064 ;
  assign n40231 = n9461 & ~n30946 ;
  assign n40232 = ~n36066 & n40231 ;
  assign n40233 = n36655 ^ n19506 ^ 1'b0 ;
  assign n40234 = n40019 ^ n29553 ^ n8828 ;
  assign n40235 = n19796 ^ n5584 ^ 1'b0 ;
  assign n40236 = n30974 | n40235 ;
  assign n40237 = n40236 ^ n15203 ^ n12094 ;
  assign n40238 = n6634 & n15389 ;
  assign n40239 = n29685 & n40238 ;
  assign n40240 = n20647 ^ n5859 ^ 1'b0 ;
  assign n40241 = n40239 | n40240 ;
  assign n40242 = n982 & ~n2183 ;
  assign n40243 = n40242 ^ n3724 ^ 1'b0 ;
  assign n40244 = n40243 ^ n358 ^ 1'b0 ;
  assign n40245 = n15526 ^ n3052 ^ 1'b0 ;
  assign n40246 = n9885 | n21419 ;
  assign n40247 = ( n3159 & ~n19228 ) | ( n3159 & n38701 ) | ( ~n19228 & n38701 ) ;
  assign n40250 = n27015 ^ n18335 ^ 1'b0 ;
  assign n40248 = n8748 | n17511 ;
  assign n40249 = n14892 | n40248 ;
  assign n40251 = n40250 ^ n40249 ^ n13356 ;
  assign n40252 = n40251 ^ n16083 ^ 1'b0 ;
  assign n40253 = n20131 & ~n28133 ;
  assign n40254 = n40253 ^ n23100 ^ 1'b0 ;
  assign n40255 = n40254 ^ n7627 ^ 1'b0 ;
  assign n40256 = n21029 ^ n5389 ^ 1'b0 ;
  assign n40257 = n3192 & n40256 ;
  assign n40258 = ( ~n11979 & n17447 ) | ( ~n11979 & n26840 ) | ( n17447 & n26840 ) ;
  assign n40259 = n40258 ^ n7325 ^ 1'b0 ;
  assign n40260 = n1701 | n40259 ;
  assign n40261 = n21651 & ~n37832 ;
  assign n40262 = ~n5519 & n40261 ;
  assign n40263 = n17574 & ~n33367 ;
  assign n40264 = n21299 & n40263 ;
  assign n40265 = n40264 ^ n26177 ^ 1'b0 ;
  assign n40266 = n15002 | n20265 ;
  assign n40267 = n40266 ^ n30664 ^ 1'b0 ;
  assign n40269 = n6791 ^ n6710 ^ 1'b0 ;
  assign n40268 = n21163 | n37424 ;
  assign n40270 = n40269 ^ n40268 ^ 1'b0 ;
  assign n40271 = ( n16430 & n40267 ) | ( n16430 & n40270 ) | ( n40267 & n40270 ) ;
  assign n40272 = n8073 | n35667 ;
  assign n40273 = n27167 ^ n23884 ^ 1'b0 ;
  assign n40274 = n27989 ^ n22940 ^ n7814 ;
  assign n40275 = n40274 ^ n33233 ^ 1'b0 ;
  assign n40276 = n25306 ^ n9924 ^ n6283 ;
  assign n40277 = n40276 ^ n29852 ^ n6157 ;
  assign n40278 = n40277 ^ n20745 ^ n10223 ;
  assign n40279 = n12138 ^ n2571 ^ 1'b0 ;
  assign n40280 = ( n1415 & n8842 ) | ( n1415 & n40279 ) | ( n8842 & n40279 ) ;
  assign n40281 = x237 & n4136 ;
  assign n40282 = ( n11982 & n40280 ) | ( n11982 & ~n40281 ) | ( n40280 & ~n40281 ) ;
  assign n40283 = n15661 ^ n672 ^ 1'b0 ;
  assign n40284 = n29520 ^ n10522 ^ n4901 ;
  assign n40285 = ( n7745 & n40283 ) | ( n7745 & ~n40284 ) | ( n40283 & ~n40284 ) ;
  assign n40286 = ~n1829 & n11806 ;
  assign n40287 = n40286 ^ n31364 ^ 1'b0 ;
  assign n40288 = n15689 ^ n15669 ^ 1'b0 ;
  assign n40289 = ~n6551 & n40288 ;
  assign n40290 = n4333 & ~n17607 ;
  assign n40291 = n4147 & n40290 ;
  assign n40292 = n20559 ^ n3612 ^ 1'b0 ;
  assign n40293 = n33097 | n40292 ;
  assign n40294 = n3257 | n40293 ;
  assign n40295 = n26483 & n40294 ;
  assign n40296 = n40295 ^ n13377 ^ 1'b0 ;
  assign n40297 = n40148 ^ n17422 ^ 1'b0 ;
  assign n40298 = n8368 & n16966 ;
  assign n40299 = n40298 ^ n16607 ^ 1'b0 ;
  assign n40300 = n11262 ^ n9164 ^ 1'b0 ;
  assign n40301 = n12440 ^ n8975 ^ x113 ;
  assign n40302 = n28344 ^ n16452 ^ n16060 ;
  assign n40305 = n4329 | n27251 ;
  assign n40303 = ~n10201 & n33722 ;
  assign n40304 = n23032 & n40303 ;
  assign n40306 = n40305 ^ n40304 ^ n5974 ;
  assign n40307 = ~n3550 & n17094 ;
  assign n40308 = n40307 ^ n22179 ^ 1'b0 ;
  assign n40309 = ~n17333 & n25100 ;
  assign n40310 = n25199 & ~n29042 ;
  assign n40311 = n40310 ^ n18693 ^ 1'b0 ;
  assign n40312 = n13560 & ~n38439 ;
  assign n40313 = n527 & n40312 ;
  assign n40314 = n6767 ^ n961 ^ 1'b0 ;
  assign n40315 = ~n17732 & n40314 ;
  assign n40316 = ~n10052 & n40315 ;
  assign n40317 = ~n6168 & n22160 ;
  assign n40318 = n14800 & n23606 ;
  assign n40319 = n14751 ^ n10304 ^ 1'b0 ;
  assign n40320 = ~n14480 & n40319 ;
  assign n40321 = n40320 ^ n32404 ^ 1'b0 ;
  assign n40322 = n40321 ^ n28462 ^ 1'b0 ;
  assign n40323 = ( n3053 & ~n3922 ) | ( n3053 & n40322 ) | ( ~n3922 & n40322 ) ;
  assign n40324 = n19624 ^ n2454 ^ 1'b0 ;
  assign n40325 = n28370 & ~n40324 ;
  assign n40326 = n40325 ^ n6159 ^ 1'b0 ;
  assign n40327 = n11261 & ~n40326 ;
  assign n40328 = n36300 ^ n2332 ^ 1'b0 ;
  assign n40329 = ( ~n8707 & n15586 ) | ( ~n8707 & n40328 ) | ( n15586 & n40328 ) ;
  assign n40330 = n22610 | n40329 ;
  assign n40331 = n7354 | n8293 ;
  assign n40332 = n1081 & ~n40331 ;
  assign n40333 = n40332 ^ n7124 ^ 1'b0 ;
  assign n40334 = n18994 ^ n8606 ^ 1'b0 ;
  assign n40335 = n1814 ^ n1511 ^ 1'b0 ;
  assign n40336 = n40335 ^ n27933 ^ n542 ;
  assign n40337 = n40336 ^ n5518 ^ 1'b0 ;
  assign n40338 = ~n22319 & n40337 ;
  assign n40339 = ~n14081 & n14242 ;
  assign n40340 = n40339 ^ n35892 ^ 1'b0 ;
  assign n40341 = n21153 ^ n17194 ^ 1'b0 ;
  assign n40342 = n16062 ^ n2916 ^ 1'b0 ;
  assign n40343 = ( n5603 & ~n22486 ) | ( n5603 & n24921 ) | ( ~n22486 & n24921 ) ;
  assign n40344 = n14490 & ~n37729 ;
  assign n40345 = ~n29431 & n40344 ;
  assign n40346 = n23271 ^ n22362 ^ 1'b0 ;
  assign n40347 = n35905 & ~n40346 ;
  assign n40348 = n4895 & n15867 ;
  assign n40349 = n40348 ^ n11257 ^ 1'b0 ;
  assign n40350 = n40349 ^ n6078 ^ 1'b0 ;
  assign n40351 = n40347 & n40350 ;
  assign n40352 = n16746 | n32398 ;
  assign n40353 = n7537 | n40352 ;
  assign n40354 = n38906 ^ n29945 ^ 1'b0 ;
  assign n40355 = n16044 | n31609 ;
  assign n40356 = n17460 ^ n302 ^ 1'b0 ;
  assign n40357 = n40355 & ~n40356 ;
  assign n40358 = n8372 | n23467 ;
  assign n40359 = ~n15833 & n23106 ;
  assign n40360 = n7515 & n25883 ;
  assign n40361 = n28677 ^ n22162 ^ 1'b0 ;
  assign n40362 = n25341 & ~n31578 ;
  assign n40363 = n5499 ^ n4619 ^ 1'b0 ;
  assign n40364 = n20714 & n40363 ;
  assign n40365 = n40364 ^ n20987 ^ n13949 ;
  assign n40366 = ( n2256 & n14422 ) | ( n2256 & n35576 ) | ( n14422 & n35576 ) ;
  assign n40367 = ( n2746 & n40365 ) | ( n2746 & n40366 ) | ( n40365 & n40366 ) ;
  assign n40368 = n14531 ^ n5975 ^ n1874 ;
  assign n40369 = ( n8657 & n13710 ) | ( n8657 & n40368 ) | ( n13710 & n40368 ) ;
  assign n40370 = n38826 | n40369 ;
  assign n40371 = n22681 & ~n40370 ;
  assign n40372 = ~n3970 & n12299 ;
  assign n40373 = ~n39778 & n40372 ;
  assign n40374 = n4090 & n8440 ;
  assign n40375 = n7173 ^ n5777 ^ n1755 ;
  assign n40376 = n40375 ^ n38811 ^ n15546 ;
  assign n40377 = n25097 ^ n12850 ^ n8051 ;
  assign n40378 = n13340 ^ n11301 ^ n7299 ;
  assign n40379 = ( ~n522 & n6926 ) | ( ~n522 & n28241 ) | ( n6926 & n28241 ) ;
  assign n40380 = ( n20335 & ~n40378 ) | ( n20335 & n40379 ) | ( ~n40378 & n40379 ) ;
  assign n40381 = n13158 ^ n8769 ^ 1'b0 ;
  assign n40384 = ~n509 & n10900 ;
  assign n40385 = n40384 ^ n12458 ^ 1'b0 ;
  assign n40382 = n1701 ^ n881 ^ 1'b0 ;
  assign n40383 = n37971 & ~n40382 ;
  assign n40386 = n40385 ^ n40383 ^ n23847 ;
  assign n40387 = ~n29961 & n32001 ;
  assign n40388 = ~n40386 & n40387 ;
  assign n40389 = n16294 | n18353 ;
  assign n40390 = n12120 & n40389 ;
  assign n40391 = n27321 & ~n40390 ;
  assign n40392 = n16688 & ~n22062 ;
  assign n40393 = n40392 ^ n26437 ^ 1'b0 ;
  assign n40394 = n31824 & n40393 ;
  assign n40395 = ~n8991 & n40394 ;
  assign n40396 = ( n7739 & n31796 ) | ( n7739 & ~n40395 ) | ( n31796 & ~n40395 ) ;
  assign n40398 = ~n11202 & n29742 ;
  assign n40399 = n11202 & n40398 ;
  assign n40397 = n28754 | n31193 ;
  assign n40400 = n40399 ^ n40397 ^ n14721 ;
  assign n40401 = n40396 & n40400 ;
  assign n40402 = n6191 | n12638 ;
  assign n40403 = n37891 ^ n35234 ^ n34751 ;
  assign n40404 = n10662 ^ n9296 ^ 1'b0 ;
  assign n40405 = n9181 & n40404 ;
  assign n40406 = n40405 ^ n3640 ^ 1'b0 ;
  assign n40407 = ( n8381 & ~n20702 ) | ( n8381 & n40406 ) | ( ~n20702 & n40406 ) ;
  assign n40408 = n10888 | n20719 ;
  assign n40409 = n2374 & ~n40408 ;
  assign n40410 = n29921 & ~n40409 ;
  assign n40411 = n3960 & n12975 ;
  assign n40412 = ~n8930 & n40411 ;
  assign n40413 = ~n25316 & n40412 ;
  assign n40414 = ~n34479 & n38358 ;
  assign n40415 = n19078 | n39243 ;
  assign n40416 = n6667 | n40415 ;
  assign n40417 = ~n26749 & n32719 ;
  assign n40418 = n17820 & ~n25894 ;
  assign n40419 = ( n3607 & n23310 ) | ( n3607 & ~n40418 ) | ( n23310 & ~n40418 ) ;
  assign n40420 = n40419 ^ n10060 ^ n6976 ;
  assign n40421 = n25924 & n27727 ;
  assign n40422 = n40421 ^ n537 ^ 1'b0 ;
  assign n40423 = n7578 ^ n4203 ^ 1'b0 ;
  assign n40424 = ~n13635 & n19523 ;
  assign n40425 = n40424 ^ n10201 ^ 1'b0 ;
  assign n40426 = ( n9939 & n40423 ) | ( n9939 & ~n40425 ) | ( n40423 & ~n40425 ) ;
  assign n40427 = n19848 | n32904 ;
  assign n40428 = n21238 & ~n40427 ;
  assign n40429 = n9887 & n35858 ;
  assign n40430 = n40429 ^ n31081 ^ 1'b0 ;
  assign n40431 = ~n17885 & n40430 ;
  assign n40432 = n30019 ^ n29660 ^ n1142 ;
  assign n40433 = n32349 ^ n10055 ^ n6305 ;
  assign n40436 = ( x213 & ~n1732 ) | ( x213 & n4214 ) | ( ~n1732 & n4214 ) ;
  assign n40434 = ~n18809 & n24911 ;
  assign n40435 = n40434 ^ n32182 ^ 1'b0 ;
  assign n40437 = n40436 ^ n40435 ^ n6339 ;
  assign n40438 = n6533 & ~n12718 ;
  assign n40439 = n40438 ^ n10232 ^ 1'b0 ;
  assign n40440 = n13559 & n40439 ;
  assign n40441 = n40440 ^ n28767 ^ n16548 ;
  assign n40445 = n18785 ^ n3316 ^ 1'b0 ;
  assign n40446 = n9358 & n40445 ;
  assign n40447 = n24362 & n40446 ;
  assign n40442 = n14758 & n29083 ;
  assign n40443 = ~n18805 & n40442 ;
  assign n40444 = n7668 & ~n40443 ;
  assign n40448 = n40447 ^ n40444 ^ 1'b0 ;
  assign n40449 = n898 | n13754 ;
  assign n40450 = n25078 | n40449 ;
  assign n40451 = ( ~n17035 & n21506 ) | ( ~n17035 & n36248 ) | ( n21506 & n36248 ) ;
  assign n40452 = ( n3247 & n36128 ) | ( n3247 & n37549 ) | ( n36128 & n37549 ) ;
  assign n40453 = n26289 ^ n4024 ^ 1'b0 ;
  assign n40456 = n14651 ^ n12587 ^ 1'b0 ;
  assign n40454 = n10360 & n21474 ;
  assign n40455 = ~n7296 & n40454 ;
  assign n40457 = n40456 ^ n40455 ^ n15183 ;
  assign n40458 = n22459 ^ n1626 ^ 1'b0 ;
  assign n40459 = ~n28494 & n40458 ;
  assign n40460 = n40459 ^ n10366 ^ 1'b0 ;
  assign n40461 = n27602 | n40460 ;
  assign n40462 = n39102 ^ n16929 ^ 1'b0 ;
  assign n40463 = ~n40461 & n40462 ;
  assign n40464 = n2311 & n2391 ;
  assign n40465 = ~n26953 & n40464 ;
  assign n40466 = n16193 ^ n1638 ^ 1'b0 ;
  assign n40467 = n2441 | n40466 ;
  assign n40468 = n8407 | n40467 ;
  assign n40470 = n17030 ^ n6082 ^ 1'b0 ;
  assign n40471 = n28502 | n40470 ;
  assign n40469 = ( n11184 & ~n13478 ) | ( n11184 & n36125 ) | ( ~n13478 & n36125 ) ;
  assign n40472 = n40471 ^ n40469 ^ n8183 ;
  assign n40473 = n844 & ~n12792 ;
  assign n40474 = n40473 ^ n5050 ^ 1'b0 ;
  assign n40475 = n20157 | n40474 ;
  assign n40476 = n40475 ^ n15493 ^ n8559 ;
  assign n40477 = n40476 ^ n8744 ^ 1'b0 ;
  assign n40478 = ~n33778 & n40264 ;
  assign n40479 = n11017 & n16032 ;
  assign n40480 = ~n21206 & n40479 ;
  assign n40481 = ( n263 & n16071 ) | ( n263 & ~n23455 ) | ( n16071 & ~n23455 ) ;
  assign n40482 = n40481 ^ n10825 ^ n9783 ;
  assign n40483 = n40482 ^ n10511 ^ 1'b0 ;
  assign n40484 = n18312 & n40483 ;
  assign n40485 = n27217 ^ n9746 ^ 1'b0 ;
  assign n40486 = ~x209 & n40485 ;
  assign n40487 = n4157 & ~n8177 ;
  assign n40488 = n40487 ^ n18748 ^ 1'b0 ;
  assign n40489 = x250 & ~n40488 ;
  assign n40490 = n40489 ^ n19737 ^ n5230 ;
  assign n40491 = n29831 ^ n17912 ^ 1'b0 ;
  assign n40492 = n5681 & n40491 ;
  assign n40493 = n40490 & n40492 ;
  assign n40494 = n27617 ^ n8937 ^ n6147 ;
  assign n40495 = n1877 | n30982 ;
  assign n40496 = n38892 & ~n40027 ;
  assign n40497 = n40496 ^ n3766 ^ 1'b0 ;
  assign n40498 = n1243 | n34602 ;
  assign n40499 = n9086 | n40498 ;
  assign n40500 = n40499 ^ n18486 ^ n10886 ;
  assign n40501 = n7001 & n40500 ;
  assign n40502 = n40501 ^ n1365 ^ 1'b0 ;
  assign n40503 = n2064 & n9902 ;
  assign n40504 = n27810 ^ n22624 ^ n4824 ;
  assign n40505 = n40027 & n40504 ;
  assign n40506 = n38907 ^ n10067 ^ 1'b0 ;
  assign n40507 = n15520 & ~n40506 ;
  assign n40508 = x109 & ~n22918 ;
  assign n40509 = n40508 ^ n599 ^ 1'b0 ;
  assign n40510 = ~n15654 & n40022 ;
  assign n40511 = n40510 ^ n26546 ^ 1'b0 ;
  assign n40512 = ~n17355 & n40511 ;
  assign n40513 = n40512 ^ n38978 ^ n32908 ;
  assign n40514 = ~n8460 & n19587 ;
  assign n40515 = n40514 ^ n27387 ^ 1'b0 ;
  assign n40516 = ( ~n7546 & n13685 ) | ( ~n7546 & n40515 ) | ( n13685 & n40515 ) ;
  assign n40517 = ( n1965 & n22728 ) | ( n1965 & ~n40516 ) | ( n22728 & ~n40516 ) ;
  assign n40518 = n30891 | n33752 ;
  assign n40519 = n14760 & ~n28643 ;
  assign n40520 = n14600 & n40519 ;
  assign n40521 = n407 & ~n37337 ;
  assign n40522 = n34099 & n40521 ;
  assign n40524 = ( ~n6549 & n21202 ) | ( ~n6549 & n30427 ) | ( n21202 & n30427 ) ;
  assign n40525 = n35056 | n40524 ;
  assign n40523 = n22387 | n25606 ;
  assign n40526 = n40525 ^ n40523 ^ 1'b0 ;
  assign n40527 = ( ~n11410 & n28379 ) | ( ~n11410 & n33070 ) | ( n28379 & n33070 ) ;
  assign n40528 = n40527 ^ n37051 ^ n37015 ;
  assign n40529 = n33823 & n40528 ;
  assign n40530 = ( ~n12196 & n13920 ) | ( ~n12196 & n31278 ) | ( n13920 & n31278 ) ;
  assign n40531 = ~n27774 & n40530 ;
  assign n40532 = n13411 & n40531 ;
  assign n40533 = n576 | n14654 ;
  assign n40534 = n36824 & n40533 ;
  assign n40535 = ~n23469 & n40534 ;
  assign n40536 = ( n37586 & n40532 ) | ( n37586 & ~n40535 ) | ( n40532 & ~n40535 ) ;
  assign n40537 = ~n25296 & n28412 ;
  assign n40538 = ~n29983 & n40537 ;
  assign n40539 = ( ~n2685 & n13513 ) | ( ~n2685 & n18824 ) | ( n13513 & n18824 ) ;
  assign n40540 = n23905 & n40539 ;
  assign n40541 = ( n892 & n17002 ) | ( n892 & n40540 ) | ( n17002 & n40540 ) ;
  assign n40542 = n31768 ^ n19484 ^ 1'b0 ;
  assign n40543 = n40542 ^ n22523 ^ n8322 ;
  assign n40544 = ~n3175 & n26499 ;
  assign n40545 = n40544 ^ n16521 ^ 1'b0 ;
  assign n40546 = n11056 | n27328 ;
  assign n40547 = n1733 & ~n40546 ;
  assign n40548 = n18190 | n40547 ;
  assign n40549 = n27222 ^ n2083 ^ 1'b0 ;
  assign n40550 = ~n5106 & n40549 ;
  assign n40551 = n40548 & n40550 ;
  assign n40552 = n40551 ^ n13040 ^ 1'b0 ;
  assign n40553 = n9653 | n11146 ;
  assign n40554 = n4844 | n40553 ;
  assign n40555 = ( ~n7985 & n15179 ) | ( ~n7985 & n40554 ) | ( n15179 & n40554 ) ;
  assign n40556 = n40555 ^ n33557 ^ 1'b0 ;
  assign n40557 = n13779 | n40556 ;
  assign n40558 = n31141 ^ n15694 ^ n868 ;
  assign n40559 = ( n2106 & n7005 ) | ( n2106 & ~n15986 ) | ( n7005 & ~n15986 ) ;
  assign n40560 = n5601 ^ n2125 ^ 1'b0 ;
  assign n40561 = n1329 & n40560 ;
  assign n40562 = n40561 ^ n21971 ^ n1818 ;
  assign n40563 = ( n12094 & ~n26657 ) | ( n12094 & n40562 ) | ( ~n26657 & n40562 ) ;
  assign n40564 = n561 | n3142 ;
  assign n40565 = n40564 ^ n29898 ^ n13618 ;
  assign n40566 = n3447 | n20671 ;
  assign n40567 = ( n9879 & n19004 ) | ( n9879 & n40566 ) | ( n19004 & n40566 ) ;
  assign n40568 = n7130 & ~n21897 ;
  assign n40569 = ~n7494 & n28133 ;
  assign n40570 = n40569 ^ n8887 ^ 1'b0 ;
  assign n40571 = ( ~n2208 & n3777 ) | ( ~n2208 & n36926 ) | ( n3777 & n36926 ) ;
  assign n40572 = n279 | n40571 ;
  assign n40573 = ~n6353 & n18229 ;
  assign n40574 = ~n40572 & n40573 ;
  assign n40575 = n7496 & n23841 ;
  assign n40576 = n21156 & ~n38230 ;
  assign n40577 = n5586 | n21834 ;
  assign n40578 = n3154 & ~n40577 ;
  assign n40580 = n27119 ^ n15273 ^ 1'b0 ;
  assign n40581 = ~n38368 & n40580 ;
  assign n40579 = n1744 | n24770 ;
  assign n40582 = n40581 ^ n40579 ^ 1'b0 ;
  assign n40583 = n14148 ^ n7566 ^ n2255 ;
  assign n40584 = n40583 ^ n1781 ^ 1'b0 ;
  assign n40585 = n4625 & ~n13943 ;
  assign n40586 = n40585 ^ n21349 ^ 1'b0 ;
  assign n40589 = n26415 ^ n5766 ^ 1'b0 ;
  assign n40587 = n4039 | n15610 ;
  assign n40588 = n5904 | n40587 ;
  assign n40590 = n40589 ^ n40588 ^ n8667 ;
  assign n40591 = n13857 | n16473 ;
  assign n40592 = ( n2690 & n9207 ) | ( n2690 & n9419 ) | ( n9207 & n9419 ) ;
  assign n40593 = n385 & ~n538 ;
  assign n40594 = n40593 ^ n8382 ^ 1'b0 ;
  assign n40595 = n8871 ^ n8746 ^ 1'b0 ;
  assign n40596 = ( n6669 & ~n29630 ) | ( n6669 & n40595 ) | ( ~n29630 & n40595 ) ;
  assign n40597 = n40596 ^ n39484 ^ 1'b0 ;
  assign n40598 = n17853 & ~n40597 ;
  assign n40599 = n699 & ~n1182 ;
  assign n40600 = n16409 & n30243 ;
  assign n40601 = n18010 ^ n12962 ^ 1'b0 ;
  assign n40602 = ( n11995 & ~n16478 ) | ( n11995 & n37861 ) | ( ~n16478 & n37861 ) ;
  assign n40604 = n2984 & n11791 ;
  assign n40605 = n40604 ^ n1283 ^ 1'b0 ;
  assign n40603 = n2974 & n24948 ;
  assign n40606 = n40605 ^ n40603 ^ 1'b0 ;
  assign n40607 = n40606 ^ n20836 ^ 1'b0 ;
  assign n40608 = n14672 & ~n30725 ;
  assign n40609 = n845 | n5578 ;
  assign n40610 = n16731 & ~n40609 ;
  assign n40611 = n9000 ^ n7779 ^ 1'b0 ;
  assign n40612 = n25304 & n39515 ;
  assign n40613 = n23340 ^ n500 ^ 1'b0 ;
  assign n40614 = n23893 & n40613 ;
  assign n40615 = n22309 ^ n18565 ^ n12716 ;
  assign n40616 = n40615 ^ n34214 ^ n21444 ;
  assign n40617 = n31286 & n40616 ;
  assign n40618 = ~n21717 & n26889 ;
  assign n40619 = n17452 ^ n13370 ^ n2403 ;
  assign n40620 = ( n32031 & n38450 ) | ( n32031 & ~n40619 ) | ( n38450 & ~n40619 ) ;
  assign n40621 = n19780 ^ n6771 ^ 1'b0 ;
  assign n40622 = n35087 & n40621 ;
  assign n40623 = n40622 ^ n3609 ^ 1'b0 ;
  assign n40624 = ( n2419 & ~n24088 ) | ( n2419 & n40623 ) | ( ~n24088 & n40623 ) ;
  assign n40625 = ~n23636 & n40624 ;
  assign n40626 = n25765 ^ n11390 ^ 1'b0 ;
  assign n40627 = n7901 & ~n40626 ;
  assign n40628 = n295 & n2833 ;
  assign n40629 = n40628 ^ n40044 ^ 1'b0 ;
  assign n40630 = n13770 ^ n6845 ^ 1'b0 ;
  assign n40631 = n24796 ^ n10134 ^ 1'b0 ;
  assign n40632 = ( n7161 & ~n11838 ) | ( n7161 & n14556 ) | ( ~n11838 & n14556 ) ;
  assign n40633 = x253 & n12807 ;
  assign n40634 = n40633 ^ n10782 ^ 1'b0 ;
  assign n40635 = ( n362 & n26718 ) | ( n362 & n40634 ) | ( n26718 & n40634 ) ;
  assign n40636 = n20386 ^ n18034 ^ n5141 ;
  assign n40637 = n40636 ^ n36182 ^ n33342 ;
  assign n40638 = n3379 | n7855 ;
  assign n40639 = n9312 | n40638 ;
  assign n40640 = n40639 ^ n496 ^ 1'b0 ;
  assign n40642 = ~n4371 & n23447 ;
  assign n40641 = n6268 & n17288 ;
  assign n40643 = n40642 ^ n40641 ^ 1'b0 ;
  assign n40645 = n9253 ^ n2911 ^ 1'b0 ;
  assign n40644 = n7296 & ~n31167 ;
  assign n40646 = n40645 ^ n40644 ^ 1'b0 ;
  assign n40647 = ( n8679 & ~n18683 ) | ( n8679 & n25319 ) | ( ~n18683 & n25319 ) ;
  assign n40648 = n13796 | n20403 ;
  assign n40649 = n40648 ^ n11822 ^ 1'b0 ;
  assign n40650 = ~n7402 & n19587 ;
  assign n40651 = ~n7210 & n40650 ;
  assign n40652 = n9485 ^ n3900 ^ 1'b0 ;
  assign n40653 = n40651 | n40652 ;
  assign n40654 = ( n12971 & ~n40649 ) | ( n12971 & n40653 ) | ( ~n40649 & n40653 ) ;
  assign n40655 = n11940 ^ n3937 ^ 1'b0 ;
  assign n40656 = ~n19421 & n40655 ;
  assign n40657 = ( n19302 & n33848 ) | ( n19302 & ~n40656 ) | ( n33848 & ~n40656 ) ;
  assign n40658 = n27895 & ~n36116 ;
  assign n40659 = n19017 ^ n2830 ^ 1'b0 ;
  assign n40660 = n18897 | n40659 ;
  assign n40661 = n33138 & ~n40660 ;
  assign n40662 = n1028 | n32166 ;
  assign n40663 = ~n12779 & n40662 ;
  assign n40664 = n6438 ^ n3693 ^ 1'b0 ;
  assign n40665 = n17894 | n40664 ;
  assign n40668 = n25258 ^ n2262 ^ 1'b0 ;
  assign n40669 = n9806 & ~n40668 ;
  assign n40667 = n27740 ^ n27672 ^ 1'b0 ;
  assign n40666 = n31978 ^ n22015 ^ 1'b0 ;
  assign n40670 = n40669 ^ n40667 ^ n40666 ;
  assign n40671 = n1194 & ~n40670 ;
  assign n40672 = n13310 & n40671 ;
  assign n40673 = n1083 & ~n6337 ;
  assign n40674 = ( ~n17072 & n25718 ) | ( ~n17072 & n40673 ) | ( n25718 & n40673 ) ;
  assign n40675 = ( n1060 & n6619 ) | ( n1060 & ~n40674 ) | ( n6619 & ~n40674 ) ;
  assign n40676 = n14193 & n30356 ;
  assign n40677 = n20874 ^ n9485 ^ 1'b0 ;
  assign n40678 = n27783 | n40677 ;
  assign n40679 = n40678 ^ n12993 ^ n2786 ;
  assign n40680 = ~n3666 & n10096 ;
  assign n40681 = n40680 ^ n4111 ^ 1'b0 ;
  assign n40682 = ~n4117 & n5144 ;
  assign n40683 = n30542 & ~n40682 ;
  assign n40685 = n23992 ^ n15964 ^ 1'b0 ;
  assign n40686 = ~n3391 & n40685 ;
  assign n40684 = n3053 | n22483 ;
  assign n40687 = n40686 ^ n40684 ^ 1'b0 ;
  assign n40689 = ~n7417 & n14309 ;
  assign n40690 = ~n5475 & n40689 ;
  assign n40688 = n3798 ^ n2724 ^ 1'b0 ;
  assign n40691 = n40690 ^ n40688 ^ n14726 ;
  assign n40692 = n6468 | n21822 ;
  assign n40693 = n40692 ^ n15304 ^ 1'b0 ;
  assign n40694 = n30124 ^ n6008 ^ 1'b0 ;
  assign n40695 = n13505 | n40694 ;
  assign n40696 = n991 & ~n33026 ;
  assign n40697 = ~n40695 & n40696 ;
  assign n40698 = ( ~n8545 & n40693 ) | ( ~n8545 & n40697 ) | ( n40693 & n40697 ) ;
  assign n40699 = n33929 ^ n23534 ^ 1'b0 ;
  assign n40700 = ( n14358 & n31309 ) | ( n14358 & ~n40699 ) | ( n31309 & ~n40699 ) ;
  assign n40701 = n8955 ^ x233 ^ 1'b0 ;
  assign n40702 = n4653 | n14646 ;
  assign n40703 = n9316 & ~n28733 ;
  assign n40704 = ~x15 & n40703 ;
  assign n40705 = n40088 ^ n38726 ^ 1'b0 ;
  assign n40706 = n30874 & n40705 ;
  assign n40707 = x90 & ~n8713 ;
  assign n40708 = n40707 ^ n22720 ^ 1'b0 ;
  assign n40709 = n21692 & n27291 ;
  assign n40710 = ~n40708 & n40709 ;
  assign n40711 = n40710 ^ n7880 ^ n1999 ;
  assign n40712 = n10094 & ~n27902 ;
  assign n40713 = n4347 ^ n1781 ^ 1'b0 ;
  assign n40714 = n14277 & ~n40713 ;
  assign n40715 = n40714 ^ n13481 ^ n2021 ;
  assign n40716 = n13513 ^ n5359 ^ 1'b0 ;
  assign n40717 = ~n30498 & n40716 ;
  assign n40718 = ~n2650 & n40717 ;
  assign n40719 = ~n2352 & n30557 ;
  assign n40720 = ~n14775 & n30476 ;
  assign n40721 = x134 ^ x90 ^ 1'b0 ;
  assign n40722 = n40721 ^ n10030 ^ n8057 ;
  assign n40723 = ( n4197 & ~n6783 ) | ( n4197 & n21711 ) | ( ~n6783 & n21711 ) ;
  assign n40724 = n20588 ^ n13310 ^ 1'b0 ;
  assign n40725 = n10597 | n40724 ;
  assign n40726 = ( n27509 & n37852 ) | ( n27509 & n38386 ) | ( n37852 & n38386 ) ;
  assign n40727 = n27075 ^ n2461 ^ n1496 ;
  assign n40728 = ( ~x183 & n3107 ) | ( ~x183 & n21875 ) | ( n3107 & n21875 ) ;
  assign n40729 = n2479 & ~n40728 ;
  assign n40730 = n40727 & n40729 ;
  assign n40731 = n15346 | n35659 ;
  assign n40732 = n40731 ^ n3945 ^ 1'b0 ;
  assign n40733 = n24953 ^ n3854 ^ 1'b0 ;
  assign n40734 = n36876 ^ n29218 ^ 1'b0 ;
  assign n40736 = n545 ^ x180 ^ 1'b0 ;
  assign n40737 = n40736 ^ n7431 ^ 1'b0 ;
  assign n40738 = n14670 & ~n40737 ;
  assign n40735 = n5685 | n17161 ;
  assign n40739 = n40738 ^ n40735 ^ n12252 ;
  assign n40740 = ( n2412 & n25688 ) | ( n2412 & ~n32125 ) | ( n25688 & ~n32125 ) ;
  assign n40741 = n40740 ^ n6351 ^ n1638 ;
  assign n40742 = n19821 ^ n6513 ^ n384 ;
  assign n40743 = n9764 | n40742 ;
  assign n40744 = n40743 ^ n11723 ^ 1'b0 ;
  assign n40745 = n29717 & ~n35967 ;
  assign n40746 = ( n1040 & ~n6430 ) | ( n1040 & n21343 ) | ( ~n6430 & n21343 ) ;
  assign n40747 = ( n1987 & n7813 ) | ( n1987 & n13515 ) | ( n7813 & n13515 ) ;
  assign n40748 = n40747 ^ n12897 ^ n1722 ;
  assign n40749 = n21146 | n33995 ;
  assign n40750 = n3210 & ~n40749 ;
  assign n40751 = n25719 ^ n15615 ^ 1'b0 ;
  assign n40752 = n10754 & n40751 ;
  assign n40753 = n12024 & ~n21595 ;
  assign n40754 = ~n7803 & n27415 ;
  assign n40755 = n40753 & n40754 ;
  assign n40756 = n12487 ^ n12131 ^ 1'b0 ;
  assign n40757 = n40756 ^ n32947 ^ 1'b0 ;
  assign n40758 = n20755 & ~n23647 ;
  assign n40759 = ~n34225 & n40758 ;
  assign n40760 = n8650 | n40759 ;
  assign n40761 = n425 & n5269 ;
  assign n40762 = n40761 ^ n24768 ^ 1'b0 ;
  assign n40763 = ( ~n3024 & n10992 ) | ( ~n3024 & n40762 ) | ( n10992 & n40762 ) ;
  assign n40764 = n15329 & ~n22430 ;
  assign n40765 = n40764 ^ n29802 ^ 1'b0 ;
  assign n40766 = n40765 ^ n15686 ^ n15168 ;
  assign n40767 = n38577 ^ n38204 ^ 1'b0 ;
  assign n40768 = n40766 & ~n40767 ;
  assign n40769 = n40768 ^ n26265 ^ 1'b0 ;
  assign n40770 = n3333 & n8774 ;
  assign n40771 = n40770 ^ n33742 ^ 1'b0 ;
  assign n40772 = n17847 ^ n14929 ^ 1'b0 ;
  assign n40773 = n16824 & n40772 ;
  assign n40774 = ~n30058 & n40773 ;
  assign n40775 = ~n37517 & n40774 ;
  assign n40776 = n4678 & n24223 ;
  assign n40777 = n16236 | n19843 ;
  assign n40778 = ( n5174 & n19568 ) | ( n5174 & n38192 ) | ( n19568 & n38192 ) ;
  assign n40779 = ~n11000 & n15787 ;
  assign n40780 = n15508 & ~n15901 ;
  assign n40781 = ~n13885 & n40780 ;
  assign n40782 = ~n4237 & n20535 ;
  assign n40783 = n8597 & n40782 ;
  assign n40784 = ~n11286 & n30431 ;
  assign n40785 = n40783 & n40784 ;
  assign n40786 = n30472 ^ n19688 ^ 1'b0 ;
  assign n40787 = n6284 & ~n40786 ;
  assign n40788 = n10053 & n20643 ;
  assign n40789 = n3080 | n4817 ;
  assign n40790 = n28727 ^ n14845 ^ 1'b0 ;
  assign n40791 = ~n40789 & n40790 ;
  assign n40792 = n6898 & ~n17390 ;
  assign n40793 = ( ~n9644 & n28678 ) | ( ~n9644 & n33461 ) | ( n28678 & n33461 ) ;
  assign n40794 = n35167 ^ n5112 ^ 1'b0 ;
  assign n40795 = ~n5359 & n10193 ;
  assign n40796 = n8047 & n26202 ;
  assign n40797 = n40796 ^ n27984 ^ 1'b0 ;
  assign n40798 = n1080 & n2317 ;
  assign n40799 = ~n6752 & n8431 ;
  assign n40800 = n40799 ^ n24872 ^ 1'b0 ;
  assign n40801 = n40798 & n40800 ;
  assign n40802 = n39816 ^ n39271 ^ 1'b0 ;
  assign n40803 = ( ~n1701 & n5078 ) | ( ~n1701 & n14473 ) | ( n5078 & n14473 ) ;
  assign n40804 = ~n25927 & n40803 ;
  assign n40805 = n31061 ^ n12265 ^ 1'b0 ;
  assign n40806 = n21835 ^ n14726 ^ n12997 ;
  assign n40807 = ( ~n17740 & n40805 ) | ( ~n17740 & n40806 ) | ( n40805 & n40806 ) ;
  assign n40808 = n15921 ^ n4444 ^ 1'b0 ;
  assign n40809 = n3047 ^ n1780 ^ 1'b0 ;
  assign n40810 = n26993 & ~n40809 ;
  assign n40811 = n19869 ^ n968 ^ 1'b0 ;
  assign n40812 = n3011 | n40811 ;
  assign n40813 = n40810 | n40812 ;
  assign n40814 = n7326 & ~n32622 ;
  assign n40815 = ~n40813 & n40814 ;
  assign n40816 = n34503 ^ n27842 ^ 1'b0 ;
  assign n40817 = n17665 & ~n40816 ;
  assign n40818 = ~n19540 & n40817 ;
  assign n40819 = ( n9266 & n17338 ) | ( n9266 & ~n29339 ) | ( n17338 & ~n29339 ) ;
  assign n40820 = n5387 & n12138 ;
  assign n40821 = n21365 & n33926 ;
  assign n40822 = n23412 & ~n40821 ;
  assign n40823 = n40822 ^ n6960 ^ 1'b0 ;
  assign n40824 = n33352 & n38539 ;
  assign n40825 = ~n8117 & n40824 ;
  assign n40826 = n17825 ^ n16406 ^ 1'b0 ;
  assign n40827 = n18335 | n40826 ;
  assign n40828 = n40827 ^ n14286 ^ x116 ;
  assign n40829 = n5374 & ~n40828 ;
  assign n40830 = n15893 & n37410 ;
  assign n40831 = n40830 ^ n12297 ^ n2095 ;
  assign n40832 = ~n905 & n10194 ;
  assign n40833 = n375 & n40832 ;
  assign n40834 = n6747 & ~n40833 ;
  assign n40835 = ~n19138 & n40834 ;
  assign n40836 = n40835 ^ n13949 ^ 1'b0 ;
  assign n40837 = n40831 & n40836 ;
  assign n40838 = x230 & ~n30267 ;
  assign n40839 = n40838 ^ n17452 ^ 1'b0 ;
  assign n40840 = n40839 ^ n18994 ^ 1'b0 ;
  assign n40844 = ~n6619 & n9586 ;
  assign n40845 = n40844 ^ n13398 ^ 1'b0 ;
  assign n40846 = n40845 ^ n30221 ^ n4493 ;
  assign n40841 = n3161 ^ n966 ^ 1'b0 ;
  assign n40842 = n36552 & n40841 ;
  assign n40843 = n21101 | n40842 ;
  assign n40847 = n40846 ^ n40843 ^ n5014 ;
  assign n40848 = ( ~n4314 & n26152 ) | ( ~n4314 & n40847 ) | ( n26152 & n40847 ) ;
  assign n40849 = n8043 | n15826 ;
  assign n40850 = n6256 & ~n40849 ;
  assign n40851 = n3115 & ~n40850 ;
  assign n40852 = n40851 ^ n37864 ^ 1'b0 ;
  assign n40853 = ~n2859 & n10738 ;
  assign n40854 = ~n40852 & n40853 ;
  assign n40856 = n6645 & ~n8939 ;
  assign n40857 = n40856 ^ n32349 ^ 1'b0 ;
  assign n40855 = n7308 & ~n17319 ;
  assign n40858 = n40857 ^ n40855 ^ 1'b0 ;
  assign n40859 = ~n29118 & n29415 ;
  assign n40860 = ~n2744 & n40859 ;
  assign n40861 = n17076 ^ n10934 ^ 1'b0 ;
  assign n40863 = n7720 ^ n6732 ^ 1'b0 ;
  assign n40862 = n14722 | n23403 ;
  assign n40864 = n40863 ^ n40862 ^ 1'b0 ;
  assign n40865 = n12249 ^ n11426 ^ 1'b0 ;
  assign n40866 = n4313 & ~n40865 ;
  assign n40867 = ( n40861 & ~n40864 ) | ( n40861 & n40866 ) | ( ~n40864 & n40866 ) ;
  assign n40868 = n25386 ^ n15734 ^ 1'b0 ;
  assign n40869 = ~n38670 & n40868 ;
  assign n40870 = ( n1701 & n29562 ) | ( n1701 & ~n40869 ) | ( n29562 & ~n40869 ) ;
  assign n40871 = n40870 ^ n37944 ^ 1'b0 ;
  assign n40872 = ( ~n1275 & n2680 ) | ( ~n1275 & n40871 ) | ( n2680 & n40871 ) ;
  assign n40873 = n22513 & ~n31378 ;
  assign n40874 = n19760 ^ n11266 ^ n4939 ;
  assign n40875 = n30518 ^ n29319 ^ 1'b0 ;
  assign n40876 = ~n24968 & n40875 ;
  assign n40877 = n40874 & n40876 ;
  assign n40878 = n40877 ^ n11805 ^ 1'b0 ;
  assign n40879 = n7521 | n40878 ;
  assign n40880 = ( n287 & n5798 ) | ( n287 & n15348 ) | ( n5798 & n15348 ) ;
  assign n40881 = n40880 ^ n26103 ^ n15436 ;
  assign n40882 = n22128 ^ n19258 ^ n5935 ;
  assign n40883 = n40882 ^ n11984 ^ 1'b0 ;
  assign n40884 = n22132 | n38668 ;
  assign n40885 = n3768 & ~n28136 ;
  assign n40886 = n2906 | n40885 ;
  assign n40887 = ( ~n1962 & n16363 ) | ( ~n1962 & n34447 ) | ( n16363 & n34447 ) ;
  assign n40888 = n40887 ^ n30377 ^ 1'b0 ;
  assign n40889 = n31877 & ~n40888 ;
  assign n40890 = n23106 ^ n6041 ^ 1'b0 ;
  assign n40891 = n11135 & n40890 ;
  assign n40892 = ~n10259 & n13643 ;
  assign n40893 = n36031 & ~n40892 ;
  assign n40894 = n40893 ^ n22297 ^ 1'b0 ;
  assign n40895 = n11169 & ~n11363 ;
  assign n40896 = n23040 & n37075 ;
  assign n40897 = ( n30284 & ~n40895 ) | ( n30284 & n40896 ) | ( ~n40895 & n40896 ) ;
  assign n40900 = n15881 ^ n10830 ^ 1'b0 ;
  assign n40898 = ~n3379 & n28735 ;
  assign n40899 = n40898 ^ n24685 ^ 1'b0 ;
  assign n40901 = n40900 ^ n40899 ^ n15746 ;
  assign n40902 = ~n1063 & n32688 ;
  assign n40903 = n23073 & n40902 ;
  assign n40904 = n1899 & n40903 ;
  assign n40905 = n31209 ^ n4371 ^ 1'b0 ;
  assign n40906 = n1720 & ~n7364 ;
  assign n40907 = n40906 ^ n7282 ^ 1'b0 ;
  assign n40909 = n5780 ^ n5012 ^ 1'b0 ;
  assign n40910 = n5287 & n40909 ;
  assign n40908 = n24053 ^ n20546 ^ n7358 ;
  assign n40911 = n40910 ^ n40908 ^ 1'b0 ;
  assign n40912 = x242 & n17372 ;
  assign n40913 = ~n7347 & n40912 ;
  assign n40914 = ( n13677 & ~n20271 ) | ( n13677 & n40913 ) | ( ~n20271 & n40913 ) ;
  assign n40915 = n36574 & ~n40914 ;
  assign n40916 = n15613 & n40915 ;
  assign n40917 = x225 & n16159 ;
  assign n40918 = n26509 ^ n5744 ^ 1'b0 ;
  assign n40919 = n26885 | n40918 ;
  assign n40920 = n11990 ^ n6958 ^ 1'b0 ;
  assign n40921 = ~n40919 & n40920 ;
  assign n40922 = n16066 & n19499 ;
  assign n40923 = ( n1906 & ~n9605 ) | ( n1906 & n24984 ) | ( ~n9605 & n24984 ) ;
  assign n40924 = n8498 & n10680 ;
  assign n40925 = n40924 ^ n9357 ^ 1'b0 ;
  assign n40926 = n40925 ^ n23900 ^ n3023 ;
  assign n40927 = n11470 & ~n40926 ;
  assign n40930 = n4489 & n16338 ;
  assign n40928 = n21875 ^ n4592 ^ 1'b0 ;
  assign n40929 = n28462 & n40928 ;
  assign n40931 = n40930 ^ n40929 ^ n20819 ;
  assign n40932 = n21676 | n34963 ;
  assign n40933 = n40932 ^ n9255 ^ 1'b0 ;
  assign n40934 = n17300 ^ n8303 ^ n5952 ;
  assign n40935 = n40934 ^ n33931 ^ n16679 ;
  assign n40936 = n10753 ^ n10636 ^ 1'b0 ;
  assign n40937 = n1399 & ~n8042 ;
  assign n40938 = n40937 ^ n21059 ^ 1'b0 ;
  assign n40939 = n15774 & ~n40938 ;
  assign n40940 = n522 & n794 ;
  assign n40941 = n40940 ^ n3726 ^ 1'b0 ;
  assign n40942 = n14176 ^ n11934 ^ 1'b0 ;
  assign n40943 = n28105 ^ n3181 ^ 1'b0 ;
  assign n40944 = n40943 ^ n40456 ^ 1'b0 ;
  assign n40945 = ~n8296 & n10190 ;
  assign n40946 = n6967 & n40945 ;
  assign n40947 = ( ~n4654 & n4835 ) | ( ~n4654 & n18463 ) | ( n4835 & n18463 ) ;
  assign n40948 = n40947 ^ n21473 ^ 1'b0 ;
  assign n40949 = n9622 ^ x196 ^ 1'b0 ;
  assign n40950 = n40949 ^ n11664 ^ 1'b0 ;
  assign n40951 = ~n15338 & n40950 ;
  assign n40952 = n5469 ^ n1047 ^ 1'b0 ;
  assign n40953 = n8348 & n40952 ;
  assign n40954 = ~n35170 & n40953 ;
  assign n40955 = ~n15174 & n40954 ;
  assign n40956 = ( n35587 & n40951 ) | ( n35587 & ~n40955 ) | ( n40951 & ~n40955 ) ;
  assign n40957 = n5578 | n7288 ;
  assign n40958 = n4950 & ~n40957 ;
  assign n40959 = n33977 & n40958 ;
  assign n40960 = n40959 ^ n4329 ^ 1'b0 ;
  assign n40961 = n22771 & n37241 ;
  assign n40962 = n28245 ^ n4947 ^ 1'b0 ;
  assign n40963 = n3318 | n40962 ;
  assign n40964 = n40963 ^ n2003 ^ 1'b0 ;
  assign n40965 = n2333 | n40964 ;
  assign n40966 = n35218 & ~n40965 ;
  assign n40967 = n16171 ^ n8980 ^ n8345 ;
  assign n40968 = n24370 ^ n15942 ^ n7639 ;
  assign n40969 = n3440 & n40968 ;
  assign n40970 = n40969 ^ n34760 ^ 1'b0 ;
  assign n40971 = ( n26808 & n36766 ) | ( n26808 & ~n40970 ) | ( n36766 & ~n40970 ) ;
  assign n40972 = ~n5165 & n9470 ;
  assign n40973 = n11910 & n40972 ;
  assign n40974 = ( n1671 & n15887 ) | ( n1671 & n40973 ) | ( n15887 & n40973 ) ;
  assign n40975 = ( n27970 & n34680 ) | ( n27970 & ~n40974 ) | ( n34680 & ~n40974 ) ;
  assign n40976 = n19728 ^ n13006 ^ 1'b0 ;
  assign n40977 = ~n9754 & n36031 ;
  assign n40978 = n3512 & ~n40977 ;
  assign n40979 = ~n9568 & n40978 ;
  assign n40980 = n19864 ^ n10675 ^ 1'b0 ;
  assign n40981 = n21135 | n40980 ;
  assign n40982 = ( ~n9687 & n27045 ) | ( ~n9687 & n30134 ) | ( n27045 & n30134 ) ;
  assign n40983 = ~n1012 & n33034 ;
  assign n40984 = n40983 ^ n35059 ^ n17401 ;
  assign n40985 = n30826 & n39825 ;
  assign n40986 = ~n33041 & n34722 ;
  assign n40987 = n13835 & n40760 ;
  assign n40988 = n19555 ^ n5108 ^ 1'b0 ;
  assign n40989 = n36693 | n40988 ;
  assign n40990 = n4618 ^ n4617 ^ 1'b0 ;
  assign n40991 = ~n1452 & n13810 ;
  assign n40992 = n5922 ^ n4858 ^ 1'b0 ;
  assign n40993 = ~n8247 & n40992 ;
  assign n40994 = ~n19501 & n40993 ;
  assign n40995 = n40994 ^ n17236 ^ n10123 ;
  assign n40996 = n12425 & n35246 ;
  assign n40997 = n40996 ^ n4118 ^ 1'b0 ;
  assign n40998 = n40997 ^ n32103 ^ 1'b0 ;
  assign n40999 = n13678 & ~n23290 ;
  assign n41000 = ( n2258 & n10060 ) | ( n2258 & n11279 ) | ( n10060 & n11279 ) ;
  assign n41006 = n18266 | n19864 ;
  assign n41003 = n1541 & n18764 ;
  assign n41004 = n16409 ^ n5436 ^ 1'b0 ;
  assign n41005 = n41003 & ~n41004 ;
  assign n41001 = n2342 | n5213 ;
  assign n41002 = n41001 ^ n15015 ^ n12906 ;
  assign n41007 = n41006 ^ n41005 ^ n41002 ;
  assign n41008 = n30118 ^ n10551 ^ 1'b0 ;
  assign n41009 = n9676 ^ n9515 ^ 1'b0 ;
  assign n41010 = ~n26907 & n41009 ;
  assign n41011 = n425 & ~n31047 ;
  assign n41012 = ~n41010 & n41011 ;
  assign n41013 = n17099 ^ n13388 ^ 1'b0 ;
  assign n41014 = n13500 & n41013 ;
  assign n41015 = ~n38187 & n41014 ;
  assign n41016 = n41012 & n41015 ;
  assign n41017 = n5119 & n38733 ;
  assign n41018 = n41017 ^ n23012 ^ 1'b0 ;
  assign n41019 = n28125 ^ n10298 ^ 1'b0 ;
  assign n41020 = n4228 & ~n41019 ;
  assign n41021 = n12244 ^ n939 ^ 1'b0 ;
  assign n41022 = n763 | n41021 ;
  assign n41023 = ( n2680 & n26986 ) | ( n2680 & n41022 ) | ( n26986 & n41022 ) ;
  assign n41024 = n9627 & n17242 ;
  assign n41025 = n41024 ^ n34474 ^ n547 ;
  assign n41026 = n10409 | n12624 ;
  assign n41027 = n41026 ^ n18735 ^ 1'b0 ;
  assign n41028 = n5011 ^ n3328 ^ 1'b0 ;
  assign n41029 = ~n41027 & n41028 ;
  assign n41030 = n12292 & n25279 ;
  assign n41031 = n41030 ^ n35142 ^ 1'b0 ;
  assign n41032 = n3180 & n16617 ;
  assign n41033 = ( ~n2349 & n5373 ) | ( ~n2349 & n7390 ) | ( n5373 & n7390 ) ;
  assign n41034 = n7784 ^ x200 ^ 1'b0 ;
  assign n41035 = n41034 ^ n39778 ^ n32049 ;
  assign n41036 = n547 & n4805 ;
  assign n41037 = n5551 & ~n10854 ;
  assign n41038 = n39738 ^ n8812 ^ 1'b0 ;
  assign n41039 = n41037 & n41038 ;
  assign n41040 = n10938 | n29647 ;
  assign n41041 = n37396 & ~n41040 ;
  assign n41042 = n19159 ^ n16964 ^ n2590 ;
  assign n41043 = n24318 ^ n14223 ^ 1'b0 ;
  assign n41044 = ~n41042 & n41043 ;
  assign n41046 = n8323 & ~n26334 ;
  assign n41045 = ~n2347 & n31619 ;
  assign n41047 = n41046 ^ n41045 ^ 1'b0 ;
  assign n41048 = n14200 & ~n34511 ;
  assign n41049 = n41048 ^ n10203 ^ 1'b0 ;
  assign n41050 = ( ~n10182 & n14761 ) | ( ~n10182 & n19390 ) | ( n14761 & n19390 ) ;
  assign n41051 = ( ~n15068 & n21333 ) | ( ~n15068 & n41050 ) | ( n21333 & n41050 ) ;
  assign n41052 = n41051 ^ n11469 ^ 1'b0 ;
  assign n41053 = ( ~n1690 & n2937 ) | ( ~n1690 & n16556 ) | ( n2937 & n16556 ) ;
  assign n41054 = n41053 ^ n34089 ^ n11380 ;
  assign n41055 = n4107 & n6418 ;
  assign n41056 = ~n30669 & n41055 ;
  assign n41057 = n41056 ^ n16140 ^ 1'b0 ;
  assign n41058 = ~n31993 & n41057 ;
  assign n41059 = n1882 & n24845 ;
  assign n41060 = n41059 ^ n10157 ^ 1'b0 ;
  assign n41061 = n16761 & n19393 ;
  assign n41062 = n17007 & n41061 ;
  assign n41063 = n41062 ^ n18858 ^ 1'b0 ;
  assign n41064 = n1671 & n41063 ;
  assign n41065 = ~n12562 & n18915 ;
  assign n41066 = ~n38031 & n41065 ;
  assign n41067 = ( n2622 & n41064 ) | ( n2622 & n41066 ) | ( n41064 & n41066 ) ;
  assign n41068 = n39203 & ~n41067 ;
  assign n41069 = n41068 ^ n33252 ^ 1'b0 ;
  assign n41070 = n22117 | n23551 ;
  assign n41071 = n13065 ^ n4260 ^ 1'b0 ;
  assign n41072 = n41071 ^ n15988 ^ 1'b0 ;
  assign n41073 = n29202 & n40440 ;
  assign n41074 = ~n405 & n41073 ;
  assign n41075 = n41072 & ~n41074 ;
  assign n41076 = n10645 & n36709 ;
  assign n41077 = ( n10514 & n23298 ) | ( n10514 & ~n41076 ) | ( n23298 & ~n41076 ) ;
  assign n41078 = ( n2619 & ~n8961 ) | ( n2619 & n17571 ) | ( ~n8961 & n17571 ) ;
  assign n41079 = n15342 & n34596 ;
  assign n41080 = n9928 & n10289 ;
  assign n41081 = n24928 & n41080 ;
  assign n41082 = n34529 | n41081 ;
  assign n41083 = n41082 ^ n5973 ^ 1'b0 ;
  assign n41084 = n20585 & n41083 ;
  assign n41085 = ( n4756 & n11982 ) | ( n4756 & n27783 ) | ( n11982 & n27783 ) ;
  assign n41086 = n9533 | n38904 ;
  assign n41087 = n3279 & n20554 ;
  assign n41088 = ~n5814 & n38015 ;
  assign n41089 = n41087 & n41088 ;
  assign n41090 = ( n16016 & n41086 ) | ( n16016 & n41089 ) | ( n41086 & n41089 ) ;
  assign n41091 = n38699 ^ n11412 ^ 1'b0 ;
  assign n41092 = ~n12587 & n41091 ;
  assign n41093 = n41092 ^ n1310 ^ 1'b0 ;
  assign n41094 = ~n41090 & n41093 ;
  assign n41095 = n12943 & n41094 ;
  assign n41096 = ( n18919 & n24473 ) | ( n18919 & n27667 ) | ( n24473 & n27667 ) ;
  assign n41097 = n29101 ^ n17275 ^ n5631 ;
  assign n41098 = n6411 | n41097 ;
  assign n41099 = n17311 | n28600 ;
  assign n41100 = n39644 | n41099 ;
  assign n41101 = n25819 & n32855 ;
  assign n41102 = n41101 ^ n30196 ^ 1'b0 ;
  assign n41103 = n24373 | n29401 ;
  assign n41104 = n17952 | n41103 ;
  assign n41105 = ( ~n19156 & n34235 ) | ( ~n19156 & n41104 ) | ( n34235 & n41104 ) ;
  assign n41106 = n36518 ^ n936 ^ 1'b0 ;
  assign n41107 = n41105 & ~n41106 ;
  assign n41108 = ~n9538 & n13035 ;
  assign n41109 = n20890 & n41108 ;
  assign n41110 = n28672 ^ n13380 ^ 1'b0 ;
  assign n41111 = n1613 & ~n41110 ;
  assign n41112 = n12476 & ~n16590 ;
  assign n41113 = n16874 ^ n15669 ^ 1'b0 ;
  assign n41114 = ~n41112 & n41113 ;
  assign n41115 = n26094 & n41114 ;
  assign n41116 = n22550 ^ n19943 ^ 1'b0 ;
  assign n41117 = n14490 & n20915 ;
  assign n41118 = n35649 & n41117 ;
  assign n41119 = n13335 & n29673 ;
  assign n41120 = ( n9431 & ~n10408 ) | ( n9431 & n11256 ) | ( ~n10408 & n11256 ) ;
  assign n41121 = n13765 ^ n13281 ^ 1'b0 ;
  assign n41122 = n41120 | n41121 ;
  assign n41124 = n14630 | n16699 ;
  assign n41123 = n25195 & n35726 ;
  assign n41125 = n41124 ^ n41123 ^ 1'b0 ;
  assign n41127 = n14386 & n14898 ;
  assign n41126 = ~n335 & n4156 ;
  assign n41128 = n41127 ^ n41126 ^ 1'b0 ;
  assign n41129 = ( ~n11032 & n20899 ) | ( ~n11032 & n22488 ) | ( n20899 & n22488 ) ;
  assign n41130 = n4546 ^ n1842 ^ 1'b0 ;
  assign n41131 = n41130 ^ n22886 ^ 1'b0 ;
  assign n41133 = n23858 ^ n19144 ^ 1'b0 ;
  assign n41132 = n35272 ^ n25280 ^ 1'b0 ;
  assign n41134 = n41133 ^ n41132 ^ n34174 ;
  assign n41135 = n10531 | n28465 ;
  assign n41136 = n23613 | n39521 ;
  assign n41137 = n41136 ^ n31708 ^ 1'b0 ;
  assign n41138 = n4955 | n24738 ;
  assign n41139 = ~n13897 & n27475 ;
  assign n41140 = n41139 ^ n19006 ^ 1'b0 ;
  assign n41141 = n27101 & n41140 ;
  assign n41143 = ~n15680 & n28727 ;
  assign n41142 = n14008 ^ n5279 ^ 1'b0 ;
  assign n41144 = n41143 ^ n41142 ^ n6216 ;
  assign n41145 = n29883 ^ n12126 ^ n3123 ;
  assign n41146 = n41145 ^ n14760 ^ 1'b0 ;
  assign n41147 = n20725 | n41146 ;
  assign n41148 = n41147 ^ n17169 ^ n13568 ;
  assign n41149 = n35696 ^ n10963 ^ 1'b0 ;
  assign n41150 = n41149 ^ n4612 ^ 1'b0 ;
  assign n41151 = n41148 & n41150 ;
  assign n41152 = n30886 & n41151 ;
  assign n41153 = n40690 ^ n39935 ^ n39050 ;
  assign n41154 = ( ~n1508 & n1766 ) | ( ~n1508 & n20316 ) | ( n1766 & n20316 ) ;
  assign n41155 = n25892 ^ n20119 ^ 1'b0 ;
  assign n41156 = ~n41154 & n41155 ;
  assign n41157 = n4635 ^ n1034 ^ 1'b0 ;
  assign n41158 = ( n18148 & n25988 ) | ( n18148 & ~n41157 ) | ( n25988 & ~n41157 ) ;
  assign n41159 = n11733 & ~n16892 ;
  assign n41160 = n41159 ^ n31768 ^ 1'b0 ;
  assign n41161 = n15660 | n41160 ;
  assign n41162 = n28948 | n41161 ;
  assign n41163 = ( n41156 & n41158 ) | ( n41156 & ~n41162 ) | ( n41158 & ~n41162 ) ;
  assign n41164 = n34486 ^ n7818 ^ 1'b0 ;
  assign n41165 = n19765 & n41164 ;
  assign n41166 = ~n888 & n14479 ;
  assign n41167 = n35019 ^ n25877 ^ 1'b0 ;
  assign n41168 = n809 ^ n717 ^ 1'b0 ;
  assign n41169 = n1729 & ~n41168 ;
  assign n41170 = ~n8572 & n41169 ;
  assign n41171 = ~x101 & n41170 ;
  assign n41172 = n1594 & ~n1600 ;
  assign n41173 = ~n41171 & n41172 ;
  assign n41174 = n8478 | n21421 ;
  assign n41175 = n1046 | n1893 ;
  assign n41176 = n6728 & ~n41175 ;
  assign n41177 = n2469 | n41176 ;
  assign n41178 = ( n2532 & ~n17333 ) | ( n2532 & n41177 ) | ( ~n17333 & n41177 ) ;
  assign n41179 = n33678 ^ n11764 ^ 1'b0 ;
  assign n41180 = n4298 | n30901 ;
  assign n41181 = n29392 ^ n24446 ^ 1'b0 ;
  assign n41182 = n7028 & ~n41181 ;
  assign n41183 = n23840 ^ n14346 ^ 1'b0 ;
  assign n41184 = n7638 | n41183 ;
  assign n41185 = n22031 & ~n34489 ;
  assign n41186 = ~n36552 & n41185 ;
  assign n41187 = ~n14563 & n34226 ;
  assign n41188 = n41187 ^ n39280 ^ 1'b0 ;
  assign n41189 = n5779 | n14929 ;
  assign n41190 = n41189 ^ n10563 ^ 1'b0 ;
  assign n41191 = n6436 | n34720 ;
  assign n41192 = n20918 & n22229 ;
  assign n41193 = n41192 ^ n13420 ^ 1'b0 ;
  assign n41194 = n4136 | n4770 ;
  assign n41195 = n41194 ^ n6812 ^ 1'b0 ;
  assign n41196 = n36613 ^ n834 ^ 1'b0 ;
  assign n41197 = n41196 ^ n25340 ^ n1907 ;
  assign n41198 = n41195 | n41197 ;
  assign n41199 = n4552 & ~n41198 ;
  assign n41200 = n11104 & ~n12042 ;
  assign n41201 = n1015 & n41200 ;
  assign n41202 = n41201 ^ n18850 ^ 1'b0 ;
  assign n41203 = n11338 | n32839 ;
  assign n41204 = x38 | n31330 ;
  assign n41205 = n41204 ^ n2547 ^ n2141 ;
  assign n41206 = ~n2162 & n31853 ;
  assign n41213 = n8955 ^ n3966 ^ n1852 ;
  assign n41207 = n586 & n40383 ;
  assign n41208 = ~x182 & n41207 ;
  assign n41209 = ~n9685 & n14004 ;
  assign n41210 = n41209 ^ n4979 ^ 1'b0 ;
  assign n41211 = n12642 | n41210 ;
  assign n41212 = n41208 & ~n41211 ;
  assign n41214 = n41213 ^ n41212 ^ n2453 ;
  assign n41215 = ~n5964 & n26633 ;
  assign n41216 = n39128 & n41215 ;
  assign n41219 = n11419 & n18488 ;
  assign n41220 = n7451 & n41219 ;
  assign n41217 = n31488 & n35561 ;
  assign n41218 = n41217 ^ n7151 ^ 1'b0 ;
  assign n41221 = n41220 ^ n41218 ^ 1'b0 ;
  assign n41222 = n17418 & ~n41221 ;
  assign n41223 = ~n31219 & n41222 ;
  assign n41224 = ~n16763 & n31418 ;
  assign n41225 = ~n17889 & n41224 ;
  assign n41226 = n35764 ^ n20414 ^ n1813 ;
  assign n41227 = n8197 & n38949 ;
  assign n41228 = n18944 | n41227 ;
  assign n41229 = n41226 | n41228 ;
  assign n41230 = n41229 ^ n20491 ^ 1'b0 ;
  assign n41231 = ~n41225 & n41230 ;
  assign n41232 = n38709 ^ n22061 ^ 1'b0 ;
  assign n41233 = n9736 & n41232 ;
  assign n41234 = n16267 | n17550 ;
  assign n41235 = ~n6153 & n41234 ;
  assign n41236 = ( n4376 & ~n23353 ) | ( n4376 & n28574 ) | ( ~n23353 & n28574 ) ;
  assign n41237 = ( n10976 & ~n16606 ) | ( n10976 & n41236 ) | ( ~n16606 & n41236 ) ;
  assign n41238 = ~n4404 & n19407 ;
  assign n41239 = ~n9187 & n41238 ;
  assign n41240 = ( n22315 & n33473 ) | ( n22315 & n41239 ) | ( n33473 & n41239 ) ;
  assign n41242 = n22999 ^ x54 ^ 1'b0 ;
  assign n41243 = n13130 & n41242 ;
  assign n41244 = ~n11373 & n41243 ;
  assign n41245 = n10945 & n41244 ;
  assign n41241 = n15529 & n37801 ;
  assign n41246 = n41245 ^ n41241 ^ 1'b0 ;
  assign n41247 = n27643 ^ n12294 ^ 1'b0 ;
  assign n41248 = n41246 & ~n41247 ;
  assign n41249 = n13863 ^ n8659 ^ 1'b0 ;
  assign n41250 = ~n38621 & n41249 ;
  assign n41251 = n11806 & n36593 ;
  assign n41252 = n41251 ^ n31883 ^ 1'b0 ;
  assign n41253 = n18004 ^ n14075 ^ 1'b0 ;
  assign n41254 = ~n11388 & n41253 ;
  assign n41255 = n39196 ^ n10395 ^ 1'b0 ;
  assign n41256 = n20554 & n41255 ;
  assign n41257 = n15410 ^ n15142 ^ 1'b0 ;
  assign n41258 = ( ~n12157 & n41256 ) | ( ~n12157 & n41257 ) | ( n41256 & n41257 ) ;
  assign n41259 = n24216 & n41258 ;
  assign n41260 = ( ~n2342 & n15989 ) | ( ~n2342 & n27319 ) | ( n15989 & n27319 ) ;
  assign n41261 = ( ~n11588 & n39039 ) | ( ~n11588 & n41260 ) | ( n39039 & n41260 ) ;
  assign n41262 = n4395 | n34090 ;
  assign n41263 = n4395 & ~n41262 ;
  assign n41264 = n41263 ^ n26712 ^ n18387 ;
  assign n41265 = n1044 | n40740 ;
  assign n41266 = n37931 ^ n20429 ^ 1'b0 ;
  assign n41267 = n41265 & ~n41266 ;
  assign n41268 = n1108 ^ n703 ^ 1'b0 ;
  assign n41269 = ~n34780 & n41268 ;
  assign n41270 = n15885 & n41269 ;
  assign n41271 = n24742 ^ n15195 ^ 1'b0 ;
  assign n41272 = n22967 ^ n4388 ^ 1'b0 ;
  assign n41273 = n15257 & ~n41272 ;
  assign n41274 = n41273 ^ n2349 ^ 1'b0 ;
  assign n41275 = n31685 ^ n4824 ^ 1'b0 ;
  assign n41276 = n8919 & ~n9906 ;
  assign n41277 = n3800 | n9764 ;
  assign n41278 = n6504 & n40910 ;
  assign n41279 = n41278 ^ n14927 ^ 1'b0 ;
  assign n41280 = n31252 & n41279 ;
  assign n41281 = n27400 ^ n1054 ^ 1'b0 ;
  assign n41282 = ( ~n5139 & n8301 ) | ( ~n5139 & n12486 ) | ( n8301 & n12486 ) ;
  assign n41283 = n5107 | n41282 ;
  assign n41284 = n21769 & ~n26920 ;
  assign n41285 = n41284 ^ n17596 ^ 1'b0 ;
  assign n41286 = n18617 | n30474 ;
  assign n41287 = n6997 & n38624 ;
  assign n41288 = ~n41286 & n41287 ;
  assign n41289 = n41285 & n41288 ;
  assign n41290 = n2828 ^ n2505 ^ n1441 ;
  assign n41291 = n18426 ^ n2925 ^ 1'b0 ;
  assign n41292 = n41290 & n41291 ;
  assign n41293 = n41292 ^ n18938 ^ n973 ;
  assign n41294 = n31409 ^ x29 ^ 1'b0 ;
  assign n41295 = n3490 | n22481 ;
  assign n41296 = n1769 & ~n39806 ;
  assign n41297 = n1030 | n27328 ;
  assign n41298 = n11709 & ~n27271 ;
  assign n41299 = n41298 ^ n30333 ^ n19154 ;
  assign n41300 = n9138 & ~n15832 ;
  assign n41301 = n41300 ^ n29876 ^ n3504 ;
  assign n41302 = n3467 & ~n23788 ;
  assign n41303 = n41302 ^ n10771 ^ 1'b0 ;
  assign n41304 = ~n1961 & n2671 ;
  assign n41305 = n41304 ^ n6858 ^ 1'b0 ;
  assign n41306 = n41305 ^ n18596 ^ 1'b0 ;
  assign n41307 = n29476 & ~n41306 ;
  assign n41308 = n428 & n39911 ;
  assign n41309 = n41308 ^ n37626 ^ 1'b0 ;
  assign n41310 = n2369 & ~n4516 ;
  assign n41311 = ( x71 & x218 ) | ( x71 & ~n2796 ) | ( x218 & ~n2796 ) ;
  assign n41312 = n12664 ^ n1448 ^ 1'b0 ;
  assign n41313 = n10959 | n41312 ;
  assign n41314 = n19610 & n21239 ;
  assign n41315 = n41313 & ~n41314 ;
  assign n41316 = n26181 | n41315 ;
  assign n41317 = n41316 ^ n26655 ^ 1'b0 ;
  assign n41318 = n1010 | n41317 ;
  assign n41319 = n41318 ^ n36232 ^ 1'b0 ;
  assign n41321 = n8771 | n10067 ;
  assign n41322 = n41321 ^ n20605 ^ 1'b0 ;
  assign n41320 = n15363 & ~n29650 ;
  assign n41323 = n41322 ^ n41320 ^ 1'b0 ;
  assign n41324 = n10191 & ~n22269 ;
  assign n41325 = n41324 ^ n6284 ^ 1'b0 ;
  assign n41326 = n10837 & n36329 ;
  assign n41327 = n35109 ^ n4334 ^ 1'b0 ;
  assign n41328 = n41327 ^ n3919 ^ 1'b0 ;
  assign n41329 = ~n25841 & n41328 ;
  assign n41330 = n41329 ^ n31205 ^ 1'b0 ;
  assign n41331 = n35919 | n36127 ;
  assign n41332 = n6135 | n20234 ;
  assign n41333 = n41332 ^ x144 ^ 1'b0 ;
  assign n41334 = n41333 ^ n12513 ^ 1'b0 ;
  assign n41335 = n41334 ^ n18416 ^ n939 ;
  assign n41336 = n13554 & ~n17108 ;
  assign n41337 = n8940 & n41336 ;
  assign n41338 = n3674 ^ n831 ^ 1'b0 ;
  assign n41339 = n41337 | n41338 ;
  assign n41340 = n9764 ^ n6254 ^ n4760 ;
  assign n41341 = n6157 | n41340 ;
  assign n41342 = n41339 & ~n41341 ;
  assign n41343 = ( n10585 & ~n10663 ) | ( n10585 & n12151 ) | ( ~n10663 & n12151 ) ;
  assign n41344 = n15803 ^ n6571 ^ 1'b0 ;
  assign n41345 = ~n24434 & n41344 ;
  assign n41346 = n41343 & ~n41345 ;
  assign n41347 = n34825 | n40000 ;
  assign n41348 = ( n686 & n12037 ) | ( n686 & ~n17030 ) | ( n12037 & ~n17030 ) ;
  assign n41349 = n2030 & ~n29260 ;
  assign n41350 = n41349 ^ n5530 ^ 1'b0 ;
  assign n41351 = ( ~n8572 & n31013 ) | ( ~n8572 & n41350 ) | ( n31013 & n41350 ) ;
  assign n41352 = n22131 ^ n13543 ^ 1'b0 ;
  assign n41353 = ~n19353 & n41352 ;
  assign n41354 = n7285 & ~n24019 ;
  assign n41355 = ( ~n25666 & n41353 ) | ( ~n25666 & n41354 ) | ( n41353 & n41354 ) ;
  assign n41356 = n8500 | n10262 ;
  assign n41357 = n6903 & n41356 ;
  assign n41358 = ~n23039 & n41357 ;
  assign n41359 = n6074 | n35857 ;
  assign n41360 = n15397 & ~n41359 ;
  assign n41361 = n4046 | n22717 ;
  assign n41362 = n41361 ^ n14832 ^ 1'b0 ;
  assign n41363 = n23245 ^ n5889 ^ n2738 ;
  assign n41364 = ( ~n20323 & n26228 ) | ( ~n20323 & n41363 ) | ( n26228 & n41363 ) ;
  assign n41365 = n35849 ^ n25870 ^ n8986 ;
  assign n41366 = n1602 & ~n4114 ;
  assign n41367 = ( n3767 & n35658 ) | ( n3767 & ~n41366 ) | ( n35658 & ~n41366 ) ;
  assign n41368 = n29255 ^ n10081 ^ 1'b0 ;
  assign n41369 = ~n27142 & n41368 ;
  assign n41370 = ~n631 & n26097 ;
  assign n41371 = n2489 & n41370 ;
  assign n41372 = n41371 ^ n31925 ^ n1626 ;
  assign n41373 = ( n35390 & n41369 ) | ( n35390 & n41372 ) | ( n41369 & n41372 ) ;
  assign n41374 = n15544 & n36679 ;
  assign n41375 = n20593 ^ n3275 ^ 1'b0 ;
  assign n41376 = n17044 & ~n41375 ;
  assign n41377 = ~n41374 & n41376 ;
  assign n41378 = n8778 & n25137 ;
  assign n41379 = n14508 | n37339 ;
  assign n41380 = n41379 ^ n7376 ^ 1'b0 ;
  assign n41381 = n2024 | n41380 ;
  assign n41382 = n10427 & ~n41381 ;
  assign n41383 = n40491 ^ n15961 ^ 1'b0 ;
  assign n41384 = n26692 ^ n15927 ^ n15486 ;
  assign n41385 = n6516 & ~n13429 ;
  assign n41386 = n41385 ^ n10017 ^ 1'b0 ;
  assign n41387 = n41386 ^ n5810 ^ 1'b0 ;
  assign n41388 = ~n2549 & n12870 ;
  assign n41389 = n41388 ^ n19993 ^ 1'b0 ;
  assign n41390 = n7740 & ~n41389 ;
  assign n41391 = n27391 ^ n18312 ^ n10793 ;
  assign n41392 = n34909 | n41391 ;
  assign n41393 = n41392 ^ n5359 ^ 1'b0 ;
  assign n41397 = n13579 ^ n2752 ^ 1'b0 ;
  assign n41398 = n5078 & ~n41397 ;
  assign n41394 = n14179 | n22891 ;
  assign n41395 = n41394 ^ n3100 ^ 1'b0 ;
  assign n41396 = n28067 & ~n41395 ;
  assign n41399 = n41398 ^ n41396 ^ 1'b0 ;
  assign n41408 = n17081 ^ n7448 ^ 1'b0 ;
  assign n41409 = n11704 & n41408 ;
  assign n41400 = ( ~n1910 & n4439 ) | ( ~n1910 & n9952 ) | ( n4439 & n9952 ) ;
  assign n41401 = n24261 ^ n13443 ^ 1'b0 ;
  assign n41402 = n41400 & n41401 ;
  assign n41403 = n22673 & n34287 ;
  assign n41404 = n41403 ^ n5919 ^ 1'b0 ;
  assign n41405 = n41404 ^ n2264 ^ 1'b0 ;
  assign n41406 = n41402 & ~n41405 ;
  assign n41407 = n10857 & n41406 ;
  assign n41410 = n41409 ^ n41407 ^ 1'b0 ;
  assign n41413 = n2350 | n15961 ;
  assign n41411 = n8737 | n12524 ;
  assign n41412 = n41411 ^ n8345 ^ 1'b0 ;
  assign n41414 = n41413 ^ n41412 ^ n10053 ;
  assign n41415 = n9154 & n31937 ;
  assign n41416 = ( n19607 & ~n25546 ) | ( n19607 & n41415 ) | ( ~n25546 & n41415 ) ;
  assign n41417 = ~n22004 & n38476 ;
  assign n41418 = n25876 & ~n34102 ;
  assign n41419 = n18546 & n41418 ;
  assign n41420 = n682 | n7637 ;
  assign n41421 = n36431 & n41420 ;
  assign n41422 = n26269 ^ n7382 ^ 1'b0 ;
  assign n41423 = n20334 | n41422 ;
  assign n41424 = ~n7895 & n13887 ;
  assign n41425 = ( n15224 & n16677 ) | ( n15224 & ~n41424 ) | ( n16677 & ~n41424 ) ;
  assign n41426 = n16691 & n41425 ;
  assign n41427 = ~n23397 & n41426 ;
  assign n41428 = n41427 ^ n24577 ^ 1'b0 ;
  assign n41429 = ~n41423 & n41428 ;
  assign n41430 = n2482 & n41029 ;
  assign n41431 = n41430 ^ n30197 ^ 1'b0 ;
  assign n41432 = n33306 ^ n27380 ^ 1'b0 ;
  assign n41433 = n38408 ^ n5889 ^ n3181 ;
  assign n41434 = n1948 | n2152 ;
  assign n41435 = n41434 ^ n19213 ^ 1'b0 ;
  assign n41436 = n12476 & n17921 ;
  assign n41437 = n12701 & n41436 ;
  assign n41438 = n16012 & ~n41437 ;
  assign n41439 = n4769 ^ n4419 ^ 1'b0 ;
  assign n41440 = n12499 | n41439 ;
  assign n41441 = n36293 | n41440 ;
  assign n41442 = n41441 ^ n28862 ^ 1'b0 ;
  assign n41443 = ( n3088 & ~n7728 ) | ( n3088 & n16241 ) | ( ~n7728 & n16241 ) ;
  assign n41444 = n11834 & n12445 ;
  assign n41445 = n4944 & n16607 ;
  assign n41446 = n32681 | n41445 ;
  assign n41447 = ( n385 & n3107 ) | ( n385 & n6020 ) | ( n3107 & n6020 ) ;
  assign n41448 = n18856 & n41447 ;
  assign n41449 = n4862 & n41448 ;
  assign n41450 = n41449 ^ n41076 ^ n36103 ;
  assign n41451 = n17187 ^ n7577 ^ 1'b0 ;
  assign n41452 = ( n16774 & n41450 ) | ( n16774 & n41451 ) | ( n41450 & n41451 ) ;
  assign n41453 = ~n4589 & n38615 ;
  assign n41454 = n41453 ^ n35310 ^ 1'b0 ;
  assign n41455 = n16522 ^ n11017 ^ 1'b0 ;
  assign n41456 = n26606 & n41455 ;
  assign n41457 = n6710 & ~n10180 ;
  assign n41458 = ~n23503 & n41457 ;
  assign n41459 = n17848 & ~n33678 ;
  assign n41460 = n30728 ^ n9943 ^ n2779 ;
  assign n41461 = ( n2230 & n26550 ) | ( n2230 & n37113 ) | ( n26550 & n37113 ) ;
  assign n41462 = ( ~n16166 & n18969 ) | ( ~n16166 & n26585 ) | ( n18969 & n26585 ) ;
  assign n41463 = n6960 & ~n41462 ;
  assign n41464 = n5244 & ~n14487 ;
  assign n41465 = n21360 & ~n21612 ;
  assign n41466 = n2586 | n41465 ;
  assign n41467 = ( n29465 & ~n41464 ) | ( n29465 & n41466 ) | ( ~n41464 & n41466 ) ;
  assign n41468 = ~n2954 & n41467 ;
  assign n41469 = n1613 & ~n20803 ;
  assign n41471 = ~n9035 & n11026 ;
  assign n41470 = n8422 & ~n18200 ;
  assign n41472 = n41471 ^ n41470 ^ 1'b0 ;
  assign n41473 = n813 | n36430 ;
  assign n41474 = n37155 ^ n5291 ^ 1'b0 ;
  assign n41475 = ~n5621 & n36865 ;
  assign n41476 = n39712 ^ n22852 ^ 1'b0 ;
  assign n41482 = n2427 | n15168 ;
  assign n41483 = n5578 & ~n41482 ;
  assign n41484 = n15074 | n41483 ;
  assign n41477 = n3029 & n25969 ;
  assign n41478 = n41422 ^ n29014 ^ 1'b0 ;
  assign n41479 = n23973 | n41478 ;
  assign n41480 = n36175 & ~n41479 ;
  assign n41481 = n41477 | n41480 ;
  assign n41485 = n41484 ^ n41481 ^ 1'b0 ;
  assign n41486 = n1399 | n39290 ;
  assign n41487 = n24504 & n29339 ;
  assign n41488 = ~n28919 & n41487 ;
  assign n41489 = n10185 & n11221 ;
  assign n41490 = n41489 ^ n18377 ^ 1'b0 ;
  assign n41491 = n29575 ^ n24803 ^ 1'b0 ;
  assign n41492 = n8887 & n22880 ;
  assign n41493 = ~n9188 & n41492 ;
  assign n41494 = n9660 ^ n1016 ^ 1'b0 ;
  assign n41495 = ~n31694 & n41494 ;
  assign n41496 = n41495 ^ n24874 ^ n9350 ;
  assign n41497 = ~n631 & n7113 ;
  assign n41498 = n41497 ^ n6016 ^ 1'b0 ;
  assign n41499 = ~n7989 & n41498 ;
  assign n41500 = n41499 ^ n5542 ^ n2800 ;
  assign n41501 = n33721 & ~n41500 ;
  assign n41502 = n19993 | n24342 ;
  assign n41503 = n41502 ^ n17618 ^ 1'b0 ;
  assign n41504 = ( n10003 & n34484 ) | ( n10003 & ~n41503 ) | ( n34484 & ~n41503 ) ;
  assign n41505 = n27141 ^ n22152 ^ 1'b0 ;
  assign n41506 = ~n485 & n41505 ;
  assign n41507 = n6847 & n36241 ;
  assign n41508 = n23955 & n41507 ;
  assign n41509 = n25742 ^ n7944 ^ n1941 ;
  assign n41510 = ~n11762 & n41509 ;
  assign n41511 = ~n12722 & n41510 ;
  assign n41512 = n3789 & ~n41511 ;
  assign n41513 = n31685 ^ n26448 ^ 1'b0 ;
  assign n41514 = n6914 & n12584 ;
  assign n41515 = n41514 ^ n18220 ^ 1'b0 ;
  assign n41516 = n41515 ^ n12742 ^ 1'b0 ;
  assign n41523 = n25909 & n26303 ;
  assign n41524 = n41523 ^ n1698 ^ 1'b0 ;
  assign n41517 = n25604 ^ n7439 ^ 1'b0 ;
  assign n41518 = n41517 ^ n20669 ^ n6261 ;
  assign n41519 = n17186 | n41518 ;
  assign n41520 = n41519 ^ n30440 ^ 1'b0 ;
  assign n41521 = n18335 ^ n3150 ^ 1'b0 ;
  assign n41522 = n41520 & ~n41521 ;
  assign n41525 = n41524 ^ n41522 ^ 1'b0 ;
  assign n41526 = n35070 & ~n41525 ;
  assign n41527 = n38824 ^ n32740 ^ 1'b0 ;
  assign n41528 = x57 & n41527 ;
  assign n41529 = n41528 ^ n1787 ^ 1'b0 ;
  assign n41530 = ( ~n12011 & n16344 ) | ( ~n12011 & n30605 ) | ( n16344 & n30605 ) ;
  assign n41531 = n41530 ^ n18318 ^ 1'b0 ;
  assign n41532 = ~n12743 & n25783 ;
  assign n41533 = ( ~n29540 & n38943 ) | ( ~n29540 & n41532 ) | ( n38943 & n41532 ) ;
  assign n41534 = n41533 ^ n2251 ^ 1'b0 ;
  assign n41535 = n25119 ^ n13721 ^ 1'b0 ;
  assign n41536 = n22365 ^ n14518 ^ 1'b0 ;
  assign n41537 = n4928 & n41536 ;
  assign n41538 = n41537 ^ n13603 ^ n956 ;
  assign n41539 = n41538 ^ x49 ^ 1'b0 ;
  assign n41540 = n1347 & ~n3523 ;
  assign n41541 = n41539 & ~n41540 ;
  assign n41542 = n16413 ^ n12434 ^ 1'b0 ;
  assign n41543 = n6111 | n41542 ;
  assign n41544 = n5594 & n16857 ;
  assign n41545 = n41543 & n41544 ;
  assign n41546 = n17805 ^ n14919 ^ 1'b0 ;
  assign n41547 = n26045 & n41546 ;
  assign n41548 = n27716 ^ n26274 ^ n17203 ;
  assign n41549 = n40769 ^ n4602 ^ 1'b0 ;
  assign n41551 = n28690 ^ n25875 ^ n15325 ;
  assign n41550 = n2401 & ~n34853 ;
  assign n41552 = n41551 ^ n41550 ^ 1'b0 ;
  assign n41553 = n37628 | n41552 ;
  assign n41554 = n35245 ^ n971 ^ 1'b0 ;
  assign n41555 = n5475 & ~n37264 ;
  assign n41556 = n41554 & n41555 ;
  assign n41558 = n28713 ^ n19513 ^ 1'b0 ;
  assign n41559 = n41558 ^ n10045 ^ 1'b0 ;
  assign n41560 = ~n28262 & n41559 ;
  assign n41557 = n7810 | n23844 ;
  assign n41561 = n41560 ^ n41557 ^ 1'b0 ;
  assign n41562 = n1962 & n3148 ;
  assign n41563 = n41562 ^ n763 ^ 1'b0 ;
  assign n41564 = n6891 & n21542 ;
  assign n41565 = n41564 ^ n33017 ^ 1'b0 ;
  assign n41567 = n13420 ^ n7466 ^ n4334 ;
  assign n41566 = n26552 & n32375 ;
  assign n41568 = n41567 ^ n41566 ^ 1'b0 ;
  assign n41569 = ~n3203 & n36420 ;
  assign n41570 = n11078 ^ n1800 ^ 1'b0 ;
  assign n41571 = ( ~n4775 & n13625 ) | ( ~n4775 & n17513 ) | ( n13625 & n17513 ) ;
  assign n41572 = x11 & n37012 ;
  assign n41573 = n14304 & n41572 ;
  assign n41574 = ( n21085 & ~n41571 ) | ( n21085 & n41573 ) | ( ~n41571 & n41573 ) ;
  assign n41575 = n5752 & ~n41574 ;
  assign n41576 = ( n5926 & ~n26946 ) | ( n5926 & n41575 ) | ( ~n26946 & n41575 ) ;
  assign n41577 = n11570 & ~n41427 ;
  assign n41578 = n41577 ^ n30650 ^ 1'b0 ;
  assign n41579 = n11170 & ~n25562 ;
  assign n41580 = ~n12679 & n41579 ;
  assign n41581 = n27646 ^ n10255 ^ 1'b0 ;
  assign n41582 = ~n41580 & n41581 ;
  assign n41583 = n17403 & n20366 ;
  assign n41584 = n9916 & ~n19027 ;
  assign n41585 = n22829 & n41584 ;
  assign n41586 = n32226 ^ n16489 ^ n11007 ;
  assign n41587 = ( n1975 & n4855 ) | ( n1975 & ~n15838 ) | ( n4855 & ~n15838 ) ;
  assign n41588 = n34145 | n41587 ;
  assign n41589 = n41586 & ~n41588 ;
  assign n41590 = ( ~n40839 & n41585 ) | ( ~n40839 & n41589 ) | ( n41585 & n41589 ) ;
  assign n41591 = ( n941 & ~n6665 ) | ( n941 & n31359 ) | ( ~n6665 & n31359 ) ;
  assign n41592 = n40968 ^ n13142 ^ 1'b0 ;
  assign n41593 = n18432 | n41592 ;
  assign n41594 = n7715 & n17306 ;
  assign n41595 = n41594 ^ n34313 ^ 1'b0 ;
  assign n41596 = n36097 ^ n17990 ^ 1'b0 ;
  assign n41597 = ~n40879 & n41596 ;
  assign n41598 = n41597 ^ n10436 ^ 1'b0 ;
  assign n41599 = n25631 ^ n3065 ^ 1'b0 ;
  assign n41600 = n7957 & ~n39001 ;
  assign n41601 = ~n19812 & n41600 ;
  assign n41602 = n5345 | n37400 ;
  assign n41603 = n41602 ^ n35273 ^ 1'b0 ;
  assign n41604 = n34750 ^ n25648 ^ n7697 ;
  assign n41605 = n7490 & n41604 ;
  assign n41606 = ( ~n1073 & n5942 ) | ( ~n1073 & n17794 ) | ( n5942 & n17794 ) ;
  assign n41607 = ( ~n4136 & n28873 ) | ( ~n4136 & n41606 ) | ( n28873 & n41606 ) ;
  assign n41608 = n18508 ^ n3463 ^ 1'b0 ;
  assign n41609 = ~n7836 & n41608 ;
  assign n41610 = n41609 ^ n18866 ^ n1578 ;
  assign n41611 = x110 & ~n17119 ;
  assign n41612 = n41611 ^ n27632 ^ 1'b0 ;
  assign n41613 = n40982 ^ n2814 ^ 1'b0 ;
  assign n41614 = n2313 & n11389 ;
  assign n41615 = n41614 ^ n36498 ^ 1'b0 ;
  assign n41616 = n20977 & ~n27403 ;
  assign n41617 = n41615 & n41616 ;
  assign n41618 = n16757 ^ n993 ^ 1'b0 ;
  assign n41619 = n40071 ^ n27702 ^ 1'b0 ;
  assign n41620 = n24265 | n41619 ;
  assign n41621 = n17317 & ~n23876 ;
  assign n41622 = n41620 & n41621 ;
  assign n41623 = n26928 ^ n5023 ^ 1'b0 ;
  assign n41624 = n24319 | n41623 ;
  assign n41625 = n12035 ^ n3229 ^ 1'b0 ;
  assign n41626 = n41624 & ~n41625 ;
  assign n41627 = n9398 ^ n6992 ^ n4307 ;
  assign n41628 = n41627 ^ n3223 ^ 1'b0 ;
  assign n41629 = n6110 | n41628 ;
  assign n41630 = ( n14905 & n17761 ) | ( n14905 & n31287 ) | ( n17761 & n31287 ) ;
  assign n41631 = n30547 ^ n3910 ^ 1'b0 ;
  assign n41632 = ~n14073 & n30695 ;
  assign n41633 = n40355 ^ n20971 ^ 1'b0 ;
  assign n41634 = ~n32474 & n41633 ;
  assign n41635 = ( n472 & n14403 ) | ( n472 & ~n23504 ) | ( n14403 & ~n23504 ) ;
  assign n41636 = n41635 ^ n22937 ^ n8631 ;
  assign n41637 = ~n490 & n41636 ;
  assign n41638 = n28190 ^ n901 ^ 1'b0 ;
  assign n41639 = n16366 | n25131 ;
  assign n41640 = n18350 | n41639 ;
  assign n41641 = n5934 & n41640 ;
  assign n41642 = n41641 ^ n28687 ^ 1'b0 ;
  assign n41643 = ~n25727 & n41642 ;
  assign n41644 = n5732 & n41643 ;
  assign n41646 = n25677 ^ n10669 ^ 1'b0 ;
  assign n41645 = n11349 | n41606 ;
  assign n41647 = n41646 ^ n41645 ^ 1'b0 ;
  assign n41648 = n6889 & n20257 ;
  assign n41649 = n7063 ^ n4016 ^ 1'b0 ;
  assign n41650 = n11497 & ~n13854 ;
  assign n41652 = n3510 & ~n33413 ;
  assign n41653 = n19964 & n41652 ;
  assign n41651 = n4474 & ~n7214 ;
  assign n41654 = n41653 ^ n41651 ^ 1'b0 ;
  assign n41660 = n5710 & ~n9047 ;
  assign n41659 = n16681 ^ n6583 ^ 1'b0 ;
  assign n41655 = n16436 & n17758 ;
  assign n41656 = ~n19546 & n41655 ;
  assign n41657 = n40254 | n41656 ;
  assign n41658 = n28917 | n41657 ;
  assign n41661 = n41660 ^ n41659 ^ n41658 ;
  assign n41662 = n16256 & n41661 ;
  assign n41663 = n41662 ^ n32190 ^ 1'b0 ;
  assign n41664 = n35634 ^ n23753 ^ n4770 ;
  assign n41665 = n3100 & n14134 ;
  assign n41666 = n9803 | n11998 ;
  assign n41667 = n11010 | n41666 ;
  assign n41668 = ( n5839 & n39689 ) | ( n5839 & ~n41667 ) | ( n39689 & ~n41667 ) ;
  assign n41669 = n41668 ^ n13614 ^ 1'b0 ;
  assign n41670 = n25927 & n37207 ;
  assign n41675 = n1579 | n20996 ;
  assign n41672 = ( n2459 & ~n9217 ) | ( n2459 & n15300 ) | ( ~n9217 & n15300 ) ;
  assign n41673 = n27563 | n41672 ;
  assign n41674 = n39424 | n41673 ;
  assign n41676 = n41675 ^ n41674 ^ 1'b0 ;
  assign n41677 = n21188 & n41676 ;
  assign n41671 = n15568 | n26008 ;
  assign n41678 = n41677 ^ n41671 ^ 1'b0 ;
  assign n41679 = ~n9300 & n12112 ;
  assign n41680 = n41679 ^ n8595 ^ 1'b0 ;
  assign n41681 = n32599 | n36427 ;
  assign n41682 = n41680 | n41681 ;
  assign n41683 = n3667 & ~n41022 ;
  assign n41684 = n35207 & n41683 ;
  assign n41685 = n36497 ^ n4033 ^ 1'b0 ;
  assign n41686 = n9530 ^ n8357 ^ 1'b0 ;
  assign n41687 = ( n15808 & n24921 ) | ( n15808 & ~n41686 ) | ( n24921 & ~n41686 ) ;
  assign n41689 = n6345 | n10910 ;
  assign n41688 = n30836 ^ n16165 ^ n9184 ;
  assign n41690 = n41689 ^ n41688 ^ 1'b0 ;
  assign n41691 = n15974 ^ n6117 ^ 1'b0 ;
  assign n41692 = n15950 & ~n41691 ;
  assign n41693 = ~n27754 & n41692 ;
  assign n41694 = n3440 & n28840 ;
  assign n41698 = ( n2598 & n3774 ) | ( n2598 & ~n31778 ) | ( n3774 & ~n31778 ) ;
  assign n41699 = n41698 ^ n12351 ^ 1'b0 ;
  assign n41700 = n37286 & ~n41699 ;
  assign n41695 = ~n33845 & n41406 ;
  assign n41696 = ~n13779 & n40474 ;
  assign n41697 = n41695 | n41696 ;
  assign n41701 = n41700 ^ n41697 ^ 1'b0 ;
  assign n41702 = n16609 ^ n15885 ^ 1'b0 ;
  assign n41703 = n38626 & ~n41702 ;
  assign n41704 = n36507 & n41703 ;
  assign n41705 = n12362 ^ n2107 ^ n2054 ;
  assign n41706 = n41705 ^ n3305 ^ 1'b0 ;
  assign n41707 = ~n36199 & n41706 ;
  assign n41708 = n19083 ^ n9319 ^ 1'b0 ;
  assign n41709 = n19350 | n41708 ;
  assign n41710 = ~n34214 & n38943 ;
  assign n41711 = n41710 ^ n27017 ^ 1'b0 ;
  assign n41712 = n41711 ^ n6556 ^ 1'b0 ;
  assign n41713 = n15431 | n41712 ;
  assign n41714 = n30163 ^ n22836 ^ 1'b0 ;
  assign n41715 = n14652 & n41714 ;
  assign n41716 = ( n19577 & ~n41713 ) | ( n19577 & n41715 ) | ( ~n41713 & n41715 ) ;
  assign n41717 = n17261 | n22783 ;
  assign n41718 = n41717 ^ n9899 ^ 1'b0 ;
  assign n41719 = n16891 & ~n41718 ;
  assign n41720 = n41719 ^ n29293 ^ n11557 ;
  assign n41721 = n17134 ^ n13622 ^ 1'b0 ;
  assign n41722 = n22608 & ~n41721 ;
  assign n41724 = n2518 | n2577 ;
  assign n41723 = n24907 ^ n8858 ^ 1'b0 ;
  assign n41725 = n41724 ^ n41723 ^ n34182 ;
  assign n41726 = n37439 ^ n25147 ^ n8999 ;
  assign n41727 = ( n9341 & ~n9731 ) | ( n9341 & n20473 ) | ( ~n9731 & n20473 ) ;
  assign n41728 = n37601 ^ n24012 ^ 1'b0 ;
  assign n41729 = n3878 | n41728 ;
  assign n41730 = n39918 ^ n24867 ^ 1'b0 ;
  assign n41731 = n6102 ^ n1107 ^ 1'b0 ;
  assign n41732 = n41731 ^ n22795 ^ 1'b0 ;
  assign n41733 = n30284 & ~n41732 ;
  assign n41734 = n12781 | n23391 ;
  assign n41735 = n41734 ^ n10850 ^ 1'b0 ;
  assign n41736 = n5764 & n18683 ;
  assign n41737 = n31761 ^ n5131 ^ 1'b0 ;
  assign n41738 = n41737 ^ n1337 ^ 1'b0 ;
  assign n41739 = n22491 | n41738 ;
  assign n41742 = n29402 ^ n24603 ^ 1'b0 ;
  assign n41740 = ( ~n10919 & n16249 ) | ( ~n10919 & n30685 ) | ( n16249 & n30685 ) ;
  assign n41741 = ( ~n8696 & n15214 ) | ( ~n8696 & n41740 ) | ( n15214 & n41740 ) ;
  assign n41743 = n41742 ^ n41741 ^ n18292 ;
  assign n41744 = n16140 ^ n1021 ^ 1'b0 ;
  assign n41745 = n16149 ^ n6276 ^ 1'b0 ;
  assign n41746 = n41744 & n41745 ;
  assign n41747 = n41746 ^ n20727 ^ 1'b0 ;
  assign n41748 = n30941 ^ n6471 ^ 1'b0 ;
  assign n41749 = n10600 ^ n9340 ^ 1'b0 ;
  assign n41750 = n7142 & ~n41749 ;
  assign n41751 = n41750 ^ n4258 ^ 1'b0 ;
  assign n41752 = x103 & n41751 ;
  assign n41753 = n41752 ^ n17004 ^ 1'b0 ;
  assign n41754 = n23929 & ~n33112 ;
  assign n41755 = n12197 & n41754 ;
  assign n41756 = n27582 ^ n21739 ^ 1'b0 ;
  assign n41757 = n3723 & ~n7197 ;
  assign n41758 = ~n9552 & n41757 ;
  assign n41759 = n7580 & ~n41758 ;
  assign n41760 = n41756 & n41759 ;
  assign n41761 = n30160 ^ n10147 ^ 1'b0 ;
  assign n41762 = n3605 & n41761 ;
  assign n41763 = n31463 ^ n692 ^ 1'b0 ;
  assign n41764 = n13848 & ~n15157 ;
  assign n41765 = n41763 & n41764 ;
  assign n41766 = n24088 ^ n12888 ^ n8781 ;
  assign n41767 = n1514 | n23636 ;
  assign n41768 = ( ~n15085 & n33401 ) | ( ~n15085 & n41767 ) | ( n33401 & n41767 ) ;
  assign n41769 = ~x187 & n23149 ;
  assign n41770 = ~n13678 & n17279 ;
  assign n41771 = n41770 ^ n19445 ^ n2779 ;
  assign n41772 = ( n2769 & n41769 ) | ( n2769 & ~n41771 ) | ( n41769 & ~n41771 ) ;
  assign n41773 = ~n14667 & n25618 ;
  assign n41774 = n41773 ^ n3631 ^ 1'b0 ;
  assign n41775 = n41774 ^ n1925 ^ 1'b0 ;
  assign n41776 = n25486 & ~n41775 ;
  assign n41777 = n1538 & n11091 ;
  assign n41778 = n3052 & n41777 ;
  assign n41779 = n41778 ^ n18321 ^ n8693 ;
  assign n41780 = n8521 & n34907 ;
  assign n41781 = ~n41779 & n41780 ;
  assign n41782 = n38875 ^ n6227 ^ 1'b0 ;
  assign n41786 = ~n18841 & n36890 ;
  assign n41783 = n10704 | n16699 ;
  assign n41784 = ~n19268 & n41783 ;
  assign n41785 = n6562 & n41784 ;
  assign n41787 = n41786 ^ n41785 ^ n7298 ;
  assign n41788 = n3222 & ~n41787 ;
  assign n41789 = n12513 | n21716 ;
  assign n41790 = n41789 ^ n25453 ^ 1'b0 ;
  assign n41791 = n27396 ^ n8076 ^ 1'b0 ;
  assign n41792 = n7694 ^ n6386 ^ 1'b0 ;
  assign n41793 = n8422 & ~n19025 ;
  assign n41794 = n41793 ^ n1634 ^ 1'b0 ;
  assign n41795 = n8887 & ~n32696 ;
  assign n41796 = ~n33640 & n41795 ;
  assign n41797 = n37879 & ~n41796 ;
  assign n41798 = n41797 ^ n4153 ^ 1'b0 ;
  assign n41799 = n26755 ^ n18126 ^ 1'b0 ;
  assign n41800 = ( n19349 & n24169 ) | ( n19349 & n39369 ) | ( n24169 & n39369 ) ;
  assign n41804 = n22853 ^ n21078 ^ n9933 ;
  assign n41805 = n7070 & ~n41804 ;
  assign n41801 = n13180 & n27904 ;
  assign n41802 = n2019 & n41801 ;
  assign n41803 = n10515 & ~n41802 ;
  assign n41806 = n41805 ^ n41803 ^ 1'b0 ;
  assign n41807 = n23067 ^ n18275 ^ 1'b0 ;
  assign n41808 = n38922 ^ n21533 ^ n19709 ;
  assign n41809 = n41808 ^ n26309 ^ n13216 ;
  assign n41810 = n41809 ^ n23139 ^ 1'b0 ;
  assign n41811 = ( n11186 & n19118 ) | ( n11186 & n21616 ) | ( n19118 & n21616 ) ;
  assign n41812 = n41811 ^ n6074 ^ 1'b0 ;
  assign n41813 = n14306 | n28531 ;
  assign n41814 = n27538 & n41813 ;
  assign n41815 = n9232 & ~n25271 ;
  assign n41816 = ~n18362 & n41815 ;
  assign n41817 = ( n10531 & n30764 ) | ( n10531 & n37974 ) | ( n30764 & n37974 ) ;
  assign n41818 = n41817 ^ n8838 ^ 1'b0 ;
  assign n41819 = n12602 ^ n1786 ^ 1'b0 ;
  assign n41820 = n33592 | n41819 ;
  assign n41821 = n2019 | n37874 ;
  assign n41822 = ( n27852 & n41820 ) | ( n27852 & ~n41821 ) | ( n41820 & ~n41821 ) ;
  assign n41823 = ( n11937 & n12234 ) | ( n11937 & n13280 ) | ( n12234 & n13280 ) ;
  assign n41824 = n30901 ^ n21192 ^ n9186 ;
  assign n41825 = ( n22741 & n27933 ) | ( n22741 & n41824 ) | ( n27933 & n41824 ) ;
  assign n41826 = n1994 & n17664 ;
  assign n41827 = n23116 & n41826 ;
  assign n41828 = n1319 & n6036 ;
  assign n41829 = n10026 | n24118 ;
  assign n41830 = n12508 & ~n41829 ;
  assign n41831 = n3121 | n41830 ;
  assign n41832 = n13525 | n28925 ;
  assign n41833 = n39557 & ~n41832 ;
  assign n41834 = ~n36225 & n41833 ;
  assign n41835 = n39515 ^ n15373 ^ 1'b0 ;
  assign n41836 = n9761 | n41835 ;
  assign n41837 = n14578 & n18919 ;
  assign n41838 = n41836 & n41837 ;
  assign n41839 = n11013 & ~n11401 ;
  assign n41840 = ~n4243 & n8709 ;
  assign n41841 = n12514 & n41840 ;
  assign n41842 = n41841 ^ n33184 ^ n13039 ;
  assign n41843 = n11403 ^ n5456 ^ 1'b0 ;
  assign n41844 = n11010 & n41843 ;
  assign n41845 = n6944 ^ n2924 ^ 1'b0 ;
  assign n41846 = n11930 & n41845 ;
  assign n41847 = n41846 ^ n5891 ^ 1'b0 ;
  assign n41848 = n41844 | n41847 ;
  assign n41849 = n15213 ^ n11257 ^ 1'b0 ;
  assign n41850 = n6945 & ~n8332 ;
  assign n41851 = n23148 ^ n16601 ^ 1'b0 ;
  assign n41852 = n11988 ^ n10639 ^ 1'b0 ;
  assign n41853 = n14496 & ~n41852 ;
  assign n41854 = n41851 & n41853 ;
  assign n41855 = n5739 & n14257 ;
  assign n41856 = n41855 ^ n39056 ^ 1'b0 ;
  assign n41857 = ~n13680 & n19689 ;
  assign n41858 = n6636 & n41857 ;
  assign n41862 = n10794 ^ n10603 ^ n515 ;
  assign n41859 = n10371 & n35525 ;
  assign n41860 = n41859 ^ n36300 ^ 1'b0 ;
  assign n41861 = ~n22968 & n41860 ;
  assign n41863 = n41862 ^ n41861 ^ 1'b0 ;
  assign n41864 = n34558 & ~n41863 ;
  assign n41866 = n39608 ^ n22940 ^ 1'b0 ;
  assign n41865 = n1749 & ~n10176 ;
  assign n41867 = n41866 ^ n41865 ^ 1'b0 ;
  assign n41868 = n22777 ^ n10832 ^ n3974 ;
  assign n41869 = ( n8181 & n8411 ) | ( n8181 & n40590 ) | ( n8411 & n40590 ) ;
  assign n41870 = n4141 & ~n4754 ;
  assign n41871 = n5840 & n41870 ;
  assign n41872 = n32029 & ~n41871 ;
  assign n41873 = n2840 & n41872 ;
  assign n41874 = ( n3803 & n16478 ) | ( n3803 & n41873 ) | ( n16478 & n41873 ) ;
  assign n41877 = ~n13314 & n22940 ;
  assign n41878 = ~n23123 & n41877 ;
  assign n41879 = n32832 ^ n13717 ^ 1'b0 ;
  assign n41880 = n41878 | n41879 ;
  assign n41875 = n7128 | n24747 ;
  assign n41876 = n18475 | n41875 ;
  assign n41881 = n41880 ^ n41876 ^ 1'b0 ;
  assign n41882 = n35574 ^ n22629 ^ 1'b0 ;
  assign n41883 = n7435 & n15044 ;
  assign n41884 = n41883 ^ n1310 ^ 1'b0 ;
  assign n41885 = n27345 | n39795 ;
  assign n41886 = n41885 ^ n16435 ^ 1'b0 ;
  assign n41887 = n1849 & ~n6480 ;
  assign n41888 = ~n28863 & n41887 ;
  assign n41889 = ( n9390 & n27850 ) | ( n9390 & ~n30710 ) | ( n27850 & ~n30710 ) ;
  assign n41890 = n6851 & ~n7208 ;
  assign n41891 = ( n4522 & n20518 ) | ( n4522 & ~n41890 ) | ( n20518 & ~n41890 ) ;
  assign n41892 = n36189 ^ n16031 ^ 1'b0 ;
  assign n41893 = x175 & n41892 ;
  assign n41894 = n5550 & ~n15665 ;
  assign n41895 = ~n41893 & n41894 ;
  assign n41896 = n25029 ^ n11509 ^ 1'b0 ;
  assign n41897 = n23710 & n41896 ;
  assign n41898 = ( ~n9457 & n40173 ) | ( ~n9457 & n41897 ) | ( n40173 & n41897 ) ;
  assign n41899 = n41895 | n41898 ;
  assign n41900 = n2110 & ~n6231 ;
  assign n41901 = n15794 | n27240 ;
  assign n41902 = n41901 ^ n7115 ^ 1'b0 ;
  assign n41903 = n37882 | n40863 ;
  assign n41904 = ~n5417 & n16325 ;
  assign n41905 = n41904 ^ n6293 ^ 1'b0 ;
  assign n41906 = n41905 ^ n5229 ^ 1'b0 ;
  assign n41907 = n37840 | n41906 ;
  assign n41908 = n41907 ^ n41811 ^ 1'b0 ;
  assign n41909 = ( n1126 & ~n40222 ) | ( n1126 & n41908 ) | ( ~n40222 & n41908 ) ;
  assign n41912 = n4823 & ~n19430 ;
  assign n41913 = ~n24759 & n41912 ;
  assign n41910 = n19029 ^ n18969 ^ 1'b0 ;
  assign n41911 = ~n1769 & n41910 ;
  assign n41914 = n41913 ^ n41911 ^ n21108 ;
  assign n41915 = n21679 ^ n15887 ^ 1'b0 ;
  assign n41916 = n28292 | n41915 ;
  assign n41917 = ( ~n12493 & n15445 ) | ( ~n12493 & n41916 ) | ( n15445 & n41916 ) ;
  assign n41918 = n12396 | n24530 ;
  assign n41919 = n5303 & ~n41918 ;
  assign n41920 = n23096 ^ n2742 ^ 1'b0 ;
  assign n41921 = n41919 | n41920 ;
  assign n41922 = x103 & n29047 ;
  assign n41923 = n5639 | n7661 ;
  assign n41924 = n7466 & ~n41923 ;
  assign n41925 = n9837 & ~n41924 ;
  assign n41926 = n7772 & ~n7974 ;
  assign n41927 = n3869 & n41926 ;
  assign n41928 = n41927 ^ n32476 ^ n26779 ;
  assign n41929 = n24191 & n41928 ;
  assign n41930 = n2769 & n41929 ;
  assign n41931 = ~n8545 & n31201 ;
  assign n41932 = n41931 ^ n9223 ^ 1'b0 ;
  assign n41933 = n41149 ^ n28711 ^ n11185 ;
  assign n41934 = n18833 | n40957 ;
  assign n41935 = n41934 ^ n8223 ^ 1'b0 ;
  assign n41936 = n41935 ^ n38011 ^ n29983 ;
  assign n41937 = n36098 ^ n35359 ^ n28607 ;
  assign n41941 = n5226 & ~n18944 ;
  assign n41942 = n41941 ^ n23705 ^ 1'b0 ;
  assign n41938 = n27178 & ~n34434 ;
  assign n41939 = ~n14076 & n41938 ;
  assign n41940 = n18737 & ~n41939 ;
  assign n41943 = n41942 ^ n41940 ^ 1'b0 ;
  assign n41944 = n4232 | n11903 ;
  assign n41946 = ~n14380 & n21578 ;
  assign n41947 = n41946 ^ n36960 ^ 1'b0 ;
  assign n41948 = ( n6965 & ~n11415 ) | ( n6965 & n41947 ) | ( ~n11415 & n41947 ) ;
  assign n41945 = n11493 | n41138 ;
  assign n41949 = n41948 ^ n41945 ^ 1'b0 ;
  assign n41950 = n10321 & ~n17469 ;
  assign n41951 = n41950 ^ n28053 ^ 1'b0 ;
  assign n41952 = n28558 ^ n27345 ^ 1'b0 ;
  assign n41953 = ( ~n12060 & n24940 ) | ( ~n12060 & n41952 ) | ( n24940 & n41952 ) ;
  assign n41954 = n1283 & n6080 ;
  assign n41955 = n41954 ^ n20019 ^ 1'b0 ;
  assign n41956 = n41955 ^ n5834 ^ 1'b0 ;
  assign n41957 = ~n1636 & n41956 ;
  assign n41958 = ( n981 & ~n9866 ) | ( n981 & n11663 ) | ( ~n9866 & n11663 ) ;
  assign n41959 = n41958 ^ n21624 ^ n13572 ;
  assign n41960 = ( ~n30202 & n41957 ) | ( ~n30202 & n41959 ) | ( n41957 & n41959 ) ;
  assign n41961 = n41960 ^ n26133 ^ n25079 ;
  assign n41962 = x25 & ~n34223 ;
  assign n41963 = n19634 & n41962 ;
  assign n41964 = n41963 ^ n12096 ^ 1'b0 ;
  assign n41965 = n41612 ^ n36484 ^ 1'b0 ;
  assign n41966 = n37393 & ~n41965 ;
  assign n41967 = ( n3679 & ~n10053 ) | ( n3679 & n11186 ) | ( ~n10053 & n11186 ) ;
  assign n41968 = n41967 ^ n19268 ^ 1'b0 ;
  assign n41969 = n22492 ^ n10274 ^ 1'b0 ;
  assign n41970 = n32885 ^ n9611 ^ 1'b0 ;
  assign n41971 = n8951 | n41970 ;
  assign n41972 = n41971 ^ n21097 ^ n16094 ;
  assign n41973 = n41972 ^ n15250 ^ n7568 ;
  assign n41974 = n41947 ^ n21761 ^ n895 ;
  assign n41975 = ( n9104 & ~n19551 ) | ( n9104 & n19740 ) | ( ~n19551 & n19740 ) ;
  assign n41976 = n41975 ^ n27941 ^ n5379 ;
  assign n41977 = ( n2458 & n3237 ) | ( n2458 & n41976 ) | ( n3237 & n41976 ) ;
  assign n41978 = n10068 | n26303 ;
  assign n41979 = ( x166 & n3581 ) | ( x166 & n17463 ) | ( n3581 & n17463 ) ;
  assign n41980 = n23016 ^ n7848 ^ 1'b0 ;
  assign n41981 = ~n41979 & n41980 ;
  assign n41982 = ~n41978 & n41981 ;
  assign n41983 = n6413 ^ n1576 ^ 1'b0 ;
  assign n41984 = ~n13734 & n41983 ;
  assign n41985 = n16403 | n35154 ;
  assign n41986 = n7081 ^ n2951 ^ n2780 ;
  assign n41987 = n34374 ^ n23665 ^ 1'b0 ;
  assign n41988 = n13214 & ~n33106 ;
  assign n41989 = ~n12476 & n41988 ;
  assign n41990 = n29872 & n32442 ;
  assign n41991 = ( x100 & n40082 ) | ( x100 & n41990 ) | ( n40082 & n41990 ) ;
  assign n41992 = ( ~n8895 & n11882 ) | ( ~n8895 & n17412 ) | ( n11882 & n17412 ) ;
  assign n41993 = n41992 ^ n33511 ^ 1'b0 ;
  assign n41994 = ~n41991 & n41993 ;
  assign n41995 = n3297 & n8311 ;
  assign n41996 = n41995 ^ n33517 ^ 1'b0 ;
  assign n41997 = n14775 | n25151 ;
  assign n41998 = n23844 ^ n21573 ^ n13846 ;
  assign n41999 = ( n19709 & n40564 ) | ( n19709 & n41998 ) | ( n40564 & n41998 ) ;
  assign n42000 = ( n20699 & ~n34982 ) | ( n20699 & n41999 ) | ( ~n34982 & n41999 ) ;
  assign n42001 = n8237 ^ n2936 ^ 1'b0 ;
  assign n42002 = ~n7032 & n42001 ;
  assign n42003 = n42000 | n42002 ;
  assign n42004 = n4670 & n11114 ;
  assign n42005 = n42004 ^ n29195 ^ 1'b0 ;
  assign n42006 = ( n22775 & n23933 ) | ( n22775 & ~n28554 ) | ( n23933 & ~n28554 ) ;
  assign n42007 = n4447 & n30892 ;
  assign n42008 = n42007 ^ n41880 ^ 1'b0 ;
  assign n42009 = n19484 ^ n7182 ^ 1'b0 ;
  assign n42010 = ~n11219 & n42009 ;
  assign n42011 = n42010 ^ n34206 ^ n9390 ;
  assign n42012 = ( n15929 & n26321 ) | ( n15929 & ~n42011 ) | ( n26321 & ~n42011 ) ;
  assign n42013 = n11018 & ~n19261 ;
  assign n42014 = n22737 ^ n7982 ^ 1'b0 ;
  assign n42015 = ~n19294 & n42014 ;
  assign n42016 = n4129 & n34576 ;
  assign n42017 = n11511 ^ n5589 ^ n2188 ;
  assign n42018 = n21520 & ~n42017 ;
  assign n42019 = ~n36577 & n42018 ;
  assign n42020 = n28941 ^ n19094 ^ 1'b0 ;
  assign n42021 = n9011 & ~n42020 ;
  assign n42022 = n2095 & ~n13138 ;
  assign n42023 = n42022 ^ n15200 ^ 1'b0 ;
  assign n42028 = ( n4690 & n5530 ) | ( n4690 & ~n39938 ) | ( n5530 & ~n39938 ) ;
  assign n42029 = n20941 ^ n13768 ^ n8411 ;
  assign n42030 = ~n42028 & n42029 ;
  assign n42024 = n6316 ^ n1326 ^ 1'b0 ;
  assign n42025 = n6040 | n42024 ;
  assign n42026 = n34536 ^ n31591 ^ n24088 ;
  assign n42027 = ~n42025 & n42026 ;
  assign n42031 = n42030 ^ n42027 ^ n17429 ;
  assign n42032 = n34875 ^ n21870 ^ n8942 ;
  assign n42036 = n26602 | n41226 ;
  assign n42033 = n5386 | n14978 ;
  assign n42034 = n6514 & ~n42033 ;
  assign n42035 = n32013 | n42034 ;
  assign n42037 = n42036 ^ n42035 ^ 1'b0 ;
  assign n42038 = n22246 ^ n1158 ^ 1'b0 ;
  assign n42039 = n619 | n8393 ;
  assign n42040 = n42039 ^ n6424 ^ 1'b0 ;
  assign n42043 = n8098 ^ x108 ^ 1'b0 ;
  assign n42044 = n3240 & n11037 ;
  assign n42045 = n42043 & n42044 ;
  assign n42041 = n17838 | n27644 ;
  assign n42042 = ( ~n5162 & n19227 ) | ( ~n5162 & n42041 ) | ( n19227 & n42041 ) ;
  assign n42046 = n42045 ^ n42042 ^ 1'b0 ;
  assign n42047 = n14670 ^ n6499 ^ n1928 ;
  assign n42048 = ~n16354 & n17429 ;
  assign n42049 = ( ~n9296 & n14120 ) | ( ~n9296 & n20428 ) | ( n14120 & n20428 ) ;
  assign n42050 = n15142 & ~n42049 ;
  assign n42051 = n10621 & ~n42050 ;
  assign n42052 = n41290 ^ n28333 ^ n15114 ;
  assign n42053 = n35179 & n42052 ;
  assign n42054 = n2373 ^ n550 ^ 1'b0 ;
  assign n42055 = n29917 & ~n42054 ;
  assign n42056 = ~n16003 & n42055 ;
  assign n42057 = n42056 ^ n30376 ^ 1'b0 ;
  assign n42058 = n42057 ^ n33433 ^ n26944 ;
  assign n42059 = n8193 & ~n33563 ;
  assign n42060 = n20459 & n42059 ;
  assign n42061 = n42060 ^ n20412 ^ 1'b0 ;
  assign n42063 = n986 & ~n11626 ;
  assign n42064 = n42063 ^ n7220 ^ 1'b0 ;
  assign n42062 = n40857 ^ n38183 ^ 1'b0 ;
  assign n42065 = n42064 ^ n42062 ^ n12681 ;
  assign n42066 = n39542 ^ n32363 ^ n11733 ;
  assign n42067 = n37078 & n42066 ;
  assign n42068 = n6826 & n26246 ;
  assign n42069 = n8364 & ~n16911 ;
  assign n42071 = n28157 ^ n7098 ^ 1'b0 ;
  assign n42072 = n7796 & n42071 ;
  assign n42070 = n3394 & n19285 ;
  assign n42073 = n42072 ^ n42070 ^ 1'b0 ;
  assign n42074 = n6433 & ~n16415 ;
  assign n42075 = n280 | n8077 ;
  assign n42076 = n42074 | n42075 ;
  assign n42077 = n42076 ^ n21321 ^ 1'b0 ;
  assign n42078 = n20591 ^ n20200 ^ n16445 ;
  assign n42079 = n42078 ^ n33124 ^ n4260 ;
  assign n42081 = n22476 ^ n3264 ^ 1'b0 ;
  assign n42082 = n21333 | n42081 ;
  assign n42080 = n24890 ^ n5996 ^ 1'b0 ;
  assign n42083 = n42082 ^ n42080 ^ 1'b0 ;
  assign n42084 = n21500 | n35447 ;
  assign n42085 = n42084 ^ n23797 ^ 1'b0 ;
  assign n42086 = n8288 ^ n7396 ^ n623 ;
  assign n42087 = ( n9837 & ~n33310 ) | ( n9837 & n42086 ) | ( ~n33310 & n42086 ) ;
  assign n42088 = n38345 ^ n23955 ^ 1'b0 ;
  assign n42089 = n42087 | n42088 ;
  assign n42090 = n25179 ^ n18602 ^ n13407 ;
  assign n42091 = n42090 ^ n30886 ^ n22513 ;
  assign n42092 = n42091 ^ n39746 ^ n35878 ;
  assign n42093 = n3247 & n9939 ;
  assign n42099 = n901 & n6137 ;
  assign n42100 = n6727 & n42099 ;
  assign n42094 = n29965 ^ n10685 ^ 1'b0 ;
  assign n42095 = ~n7562 & n28820 ;
  assign n42096 = n23091 & n42095 ;
  assign n42097 = n42094 & ~n42096 ;
  assign n42098 = n42097 ^ n10013 ^ 1'b0 ;
  assign n42101 = n42100 ^ n42098 ^ 1'b0 ;
  assign n42102 = n15810 | n16197 ;
  assign n42103 = ~n9853 & n20895 ;
  assign n42104 = n42103 ^ n23729 ^ n10251 ;
  assign n42105 = n13121 ^ x210 ^ 1'b0 ;
  assign n42106 = ~n9115 & n42105 ;
  assign n42107 = ( n28863 & n42104 ) | ( n28863 & ~n42106 ) | ( n42104 & ~n42106 ) ;
  assign n42108 = n38494 ^ n4303 ^ 1'b0 ;
  assign n42109 = ~n30648 & n42108 ;
  assign n42110 = ( n567 & ~n22132 ) | ( n567 & n42109 ) | ( ~n22132 & n42109 ) ;
  assign n42111 = n39846 ^ n20437 ^ 1'b0 ;
  assign n42112 = n12071 & n12400 ;
  assign n42113 = ~n20973 & n42112 ;
  assign n42114 = n42113 ^ n24767 ^ n24312 ;
  assign n42115 = n10090 | n13007 ;
  assign n42116 = n42115 ^ n40040 ^ 1'b0 ;
  assign n42117 = ( n1685 & ~n12034 ) | ( n1685 & n42116 ) | ( ~n12034 & n42116 ) ;
  assign n42118 = n32610 ^ n13081 ^ 1'b0 ;
  assign n42119 = n42118 ^ n33044 ^ 1'b0 ;
  assign n42120 = ~n4927 & n7079 ;
  assign n42121 = n42120 ^ n9461 ^ 1'b0 ;
  assign n42122 = ~n12401 & n23818 ;
  assign n42123 = n42121 & n42122 ;
  assign n42124 = n27640 ^ n2850 ^ 1'b0 ;
  assign n42125 = ~n14809 & n42124 ;
  assign n42126 = n10474 & ~n17817 ;
  assign n42127 = n17817 & n42126 ;
  assign n42128 = n8307 | n9897 ;
  assign n42129 = n42127 & ~n42128 ;
  assign n42130 = n27295 ^ n6788 ^ 1'b0 ;
  assign n42131 = n3866 | n42130 ;
  assign n42132 = n42131 ^ n7395 ^ 1'b0 ;
  assign n42133 = n2567 & ~n42132 ;
  assign n42134 = n36252 & ~n42133 ;
  assign n42135 = ( n36710 & ~n42129 ) | ( n36710 & n42134 ) | ( ~n42129 & n42134 ) ;
  assign n42136 = ( n5879 & ~n7740 ) | ( n5879 & n9332 ) | ( ~n7740 & n9332 ) ;
  assign n42137 = x76 & n42136 ;
  assign n42138 = n42137 ^ n14689 ^ 1'b0 ;
  assign n42139 = n22335 & n42138 ;
  assign n42140 = n9266 & ~n9736 ;
  assign n42141 = ~n19970 & n42140 ;
  assign n42142 = x202 | n24631 ;
  assign n42143 = n28494 ^ n20998 ^ n14427 ;
  assign n42144 = n22371 ^ n7037 ^ n704 ;
  assign n42145 = n21209 | n42144 ;
  assign n42146 = n42143 & ~n42145 ;
  assign n42147 = n30147 & ~n35245 ;
  assign n42148 = n31087 ^ n29000 ^ 1'b0 ;
  assign n42149 = ~n7214 & n42148 ;
  assign n42150 = n22510 ^ n1564 ^ 1'b0 ;
  assign n42151 = n42149 & ~n42150 ;
  assign n42153 = n8415 & ~n40253 ;
  assign n42154 = n42153 ^ n6428 ^ 1'b0 ;
  assign n42152 = n1463 & ~n18911 ;
  assign n42155 = n42154 ^ n42152 ^ 1'b0 ;
  assign n42156 = ( n15487 & n39754 ) | ( n15487 & ~n41532 ) | ( n39754 & ~n41532 ) ;
  assign n42157 = n3597 & ~n4913 ;
  assign n42158 = n2256 & n29741 ;
  assign n42159 = ~n4745 & n42158 ;
  assign n42160 = ( n7644 & ~n11259 ) | ( n7644 & n42159 ) | ( ~n11259 & n42159 ) ;
  assign n42161 = n41109 | n42160 ;
  assign n42162 = n30647 & ~n42161 ;
  assign n42163 = n22832 ^ n21980 ^ n17456 ;
  assign n42164 = ~n26115 & n42163 ;
  assign n42165 = ~n654 & n42164 ;
  assign n42166 = n15836 ^ n3939 ^ 1'b0 ;
  assign n42167 = n2816 & n42166 ;
  assign n42168 = n11231 & n42167 ;
  assign n42169 = n42165 & n42168 ;
  assign n42170 = n7015 & ~n33724 ;
  assign n42171 = ~n25171 & n42170 ;
  assign n42172 = n36141 ^ n6075 ^ x196 ;
  assign n42173 = n42172 ^ n12743 ^ 1'b0 ;
  assign n42174 = ( n1138 & n24423 ) | ( n1138 & ~n37903 ) | ( n24423 & ~n37903 ) ;
  assign n42175 = n14276 | n17607 ;
  assign n42176 = n13384 ^ n3547 ^ 1'b0 ;
  assign n42177 = n16157 & n42176 ;
  assign n42178 = n8962 | n24667 ;
  assign n42179 = n42177 | n42178 ;
  assign n42180 = n33075 ^ n11214 ^ 1'b0 ;
  assign n42181 = n42180 ^ n30758 ^ 1'b0 ;
  assign n42182 = n15732 | n42181 ;
  assign n42183 = x175 | n42182 ;
  assign n42184 = n16545 ^ n3893 ^ 1'b0 ;
  assign n42185 = n9785 ^ n7851 ^ 1'b0 ;
  assign n42186 = ( n4251 & n34685 ) | ( n4251 & ~n42185 ) | ( n34685 & ~n42185 ) ;
  assign n42187 = n42186 ^ n26531 ^ 1'b0 ;
  assign n42188 = n30366 ^ n1629 ^ n616 ;
  assign n42191 = n16073 | n39573 ;
  assign n42192 = n42191 ^ n26107 ^ 1'b0 ;
  assign n42189 = n11535 ^ n2165 ^ n457 ;
  assign n42190 = ( n19629 & ~n23900 ) | ( n19629 & n42189 ) | ( ~n23900 & n42189 ) ;
  assign n42193 = n42192 ^ n42190 ^ n17343 ;
  assign n42194 = n22580 | n24890 ;
  assign n42195 = n42194 ^ n35229 ^ 1'b0 ;
  assign n42196 = ~n5582 & n35138 ;
  assign n42197 = n24048 & ~n42196 ;
  assign n42198 = n42195 & n42197 ;
  assign n42199 = n427 | n16106 ;
  assign n42200 = n19431 & ~n42199 ;
  assign n42201 = n42200 ^ n18780 ^ n7893 ;
  assign n42202 = n31956 ^ n3219 ^ 1'b0 ;
  assign n42203 = n25023 | n27614 ;
  assign n42204 = n19759 & n32695 ;
  assign n42205 = n42204 ^ n6850 ^ 1'b0 ;
  assign n42206 = n10654 & ~n12110 ;
  assign n42208 = n3437 | n5803 ;
  assign n42209 = n42208 ^ n26329 ^ n3983 ;
  assign n42207 = ( n8932 & ~n10954 ) | ( n8932 & n32881 ) | ( ~n10954 & n32881 ) ;
  assign n42210 = n42209 ^ n42207 ^ 1'b0 ;
  assign n42211 = n8358 & n42210 ;
  assign n42212 = ( n11276 & ~n28214 ) | ( n11276 & n42211 ) | ( ~n28214 & n42211 ) ;
  assign n42213 = n40349 ^ n35598 ^ 1'b0 ;
  assign n42214 = n10038 & ~n16767 ;
  assign n42215 = n42214 ^ n30325 ^ 1'b0 ;
  assign n42216 = n42215 ^ n19490 ^ 1'b0 ;
  assign n42217 = n42216 ^ n5701 ^ 1'b0 ;
  assign n42218 = n10251 | n27478 ;
  assign n42220 = n19484 ^ n3573 ^ n1951 ;
  assign n42219 = n25632 ^ n1082 ^ 1'b0 ;
  assign n42221 = n42220 ^ n42219 ^ 1'b0 ;
  assign n42222 = n1243 | n36303 ;
  assign n42223 = n2760 & ~n42222 ;
  assign n42224 = n11351 | n38601 ;
  assign n42225 = n18116 & ~n42224 ;
  assign n42226 = n42225 ^ n8477 ^ 1'b0 ;
  assign n42227 = n34576 & ~n42226 ;
  assign n42228 = n31608 ^ n6174 ^ 1'b0 ;
  assign n42229 = n11774 & n31285 ;
  assign n42230 = n24220 & ~n42229 ;
  assign n42231 = n42228 & n42230 ;
  assign n42233 = n3940 | n16923 ;
  assign n42232 = ~n675 & n5858 ;
  assign n42234 = n42233 ^ n42232 ^ n23188 ;
  assign n42235 = n13070 ^ n13033 ^ 1'b0 ;
  assign n42236 = n39557 ^ n2922 ^ 1'b0 ;
  assign n42237 = ~n30824 & n42236 ;
  assign n42238 = n6420 & n6594 ;
  assign n42239 = n42238 ^ n9484 ^ 1'b0 ;
  assign n42240 = n379 & n42239 ;
  assign n42241 = n7638 | n32383 ;
  assign n42242 = n6875 & ~n7754 ;
  assign n42243 = n42242 ^ n13357 ^ 1'b0 ;
  assign n42244 = ( n11989 & n12968 ) | ( n11989 & ~n33116 ) | ( n12968 & ~n33116 ) ;
  assign n42245 = n34850 ^ n31825 ^ n19980 ;
  assign n42247 = n38441 ^ n15917 ^ n9685 ;
  assign n42246 = ~n15392 & n37462 ;
  assign n42248 = n42247 ^ n42246 ^ 1'b0 ;
  assign n42249 = ~n1051 & n2280 ;
  assign n42250 = n42249 ^ n12504 ^ 1'b0 ;
  assign n42251 = ( x43 & ~n21113 ) | ( x43 & n25451 ) | ( ~n21113 & n25451 ) ;
  assign n42252 = n42250 | n42251 ;
  assign n42253 = n672 | n14275 ;
  assign n42254 = n42253 ^ n28803 ^ 1'b0 ;
  assign n42255 = n31209 & ~n38832 ;
  assign n42256 = ( ~n1406 & n1780 ) | ( ~n1406 & n15892 ) | ( n1780 & n15892 ) ;
  assign n42257 = x250 & n14189 ;
  assign n42258 = n5592 & n42257 ;
  assign n42259 = n16499 ^ n2690 ^ 1'b0 ;
  assign n42260 = ~n42258 & n42259 ;
  assign n42261 = n13404 & ~n25402 ;
  assign n42262 = n8018 | n42261 ;
  assign n42263 = n42260 | n42262 ;
  assign n42264 = ~n4893 & n11550 ;
  assign n42265 = ~n5855 & n42264 ;
  assign n42266 = n30809 ^ n15130 ^ 1'b0 ;
  assign n42267 = n4857 | n42266 ;
  assign n42268 = n42267 ^ n36087 ^ n31967 ;
  assign n42269 = n5841 | n38575 ;
  assign n42270 = n32744 & ~n42269 ;
  assign n42271 = n25786 & ~n42270 ;
  assign n42272 = n697 | n28923 ;
  assign n42273 = n17353 ^ n2412 ^ 1'b0 ;
  assign n42274 = ~n17558 & n33457 ;
  assign n42275 = n42274 ^ n6881 ^ 1'b0 ;
  assign n42276 = n30699 & ~n42275 ;
  assign n42277 = ~n42273 & n42276 ;
  assign n42278 = n38247 & n42277 ;
  assign n42279 = n16872 ^ n12544 ^ n9641 ;
  assign n42280 = ~n13954 & n42279 ;
  assign n42281 = n37701 ^ n24432 ^ 1'b0 ;
  assign n42282 = ~n9986 & n42281 ;
  assign n42283 = n20862 & ~n28339 ;
  assign n42284 = n42283 ^ n11670 ^ 1'b0 ;
  assign n42285 = n2263 | n42284 ;
  assign n42286 = n6218 & ~n42285 ;
  assign n42287 = n42286 ^ n29772 ^ 1'b0 ;
  assign n42288 = n32975 | n42287 ;
  assign n42289 = n42282 & ~n42288 ;
  assign n42290 = n42280 & n42289 ;
  assign n42291 = n42288 ^ n13810 ^ 1'b0 ;
  assign n42292 = n41515 ^ n1727 ^ 1'b0 ;
  assign n42293 = n42292 ^ n9461 ^ n2603 ;
  assign n42294 = n42293 ^ n24933 ^ 1'b0 ;
  assign n42295 = n23884 ^ n15522 ^ 1'b0 ;
  assign n42296 = ( ~n2427 & n10854 ) | ( ~n2427 & n36796 ) | ( n10854 & n36796 ) ;
  assign n42297 = n42296 ^ x120 ^ 1'b0 ;
  assign n42298 = n42297 ^ n3731 ^ 1'b0 ;
  assign n42299 = n30734 & ~n42298 ;
  assign n42300 = n4811 ^ n3396 ^ 1'b0 ;
  assign n42301 = n42299 & ~n42300 ;
  assign n42302 = n6075 | n31467 ;
  assign n42303 = n25977 ^ n11882 ^ n10847 ;
  assign n42304 = n19871 ^ n15584 ^ 1'b0 ;
  assign n42305 = n8486 & n16591 ;
  assign n42306 = ~n28634 & n42305 ;
  assign n42307 = n42306 ^ n24164 ^ 1'b0 ;
  assign n42308 = n42307 ^ n5715 ^ n2452 ;
  assign n42309 = n8286 & n25220 ;
  assign n42310 = ~n6996 & n42309 ;
  assign n42311 = n42310 ^ n14186 ^ 1'b0 ;
  assign n42312 = ~n3669 & n37717 ;
  assign n42313 = n42312 ^ n39709 ^ n5926 ;
  assign n42314 = n10450 | n42077 ;
  assign n42315 = n12158 | n42314 ;
  assign n42318 = n2823 | n19199 ;
  assign n42316 = n1179 & ~n29985 ;
  assign n42317 = ( n1637 & ~n7570 ) | ( n1637 & n42316 ) | ( ~n7570 & n42316 ) ;
  assign n42319 = n42318 ^ n42317 ^ 1'b0 ;
  assign n42320 = n12390 & ~n31074 ;
  assign n42321 = n9527 ^ n9518 ^ 1'b0 ;
  assign n42322 = n11474 | n42321 ;
  assign n42323 = ( ~n1162 & n13986 ) | ( ~n1162 & n42322 ) | ( n13986 & n42322 ) ;
  assign n42324 = n28239 | n42323 ;
  assign n42325 = ( n16376 & ~n21604 ) | ( n16376 & n42324 ) | ( ~n21604 & n42324 ) ;
  assign n42326 = n5181 & n14985 ;
  assign n42327 = n6772 ^ n4662 ^ 1'b0 ;
  assign n42328 = n9929 & n20602 ;
  assign n42329 = n31552 ^ n23775 ^ 1'b0 ;
  assign n42330 = n6618 & ~n11168 ;
  assign n42331 = n42330 ^ n4122 ^ 1'b0 ;
  assign n42332 = n7578 ^ n805 ^ 1'b0 ;
  assign n42333 = n9622 & n42332 ;
  assign n42334 = n42333 ^ n28937 ^ n23877 ;
  assign n42335 = ( ~n4525 & n5495 ) | ( ~n4525 & n27280 ) | ( n5495 & n27280 ) ;
  assign n42336 = n3030 & ~n42335 ;
  assign n42337 = n4707 | n16653 ;
  assign n42338 = n15210 ^ n8846 ^ 1'b0 ;
  assign n42339 = n42337 & n42338 ;
  assign n42340 = n32551 & n42339 ;
  assign n42341 = n4490 | n38802 ;
  assign n42342 = ~n12754 & n28914 ;
  assign n42343 = n29819 & n42342 ;
  assign n42344 = n11025 & n11693 ;
  assign n42345 = n42344 ^ n22476 ^ 1'b0 ;
  assign n42346 = n42345 ^ n26244 ^ n17282 ;
  assign n42348 = n10257 ^ n3694 ^ 1'b0 ;
  assign n42349 = ~n12375 & n42348 ;
  assign n42347 = n4138 & ~n9153 ;
  assign n42350 = n42349 ^ n42347 ^ 1'b0 ;
  assign n42351 = ( ~n21059 & n24143 ) | ( ~n21059 & n42350 ) | ( n24143 & n42350 ) ;
  assign n42352 = n8404 | n25865 ;
  assign n42353 = n42352 ^ n37879 ^ 1'b0 ;
  assign n42354 = n29776 ^ n27476 ^ 1'b0 ;
  assign n42355 = n42353 & ~n42354 ;
  assign n42356 = n7132 | n24157 ;
  assign n42357 = n19797 & ~n42356 ;
  assign n42358 = n28419 ^ n3282 ^ 1'b0 ;
  assign n42359 = ~n42357 & n42358 ;
  assign n42360 = n20952 ^ n19529 ^ n7030 ;
  assign n42361 = n14234 ^ n13348 ^ 1'b0 ;
  assign n42362 = n7586 & ~n42361 ;
  assign n42363 = n12778 & n31091 ;
  assign n42364 = n42363 ^ n21838 ^ 1'b0 ;
  assign n42365 = n14779 | n34442 ;
  assign n42366 = n27190 | n42365 ;
  assign n42367 = ~n19190 & n42366 ;
  assign n42368 = n42367 ^ n24518 ^ 1'b0 ;
  assign n42369 = n42368 ^ n7376 ^ 1'b0 ;
  assign n42370 = n462 & n42369 ;
  assign n42371 = ~n35932 & n42370 ;
  assign n42372 = n21717 ^ n8275 ^ 1'b0 ;
  assign n42373 = n30454 & ~n39716 ;
  assign n42374 = n30792 ^ n14661 ^ n7621 ;
  assign n42375 = n24058 ^ n14731 ^ 1'b0 ;
  assign n42376 = n6968 | n42375 ;
  assign n42377 = n42376 ^ n9288 ^ 1'b0 ;
  assign n42378 = n9513 ^ n569 ^ 1'b0 ;
  assign n42379 = n5662 & n42378 ;
  assign n42380 = n8483 ^ n1633 ^ 1'b0 ;
  assign n42381 = n42379 & ~n42380 ;
  assign n42382 = n7761 ^ n7001 ^ 1'b0 ;
  assign n42383 = ~n11802 & n33079 ;
  assign n42384 = n42383 ^ n17007 ^ 1'b0 ;
  assign n42385 = n42384 ^ n30037 ^ n1760 ;
  assign n42386 = n7016 | n42385 ;
  assign n42387 = n29540 ^ n16519 ^ 1'b0 ;
  assign n42388 = n28801 ^ n14215 ^ n5963 ;
  assign n42389 = n31096 ^ n22208 ^ n5391 ;
  assign n42390 = ( n4068 & ~n42388 ) | ( n4068 & n42389 ) | ( ~n42388 & n42389 ) ;
  assign n42391 = ( n704 & n20017 ) | ( n704 & n25278 ) | ( n20017 & n25278 ) ;
  assign n42392 = n27115 ^ n7974 ^ 1'b0 ;
  assign n42393 = ~n12036 & n42392 ;
  assign n42394 = ~n28383 & n35469 ;
  assign n42395 = n28383 & n42394 ;
  assign n42396 = n42395 ^ n25371 ^ 1'b0 ;
  assign n42397 = n7481 & ~n42396 ;
  assign n42398 = n10932 & ~n23355 ;
  assign n42399 = n32116 & n42398 ;
  assign n42400 = ( ~n4874 & n23217 ) | ( ~n4874 & n42399 ) | ( n23217 & n42399 ) ;
  assign n42401 = n42397 & n42400 ;
  assign n42402 = ~n8048 & n24828 ;
  assign n42403 = n9158 & n42402 ;
  assign n42404 = n8801 | n27021 ;
  assign n42405 = n8969 ^ n5102 ^ 1'b0 ;
  assign n42406 = n30629 ^ n29988 ^ n9731 ;
  assign n42407 = n41676 & n42406 ;
  assign n42408 = n33000 ^ n11665 ^ 1'b0 ;
  assign n42411 = n7854 ^ n4219 ^ 1'b0 ;
  assign n42412 = n42411 ^ n33200 ^ 1'b0 ;
  assign n42413 = n9122 | n42412 ;
  assign n42409 = n39473 ^ n2374 ^ 1'b0 ;
  assign n42410 = n24521 | n42409 ;
  assign n42414 = n42413 ^ n42410 ^ 1'b0 ;
  assign n42415 = n17562 ^ n13204 ^ 1'b0 ;
  assign n42416 = n18091 & ~n42415 ;
  assign n42417 = n453 | n1465 ;
  assign n42418 = n9351 | n42417 ;
  assign n42419 = n4606 & ~n9885 ;
  assign n42420 = n42419 ^ n22736 ^ 1'b0 ;
  assign n42421 = n17662 & n20223 ;
  assign n42422 = n42420 & n42421 ;
  assign n42423 = n13397 & n22644 ;
  assign n42424 = n14000 & n42423 ;
  assign n42425 = n30498 & ~n42424 ;
  assign n42426 = ( n28719 & n34909 ) | ( n28719 & ~n42425 ) | ( n34909 & ~n42425 ) ;
  assign n42428 = ( n2491 & n17691 ) | ( n2491 & n29425 ) | ( n17691 & n29425 ) ;
  assign n42427 = n603 & n11428 ;
  assign n42429 = n42428 ^ n42427 ^ 1'b0 ;
  assign n42430 = n22163 ^ n1527 ^ 1'b0 ;
  assign n42431 = n11371 & ~n42430 ;
  assign n42432 = ~n8116 & n42431 ;
  assign n42433 = n16383 ^ n8634 ^ n4149 ;
  assign n42434 = n28240 & n42433 ;
  assign n42435 = n1374 | n15971 ;
  assign n42436 = n42434 & ~n42435 ;
  assign n42437 = n23893 ^ n6986 ^ 1'b0 ;
  assign n42438 = n22759 & ~n42437 ;
  assign n42439 = ~n6367 & n33919 ;
  assign n42440 = n23045 ^ n20154 ^ 1'b0 ;
  assign n42441 = n15788 ^ n13988 ^ n9292 ;
  assign n42442 = n13452 | n42441 ;
  assign n42443 = n7837 & ~n10829 ;
  assign n42444 = ~n31044 & n42443 ;
  assign n42445 = n21260 ^ n2779 ^ 1'b0 ;
  assign n42446 = n4191 & n42445 ;
  assign n42447 = n1053 & n33835 ;
  assign n42448 = n23590 | n34612 ;
  assign n42449 = n2059 & n18794 ;
  assign n42450 = n10155 & ~n32954 ;
  assign n42451 = ~n24445 & n42450 ;
  assign n42452 = ( ~n16340 & n24386 ) | ( ~n16340 & n33493 ) | ( n24386 & n33493 ) ;
  assign n42453 = n16246 | n16847 ;
  assign n42454 = n42453 ^ n19499 ^ 1'b0 ;
  assign n42455 = n42452 & ~n42454 ;
  assign n42458 = ( n6262 & n11005 ) | ( n6262 & ~n17191 ) | ( n11005 & ~n17191 ) ;
  assign n42456 = n24566 | n34196 ;
  assign n42457 = n42456 ^ n19284 ^ 1'b0 ;
  assign n42459 = n42458 ^ n42457 ^ n28669 ;
  assign n42460 = ~n8382 & n35329 ;
  assign n42461 = ~n42189 & n42460 ;
  assign n42462 = n34171 & n42461 ;
  assign n42463 = n33384 ^ n25040 ^ n4061 ;
  assign n42464 = n409 & ~n27737 ;
  assign n42465 = n28508 ^ n21098 ^ 1'b0 ;
  assign n42466 = n20649 & n42465 ;
  assign n42467 = ( n5462 & n9100 ) | ( n5462 & ~n20927 ) | ( n9100 & ~n20927 ) ;
  assign n42468 = n42467 ^ n13219 ^ 1'b0 ;
  assign n42471 = n15438 ^ n7696 ^ n3955 ;
  assign n42472 = n4416 & n42471 ;
  assign n42473 = n42472 ^ n20480 ^ 1'b0 ;
  assign n42474 = n11231 ^ n7361 ^ 1'b0 ;
  assign n42475 = n42473 | n42474 ;
  assign n42469 = n18251 ^ n7459 ^ 1'b0 ;
  assign n42470 = ( n3047 & ~n21546 ) | ( n3047 & n42469 ) | ( ~n21546 & n42469 ) ;
  assign n42476 = n42475 ^ n42470 ^ 1'b0 ;
  assign n42477 = ( n4719 & n15953 ) | ( n4719 & ~n17817 ) | ( n15953 & ~n17817 ) ;
  assign n42478 = n42477 ^ n6946 ^ 1'b0 ;
  assign n42479 = n287 & ~n10859 ;
  assign n42480 = n42479 ^ n9927 ^ n4840 ;
  assign n42481 = n42480 ^ n24780 ^ 1'b0 ;
  assign n42482 = n11200 | n21654 ;
  assign n42483 = n27141 | n42482 ;
  assign n42484 = n42483 ^ n33467 ^ 1'b0 ;
  assign n42485 = n42484 ^ n39855 ^ 1'b0 ;
  assign n42486 = ~n5460 & n22799 ;
  assign n42487 = n2921 & n42486 ;
  assign n42488 = n1265 & n2703 ;
  assign n42489 = n12526 | n42488 ;
  assign n42490 = n42487 & ~n42489 ;
  assign n42491 = n42490 ^ n19580 ^ 1'b0 ;
  assign n42492 = n33162 | n37294 ;
  assign n42493 = n26704 ^ n14712 ^ 1'b0 ;
  assign n42494 = ~n7392 & n42493 ;
  assign n42495 = n28769 ^ n3652 ^ 1'b0 ;
  assign n42496 = n41675 ^ n20250 ^ 1'b0 ;
  assign n42497 = n26330 ^ n9207 ^ 1'b0 ;
  assign n42498 = ~n29524 & n42497 ;
  assign n42499 = ( n9906 & n13527 ) | ( n9906 & n40122 ) | ( n13527 & n40122 ) ;
  assign n42500 = n12210 ^ n3859 ^ 1'b0 ;
  assign n42501 = n28611 & n42500 ;
  assign n42502 = n2245 & ~n5001 ;
  assign n42503 = n42502 ^ n9702 ^ 1'b0 ;
  assign n42504 = n23907 ^ n11963 ^ 1'b0 ;
  assign n42505 = n42503 & n42504 ;
  assign n42506 = n12787 ^ n8926 ^ n890 ;
  assign n42507 = n28033 & n42506 ;
  assign n42508 = x113 & n42507 ;
  assign n42509 = ~n15486 & n42508 ;
  assign n42510 = n7473 | n11888 ;
  assign n42511 = ( n1504 & n10189 ) | ( n1504 & n23563 ) | ( n10189 & n23563 ) ;
  assign n42516 = n18306 ^ n10483 ^ n10052 ;
  assign n42517 = ( n7486 & ~n17979 ) | ( n7486 & n42516 ) | ( ~n17979 & n42516 ) ;
  assign n42512 = n15677 ^ n11355 ^ n10201 ;
  assign n42513 = n3826 & ~n42512 ;
  assign n42514 = n42513 ^ n23068 ^ 1'b0 ;
  assign n42515 = n42514 ^ n33773 ^ n7396 ;
  assign n42518 = n42517 ^ n42515 ^ n36223 ;
  assign n42519 = ( ~n584 & n19143 ) | ( ~n584 & n19621 ) | ( n19143 & n19621 ) ;
  assign n42520 = n17473 & ~n42292 ;
  assign n42521 = n42520 ^ n41543 ^ 1'b0 ;
  assign n42522 = ~n18836 & n19569 ;
  assign n42523 = ~n11313 & n37524 ;
  assign n42526 = n38175 ^ n2250 ^ 1'b0 ;
  assign n42524 = ~n7787 & n20145 ;
  assign n42525 = n42524 ^ n14729 ^ n11157 ;
  assign n42527 = n42526 ^ n42525 ^ 1'b0 ;
  assign n42528 = n42523 | n42527 ;
  assign n42529 = n25464 ^ n19058 ^ 1'b0 ;
  assign n42530 = n13684 & ~n26184 ;
  assign n42531 = n42530 ^ n29346 ^ 1'b0 ;
  assign n42532 = n9276 | n42531 ;
  assign n42533 = n42532 ^ n10317 ^ 1'b0 ;
  assign n42534 = ~n588 & n24845 ;
  assign n42535 = n5518 & n42534 ;
  assign n42536 = n24250 & n42535 ;
  assign n42537 = n42536 ^ n32891 ^ 1'b0 ;
  assign n42538 = n40821 ^ n26912 ^ n8406 ;
  assign n42539 = n33931 ^ n8991 ^ 1'b0 ;
  assign n42540 = n10121 & n30922 ;
  assign n42541 = n42540 ^ n8065 ^ 1'b0 ;
  assign n42542 = n31779 | n42541 ;
  assign n42543 = n42512 ^ n16215 ^ 1'b0 ;
  assign n42544 = n42542 & ~n42543 ;
  assign n42545 = n5472 & ~n42544 ;
  assign n42546 = n17292 & n42545 ;
  assign n42547 = n13888 ^ n6459 ^ 1'b0 ;
  assign n42548 = n5287 ^ n4112 ^ 1'b0 ;
  assign n42549 = n42548 ^ n983 ^ 1'b0 ;
  assign n42550 = ~n42547 & n42549 ;
  assign n42551 = n1727 & n19388 ;
  assign n42552 = ~n35440 & n42551 ;
  assign n42553 = n7077 ^ n2877 ^ 1'b0 ;
  assign n42554 = n42553 ^ n19065 ^ 1'b0 ;
  assign n42555 = n2746 & ~n3029 ;
  assign n42556 = n41957 ^ n23361 ^ n9976 ;
  assign n42557 = ( n3379 & n31188 ) | ( n3379 & ~n42556 ) | ( n31188 & ~n42556 ) ;
  assign n42558 = n42557 ^ n33787 ^ 1'b0 ;
  assign n42560 = ( n15557 & n33231 ) | ( n15557 & n34829 ) | ( n33231 & n34829 ) ;
  assign n42559 = n5552 & n8406 ;
  assign n42561 = n42560 ^ n42559 ^ 1'b0 ;
  assign n42564 = n13100 ^ n6386 ^ x48 ;
  assign n42562 = ( n11934 & n16555 ) | ( n11934 & ~n28551 ) | ( n16555 & ~n28551 ) ;
  assign n42563 = ~n29511 & n42562 ;
  assign n42565 = n42564 ^ n42563 ^ 1'b0 ;
  assign n42568 = ~n13377 & n13860 ;
  assign n42569 = n42568 ^ n13177 ^ 1'b0 ;
  assign n42566 = n9737 & ~n18702 ;
  assign n42567 = ~n36346 & n42566 ;
  assign n42570 = n42569 ^ n42567 ^ 1'b0 ;
  assign n42571 = ( n2314 & n11606 ) | ( n2314 & n27099 ) | ( n11606 & n27099 ) ;
  assign n42572 = n18355 ^ n802 ^ 1'b0 ;
  assign n42573 = ( n15267 & ~n22497 ) | ( n15267 & n25224 ) | ( ~n22497 & n25224 ) ;
  assign n42574 = n8935 & ~n41138 ;
  assign n42575 = n3023 | n41160 ;
  assign n42576 = n42575 ^ n7111 ^ 1'b0 ;
  assign n42577 = n27652 ^ n22476 ^ n15252 ;
  assign n42578 = n29820 ^ n16617 ^ 1'b0 ;
  assign n42579 = n42577 & n42578 ;
  assign n42580 = n11210 & n15449 ;
  assign n42581 = n42580 ^ n25404 ^ 1'b0 ;
  assign n42582 = n5356 & ~n42581 ;
  assign n42583 = n9192 & n27449 ;
  assign n42584 = n4431 & n42583 ;
  assign n42585 = n42584 ^ n41164 ^ n25686 ;
  assign n42586 = ~n5541 & n18875 ;
  assign n42587 = ~n24104 & n42586 ;
  assign n42588 = n35952 & ~n42587 ;
  assign n42589 = n17587 & n42588 ;
  assign n42590 = ( ~n1843 & n13225 ) | ( ~n1843 & n32302 ) | ( n13225 & n32302 ) ;
  assign n42591 = ( n3328 & n42589 ) | ( n3328 & ~n42590 ) | ( n42589 & ~n42590 ) ;
  assign n42592 = n38285 ^ n4875 ^ 1'b0 ;
  assign n42593 = n37891 ^ n11308 ^ 1'b0 ;
  assign n42594 = n22611 ^ n21667 ^ 1'b0 ;
  assign n42595 = n34233 | n42594 ;
  assign n42596 = n24998 ^ n9353 ^ n5359 ;
  assign n42597 = n11268 | n42596 ;
  assign n42598 = n29904 ^ n15115 ^ n3557 ;
  assign n42599 = n5608 & ~n34175 ;
  assign n42600 = n42599 ^ n7784 ^ 1'b0 ;
  assign n42601 = n16518 | n19891 ;
  assign n42602 = n42601 ^ n22598 ^ 1'b0 ;
  assign n42603 = x8 | n22665 ;
  assign n42604 = ( ~n8424 & n12449 ) | ( ~n8424 & n40621 ) | ( n12449 & n40621 ) ;
  assign n42605 = n7983 | n42604 ;
  assign n42606 = ~n10465 & n18565 ;
  assign n42607 = n36674 ^ n28816 ^ 1'b0 ;
  assign n42608 = n16396 & ~n20127 ;
  assign n42609 = ~n4079 & n42608 ;
  assign n42610 = n42609 ^ n30597 ^ 1'b0 ;
  assign n42611 = n15875 & ~n42007 ;
  assign n42612 = n21126 ^ n12573 ^ 1'b0 ;
  assign n42613 = n42612 ^ n2440 ^ 1'b0 ;
  assign n42614 = n42611 & ~n42613 ;
  assign n42615 = ~n39429 & n42614 ;
  assign n42616 = n8674 ^ n1369 ^ n675 ;
  assign n42617 = n11857 | n42616 ;
  assign n42618 = n27652 ^ n16713 ^ 1'b0 ;
  assign n42619 = n42618 ^ n42184 ^ 1'b0 ;
  assign n42620 = n12861 & n42619 ;
  assign n42621 = n26502 ^ n9470 ^ 1'b0 ;
  assign n42622 = n26747 & ~n42621 ;
  assign n42623 = n33199 ^ n11298 ^ 1'b0 ;
  assign n42624 = ~n33967 & n42623 ;
  assign n42625 = n42624 ^ n39486 ^ n34132 ;
  assign n42626 = ~n10208 & n21184 ;
  assign n42627 = n42626 ^ n40614 ^ n17902 ;
  assign n42628 = n5881 & n16688 ;
  assign n42629 = n4311 & n42628 ;
  assign n42630 = n42629 ^ n42030 ^ n7794 ;
  assign n42631 = n29984 ^ n5934 ^ 1'b0 ;
  assign n42632 = ~n33393 & n42631 ;
  assign n42633 = n32114 ^ n5687 ^ 1'b0 ;
  assign n42634 = n3789 | n42633 ;
  assign n42635 = n10505 | n42634 ;
  assign n42636 = n35429 ^ n20168 ^ n8810 ;
  assign n42637 = ~n1653 & n42636 ;
  assign n42638 = n17301 & n19702 ;
  assign n42639 = n21633 ^ n20265 ^ n12048 ;
  assign n42640 = n9073 | n33265 ;
  assign n42641 = ( n25056 & ~n30355 ) | ( n25056 & n41420 ) | ( ~n30355 & n41420 ) ;
  assign n42642 = ~n5539 & n16565 ;
  assign n42643 = ( n1190 & n7269 ) | ( n1190 & ~n8198 ) | ( n7269 & ~n8198 ) ;
  assign n42644 = n42643 ^ n14117 ^ 1'b0 ;
  assign n42645 = n16227 | n42644 ;
  assign n42646 = n5882 & ~n24550 ;
  assign n42647 = ( n2845 & n8158 ) | ( n2845 & n39542 ) | ( n8158 & n39542 ) ;
  assign n42648 = n41063 ^ n8363 ^ 1'b0 ;
  assign n42649 = ( n39139 & n42647 ) | ( n39139 & n42648 ) | ( n42647 & n42648 ) ;
  assign n42650 = n6027 ^ n4226 ^ n1244 ;
  assign n42651 = n42650 ^ n9740 ^ n5033 ;
  assign n42652 = n42651 ^ n3934 ^ 1'b0 ;
  assign n42653 = ~n42649 & n42652 ;
  assign n42654 = n8683 ^ n3825 ^ 1'b0 ;
  assign n42655 = n8819 | n24195 ;
  assign n42656 = n42654 & ~n42655 ;
  assign n42657 = ~n4411 & n39864 ;
  assign n42658 = n42657 ^ n33135 ^ n17213 ;
  assign n42659 = n9812 & ~n21349 ;
  assign n42660 = n42659 ^ n1202 ^ 1'b0 ;
  assign n42661 = ( n8572 & n14271 ) | ( n8572 & n42660 ) | ( n14271 & n42660 ) ;
  assign n42662 = n32872 ^ n30836 ^ 1'b0 ;
  assign n42663 = n42662 ^ n42099 ^ n15712 ;
  assign n42664 = n3997 | n5996 ;
  assign n42665 = n15662 ^ n11013 ^ 1'b0 ;
  assign n42666 = ~n4419 & n42665 ;
  assign n42667 = n42666 ^ n24666 ^ 1'b0 ;
  assign n42668 = ~n1899 & n42667 ;
  assign n42669 = n1955 | n23965 ;
  assign n42670 = ~n21195 & n42669 ;
  assign n42671 = ~n42668 & n42670 ;
  assign n42672 = n24412 & ~n25079 ;
  assign n42673 = ~n15950 & n42672 ;
  assign n42674 = ~n41288 & n42673 ;
  assign n42676 = ~n18175 & n19767 ;
  assign n42677 = n42676 ^ n27980 ^ 1'b0 ;
  assign n42675 = ~n1225 & n21864 ;
  assign n42678 = n42677 ^ n42675 ^ 1'b0 ;
  assign n42679 = ~n17806 & n36259 ;
  assign n42680 = n22712 & n42679 ;
  assign n42681 = n42680 ^ n13405 ^ n12591 ;
  assign n42682 = n19728 & n42681 ;
  assign n42683 = n25906 & n42682 ;
  assign n42684 = n27827 ^ n21180 ^ 1'b0 ;
  assign n42686 = n5892 & ~n9423 ;
  assign n42685 = n28696 ^ n16555 ^ 1'b0 ;
  assign n42687 = n42686 ^ n42685 ^ n10298 ;
  assign n42688 = ( ~n6344 & n20644 ) | ( ~n6344 & n42687 ) | ( n20644 & n42687 ) ;
  assign n42689 = n1696 & n15060 ;
  assign n42690 = n14929 & n42689 ;
  assign n42691 = n42690 ^ n13256 ^ n12469 ;
  assign n42692 = n42691 ^ n30725 ^ n16781 ;
  assign n42694 = n4845 & ~n21929 ;
  assign n42695 = ~n7346 & n42694 ;
  assign n42693 = n16859 & ~n41771 ;
  assign n42696 = n42695 ^ n42693 ^ 1'b0 ;
  assign n42697 = n27716 | n42696 ;
  assign n42698 = n1664 & ~n42697 ;
  assign n42699 = n42698 ^ n10993 ^ 1'b0 ;
  assign n42700 = ~n27096 & n30287 ;
  assign n42701 = n4034 & n30479 ;
  assign n42702 = n19939 ^ n13281 ^ n13105 ;
  assign n42703 = ( ~n10755 & n42701 ) | ( ~n10755 & n42702 ) | ( n42701 & n42702 ) ;
  assign n42704 = ~n22741 & n31278 ;
  assign n42705 = n42704 ^ n37846 ^ 1'b0 ;
  assign n42706 = n42703 | n42705 ;
  assign n42707 = n12000 | n34475 ;
  assign n42708 = n40550 & ~n42707 ;
  assign n42709 = n3471 & n16809 ;
  assign n42710 = n42709 ^ n29426 ^ 1'b0 ;
  assign n42711 = n42710 ^ n28019 ^ n23758 ;
  assign n42712 = n20647 ^ n6016 ^ n5060 ;
  assign n42713 = n20707 | n30667 ;
  assign n42714 = n16346 & ~n42713 ;
  assign n42715 = n35212 ^ n14204 ^ 1'b0 ;
  assign n42716 = n25565 ^ n20857 ^ 1'b0 ;
  assign n42717 = n18794 & ~n42716 ;
  assign n42718 = n19075 & ~n37567 ;
  assign n42719 = n42718 ^ n14629 ^ n2030 ;
  assign n42720 = n31267 ^ n2596 ^ 1'b0 ;
  assign n42721 = ( x234 & ~n24537 ) | ( x234 & n42720 ) | ( ~n24537 & n42720 ) ;
  assign n42722 = n35334 ^ n34829 ^ 1'b0 ;
  assign n42723 = ~n25258 & n42722 ;
  assign n42724 = n35620 & n42507 ;
  assign n42725 = n42724 ^ n39823 ^ 1'b0 ;
  assign n42726 = n8307 | n34348 ;
  assign n42727 = ( ~n12953 & n26441 ) | ( ~n12953 & n37119 ) | ( n26441 & n37119 ) ;
  assign n42728 = n42727 ^ n26281 ^ 1'b0 ;
  assign n42729 = n22885 ^ n19369 ^ n13064 ;
  assign n42730 = n42729 ^ n25334 ^ n3510 ;
  assign n42731 = ~n533 & n24904 ;
  assign n42732 = n42731 ^ n21163 ^ 1'b0 ;
  assign n42734 = ~n3080 & n23635 ;
  assign n42733 = n18337 | n20408 ;
  assign n42735 = n42734 ^ n42733 ^ 1'b0 ;
  assign n42736 = n26840 ^ n22131 ^ n14743 ;
  assign n42737 = n6190 & ~n42736 ;
  assign n42738 = ~n490 & n42737 ;
  assign n42739 = n39169 ^ n764 ^ 1'b0 ;
  assign n42740 = ~n23675 & n42739 ;
  assign n42742 = n8824 ^ n4977 ^ 1'b0 ;
  assign n42743 = n684 | n2769 ;
  assign n42744 = n42742 & ~n42743 ;
  assign n42741 = n4026 & n31546 ;
  assign n42745 = n42744 ^ n42741 ^ 1'b0 ;
  assign n42746 = n10601 & ~n37900 ;
  assign n42747 = n28198 ^ n22252 ^ n9189 ;
  assign n42748 = n16185 ^ n9809 ^ 1'b0 ;
  assign n42749 = ~n32821 & n42748 ;
  assign n42750 = n42749 ^ n34097 ^ n20891 ;
  assign n42751 = ( n14137 & n19495 ) | ( n14137 & n21255 ) | ( n19495 & n21255 ) ;
  assign n42752 = ( ~n7233 & n34237 ) | ( ~n7233 & n35038 ) | ( n34237 & n35038 ) ;
  assign n42753 = n10740 & ~n19610 ;
  assign n42754 = n42753 ^ n18926 ^ 1'b0 ;
  assign n42755 = n36656 ^ n29975 ^ 1'b0 ;
  assign n42756 = n1557 | n3308 ;
  assign n42757 = n42756 ^ x73 ^ 1'b0 ;
  assign n42758 = n22462 ^ n18353 ^ 1'b0 ;
  assign n42759 = n42757 & ~n42758 ;
  assign n42760 = n42759 ^ n20695 ^ 1'b0 ;
  assign n42761 = ~n14663 & n42760 ;
  assign n42762 = ~n3475 & n32885 ;
  assign n42763 = n5938 & n42762 ;
  assign n42764 = n32182 | n42763 ;
  assign n42765 = n2164 & ~n42764 ;
  assign n42766 = n19701 ^ n14660 ^ 1'b0 ;
  assign n42767 = ~n26522 & n40084 ;
  assign n42768 = n1936 & ~n3254 ;
  assign n42769 = n8867 & n42768 ;
  assign n42770 = n42769 ^ n292 ^ 1'b0 ;
  assign n42771 = n9675 | n30164 ;
  assign n42772 = n42771 ^ n16911 ^ 1'b0 ;
  assign n42773 = ~n8618 & n13605 ;
  assign n42774 = n41366 ^ n11361 ^ 1'b0 ;
  assign n42775 = ~n5077 & n40799 ;
  assign n42776 = n3283 & n42775 ;
  assign n42777 = n42776 ^ n36626 ^ n19347 ;
  assign n42778 = n36995 | n39642 ;
  assign n42779 = n12360 | n27995 ;
  assign n42780 = n42779 ^ n22233 ^ 1'b0 ;
  assign n42781 = n15182 | n30529 ;
  assign n42782 = n20250 | n42781 ;
  assign n42784 = n4249 ^ n2204 ^ 1'b0 ;
  assign n42785 = n42784 ^ n6745 ^ n2379 ;
  assign n42783 = n27361 ^ n24089 ^ n10165 ;
  assign n42786 = n42785 ^ n42783 ^ 1'b0 ;
  assign n42787 = ( n22165 & ~n24474 ) | ( n22165 & n37821 ) | ( ~n24474 & n37821 ) ;
  assign n42790 = n16172 & n24164 ;
  assign n42788 = n19363 ^ n7784 ^ 1'b0 ;
  assign n42789 = n6196 & ~n42788 ;
  assign n42791 = n42790 ^ n42789 ^ 1'b0 ;
  assign n42792 = n33102 ^ n3813 ^ 1'b0 ;
  assign n42793 = ( ~n16390 & n34949 ) | ( ~n16390 & n42792 ) | ( n34949 & n42792 ) ;
  assign n42794 = n1590 ^ n866 ^ 1'b0 ;
  assign n42795 = ( n13261 & n14764 ) | ( n13261 & n21429 ) | ( n14764 & n21429 ) ;
  assign n42796 = n314 | n42795 ;
  assign n42797 = n25582 & n36470 ;
  assign n42798 = n3401 | n24706 ;
  assign n42799 = n42797 & ~n42798 ;
  assign n42800 = n4670 & ~n11747 ;
  assign n42801 = n42800 ^ n2240 ^ 1'b0 ;
  assign n42802 = n35476 ^ n9441 ^ n536 ;
  assign n42803 = ( n24195 & ~n42801 ) | ( n24195 & n42802 ) | ( ~n42801 & n42802 ) ;
  assign n42804 = n2083 | n26374 ;
  assign n42805 = ( ~n11422 & n33884 ) | ( ~n11422 & n42804 ) | ( n33884 & n42804 ) ;
  assign n42806 = n42803 & n42805 ;
  assign n42807 = n42806 ^ n28983 ^ 1'b0 ;
  assign n42808 = ( n13625 & n19367 ) | ( n13625 & ~n36612 ) | ( n19367 & ~n36612 ) ;
  assign n42809 = ~n3640 & n17639 ;
  assign n42810 = ( n9514 & n26003 ) | ( n9514 & ~n29145 ) | ( n26003 & ~n29145 ) ;
  assign n42811 = ~n26042 & n42810 ;
  assign n42812 = n22538 ^ n22146 ^ n13106 ;
  assign n42813 = ( n11221 & ~n24174 ) | ( n11221 & n42812 ) | ( ~n24174 & n42812 ) ;
  assign n42814 = n8140 | n8830 ;
  assign n42815 = n42814 ^ n9754 ^ 1'b0 ;
  assign n42816 = n38311 ^ x75 ^ 1'b0 ;
  assign n42817 = n4090 | n42816 ;
  assign n42820 = n1933 | n13100 ;
  assign n42821 = ( n21551 & n39161 ) | ( n21551 & n42820 ) | ( n39161 & n42820 ) ;
  assign n42818 = ~n1211 & n32409 ;
  assign n42819 = ~n28813 & n42818 ;
  assign n42822 = n42821 ^ n42819 ^ n8208 ;
  assign n42823 = n25471 ^ n22622 ^ 1'b0 ;
  assign n42824 = n32355 ^ n5432 ^ 1'b0 ;
  assign n42825 = ( n4952 & n5232 ) | ( n4952 & n18218 ) | ( n5232 & n18218 ) ;
  assign n42826 = n10218 | n42825 ;
  assign n42827 = n42824 | n42826 ;
  assign n42828 = n1196 & ~n13497 ;
  assign n42829 = n42828 ^ n27730 ^ 1'b0 ;
  assign n42830 = n23111 ^ n1247 ^ 1'b0 ;
  assign n42831 = n18287 ^ n8309 ^ 1'b0 ;
  assign n42832 = n14901 & ~n42831 ;
  assign n42833 = n37757 ^ n26011 ^ 1'b0 ;
  assign n42834 = n19917 | n42833 ;
  assign n42835 = n32961 ^ n30834 ^ 1'b0 ;
  assign n42836 = ( n19004 & ~n20224 ) | ( n19004 & n42835 ) | ( ~n20224 & n42835 ) ;
  assign n42837 = n29428 ^ n18247 ^ 1'b0 ;
  assign n42838 = n42836 & ~n42837 ;
  assign n42839 = n19640 ^ n3158 ^ 1'b0 ;
  assign n42840 = n4611 | n16425 ;
  assign n42844 = n27290 & ~n38207 ;
  assign n42841 = n5800 ^ n3213 ^ 1'b0 ;
  assign n42842 = n29521 & ~n42841 ;
  assign n42843 = n42842 ^ n28078 ^ 1'b0 ;
  assign n42845 = n42844 ^ n42843 ^ n4617 ;
  assign n42846 = n31038 ^ n21474 ^ 1'b0 ;
  assign n42847 = ~n8025 & n42846 ;
  assign n42848 = n13620 & n42847 ;
  assign n42849 = n42848 ^ n7943 ^ 1'b0 ;
  assign n42850 = n5178 | n11786 ;
  assign n42851 = n25490 & ~n42850 ;
  assign n42852 = n347 & n11670 ;
  assign n42853 = n42851 & n42852 ;
  assign n42854 = n3637 | n38219 ;
  assign n42855 = n7416 ^ n2504 ^ 1'b0 ;
  assign n42856 = n11376 ^ n2290 ^ 1'b0 ;
  assign n42857 = n4928 & ~n9553 ;
  assign n42858 = ~n3037 & n28939 ;
  assign n42859 = ~n7246 & n12907 ;
  assign n42860 = n42858 & n42859 ;
  assign n42861 = n28010 ^ n27380 ^ 1'b0 ;
  assign n42862 = x202 | n42861 ;
  assign n42863 = ~n1689 & n6080 ;
  assign n42864 = ~n335 & n42863 ;
  assign n42865 = ~n3420 & n42864 ;
  assign n42870 = n19104 | n34373 ;
  assign n42866 = n7643 ^ n6669 ^ 1'b0 ;
  assign n42867 = n5266 & ~n42866 ;
  assign n42868 = ( n2360 & n3391 ) | ( n2360 & n42867 ) | ( n3391 & n42867 ) ;
  assign n42869 = ~n16354 & n42868 ;
  assign n42871 = n42870 ^ n42869 ^ 1'b0 ;
  assign n42872 = n30169 | n39432 ;
  assign n42873 = n41477 ^ n31675 ^ 1'b0 ;
  assign n42874 = n27842 ^ n7317 ^ 1'b0 ;
  assign n42875 = ( n10265 & n34109 ) | ( n10265 & n42874 ) | ( n34109 & n42874 ) ;
  assign n42876 = n42875 ^ n22547 ^ n17925 ;
  assign n42877 = ( n12138 & n14665 ) | ( n12138 & ~n41990 ) | ( n14665 & ~n41990 ) ;
  assign n42878 = n42877 ^ n32499 ^ n4995 ;
  assign n42879 = n15509 ^ n639 ^ 1'b0 ;
  assign n42881 = n26233 ^ n17061 ^ n6463 ;
  assign n42880 = n17286 & ~n18801 ;
  assign n42882 = n42881 ^ n42880 ^ n23808 ;
  assign n42883 = n9976 & n42882 ;
  assign n42886 = ~n1332 & n3368 ;
  assign n42884 = n5297 | n20019 ;
  assign n42885 = n42884 ^ n8898 ^ 1'b0 ;
  assign n42887 = n42886 ^ n42885 ^ n13310 ;
  assign n42888 = n42887 ^ n4754 ^ n900 ;
  assign n42889 = n4544 ^ n3796 ^ 1'b0 ;
  assign n42890 = n42889 ^ n34385 ^ n5988 ;
  assign n42891 = n11152 ^ n5579 ^ 1'b0 ;
  assign n42892 = ( n9996 & n42890 ) | ( n9996 & n42891 ) | ( n42890 & n42891 ) ;
  assign n42893 = n16155 & ~n26307 ;
  assign n42894 = n42893 ^ n27579 ^ 1'b0 ;
  assign n42895 = ( n13039 & n13051 ) | ( n13039 & n13267 ) | ( n13051 & n13267 ) ;
  assign n42896 = n27284 ^ n11397 ^ 1'b0 ;
  assign n42897 = n4537 & n42896 ;
  assign n42899 = ~n18297 & n31977 ;
  assign n42900 = n5107 & n42899 ;
  assign n42898 = ~n3877 & n9108 ;
  assign n42901 = n42900 ^ n42898 ^ 1'b0 ;
  assign n42902 = n8117 & ~n8129 ;
  assign n42903 = n3953 & n31414 ;
  assign n42904 = n42903 ^ n25660 ^ 1'b0 ;
  assign n42905 = n6594 & ~n17771 ;
  assign n42906 = n42905 ^ n10629 ^ 1'b0 ;
  assign n42907 = ( ~n5471 & n42904 ) | ( ~n5471 & n42906 ) | ( n42904 & n42906 ) ;
  assign n42908 = n6043 | n18007 ;
  assign n42909 = n42908 ^ n5717 ^ 1'b0 ;
  assign n42910 = ~n15175 & n42909 ;
  assign n42911 = ~n40446 & n42910 ;
  assign n42912 = n20049 & ~n42911 ;
  assign n42913 = ( n11446 & n37504 ) | ( n11446 & ~n37685 ) | ( n37504 & ~n37685 ) ;
  assign n42914 = n6699 | n10821 ;
  assign n42915 = n20295 & ~n42914 ;
  assign n42916 = n318 & ~n42915 ;
  assign n42917 = n42916 ^ n39426 ^ 1'b0 ;
  assign n42918 = ~n14508 & n34405 ;
  assign n42919 = n42918 ^ n11061 ^ 1'b0 ;
  assign n42920 = n17792 & n42919 ;
  assign n42921 = ~n6050 & n42920 ;
  assign n42922 = n42921 ^ n30071 ^ 1'b0 ;
  assign n42923 = n41656 ^ n4444 ^ 1'b0 ;
  assign n42924 = n27883 ^ n7131 ^ 1'b0 ;
  assign n42925 = ~n13495 & n42924 ;
  assign n42927 = n7946 ^ n6882 ^ 1'b0 ;
  assign n42926 = n1380 | n19195 ;
  assign n42928 = n42927 ^ n42926 ^ 1'b0 ;
  assign n42929 = n7961 & n38056 ;
  assign n42930 = n22967 ^ n18365 ^ n17817 ;
  assign n42931 = ( n8386 & ~n10789 ) | ( n8386 & n42930 ) | ( ~n10789 & n42930 ) ;
  assign n42932 = n642 & ~n34730 ;
  assign n42933 = n24696 ^ n19679 ^ 1'b0 ;
  assign n42934 = ~n11000 & n42933 ;
  assign n42935 = n42934 ^ n23211 ^ 1'b0 ;
  assign n42936 = n25086 ^ n10189 ^ n2344 ;
  assign n42937 = n16388 & ~n42936 ;
  assign n42938 = n42937 ^ n9089 ^ 1'b0 ;
  assign n42939 = ( n19190 & ~n30843 ) | ( n19190 & n41832 ) | ( ~n30843 & n41832 ) ;
  assign n42940 = ( n42935 & ~n42938 ) | ( n42935 & n42939 ) | ( ~n42938 & n42939 ) ;
  assign n42941 = n21650 ^ n16726 ^ 1'b0 ;
  assign n42942 = ~n3758 & n21592 ;
  assign n42943 = ~n10031 & n24858 ;
  assign n42944 = n42943 ^ n20467 ^ 1'b0 ;
  assign n42945 = ( n20548 & n27801 ) | ( n20548 & ~n42944 ) | ( n27801 & ~n42944 ) ;
  assign n42946 = n27183 ^ n8805 ^ n8715 ;
  assign n42947 = n3188 & ~n42946 ;
  assign n42948 = n30523 ^ n20697 ^ n14901 ;
  assign n42949 = ~n30164 & n34290 ;
  assign n42950 = n42949 ^ n11977 ^ 1'b0 ;
  assign n42951 = n19037 & n42480 ;
  assign n42952 = ~n32796 & n42951 ;
  assign n42953 = n38859 ^ n35626 ^ 1'b0 ;
  assign n42954 = n21875 | n42953 ;
  assign n42956 = n22854 ^ n12788 ^ 1'b0 ;
  assign n42957 = n28592 & ~n42956 ;
  assign n42955 = n33993 & n35613 ;
  assign n42958 = n42957 ^ n42955 ^ 1'b0 ;
  assign n42963 = n3830 | n6320 ;
  assign n42959 = n11779 & n19402 ;
  assign n42960 = ( n1847 & n11631 ) | ( n1847 & ~n42959 ) | ( n11631 & ~n42959 ) ;
  assign n42961 = ~n39488 & n42960 ;
  assign n42962 = n25894 & n42961 ;
  assign n42964 = n42963 ^ n42962 ^ n19614 ;
  assign n42965 = n5901 ^ n5520 ^ 1'b0 ;
  assign n42966 = n42964 | n42965 ;
  assign n42967 = n13162 & ~n20941 ;
  assign n42968 = n39297 & n42967 ;
  assign n42969 = n18143 & ~n42968 ;
  assign n42970 = n42969 ^ n23484 ^ 1'b0 ;
  assign n42971 = n27725 ^ n13298 ^ n10099 ;
  assign n42972 = n29298 ^ n26827 ^ 1'b0 ;
  assign n42973 = ( n1076 & ~n3371 ) | ( n1076 & n42972 ) | ( ~n3371 & n42972 ) ;
  assign n42974 = n37205 ^ n8790 ^ n4094 ;
  assign n42975 = ( n42971 & ~n42973 ) | ( n42971 & n42974 ) | ( ~n42973 & n42974 ) ;
  assign n42976 = n12457 | n26394 ;
  assign n42977 = n15462 & ~n37646 ;
  assign n42978 = n42977 ^ n37988 ^ 1'b0 ;
  assign n42979 = n14400 & n20671 ;
  assign n42980 = n42979 ^ n5141 ^ 1'b0 ;
  assign n42981 = ~n18895 & n25037 ;
  assign n42982 = ~n39974 & n42981 ;
  assign n42983 = n16977 ^ n16350 ^ n13851 ;
  assign n42984 = n12582 & n35507 ;
  assign n42985 = ~n36498 & n42984 ;
  assign n42986 = ( n28611 & ~n42983 ) | ( n28611 & n42985 ) | ( ~n42983 & n42985 ) ;
  assign n42987 = ~n20335 & n42986 ;
  assign n42988 = n29790 ^ n16461 ^ 1'b0 ;
  assign n42989 = n27783 ^ n4191 ^ 1'b0 ;
  assign n42990 = n3796 | n22530 ;
  assign n42991 = ~n3358 & n35313 ;
  assign n42992 = n42991 ^ n12898 ^ 1'b0 ;
  assign n42993 = n42992 ^ n29094 ^ 1'b0 ;
  assign n42994 = ~n2507 & n42993 ;
  assign n42995 = n17696 ^ n8893 ^ 1'b0 ;
  assign n42996 = n36339 ^ n17208 ^ 1'b0 ;
  assign n42997 = n6382 & ~n10753 ;
  assign n42998 = n18488 & n42997 ;
  assign n42999 = n42998 ^ n17863 ^ n5162 ;
  assign n43000 = ~n8393 & n14533 ;
  assign n43001 = n29965 & ~n43000 ;
  assign n43002 = n43001 ^ n33584 ^ n10383 ;
  assign n43003 = ( ~n354 & n24813 ) | ( ~n354 & n40759 ) | ( n24813 & n40759 ) ;
  assign n43004 = ( n20455 & ~n41066 ) | ( n20455 & n43003 ) | ( ~n41066 & n43003 ) ;
  assign n43005 = n1702 & ~n16767 ;
  assign n43006 = n10395 & n43005 ;
  assign n43007 = n43006 ^ n37293 ^ 1'b0 ;
  assign n43008 = n2703 | n40283 ;
  assign n43009 = n43008 ^ n37699 ^ 1'b0 ;
  assign n43010 = ( n8456 & ~n11398 ) | ( n8456 & n41871 ) | ( ~n11398 & n41871 ) ;
  assign n43011 = n4824 & n8286 ;
  assign n43012 = n11325 & ~n43011 ;
  assign n43013 = n43010 & n43012 ;
  assign n43014 = ~n17263 & n23965 ;
  assign n43015 = n39958 & n43014 ;
  assign n43016 = n12046 | n43015 ;
  assign n43020 = n7586 & ~n8433 ;
  assign n43017 = n8302 ^ n7322 ^ 1'b0 ;
  assign n43018 = ~n9512 & n43017 ;
  assign n43019 = n12554 | n43018 ;
  assign n43021 = n43020 ^ n43019 ^ n4413 ;
  assign n43022 = ~n10039 & n43021 ;
  assign n43023 = n18131 & ~n43022 ;
  assign n43024 = n2136 & ~n4361 ;
  assign n43025 = n43024 ^ n5044 ^ 1'b0 ;
  assign n43026 = n43025 ^ n37722 ^ n28403 ;
  assign n43027 = n16890 & n18250 ;
  assign n43028 = n43027 ^ n14784 ^ 1'b0 ;
  assign n43029 = ~n31826 & n43028 ;
  assign n43030 = n10402 | n11449 ;
  assign n43031 = n24820 & ~n29738 ;
  assign n43032 = n43031 ^ n16773 ^ 1'b0 ;
  assign n43033 = ~n28577 & n43032 ;
  assign n43034 = n6967 & n43033 ;
  assign n43035 = n1232 & n18597 ;
  assign n43036 = n43035 ^ n31855 ^ 1'b0 ;
  assign n43037 = n1468 & ~n43036 ;
  assign n43038 = n26061 | n32815 ;
  assign n43039 = n10031 | n43038 ;
  assign n43040 = n6735 ^ n6511 ^ 1'b0 ;
  assign n43041 = n684 & n43040 ;
  assign n43042 = n29126 & n43041 ;
  assign n43043 = ~n20788 & n42881 ;
  assign n43044 = n43043 ^ n16083 ^ 1'b0 ;
  assign n43045 = n3136 | n4254 ;
  assign n43046 = n43045 ^ n26247 ^ n12491 ;
  assign n43047 = n30061 | n36135 ;
  assign n43048 = ~n5795 & n16021 ;
  assign n43049 = n43048 ^ n9033 ^ 1'b0 ;
  assign n43050 = n12470 & n35106 ;
  assign n43051 = n13765 & n43050 ;
  assign n43052 = n43051 ^ n5694 ^ n3315 ;
  assign n43053 = n32942 & n43052 ;
  assign n43054 = ( n12265 & n31759 ) | ( n12265 & n37761 ) | ( n31759 & n37761 ) ;
  assign n43055 = n30061 ^ n25079 ^ 1'b0 ;
  assign n43056 = n20255 & n43055 ;
  assign n43057 = n13069 | n40112 ;
  assign n43058 = n43057 ^ n38031 ^ 1'b0 ;
  assign n43059 = n43058 ^ n33807 ^ n2665 ;
  assign n43060 = n13691 & ~n39255 ;
  assign n43061 = ~n8025 & n43060 ;
  assign n43062 = n15204 & ~n15431 ;
  assign n43063 = ~n10892 & n43062 ;
  assign n43064 = n30958 ^ n21923 ^ 1'b0 ;
  assign n43065 = n8058 ^ n6467 ^ n2798 ;
  assign n43066 = ~n5579 & n6981 ;
  assign n43067 = n43066 ^ n37625 ^ 1'b0 ;
  assign n43068 = ( n24566 & n43065 ) | ( n24566 & n43067 ) | ( n43065 & n43067 ) ;
  assign n43069 = ( n1752 & ~n4435 ) | ( n1752 & n9445 ) | ( ~n4435 & n9445 ) ;
  assign n43070 = n43069 ^ n21856 ^ n20290 ;
  assign n43071 = n8757 & n21382 ;
  assign n43072 = ~n35469 & n43071 ;
  assign n43073 = n3515 ^ n1944 ^ 1'b0 ;
  assign n43074 = ~n9670 & n18721 ;
  assign n43075 = n16796 & n20672 ;
  assign n43076 = ~n10332 & n43075 ;
  assign n43077 = ( n10932 & ~n23282 ) | ( n10932 & n30695 ) | ( ~n23282 & n30695 ) ;
  assign n43078 = n20871 | n43077 ;
  assign n43079 = n11371 ^ n4858 ^ 1'b0 ;
  assign n43080 = n10010 & ~n28906 ;
  assign n43081 = n43079 & ~n43080 ;
  assign n43082 = x214 & n731 ;
  assign n43083 = ~x214 & n43082 ;
  assign n43084 = x98 & x214 ;
  assign n43085 = n43083 & n43084 ;
  assign n43086 = n43085 ^ n1090 ^ 1'b0 ;
  assign n43087 = n11286 ^ n10310 ^ 1'b0 ;
  assign n43088 = n43086 & ~n43087 ;
  assign n43089 = ( n17750 & ~n21949 ) | ( n17750 & n43088 ) | ( ~n21949 & n43088 ) ;
  assign n43090 = n31158 & ~n32927 ;
  assign n43091 = n43090 ^ n7434 ^ 1'b0 ;
  assign n43092 = n15703 ^ n1394 ^ 1'b0 ;
  assign n43093 = n10346 ^ n1848 ^ 1'b0 ;
  assign n43094 = n9110 ^ n1935 ^ 1'b0 ;
  assign n43095 = n7256 & ~n43094 ;
  assign n43096 = n43095 ^ n13004 ^ 1'b0 ;
  assign n43097 = n3447 & n43096 ;
  assign n43098 = n8179 ^ n6361 ^ 1'b0 ;
  assign n43099 = n16111 ^ n12870 ^ 1'b0 ;
  assign n43100 = n13064 | n43099 ;
  assign n43101 = ( n24622 & n43098 ) | ( n24622 & ~n43100 ) | ( n43098 & ~n43100 ) ;
  assign n43102 = n27247 ^ n26668 ^ n18785 ;
  assign n43103 = ~n18487 & n35891 ;
  assign n43104 = ( n3939 & n43102 ) | ( n3939 & ~n43103 ) | ( n43102 & ~n43103 ) ;
  assign n43105 = n12091 ^ n5187 ^ 1'b0 ;
  assign n43106 = ~n16573 & n43105 ;
  assign n43107 = ~n10533 & n14077 ;
  assign n43108 = n43107 ^ n8331 ^ 1'b0 ;
  assign n43109 = n43106 & ~n43108 ;
  assign n43110 = ~n9599 & n43109 ;
  assign n43111 = n21683 & n43110 ;
  assign n43112 = n34604 ^ n12826 ^ n2009 ;
  assign n43113 = n28756 ^ n11749 ^ 1'b0 ;
  assign n43114 = ~n41503 & n43113 ;
  assign n43115 = n4668 ^ x166 ^ 1'b0 ;
  assign n43116 = n19932 | n43115 ;
  assign n43117 = n43116 ^ n18619 ^ n16961 ;
  assign n43118 = n13004 & n43117 ;
  assign n43119 = n43118 ^ n4770 ^ 1'b0 ;
  assign n43120 = n5296 ^ n4672 ^ 1'b0 ;
  assign n43121 = n2390 & ~n12579 ;
  assign n43122 = n43121 ^ n326 ^ 1'b0 ;
  assign n43123 = n39087 ^ n16008 ^ 1'b0 ;
  assign n43124 = x26 & n43123 ;
  assign n43125 = n43124 ^ n17656 ^ 1'b0 ;
  assign n43126 = n16394 | n31192 ;
  assign n43127 = n30824 | n40395 ;
  assign n43128 = n43126 & ~n43127 ;
  assign n43129 = ( n28227 & ~n29681 ) | ( n28227 & n43128 ) | ( ~n29681 & n43128 ) ;
  assign n43130 = n15575 ^ n14212 ^ 1'b0 ;
  assign n43131 = ( n11493 & n26075 ) | ( n11493 & n43130 ) | ( n26075 & n43130 ) ;
  assign n43132 = n43131 ^ n38472 ^ 1'b0 ;
  assign n43133 = n42795 ^ n28185 ^ n17059 ;
  assign n43134 = n16109 & ~n22098 ;
  assign n43135 = n43133 & n43134 ;
  assign n43136 = n24424 ^ n8357 ^ 1'b0 ;
  assign n43137 = ~n7373 & n43136 ;
  assign n43138 = ~n1943 & n43137 ;
  assign n43139 = n22302 & ~n32551 ;
  assign n43140 = n43139 ^ n21318 ^ 1'b0 ;
  assign n43141 = n41382 ^ n33552 ^ 1'b0 ;
  assign n43142 = n5491 & n19523 ;
  assign n43143 = n11483 | n43142 ;
  assign n43144 = ( n10298 & n19521 ) | ( n10298 & ~n43143 ) | ( n19521 & ~n43143 ) ;
  assign n43145 = n40191 ^ n9461 ^ 1'b0 ;
  assign n43146 = ~n19109 & n19851 ;
  assign n43147 = ~n14040 & n43146 ;
  assign n43148 = n4569 & ~n22961 ;
  assign n43149 = n28874 ^ n10619 ^ 1'b0 ;
  assign n43150 = n4422 ^ n3428 ^ 1'b0 ;
  assign n43151 = n13126 & n28274 ;
  assign n43152 = ~n8028 & n43151 ;
  assign n43153 = n26091 ^ n901 ^ 1'b0 ;
  assign n43154 = n43153 ^ n25915 ^ n14634 ;
  assign n43155 = n29945 ^ n15114 ^ n481 ;
  assign n43156 = n20122 & ~n21553 ;
  assign n43157 = n26244 & n43156 ;
  assign n43158 = n23866 ^ n2841 ^ 1'b0 ;
  assign n43159 = n2440 & n43158 ;
  assign n43160 = n26835 & n38493 ;
  assign n43161 = n43160 ^ n16606 ^ 1'b0 ;
  assign n43162 = n13717 & n35866 ;
  assign n43163 = ~n7876 & n43162 ;
  assign n43164 = n43163 ^ n20821 ^ 1'b0 ;
  assign n43165 = ~n29000 & n29508 ;
  assign n43166 = n15218 & n43165 ;
  assign n43167 = n34206 ^ n29826 ^ n13637 ;
  assign n43168 = n7145 & ~n43167 ;
  assign n43169 = ~n19973 & n43168 ;
  assign n43170 = n7553 & ~n13335 ;
  assign n43171 = n43170 ^ n25433 ^ n7004 ;
  assign n43172 = ( x240 & n12165 ) | ( x240 & ~n18594 ) | ( n12165 & ~n18594 ) ;
  assign n43173 = n9189 & n10506 ;
  assign n43174 = n43173 ^ n22398 ^ 1'b0 ;
  assign n43175 = n43174 ^ n43095 ^ n42904 ;
  assign n43176 = ( n13453 & n19606 ) | ( n13453 & n39687 ) | ( n19606 & n39687 ) ;
  assign n43177 = n3095 | n12267 ;
  assign n43178 = n2331 | n43177 ;
  assign n43179 = n14137 & n27330 ;
  assign n43180 = ~n43178 & n43179 ;
  assign n43181 = n7116 & n16362 ;
  assign n43182 = n19356 ^ n4020 ^ 1'b0 ;
  assign n43183 = ~n2196 & n6804 ;
  assign n43185 = n9878 & ~n11115 ;
  assign n43184 = ~n15226 & n25179 ;
  assign n43186 = n43185 ^ n43184 ^ 1'b0 ;
  assign n43187 = ( n4351 & n13659 ) | ( n4351 & ~n27281 ) | ( n13659 & ~n27281 ) ;
  assign n43188 = ( n10750 & n12861 ) | ( n10750 & n25660 ) | ( n12861 & n25660 ) ;
  assign n43189 = n8773 & ~n31909 ;
  assign n43190 = n43188 & n43189 ;
  assign n43191 = ( n4173 & n13276 ) | ( n4173 & ~n27302 ) | ( n13276 & ~n27302 ) ;
  assign n43192 = n23773 & ~n43191 ;
  assign n43193 = ~n8991 & n43192 ;
  assign n43194 = ~n2356 & n20075 ;
  assign n43195 = n43193 & n43194 ;
  assign n43196 = n14053 ^ n5399 ^ 1'b0 ;
  assign n43197 = n8941 ^ n5416 ^ 1'b0 ;
  assign n43198 = n43196 & n43197 ;
  assign n43199 = n9853 ^ n4228 ^ n3222 ;
  assign n43200 = n11135 | n43199 ;
  assign n43201 = ~n23653 & n43200 ;
  assign n43202 = n43201 ^ n15228 ^ 1'b0 ;
  assign n43203 = ~n6698 & n13986 ;
  assign n43204 = ~n43202 & n43203 ;
  assign n43205 = n43204 ^ n4812 ^ 1'b0 ;
  assign n43206 = n1825 | n43205 ;
  assign n43209 = n12113 ^ n1289 ^ 1'b0 ;
  assign n43207 = n9734 ^ n8709 ^ x147 ;
  assign n43208 = n21195 | n43207 ;
  assign n43210 = n43209 ^ n43208 ^ 1'b0 ;
  assign n43211 = n20328 & ~n43210 ;
  assign n43212 = n1082 & n21260 ;
  assign n43213 = n43212 ^ n30633 ^ 1'b0 ;
  assign n43214 = n42072 | n43213 ;
  assign n43215 = n31769 ^ n9880 ^ 1'b0 ;
  assign n43216 = n21291 & n43215 ;
  assign n43217 = n43216 ^ n27652 ^ 1'b0 ;
  assign n43218 = x83 & ~n21040 ;
  assign n43219 = ~n6728 & n43218 ;
  assign n43220 = n43219 ^ n39629 ^ 1'b0 ;
  assign n43221 = ( n21857 & n21978 ) | ( n21857 & n43220 ) | ( n21978 & n43220 ) ;
  assign n43222 = n26829 ^ n3578 ^ 1'b0 ;
  assign n43223 = n41992 & n43222 ;
  assign n43224 = ( n29534 & n29839 ) | ( n29534 & n43223 ) | ( n29839 & n43223 ) ;
  assign n43225 = n11629 ^ n2826 ^ n1781 ;
  assign n43226 = ~n569 & n8960 ;
  assign n43227 = ( n14276 & ~n43225 ) | ( n14276 & n43226 ) | ( ~n43225 & n43226 ) ;
  assign n43228 = n4083 & n15588 ;
  assign n43229 = n43228 ^ n39211 ^ 1'b0 ;
  assign n43230 = ( n3034 & n22929 ) | ( n3034 & n43229 ) | ( n22929 & n43229 ) ;
  assign n43233 = n2577 | n23844 ;
  assign n43234 = n8941 | n43233 ;
  assign n43235 = n4098 & n43234 ;
  assign n43236 = n43235 ^ n1828 ^ 1'b0 ;
  assign n43231 = n7319 ^ n287 ^ 1'b0 ;
  assign n43232 = x39 & ~n43231 ;
  assign n43237 = n43236 ^ n43232 ^ 1'b0 ;
  assign n43238 = n9521 & n37947 ;
  assign n43239 = n43238 ^ n11535 ^ 1'b0 ;
  assign n43240 = n34207 ^ n22857 ^ n2151 ;
  assign n43241 = n10436 ^ n9818 ^ 1'b0 ;
  assign n43242 = n43241 ^ n34368 ^ 1'b0 ;
  assign n43243 = ( ~n1138 & n30725 ) | ( ~n1138 & n43242 ) | ( n30725 & n43242 ) ;
  assign n43244 = n6917 & ~n32002 ;
  assign n43245 = ~n43243 & n43244 ;
  assign n43246 = ( n11445 & n18568 ) | ( n11445 & n43245 ) | ( n18568 & n43245 ) ;
  assign n43247 = ~x53 & n25340 ;
  assign n43248 = n30865 ^ n17991 ^ 1'b0 ;
  assign n43249 = ~n43247 & n43248 ;
  assign n43250 = n43249 ^ n41412 ^ 1'b0 ;
  assign n43251 = ( n2073 & ~n3387 ) | ( n2073 & n8294 ) | ( ~n3387 & n8294 ) ;
  assign n43252 = ~n3172 & n7939 ;
  assign n43253 = ~n31852 & n43252 ;
  assign n43254 = n43253 ^ n4602 ^ 1'b0 ;
  assign n43255 = n25901 & ~n43254 ;
  assign n43256 = n654 & ~n21089 ;
  assign n43257 = ~n12413 & n43256 ;
  assign n43258 = n4330 & ~n38293 ;
  assign n43259 = n15549 & n36199 ;
  assign n43260 = n32962 ^ n3529 ^ 1'b0 ;
  assign n43261 = ~n4581 & n13032 ;
  assign n43262 = ~n10358 & n43261 ;
  assign n43263 = ( n10585 & n28403 ) | ( n10585 & ~n43262 ) | ( n28403 & ~n43262 ) ;
  assign n43264 = n14548 ^ n3297 ^ n1393 ;
  assign n43265 = ( ~n16877 & n36824 ) | ( ~n16877 & n43264 ) | ( n36824 & n43264 ) ;
  assign n43266 = ~n16402 & n23777 ;
  assign n43267 = n43266 ^ n35040 ^ 1'b0 ;
  assign n43268 = n4223 & n15795 ;
  assign n43269 = n43267 & n43268 ;
  assign n43270 = n15494 & n34032 ;
  assign n43271 = n17116 ^ n15380 ^ 1'b0 ;
  assign n43272 = n43270 | n43271 ;
  assign n43273 = n11562 & ~n43272 ;
  assign n43274 = ~n19766 & n43273 ;
  assign n43275 = n25713 ^ n13007 ^ 1'b0 ;
  assign n43277 = ~n13762 & n17473 ;
  assign n43278 = n28547 ^ n25909 ^ 1'b0 ;
  assign n43279 = n43277 & ~n43278 ;
  assign n43276 = n9803 | n18866 ;
  assign n43280 = n43279 ^ n43276 ^ 1'b0 ;
  assign n43281 = n9212 ^ n3532 ^ 1'b0 ;
  assign n43282 = ( n9628 & ~n19709 ) | ( n9628 & n43281 ) | ( ~n19709 & n43281 ) ;
  assign n43283 = n6406 ^ n4013 ^ 1'b0 ;
  assign n43284 = ( n658 & n41260 ) | ( n658 & n43283 ) | ( n41260 & n43283 ) ;
  assign n43285 = ( n6610 & n15924 ) | ( n6610 & n36572 ) | ( n15924 & n36572 ) ;
  assign n43286 = ( ~x145 & n6758 ) | ( ~x145 & n11517 ) | ( n6758 & n11517 ) ;
  assign n43287 = n38107 | n43286 ;
  assign n43288 = n493 & ~n43287 ;
  assign n43289 = n43288 ^ n3646 ^ 1'b0 ;
  assign n43290 = n15240 & n43289 ;
  assign n43291 = n32000 ^ n13320 ^ n12676 ;
  assign n43292 = n19727 ^ n288 ^ 1'b0 ;
  assign n43295 = n20360 ^ n20021 ^ 1'b0 ;
  assign n43296 = n7100 & ~n43295 ;
  assign n43297 = n43296 ^ n23358 ^ 1'b0 ;
  assign n43293 = n38239 ^ n18675 ^ n4657 ;
  assign n43294 = n30278 & n43293 ;
  assign n43298 = n43297 ^ n43294 ^ 1'b0 ;
  assign n43299 = n43011 ^ n5638 ^ 1'b0 ;
  assign n43300 = n28757 & n43299 ;
  assign n43301 = n20049 ^ n11748 ^ 1'b0 ;
  assign n43302 = ~n1700 & n43301 ;
  assign n43303 = n43302 ^ n36708 ^ 1'b0 ;
  assign n43304 = n5495 & n43303 ;
  assign n43305 = n43304 ^ x46 ^ 1'b0 ;
  assign n43306 = ~n5925 & n43305 ;
  assign n43307 = n36674 ^ n34394 ^ n8742 ;
  assign n43308 = n5081 | n8969 ;
  assign n43309 = n43308 ^ n2411 ^ 1'b0 ;
  assign n43310 = n1510 & ~n10142 ;
  assign n43311 = n43309 & n43310 ;
  assign n43312 = n35669 ^ n22209 ^ 1'b0 ;
  assign n43313 = n633 | n43312 ;
  assign n43314 = n2760 & ~n18051 ;
  assign n43315 = ( n32498 & ~n36012 ) | ( n32498 & n43314 ) | ( ~n36012 & n43314 ) ;
  assign n43316 = n24256 ^ n16673 ^ n5857 ;
  assign n43317 = n21178 ^ n10674 ^ 1'b0 ;
  assign n43318 = ~n5484 & n43317 ;
  assign n43319 = ~n1979 & n43318 ;
  assign n43321 = ~n12677 & n31340 ;
  assign n43320 = ~n9927 & n12870 ;
  assign n43322 = n43321 ^ n43320 ^ 1'b0 ;
  assign n43323 = n25169 ^ n2225 ^ 1'b0 ;
  assign n43324 = ~n923 & n6606 ;
  assign n43325 = n9996 & n43324 ;
  assign n43326 = n23279 ^ n14604 ^ 1'b0 ;
  assign n43327 = n3283 ^ n294 ^ 1'b0 ;
  assign n43328 = n19395 | n43327 ;
  assign n43329 = ~n17119 & n23907 ;
  assign n43330 = ( ~n1382 & n35154 ) | ( ~n1382 & n43329 ) | ( n35154 & n43329 ) ;
  assign n43331 = ~n7805 & n15966 ;
  assign n43332 = n945 & n5755 ;
  assign n43333 = ( n8149 & n43331 ) | ( n8149 & ~n43332 ) | ( n43331 & ~n43332 ) ;
  assign n43334 = n6315 & n22609 ;
  assign n43335 = n43334 ^ n24723 ^ 1'b0 ;
  assign n43336 = n9681 & n16181 ;
  assign n43337 = n290 & n43336 ;
  assign n43338 = ( ~n1936 & n20574 ) | ( ~n1936 & n26120 ) | ( n20574 & n26120 ) ;
  assign n43339 = n43338 ^ n7119 ^ x218 ;
  assign n43340 = n24324 ^ n6759 ^ 1'b0 ;
  assign n43341 = n43339 & n43340 ;
  assign n43342 = n43341 ^ n33079 ^ 1'b0 ;
  assign n43343 = n31133 ^ n26232 ^ n5426 ;
  assign n43344 = n43343 ^ n10518 ^ 1'b0 ;
  assign n43345 = ~n32639 & n43344 ;
  assign n43346 = n20433 ^ n2192 ^ 1'b0 ;
  assign n43347 = n13625 & n43346 ;
  assign n43348 = n38143 ^ n27752 ^ 1'b0 ;
  assign n43349 = n14469 & n43348 ;
  assign n43350 = n30208 ^ n7780 ^ n2004 ;
  assign n43351 = ~n845 & n40164 ;
  assign n43352 = n43351 ^ n21385 ^ 1'b0 ;
  assign n43353 = n43352 ^ n22962 ^ n702 ;
  assign n43354 = ~n13877 & n28498 ;
  assign n43355 = n43354 ^ n16824 ^ n7113 ;
  assign n43356 = n10470 & ~n43355 ;
  assign n43357 = n43356 ^ n30787 ^ 1'b0 ;
  assign n43358 = n26686 ^ n10003 ^ 1'b0 ;
  assign n43359 = n40736 & n43358 ;
  assign n43360 = n30382 | n43359 ;
  assign n43361 = n4912 & n10487 ;
  assign n43362 = ( n2671 & n6192 ) | ( n2671 & ~n34495 ) | ( n6192 & ~n34495 ) ;
  assign n43363 = ~n19595 & n43362 ;
  assign n43364 = ~n39598 & n43363 ;
  assign n43365 = n2205 | n9422 ;
  assign n43366 = n43365 ^ n4243 ^ 1'b0 ;
  assign n43373 = n13448 & ~n25758 ;
  assign n43374 = n43373 ^ n22590 ^ n16005 ;
  assign n43368 = ~n3947 & n8751 ;
  assign n43369 = ~n26587 & n43368 ;
  assign n43370 = n43369 ^ n25335 ^ 1'b0 ;
  assign n43371 = n43370 ^ n20616 ^ n15307 ;
  assign n43367 = n1847 & ~n29657 ;
  assign n43372 = n43371 ^ n43367 ^ 1'b0 ;
  assign n43375 = n43374 ^ n43372 ^ n933 ;
  assign n43376 = n15039 ^ n4340 ^ 1'b0 ;
  assign n43377 = ~n17765 & n43376 ;
  assign n43378 = n43377 ^ n18675 ^ n5292 ;
  assign n43379 = n30458 & ~n31924 ;
  assign n43380 = n28395 & n43379 ;
  assign n43381 = n43380 ^ n11202 ^ 1'b0 ;
  assign n43382 = n21345 & n24250 ;
  assign n43383 = ~n37919 & n43382 ;
  assign n43386 = n19701 ^ n9077 ^ 1'b0 ;
  assign n43387 = n7098 | n43386 ;
  assign n43384 = n23488 & n40830 ;
  assign n43385 = n7464 & n43384 ;
  assign n43388 = n43387 ^ n43385 ^ 1'b0 ;
  assign n43389 = n7812 & n30329 ;
  assign n43390 = n43389 ^ n33070 ^ 1'b0 ;
  assign n43391 = n18182 & n43390 ;
  assign n43392 = n18273 | n22967 ;
  assign n43393 = n36341 ^ n13994 ^ 1'b0 ;
  assign n43394 = n25442 ^ n7880 ^ 1'b0 ;
  assign n43395 = ~n10851 & n43394 ;
  assign n43396 = ( n19785 & n27359 ) | ( n19785 & ~n43395 ) | ( n27359 & ~n43395 ) ;
  assign n43397 = n13263 & ~n43396 ;
  assign n43398 = n8559 & ~n43397 ;
  assign n43399 = n11582 & n43398 ;
  assign n43400 = n24285 ^ n22134 ^ n14747 ;
  assign n43401 = n38531 ^ n7946 ^ n5160 ;
  assign n43402 = n33810 ^ n8276 ^ 1'b0 ;
  assign n43403 = n16227 ^ n15807 ^ 1'b0 ;
  assign n43404 = n610 & ~n24863 ;
  assign n43405 = ( n2567 & n7508 ) | ( n2567 & ~n12971 ) | ( n7508 & ~n12971 ) ;
  assign n43406 = n2954 ^ n1871 ^ 1'b0 ;
  assign n43407 = n994 & ~n43406 ;
  assign n43408 = ~n11082 & n43407 ;
  assign n43409 = n43405 & n43408 ;
  assign n43410 = n32793 | n43409 ;
  assign n43411 = n13982 & ~n43410 ;
  assign n43412 = n3207 & n9612 ;
  assign n43413 = n43412 ^ n20163 ^ 1'b0 ;
  assign n43414 = n4310 & n43413 ;
  assign n43415 = n43414 ^ n9041 ^ 1'b0 ;
  assign n43416 = ( n4616 & n26861 ) | ( n4616 & n38531 ) | ( n26861 & n38531 ) ;
  assign n43417 = n4350 ^ n639 ^ 1'b0 ;
  assign n43418 = ( n7242 & n25329 ) | ( n7242 & ~n33546 ) | ( n25329 & ~n33546 ) ;
  assign n43419 = n38641 & ~n42000 ;
  assign n43420 = n29047 ^ n4055 ^ 1'b0 ;
  assign n43421 = n9772 & n43420 ;
  assign n43422 = ~n24454 & n43421 ;
  assign n43423 = n43422 ^ n21139 ^ n3624 ;
  assign n43424 = n29513 ^ n15927 ^ 1'b0 ;
  assign n43425 = n16267 ^ n8420 ^ n5062 ;
  assign n43426 = n13511 ^ x220 ^ 1'b0 ;
  assign n43427 = ~n36131 & n43426 ;
  assign n43428 = n43427 ^ x108 ^ 1'b0 ;
  assign n43429 = ~n21149 & n37807 ;
  assign n43430 = ~n27743 & n43429 ;
  assign n43431 = n43430 ^ n2654 ^ 1'b0 ;
  assign n43432 = n33184 & n43431 ;
  assign n43433 = n32109 ^ n31624 ^ 1'b0 ;
  assign n43434 = n13512 & ~n32788 ;
  assign n43435 = ~n2301 & n19775 ;
  assign n43436 = ( n9764 & n33036 ) | ( n9764 & n43435 ) | ( n33036 & n43435 ) ;
  assign n43437 = n31514 ^ n7776 ^ 1'b0 ;
  assign n43438 = n40019 ^ n35252 ^ n16619 ;
  assign n43439 = n43437 & n43438 ;
  assign n43440 = n22287 ^ n16195 ^ n5276 ;
  assign n43441 = ( n2349 & n6915 ) | ( n2349 & ~n17415 ) | ( n6915 & ~n17415 ) ;
  assign n43442 = ~n10009 & n13911 ;
  assign n43443 = ( n7120 & ~n43441 ) | ( n7120 & n43442 ) | ( ~n43441 & n43442 ) ;
  assign n43444 = n3578 & n43443 ;
  assign n43445 = n43440 & n43444 ;
  assign n43446 = n18158 & n33730 ;
  assign n43447 = ~n36569 & n43446 ;
  assign n43448 = n9449 ^ n811 ^ 1'b0 ;
  assign n43449 = ~n43447 & n43448 ;
  assign n43450 = ~n2263 & n23447 ;
  assign n43451 = n14472 & n43450 ;
  assign n43452 = n43451 ^ n19188 ^ 1'b0 ;
  assign n43453 = n22330 | n25476 ;
  assign n43454 = n3836 | n20242 ;
  assign n43455 = n43454 ^ n21652 ^ 1'b0 ;
  assign n43456 = n43455 ^ n1727 ^ 1'b0 ;
  assign n43457 = ( ~n23527 & n43453 ) | ( ~n23527 & n43456 ) | ( n43453 & n43456 ) ;
  assign n43458 = n27149 ^ n24756 ^ n7532 ;
  assign n43459 = n25731 ^ n7500 ^ 1'b0 ;
  assign n43463 = n23109 ^ n21103 ^ n8930 ;
  assign n43460 = n5398 | n16080 ;
  assign n43461 = n26241 & ~n43460 ;
  assign n43462 = n43461 ^ n30571 ^ n17631 ;
  assign n43464 = n43463 ^ n43462 ^ 1'b0 ;
  assign n43465 = n12374 & n22916 ;
  assign n43466 = n3190 & n43465 ;
  assign n43467 = n25733 | n43466 ;
  assign n43468 = n43467 ^ n3262 ^ 1'b0 ;
  assign n43469 = n8836 | n9775 ;
  assign n43470 = n43469 ^ n32002 ^ 1'b0 ;
  assign n43471 = n2669 | n42444 ;
  assign n43473 = ( ~n8046 & n18218 ) | ( ~n8046 & n30479 ) | ( n18218 & n30479 ) ;
  assign n43474 = ~n23107 & n43473 ;
  assign n43475 = n43474 ^ n10339 ^ 1'b0 ;
  assign n43472 = ( ~n5527 & n23160 ) | ( ~n5527 & n32308 ) | ( n23160 & n32308 ) ;
  assign n43476 = n43475 ^ n43472 ^ n30877 ;
  assign n43477 = n6097 & n14923 ;
  assign n43478 = n43477 ^ n27280 ^ 1'b0 ;
  assign n43480 = ( n5377 & n12215 ) | ( n5377 & n16677 ) | ( n12215 & n16677 ) ;
  assign n43479 = n19696 ^ n7798 ^ n4890 ;
  assign n43481 = n43480 ^ n43479 ^ 1'b0 ;
  assign n43483 = ( ~n1004 & n10436 ) | ( ~n1004 & n20994 ) | ( n10436 & n20994 ) ;
  assign n43482 = ( n11635 & n18328 ) | ( n11635 & n18766 ) | ( n18328 & n18766 ) ;
  assign n43484 = n43483 ^ n43482 ^ 1'b0 ;
  assign n43485 = n40012 & ~n43484 ;
  assign n43486 = ~n2363 & n4398 ;
  assign n43487 = n43486 ^ n368 ^ 1'b0 ;
  assign n43494 = ~n4869 & n27984 ;
  assign n43495 = n9626 & n43494 ;
  assign n43491 = ( ~n5588 & n5759 ) | ( ~n5588 & n25562 ) | ( n5759 & n25562 ) ;
  assign n43488 = n14578 & n36878 ;
  assign n43489 = n8052 & n43488 ;
  assign n43490 = n13398 | n43489 ;
  assign n43492 = n43491 ^ n43490 ^ n21603 ;
  assign n43493 = n26529 & n43492 ;
  assign n43496 = n43495 ^ n43493 ^ 1'b0 ;
  assign n43497 = n17924 & ~n18321 ;
  assign n43498 = n43497 ^ n24370 ^ 1'b0 ;
  assign n43499 = n13788 & n30235 ;
  assign n43500 = n43499 ^ n25891 ^ 1'b0 ;
  assign n43501 = n1863 | n8017 ;
  assign n43502 = n43501 ^ n7530 ^ 1'b0 ;
  assign n43503 = n9486 | n28287 ;
  assign n43504 = n43503 ^ n37746 ^ n14759 ;
  assign n43505 = n43504 ^ n19679 ^ n16979 ;
  assign n43506 = n28753 ^ n17355 ^ 1'b0 ;
  assign n43507 = n43506 ^ n31171 ^ n1707 ;
  assign n43508 = n13647 & ~n24184 ;
  assign n43509 = n43508 ^ n31948 ^ 1'b0 ;
  assign n43510 = ~n31698 & n43509 ;
  assign n43511 = n5613 & n9460 ;
  assign n43512 = n2386 | n43511 ;
  assign n43513 = n43512 ^ n15010 ^ 1'b0 ;
  assign n43514 = n40527 ^ n11426 ^ 1'b0 ;
  assign n43515 = n17948 & ~n43514 ;
  assign n43516 = n2348 | n23403 ;
  assign n43517 = ( ~n7273 & n43515 ) | ( ~n7273 & n43516 ) | ( n43515 & n43516 ) ;
  assign n43518 = n2778 & ~n21887 ;
  assign n43519 = n2847 ^ n876 ^ 1'b0 ;
  assign n43520 = n43518 | n43519 ;
  assign n43521 = n2078 | n43520 ;
  assign n43522 = n10557 & n35707 ;
  assign n43523 = n43522 ^ n30643 ^ 1'b0 ;
  assign n43524 = n43523 ^ n12267 ^ 1'b0 ;
  assign n43525 = n13515 ^ n9082 ^ 1'b0 ;
  assign n43526 = n33240 ^ n1069 ^ 1'b0 ;
  assign n43527 = ~n35506 & n43526 ;
  assign n43528 = n26871 ^ n16945 ^ n745 ;
  assign n43529 = n43527 & n43528 ;
  assign n43530 = n15731 | n16051 ;
  assign n43531 = n13623 & n32267 ;
  assign n43532 = n43531 ^ n27787 ^ 1'b0 ;
  assign n43533 = n41420 ^ n22035 ^ 1'b0 ;
  assign n43534 = ~n14796 & n43533 ;
  assign n43535 = ~n17649 & n20506 ;
  assign n43536 = n40666 & n43535 ;
  assign n43537 = n14147 ^ n2828 ^ 1'b0 ;
  assign n43538 = n16284 & n43537 ;
  assign n43539 = n32314 & n43538 ;
  assign n43540 = n12374 & ~n34641 ;
  assign n43541 = n12353 ^ n3104 ^ 1'b0 ;
  assign n43542 = ( ~n2850 & n12091 ) | ( ~n2850 & n19375 ) | ( n12091 & n19375 ) ;
  assign n43543 = n9113 & ~n38168 ;
  assign n43544 = n38766 ^ n1100 ^ 1'b0 ;
  assign n43545 = n21729 ^ n310 ^ 1'b0 ;
  assign n43546 = n42801 ^ n6832 ^ 1'b0 ;
  assign n43547 = n20483 ^ n11251 ^ 1'b0 ;
  assign n43548 = n25917 | n43547 ;
  assign n43549 = n10326 ^ n7885 ^ n1950 ;
  assign n43550 = n43549 ^ n37559 ^ n18349 ;
  assign n43551 = n43303 ^ n7990 ^ n921 ;
  assign n43552 = n43551 ^ n21206 ^ 1'b0 ;
  assign n43553 = n16569 ^ n15870 ^ 1'b0 ;
  assign n43554 = n42972 ^ n7601 ^ 1'b0 ;
  assign n43555 = ~n13262 & n43554 ;
  assign n43556 = n9871 & n43555 ;
  assign n43557 = ~n4487 & n43556 ;
  assign n43558 = n381 | n8494 ;
  assign n43559 = n43558 ^ n26646 ^ 1'b0 ;
  assign n43560 = n14677 ^ n11790 ^ n2075 ;
  assign n43561 = n43560 ^ n18956 ^ n8835 ;
  assign n43562 = n16311 & n37495 ;
  assign n43563 = n43562 ^ n43234 ^ 1'b0 ;
  assign n43564 = n32602 | n42553 ;
  assign n43565 = n22161 ^ n9884 ^ 1'b0 ;
  assign n43566 = n18516 ^ n678 ^ 1'b0 ;
  assign n43567 = ~n43565 & n43566 ;
  assign n43568 = n32168 ^ n28643 ^ 1'b0 ;
  assign n43569 = n7966 | n43568 ;
  assign n43570 = n43569 ^ n16571 ^ 1'b0 ;
  assign n43571 = n12691 & ~n43570 ;
  assign n43572 = ( n22794 & n24914 ) | ( n22794 & n34496 ) | ( n24914 & n34496 ) ;
  assign n43574 = n18778 ^ n1179 ^ 1'b0 ;
  assign n43573 = ( ~n13268 & n17044 ) | ( ~n13268 & n26383 ) | ( n17044 & n26383 ) ;
  assign n43575 = n43574 ^ n43573 ^ n7885 ;
  assign n43576 = n35170 ^ n18416 ^ n12896 ;
  assign n43577 = ~n24446 & n43576 ;
  assign n43578 = n13420 & n25065 ;
  assign n43579 = n9277 & n43578 ;
  assign n43580 = ~n26604 & n34756 ;
  assign n43587 = ( n18602 & n22254 ) | ( n18602 & n24103 ) | ( n22254 & n24103 ) ;
  assign n43581 = n32015 ^ n14183 ^ 1'b0 ;
  assign n43582 = n30599 | n43581 ;
  assign n43583 = ~n10973 & n13067 ;
  assign n43584 = n43582 & n43583 ;
  assign n43585 = ( x53 & ~n41518 ) | ( x53 & n43584 ) | ( ~n41518 & n43584 ) ;
  assign n43586 = ~n20913 & n43585 ;
  assign n43588 = n43587 ^ n43586 ^ 1'b0 ;
  assign n43589 = n17023 ^ n11817 ^ 1'b0 ;
  assign n43590 = ( n2919 & n5317 ) | ( n2919 & n7337 ) | ( n5317 & n7337 ) ;
  assign n43591 = ( ~n5331 & n13637 ) | ( ~n5331 & n43590 ) | ( n13637 & n43590 ) ;
  assign n43592 = n18114 ^ n7900 ^ 1'b0 ;
  assign n43593 = n15591 ^ n13981 ^ 1'b0 ;
  assign n43594 = n23509 & ~n43593 ;
  assign n43595 = n11131 & ~n19122 ;
  assign n43596 = ~n43594 & n43595 ;
  assign n43597 = x247 & ~n33296 ;
  assign n43598 = ~n7037 & n43597 ;
  assign n43599 = n9675 | n43598 ;
  assign n43600 = n43599 ^ n7015 ^ 1'b0 ;
  assign n43601 = n6815 | n13250 ;
  assign n43602 = n41204 | n43601 ;
  assign n43603 = n25601 ^ n9349 ^ 1'b0 ;
  assign n43604 = n20207 ^ n15224 ^ 1'b0 ;
  assign n43605 = n24041 | n43604 ;
  assign n43606 = n13508 & ~n43605 ;
  assign n43607 = n42323 ^ n24096 ^ n2210 ;
  assign n43608 = n20369 & n27072 ;
  assign n43609 = n43608 ^ n15418 ^ 1'b0 ;
  assign n43610 = n43609 ^ n42919 ^ n7384 ;
  assign n43611 = n43610 ^ n27230 ^ n18519 ;
  assign n43612 = n18347 ^ n13102 ^ n3479 ;
  assign n43613 = n22682 ^ n17651 ^ 1'b0 ;
  assign n43614 = n7493 | n43613 ;
  assign n43615 = n43614 ^ n43101 ^ 1'b0 ;
  assign n43616 = n7805 | n43615 ;
  assign n43617 = ~n453 & n36367 ;
  assign n43618 = n43617 ^ n6322 ^ 1'b0 ;
  assign n43619 = ~n13999 & n35857 ;
  assign n43620 = n22047 ^ n21886 ^ 1'b0 ;
  assign n43621 = n43609 & n43620 ;
  assign n43622 = ( n20979 & n28374 ) | ( n20979 & n30160 ) | ( n28374 & n30160 ) ;
  assign n43623 = n32160 ^ n17367 ^ 1'b0 ;
  assign n43624 = n43067 ^ n12006 ^ 1'b0 ;
  assign n43625 = n7761 | n15086 ;
  assign n43626 = ( n27981 & n43624 ) | ( n27981 & ~n43625 ) | ( n43624 & ~n43625 ) ;
  assign n43627 = n43264 ^ n19785 ^ n11532 ;
  assign n43628 = n9296 & n17213 ;
  assign n43629 = ~n7892 & n33184 ;
  assign n43630 = n28264 & n43629 ;
  assign n43631 = n1545 ^ n917 ^ 1'b0 ;
  assign n43632 = ~n21154 & n43631 ;
  assign n43633 = n2651 | n11082 ;
  assign n43643 = ~n19558 & n23885 ;
  assign n43641 = n6839 & n9237 ;
  assign n43642 = n8928 & n43641 ;
  assign n43637 = n5416 | n5947 ;
  assign n43638 = n11800 & ~n43637 ;
  assign n43639 = ~n20219 & n43638 ;
  assign n43634 = n16067 ^ n8240 ^ 1'b0 ;
  assign n43635 = n35475 & ~n43634 ;
  assign n43636 = n8658 & n43635 ;
  assign n43640 = n43639 ^ n43636 ^ 1'b0 ;
  assign n43644 = n43643 ^ n43642 ^ n43640 ;
  assign n43645 = n17766 ^ n7028 ^ 1'b0 ;
  assign n43646 = n863 | n31502 ;
  assign n43647 = n43646 ^ n22342 ^ 1'b0 ;
  assign n43648 = n43647 ^ n24545 ^ n12010 ;
  assign n43649 = n545 | n7788 ;
  assign n43650 = n9937 | n11501 ;
  assign n43651 = n43650 ^ n29037 ^ 1'b0 ;
  assign n43652 = ~n41888 & n43651 ;
  assign n43653 = n41089 & n43652 ;
  assign n43654 = n8997 & n30957 ;
  assign n43655 = n2007 & ~n34853 ;
  assign n43656 = n38311 ^ n7393 ^ 1'b0 ;
  assign n43657 = n29600 & ~n43656 ;
  assign n43658 = ~n34976 & n39165 ;
  assign n43659 = n18803 | n38249 ;
  assign n43660 = n34646 | n43659 ;
  assign n43661 = n43660 ^ n24347 ^ 1'b0 ;
  assign n43662 = ~n7851 & n20448 ;
  assign n43663 = n43662 ^ n1367 ^ 1'b0 ;
  assign n43664 = ( ~n16474 & n16992 ) | ( ~n16474 & n43663 ) | ( n16992 & n43663 ) ;
  assign n43665 = n7242 & n12326 ;
  assign n43666 = n12944 & ~n43665 ;
  assign n43667 = n37235 ^ n23109 ^ n22611 ;
  assign n43668 = x254 | n4229 ;
  assign n43669 = ( n12593 & ~n26799 ) | ( n12593 & n43668 ) | ( ~n26799 & n43668 ) ;
  assign n43670 = n5789 & n31829 ;
  assign n43671 = n10344 & ~n25721 ;
  assign n43672 = n43671 ^ n1194 ^ 1'b0 ;
  assign n43673 = ~n815 & n9290 ;
  assign n43674 = n4200 | n12964 ;
  assign n43675 = n29453 & ~n43674 ;
  assign n43676 = ( n21365 & ~n28437 ) | ( n21365 & n33050 ) | ( ~n28437 & n33050 ) ;
  assign n43677 = x211 & n4074 ;
  assign n43678 = n43677 ^ n4050 ^ 1'b0 ;
  assign n43679 = ( x9 & ~n26756 ) | ( x9 & n43678 ) | ( ~n26756 & n43678 ) ;
  assign n43680 = n10945 & ~n15228 ;
  assign n43681 = n16785 ^ n12189 ^ 1'b0 ;
  assign n43682 = ~n41769 & n43681 ;
  assign n43683 = ~n1930 & n33784 ;
  assign n43684 = n43683 ^ n5097 ^ 1'b0 ;
  assign n43685 = n19911 ^ n15841 ^ 1'b0 ;
  assign n43686 = n12104 | n43685 ;
  assign n43687 = n39989 ^ n20223 ^ 1'b0 ;
  assign n43688 = ~n43686 & n43687 ;
  assign n43689 = n37820 ^ n9041 ^ 1'b0 ;
  assign n43690 = n9822 | n43689 ;
  assign n43691 = ( n3714 & n5215 ) | ( n3714 & ~n16599 ) | ( n5215 & ~n16599 ) ;
  assign n43692 = n3625 & ~n43691 ;
  assign n43693 = n13545 ^ n9790 ^ 1'b0 ;
  assign n43694 = ~n1339 & n43693 ;
  assign n43695 = n43694 ^ n16380 ^ 1'b0 ;
  assign n43696 = ( n3199 & n5444 ) | ( n3199 & ~n8069 ) | ( n5444 & ~n8069 ) ;
  assign n43697 = n43696 ^ x24 ^ 1'b0 ;
  assign n43698 = ~n43695 & n43697 ;
  assign n43699 = ~n35899 & n43698 ;
  assign n43700 = ( ~n9823 & n38640 ) | ( ~n9823 & n43699 ) | ( n38640 & n43699 ) ;
  assign n43701 = n29183 ^ n28086 ^ n10292 ;
  assign n43702 = n31228 ^ n23967 ^ n11966 ;
  assign n43703 = n27220 ^ n4356 ^ 1'b0 ;
  assign n43704 = n43702 | n43703 ;
  assign n43705 = ~n363 & n21616 ;
  assign n43706 = n354 ^ x182 ^ 1'b0 ;
  assign n43707 = n19180 & n43706 ;
  assign n43708 = ( n21892 & n28208 ) | ( n21892 & n43707 ) | ( n28208 & n43707 ) ;
  assign n43709 = ~n9506 & n20172 ;
  assign n43710 = ~n3528 & n43709 ;
  assign n43711 = n43710 ^ n18924 ^ n13068 ;
  assign n43712 = n9682 ^ n5670 ^ 1'b0 ;
  assign n43713 = n32572 | n43712 ;
  assign n43714 = n3080 & ~n43713 ;
  assign n43715 = n6530 & n10003 ;
  assign n43716 = n43715 ^ n14606 ^ 1'b0 ;
  assign n43717 = ( n27600 & n43714 ) | ( n27600 & ~n43716 ) | ( n43714 & ~n43716 ) ;
  assign n43718 = ( ~n7747 & n9610 ) | ( ~n7747 & n11811 ) | ( n9610 & n11811 ) ;
  assign n43719 = ~n10121 & n16106 ;
  assign n43720 = ( n28024 & n43718 ) | ( n28024 & n43719 ) | ( n43718 & n43719 ) ;
  assign n43721 = n13035 ^ n12969 ^ 1'b0 ;
  assign n43722 = n3093 & ~n43721 ;
  assign n43723 = n23086 & ~n43722 ;
  assign n43726 = ~n37553 & n41612 ;
  assign n43724 = ~n840 & n6260 ;
  assign n43725 = ~n15306 & n43724 ;
  assign n43727 = n43726 ^ n43725 ^ 1'b0 ;
  assign n43728 = n3792 & n25294 ;
  assign n43729 = ~n32529 & n43728 ;
  assign n43730 = n43729 ^ n24379 ^ 1'b0 ;
  assign n43731 = n1048 & n20945 ;
  assign n43732 = n43731 ^ n41440 ^ 1'b0 ;
  assign n43733 = n7860 & ~n37211 ;
  assign n43734 = ( n11418 & n15707 ) | ( n11418 & ~n33430 ) | ( n15707 & ~n33430 ) ;
  assign n43737 = n4730 & ~n5947 ;
  assign n43738 = ~n1393 & n43737 ;
  assign n43735 = n4033 & ~n9088 ;
  assign n43736 = n43735 ^ n18033 ^ 1'b0 ;
  assign n43739 = n43738 ^ n43736 ^ n33590 ;
  assign n43740 = n30387 ^ n29922 ^ n4933 ;
  assign n43741 = ~n32658 & n43740 ;
  assign n43742 = n8905 ^ n1962 ^ 1'b0 ;
  assign n43743 = x130 & ~n28798 ;
  assign n43744 = n43743 ^ n22513 ^ 1'b0 ;
  assign n43745 = n43742 & n43744 ;
  assign n43747 = ~n12458 & n38617 ;
  assign n43748 = n28955 & n43747 ;
  assign n43749 = ( n3356 & n19386 ) | ( n3356 & ~n43748 ) | ( n19386 & ~n43748 ) ;
  assign n43746 = x169 & ~n32433 ;
  assign n43750 = n43749 ^ n43746 ^ 1'b0 ;
  assign n43751 = n37389 ^ n36764 ^ 1'b0 ;
  assign n43752 = n41599 | n43751 ;
  assign n43753 = n14689 ^ n10939 ^ n9296 ;
  assign n43754 = n12796 | n43753 ;
  assign n43755 = n8198 & n18889 ;
  assign n43756 = n43755 ^ n13158 ^ 1'b0 ;
  assign n43757 = ( n22824 & n38386 ) | ( n22824 & ~n43756 ) | ( n38386 & ~n43756 ) ;
  assign n43758 = n5112 | n7936 ;
  assign n43759 = n34642 ^ n7814 ^ n6143 ;
  assign n43760 = n22519 & n29081 ;
  assign n43761 = n43760 ^ n29753 ^ 1'b0 ;
  assign n43762 = n12939 & n38014 ;
  assign n43763 = ~n39041 & n43762 ;
  assign n43764 = n14443 ^ n2314 ^ 1'b0 ;
  assign n43765 = n17115 & n43764 ;
  assign n43768 = ( n1971 & ~n18009 ) | ( n1971 & n37589 ) | ( ~n18009 & n37589 ) ;
  assign n43769 = n12493 & ~n24392 ;
  assign n43770 = ~n1010 & n43769 ;
  assign n43771 = ( n3166 & ~n43768 ) | ( n3166 & n43770 ) | ( ~n43768 & n43770 ) ;
  assign n43766 = n15128 & ~n32988 ;
  assign n43767 = ~n4661 & n43766 ;
  assign n43772 = n43771 ^ n43767 ^ n27314 ;
  assign n43773 = n503 & ~n38003 ;
  assign n43774 = ( n2083 & ~n9364 ) | ( n2083 & n42842 ) | ( ~n9364 & n42842 ) ;
  assign n43775 = n23387 ^ n7478 ^ 1'b0 ;
  assign n43776 = n32654 ^ n22726 ^ n2005 ;
  assign n43777 = ( n18800 & ~n43775 ) | ( n18800 & n43776 ) | ( ~n43775 & n43776 ) ;
  assign n43778 = n39297 ^ n1655 ^ 1'b0 ;
  assign n43779 = n43777 & n43778 ;
  assign n43780 = ( n7759 & n11251 ) | ( n7759 & n26441 ) | ( n11251 & n26441 ) ;
  assign n43781 = ~n8430 & n43780 ;
  assign n43782 = n7942 & n43781 ;
  assign n43784 = ~n21108 & n23544 ;
  assign n43785 = n43784 ^ n36560 ^ 1'b0 ;
  assign n43783 = n6259 | n31399 ;
  assign n43786 = n43785 ^ n43783 ^ 1'b0 ;
  assign n43787 = n11207 ^ n8521 ^ 1'b0 ;
  assign n43788 = n37891 | n43787 ;
  assign n43789 = n7995 & ~n43788 ;
  assign n43790 = n43789 ^ n21339 ^ 1'b0 ;
  assign n43791 = n22917 ^ n17358 ^ 1'b0 ;
  assign n43792 = n11228 | n43791 ;
  assign n43793 = n38158 ^ n11234 ^ 1'b0 ;
  assign n43794 = ~n5424 & n43793 ;
  assign n43798 = n25034 ^ n20631 ^ 1'b0 ;
  assign n43795 = n19186 & n40701 ;
  assign n43796 = ~n5909 & n43795 ;
  assign n43797 = n32983 | n43796 ;
  assign n43799 = n43798 ^ n43797 ^ 1'b0 ;
  assign n43800 = n1862 | n37625 ;
  assign n43801 = n1063 & ~n2937 ;
  assign n43802 = n3639 & n13743 ;
  assign n43803 = n43802 ^ n11613 ^ 1'b0 ;
  assign n43804 = n43803 ^ n12715 ^ 1'b0 ;
  assign n43806 = ( ~n8623 & n18250 ) | ( ~n8623 & n20162 ) | ( n18250 & n20162 ) ;
  assign n43805 = n6841 & n16758 ;
  assign n43807 = n43806 ^ n43805 ^ 1'b0 ;
  assign n43808 = ~n4840 & n8762 ;
  assign n43809 = n7242 & n43808 ;
  assign n43810 = n4989 & ~n43809 ;
  assign n43811 = n43807 & n43810 ;
  assign n43812 = n10266 ^ n5144 ^ 1'b0 ;
  assign n43813 = ~n6616 & n43812 ;
  assign n43814 = ( n5518 & n5842 ) | ( n5518 & n43813 ) | ( n5842 & n43813 ) ;
  assign n43815 = n40141 | n43814 ;
  assign n43816 = ~n4597 & n20875 ;
  assign n43817 = n20442 & n42002 ;
  assign n43818 = n43817 ^ n12021 ^ 1'b0 ;
  assign n43819 = n13234 ^ n2019 ^ 1'b0 ;
  assign n43820 = n22299 & n43819 ;
  assign n43821 = ( n27281 & n29986 ) | ( n27281 & ~n38187 ) | ( n29986 & ~n38187 ) ;
  assign n43822 = n23462 ^ n5106 ^ 1'b0 ;
  assign n43823 = n43822 ^ n36638 ^ n7520 ;
  assign n43824 = n15686 ^ n7168 ^ n947 ;
  assign n43825 = ~n5987 & n9059 ;
  assign n43826 = n43825 ^ n43190 ^ 1'b0 ;
  assign n43827 = n11979 & ~n17756 ;
  assign n43828 = n23784 & n43827 ;
  assign n43829 = n270 & n43828 ;
  assign n43830 = x217 & n38494 ;
  assign n43831 = n43830 ^ n11188 ^ 1'b0 ;
  assign n43832 = n21162 ^ n8250 ^ x131 ;
  assign n43833 = ~n27893 & n43832 ;
  assign n43834 = ~n23584 & n39340 ;
  assign n43835 = n27060 & ~n40053 ;
  assign n43836 = n43835 ^ n4528 ^ 1'b0 ;
  assign n43837 = n43836 ^ n35493 ^ n3475 ;
  assign n43838 = n6509 ^ n4256 ^ 1'b0 ;
  assign n43839 = n27264 & n43838 ;
  assign n43840 = n3858 & ~n20642 ;
  assign n43841 = n43840 ^ n3223 ^ 1'b0 ;
  assign n43842 = ( ~n40540 & n43839 ) | ( ~n40540 & n43841 ) | ( n43839 & n43841 ) ;
  assign n43843 = n31188 ^ n7589 ^ n7173 ;
  assign n43844 = n43843 ^ n2362 ^ 1'b0 ;
  assign n43846 = n24975 ^ n3410 ^ 1'b0 ;
  assign n43847 = n1742 | n43846 ;
  assign n43848 = n39399 & ~n43847 ;
  assign n43849 = n16978 & ~n43848 ;
  assign n43850 = n43849 ^ n16877 ^ 1'b0 ;
  assign n43845 = ~n16686 & n43161 ;
  assign n43851 = n43850 ^ n43845 ^ 1'b0 ;
  assign n43852 = ~n25732 & n33817 ;
  assign n43853 = n43852 ^ n42399 ^ 1'b0 ;
  assign n43855 = n28762 ^ n18055 ^ x148 ;
  assign n43856 = ~n9388 & n11330 ;
  assign n43857 = n43855 & n43856 ;
  assign n43854 = n25170 & ~n43190 ;
  assign n43858 = n43857 ^ n43854 ^ 1'b0 ;
  assign n43859 = n22005 & ~n42052 ;
  assign n43860 = n4296 | n20724 ;
  assign n43861 = ( n1532 & n22885 ) | ( n1532 & n43860 ) | ( n22885 & n43860 ) ;
  assign n43862 = ( ~n15081 & n24256 ) | ( ~n15081 & n43861 ) | ( n24256 & n43861 ) ;
  assign n43863 = n12902 | n26219 ;
  assign n43864 = ~x206 & n14765 ;
  assign n43865 = n43864 ^ n42533 ^ 1'b0 ;
  assign n43866 = ~n4114 & n43865 ;
  assign n43867 = ~n13629 & n15217 ;
  assign n43868 = n7653 ^ n2877 ^ 1'b0 ;
  assign n43869 = n3590 & ~n43868 ;
  assign n43870 = ( ~n3255 & n15724 ) | ( ~n3255 & n43869 ) | ( n15724 & n43869 ) ;
  assign n43871 = n43870 ^ n24120 ^ n22459 ;
  assign n43872 = n24094 ^ n18848 ^ 1'b0 ;
  assign n43873 = n15361 ^ n13172 ^ 1'b0 ;
  assign n43874 = n17294 ^ n14621 ^ 1'b0 ;
  assign n43875 = n17226 | n43874 ;
  assign n43876 = n2256 & ~n43875 ;
  assign n43877 = n4935 & n8585 ;
  assign n43878 = ~n5945 & n43877 ;
  assign n43879 = n729 | n6940 ;
  assign n43880 = n43879 ^ n5564 ^ 1'b0 ;
  assign n43881 = n43880 ^ n39340 ^ n32994 ;
  assign n43882 = n3511 & n21417 ;
  assign n43883 = ~n15654 & n43882 ;
  assign n43884 = n43883 ^ n1538 ^ 1'b0 ;
  assign n43885 = n43881 & ~n43884 ;
  assign n43886 = n24442 ^ n16213 ^ n13766 ;
  assign n43887 = n20343 ^ n2453 ^ 1'b0 ;
  assign n43888 = n31172 ^ n17851 ^ n5515 ;
  assign n43889 = n1173 & ~n23129 ;
  assign n43890 = n43889 ^ n31406 ^ 1'b0 ;
  assign n43891 = ~n23781 & n36376 ;
  assign n43892 = n16221 & n43891 ;
  assign n43893 = n5174 & ~n13584 ;
  assign n43894 = n18493 ^ n13992 ^ 1'b0 ;
  assign n43895 = n9525 & ~n43894 ;
  assign n43896 = ~n43893 & n43895 ;
  assign n43897 = n27883 ^ n3581 ^ 1'b0 ;
  assign n43898 = n12852 & ~n32084 ;
  assign n43899 = n43898 ^ n23030 ^ n21369 ;
  assign n43900 = ( ~n15630 & n28010 ) | ( ~n15630 & n42783 ) | ( n28010 & n42783 ) ;
  assign n43903 = ~n33897 & n35463 ;
  assign n43901 = n21206 ^ n9807 ^ 1'b0 ;
  assign n43902 = n9015 & n43901 ;
  assign n43904 = n43903 ^ n43902 ^ n10856 ;
  assign n43906 = n22186 & ~n43219 ;
  assign n43907 = ~n7028 & n43906 ;
  assign n43905 = ~n11296 & n14789 ;
  assign n43908 = n43907 ^ n43905 ^ 1'b0 ;
  assign n43909 = n15881 ^ n7022 ^ 1'b0 ;
  assign n43910 = n4457 & ~n43909 ;
  assign n43911 = n31793 & n43910 ;
  assign n43912 = ~n18331 & n43911 ;
  assign n43913 = n43912 ^ n13317 ^ 1'b0 ;
  assign n43914 = n27321 ^ n17649 ^ n8194 ;
  assign n43915 = n18550 & ~n22361 ;
  assign n43916 = n43915 ^ n24103 ^ 1'b0 ;
  assign n43917 = ( n19725 & n28507 ) | ( n19725 & ~n43916 ) | ( n28507 & ~n43916 ) ;
  assign n43918 = ( n13614 & ~n14324 ) | ( n13614 & n27108 ) | ( ~n14324 & n27108 ) ;
  assign n43919 = n43918 ^ n7031 ^ n2983 ;
  assign n43920 = n2831 & ~n43919 ;
  assign n43921 = n41737 ^ n7608 ^ 1'b0 ;
  assign n43922 = n11387 | n43921 ;
  assign n43923 = n43922 ^ n10722 ^ 1'b0 ;
  assign n43924 = n16725 & ~n38985 ;
  assign n43925 = n9618 & ~n25850 ;
  assign n43926 = n378 & n43925 ;
  assign n43927 = n8388 | n43926 ;
  assign n43928 = n3590 | n43927 ;
  assign n43929 = ~n19227 & n43928 ;
  assign n43931 = n28786 ^ n4715 ^ 1'b0 ;
  assign n43932 = n19766 & ~n43931 ;
  assign n43930 = n3662 & n31277 ;
  assign n43933 = n43932 ^ n43930 ^ n3100 ;
  assign n43934 = n15858 & ~n23109 ;
  assign n43935 = ~n43933 & n43934 ;
  assign n43936 = n24231 & n25546 ;
  assign n43937 = n40157 ^ n36507 ^ n20486 ;
  assign n43938 = n23370 & ~n25776 ;
  assign n43939 = n5969 & ~n20556 ;
  assign n43941 = n10122 ^ n3667 ^ 1'b0 ;
  assign n43940 = x204 & ~n32574 ;
  assign n43942 = n43941 ^ n43940 ^ 1'b0 ;
  assign n43943 = ~n16097 & n36146 ;
  assign n43944 = n43943 ^ n26996 ^ n928 ;
  assign n43945 = n25917 & ~n43944 ;
  assign n43946 = n13241 ^ n12014 ^ 1'b0 ;
  assign n43947 = ( n20752 & ~n35624 ) | ( n20752 & n36245 ) | ( ~n35624 & n36245 ) ;
  assign n43948 = n2662 & ~n22568 ;
  assign n43949 = n32673 ^ n11790 ^ n6188 ;
  assign n43950 = n12470 | n43949 ;
  assign n43951 = n11174 | n28800 ;
  assign n43952 = n43951 ^ n12598 ^ 1'b0 ;
  assign n43954 = n33763 ^ n10832 ^ 1'b0 ;
  assign n43955 = ~n40542 & n43954 ;
  assign n43953 = n34145 | n42646 ;
  assign n43956 = n43955 ^ n43953 ^ 1'b0 ;
  assign n43957 = n1401 | n13968 ;
  assign n43958 = n43957 ^ n34754 ^ n22209 ;
  assign n43959 = n6008 & ~n23604 ;
  assign n43960 = n43959 ^ n18722 ^ 1'b0 ;
  assign n43961 = n36468 ^ n26527 ^ n8580 ;
  assign n43962 = n1415 | n6165 ;
  assign n43963 = n43961 & ~n43962 ;
  assign n43964 = n43963 ^ n15385 ^ n12247 ;
  assign n43965 = ( n12694 & n21194 ) | ( n12694 & ~n43964 ) | ( n21194 & ~n43964 ) ;
  assign n43966 = n29069 | n31700 ;
  assign n43967 = n3656 & ~n43966 ;
  assign n43968 = ~n14630 & n42317 ;
  assign n43969 = n23182 ^ n7638 ^ 1'b0 ;
  assign n43970 = n593 & ~n43969 ;
  assign n43971 = n43970 ^ n35343 ^ 1'b0 ;
  assign n43972 = n25994 ^ n9759 ^ 1'b0 ;
  assign n43973 = ( n6678 & ~n11635 ) | ( n6678 & n14852 ) | ( ~n11635 & n14852 ) ;
  assign n43974 = n12122 & n43973 ;
  assign n43975 = n38813 ^ n19591 ^ n8834 ;
  assign n43976 = n9129 & n20339 ;
  assign n43977 = n43976 ^ n2117 ^ 1'b0 ;
  assign n43978 = n10154 & ~n13399 ;
  assign n43979 = n12342 & n43978 ;
  assign n43980 = ~n639 & n43979 ;
  assign n43981 = n43980 ^ n19648 ^ 1'b0 ;
  assign n43982 = n20254 ^ n14122 ^ 1'b0 ;
  assign n43983 = n8057 | n43982 ;
  assign n43984 = n12064 | n43983 ;
  assign n43985 = n43984 ^ n20505 ^ 1'b0 ;
  assign n43986 = n42233 ^ n13857 ^ n8981 ;
  assign n43987 = n43986 ^ n13667 ^ 1'b0 ;
  assign n43988 = ~n10085 & n43987 ;
  assign n43989 = n13632 & ~n20438 ;
  assign n43990 = n43989 ^ n9274 ^ 1'b0 ;
  assign n43991 = n10691 & ~n43990 ;
  assign n43992 = ( n1361 & n2769 ) | ( n1361 & n14366 ) | ( n2769 & n14366 ) ;
  assign n43993 = ~n15359 & n26993 ;
  assign n43994 = n38937 | n43993 ;
  assign n43995 = n39315 ^ n20980 ^ n8155 ;
  assign n43996 = ~n3831 & n7694 ;
  assign n43997 = n43996 ^ n15950 ^ 1'b0 ;
  assign n43998 = n270 | n43997 ;
  assign n43999 = n26545 ^ n21222 ^ n1334 ;
  assign n44000 = n16441 | n43999 ;
  assign n44001 = n2942 | n44000 ;
  assign n44002 = n20909 ^ n1831 ^ 1'b0 ;
  assign n44003 = n16600 & n44002 ;
  assign n44004 = ~n3053 & n11412 ;
  assign n44005 = ~n1152 & n44004 ;
  assign n44006 = n19648 | n19957 ;
  assign n44007 = ( n2443 & n11448 ) | ( n2443 & n44006 ) | ( n11448 & n44006 ) ;
  assign n44008 = ( ~n15478 & n44005 ) | ( ~n15478 & n44007 ) | ( n44005 & n44007 ) ;
  assign n44009 = n2840 ^ x104 ^ 1'b0 ;
  assign n44010 = ( n5779 & ~n11852 ) | ( n5779 & n40957 ) | ( ~n11852 & n40957 ) ;
  assign n44011 = n29975 ^ n6434 ^ x56 ;
  assign n44012 = n10289 & n15451 ;
  assign n44013 = n44012 ^ n4055 ^ 1'b0 ;
  assign n44014 = n8481 & ~n44013 ;
  assign n44015 = n44014 ^ n22737 ^ 1'b0 ;
  assign n44016 = n5381 ^ n1999 ^ 1'b0 ;
  assign n44017 = n9816 & ~n44016 ;
  assign n44018 = n27827 ^ n8358 ^ 1'b0 ;
  assign n44019 = n24003 | n44018 ;
  assign n44020 = n2671 & ~n18112 ;
  assign n44021 = ~x44 & n27730 ;
  assign n44022 = ( n3991 & n35903 ) | ( n3991 & n44021 ) | ( n35903 & n44021 ) ;
  assign n44029 = ( n15431 & ~n27176 ) | ( n15431 & n40164 ) | ( ~n27176 & n40164 ) ;
  assign n44024 = n1129 & ~n4039 ;
  assign n44026 = n556 & ~n20164 ;
  assign n44025 = n1733 | n11001 ;
  assign n44027 = n44026 ^ n44025 ^ 1'b0 ;
  assign n44028 = ~n44024 & n44027 ;
  assign n44023 = n10432 ^ n6551 ^ x61 ;
  assign n44030 = n44029 ^ n44028 ^ n44023 ;
  assign n44031 = ( n8894 & n34465 ) | ( n8894 & ~n41604 ) | ( n34465 & ~n41604 ) ;
  assign n44032 = n44031 ^ n25072 ^ n2464 ;
  assign n44033 = ( n19858 & n26379 ) | ( n19858 & n28791 ) | ( n26379 & n28791 ) ;
  assign n44034 = n18255 | n19533 ;
  assign n44035 = n44034 ^ n3632 ^ 1'b0 ;
  assign n44036 = ( n6603 & n11106 ) | ( n6603 & n44035 ) | ( n11106 & n44035 ) ;
  assign n44037 = ~n27029 & n44036 ;
  assign n44038 = n42275 ^ n10516 ^ 1'b0 ;
  assign n44039 = n23876 ^ n545 ^ 1'b0 ;
  assign n44040 = n18561 ^ n17365 ^ 1'b0 ;
  assign n44041 = ( n256 & n6523 ) | ( n256 & n8521 ) | ( n6523 & n8521 ) ;
  assign n44042 = ( n14171 & ~n23370 ) | ( n14171 & n44041 ) | ( ~n23370 & n44041 ) ;
  assign n44043 = n20215 ^ n12944 ^ n12435 ;
  assign n44044 = n9781 ^ n1009 ^ 1'b0 ;
  assign n44045 = ( n3529 & n44043 ) | ( n3529 & ~n44044 ) | ( n44043 & ~n44044 ) ;
  assign n44046 = ~n9264 & n24608 ;
  assign n44047 = n15305 & n44046 ;
  assign n44048 = n44047 ^ n5680 ^ 1'b0 ;
  assign n44049 = n43944 ^ n42526 ^ 1'b0 ;
  assign n44050 = n11981 ^ n6221 ^ 1'b0 ;
  assign n44051 = ~n14548 & n44050 ;
  assign n44052 = n27732 & ~n44051 ;
  assign n44053 = n44052 ^ n30369 ^ 1'b0 ;
  assign n44054 = n19197 ^ n5502 ^ 1'b0 ;
  assign n44055 = n37233 ^ n24420 ^ 1'b0 ;
  assign n44056 = n16195 ^ n14911 ^ n3275 ;
  assign n44057 = n1842 & n2828 ;
  assign n44058 = n34201 ^ n23672 ^ 1'b0 ;
  assign n44059 = n44057 | n44058 ;
  assign n44060 = n44059 ^ n34803 ^ n1266 ;
  assign n44061 = n34961 ^ n30795 ^ n11192 ;
  assign n44062 = n12231 | n12279 ;
  assign n44063 = n27385 & ~n44062 ;
  assign n44064 = n38546 ^ n19872 ^ 1'b0 ;
  assign n44065 = n25081 | n32641 ;
  assign n44066 = n11023 & ~n14314 ;
  assign n44070 = n12326 ^ n5740 ^ 1'b0 ;
  assign n44067 = n37154 ^ n1472 ^ n759 ;
  assign n44068 = n26446 ^ n16142 ^ 1'b0 ;
  assign n44069 = ( n25824 & n44067 ) | ( n25824 & ~n44068 ) | ( n44067 & ~n44068 ) ;
  assign n44071 = n44070 ^ n44069 ^ 1'b0 ;
  assign n44072 = n20614 ^ n3729 ^ n2489 ;
  assign n44073 = n24379 ^ n10357 ^ 1'b0 ;
  assign n44074 = n27489 & ~n38575 ;
  assign n44075 = ~n25994 & n44074 ;
  assign n44076 = n4756 & ~n17554 ;
  assign n44077 = n2737 | n41483 ;
  assign n44078 = n44077 ^ n2199 ^ n1048 ;
  assign n44079 = n39486 ^ n2680 ^ 1'b0 ;
  assign n44080 = ~n10181 & n44079 ;
  assign n44081 = ~n2658 & n36747 ;
  assign n44082 = ( n33121 & n44080 ) | ( n33121 & n44081 ) | ( n44080 & n44081 ) ;
  assign n44083 = n35104 ^ n31792 ^ 1'b0 ;
  assign n44084 = n18607 & ~n44083 ;
  assign n44085 = ~n19453 & n44084 ;
  assign n44086 = n33308 ^ n33053 ^ 1'b0 ;
  assign n44088 = n25796 ^ n22824 ^ n9100 ;
  assign n44089 = ( x2 & ~n2089 ) | ( x2 & n44088 ) | ( ~n2089 & n44088 ) ;
  assign n44087 = n3425 | n15239 ;
  assign n44090 = n44089 ^ n44087 ^ n21291 ;
  assign n44091 = n44086 & n44090 ;
  assign n44092 = n13359 & ~n22342 ;
  assign n44093 = n44092 ^ n36675 ^ 1'b0 ;
  assign n44095 = n26557 ^ n15010 ^ n3054 ;
  assign n44094 = ~n35290 & n35921 ;
  assign n44096 = n44095 ^ n44094 ^ 1'b0 ;
  assign n44097 = n37608 ^ n2192 ^ 1'b0 ;
  assign n44098 = n31929 ^ n12487 ^ 1'b0 ;
  assign n44099 = n12115 | n40040 ;
  assign n44100 = ~n1703 & n7222 ;
  assign n44101 = n1865 | n23366 ;
  assign n44102 = n44101 ^ n15803 ^ 1'b0 ;
  assign n44103 = ~n14133 & n42526 ;
  assign n44104 = n44103 ^ n3181 ^ 1'b0 ;
  assign n44105 = n31074 & ~n39611 ;
  assign n44106 = ~n34252 & n44105 ;
  assign n44107 = n2006 ^ n467 ^ 1'b0 ;
  assign n44108 = n7760 & ~n13099 ;
  assign n44109 = ~n7784 & n44108 ;
  assign n44111 = n5483 ^ n3000 ^ 1'b0 ;
  assign n44110 = n9577 | n14974 ;
  assign n44112 = n44111 ^ n44110 ^ n33599 ;
  assign n44113 = ( n16206 & n35209 ) | ( n16206 & ~n40511 ) | ( n35209 & ~n40511 ) ;
  assign n44114 = ~n14407 & n24921 ;
  assign n44115 = n44114 ^ n39480 ^ 1'b0 ;
  assign n44116 = n35403 ^ n12614 ^ 1'b0 ;
  assign n44117 = n874 & ~n44116 ;
  assign n44118 = n16243 & ~n44117 ;
  assign n44119 = n24076 & ~n38767 ;
  assign n44120 = ~n27852 & n44119 ;
  assign n44121 = n44120 ^ n4826 ^ 1'b0 ;
  assign n44122 = ~n4968 & n21992 ;
  assign n44123 = n3437 | n44122 ;
  assign n44124 = n2799 ^ n827 ^ 1'b0 ;
  assign n44125 = n2392 & ~n44124 ;
  assign n44126 = n44125 ^ n35263 ^ n8743 ;
  assign n44127 = n29126 ^ n16149 ^ n15788 ;
  assign n44128 = ( ~n40887 & n44126 ) | ( ~n40887 & n44127 ) | ( n44126 & n44127 ) ;
  assign n44129 = n1011 | n6889 ;
  assign n44130 = n6487 & ~n17033 ;
  assign n44131 = n44130 ^ n16081 ^ 1'b0 ;
  assign n44132 = ~n9551 & n26731 ;
  assign n44133 = n44132 ^ n25937 ^ 1'b0 ;
  assign n44134 = n25999 ^ n5649 ^ 1'b0 ;
  assign n44135 = ~n44133 & n44134 ;
  assign n44136 = n40061 ^ n30660 ^ 1'b0 ;
  assign n44137 = n15350 & n39729 ;
  assign n44138 = ~n21500 & n44137 ;
  assign n44139 = n44138 ^ n31524 ^ n21820 ;
  assign n44140 = n40107 ^ n30212 ^ 1'b0 ;
  assign n44141 = ~n17136 & n32287 ;
  assign n44142 = ~n12863 & n44141 ;
  assign n44143 = n8294 & ~n20674 ;
  assign n44144 = n44143 ^ n13065 ^ 1'b0 ;
  assign n44145 = ~n1653 & n10634 ;
  assign n44146 = n44145 ^ n2189 ^ 1'b0 ;
  assign n44147 = ( ~n3904 & n9022 ) | ( ~n3904 & n31628 ) | ( n9022 & n31628 ) ;
  assign n44148 = ~n8606 & n16220 ;
  assign n44149 = n44148 ^ n18001 ^ n5496 ;
  assign n44150 = ( n10961 & n26031 ) | ( n10961 & n44149 ) | ( n26031 & n44149 ) ;
  assign n44151 = n8277 ^ n1937 ^ 1'b0 ;
  assign n44152 = n13273 | n44151 ;
  assign n44153 = n44152 ^ n11048 ^ 1'b0 ;
  assign n44154 = ( n4592 & n6576 ) | ( n4592 & n30217 ) | ( n6576 & n30217 ) ;
  assign n44155 = n16992 & n21283 ;
  assign n44156 = ~n31373 & n44155 ;
  assign n44157 = n4121 & n9682 ;
  assign n44158 = n16049 & n44157 ;
  assign n44159 = n293 | n44158 ;
  assign n44160 = n3485 & ~n44159 ;
  assign n44161 = n26949 ^ n22413 ^ 1'b0 ;
  assign n44162 = n44161 ^ n30636 ^ 1'b0 ;
  assign n44163 = ( n32639 & n38932 ) | ( n32639 & ~n44162 ) | ( n38932 & ~n44162 ) ;
  assign n44164 = n2640 & n44163 ;
  assign n44165 = n44164 ^ n42247 ^ 1'b0 ;
  assign n44166 = n3188 & ~n9814 ;
  assign n44167 = ~n18822 & n44166 ;
  assign n44168 = n16577 | n29186 ;
  assign n44169 = n44167 & ~n44168 ;
  assign n44172 = n13493 & ~n14687 ;
  assign n44173 = n44172 ^ n2114 ^ 1'b0 ;
  assign n44174 = n44173 ^ n18778 ^ 1'b0 ;
  assign n44175 = n18092 & n44174 ;
  assign n44170 = n18233 ^ n11322 ^ 1'b0 ;
  assign n44171 = n30212 & n44170 ;
  assign n44176 = n44175 ^ n44171 ^ 1'b0 ;
  assign n44177 = n6804 ^ n1548 ^ 1'b0 ;
  assign n44178 = n9346 & n44177 ;
  assign n44179 = n44178 ^ n44175 ^ n27466 ;
  assign n44180 = n10912 & ~n42457 ;
  assign n44181 = ~n22282 & n43686 ;
  assign n44182 = n16553 ^ n7919 ^ 1'b0 ;
  assign n44183 = n9902 & ~n21198 ;
  assign n44184 = n44183 ^ n30781 ^ 1'b0 ;
  assign n44185 = n21563 | n24062 ;
  assign n44186 = n13922 | n44185 ;
  assign n44187 = n44186 ^ n10860 ^ 1'b0 ;
  assign n44188 = ( n6805 & n25942 ) | ( n6805 & ~n31339 ) | ( n25942 & ~n31339 ) ;
  assign n44189 = n44188 ^ n1849 ^ 1'b0 ;
  assign n44190 = n5807 & ~n31767 ;
  assign n44191 = ~n13484 & n44190 ;
  assign n44196 = n19889 & n25444 ;
  assign n44195 = ( n270 & n9234 ) | ( n270 & n29998 ) | ( n9234 & n29998 ) ;
  assign n44192 = n3541 & n4801 ;
  assign n44193 = ~n13081 & n44192 ;
  assign n44194 = n44193 ^ n38087 ^ 1'b0 ;
  assign n44197 = n44196 ^ n44195 ^ n44194 ;
  assign n44198 = n34084 ^ n33864 ^ n15237 ;
  assign n44199 = n40547 | n41587 ;
  assign n44200 = ( n1592 & n13262 ) | ( n1592 & ~n13499 ) | ( n13262 & ~n13499 ) ;
  assign n44201 = n44200 ^ n23131 ^ n9752 ;
  assign n44202 = n5897 | n19897 ;
  assign n44203 = n44202 ^ x212 ^ 1'b0 ;
  assign n44204 = n33831 & ~n44203 ;
  assign n44205 = n3389 ^ n1240 ^ 1'b0 ;
  assign n44206 = n25179 & n44205 ;
  assign n44207 = n43175 ^ x54 ^ 1'b0 ;
  assign n44208 = ~n24387 & n44207 ;
  assign n44209 = x110 & n14999 ;
  assign n44210 = x249 & ~n44209 ;
  assign n44211 = n44210 ^ n24784 ^ 1'b0 ;
  assign n44212 = ~n7910 & n44211 ;
  assign n44213 = ~n7995 & n39104 ;
  assign n44214 = n15292 & n44213 ;
  assign n44215 = n6718 | n44214 ;
  assign n44216 = n37118 ^ n28485 ^ 1'b0 ;
  assign n44217 = ( ~n12898 & n44215 ) | ( ~n12898 & n44216 ) | ( n44215 & n44216 ) ;
  assign n44218 = n44217 ^ n11037 ^ 1'b0 ;
  assign n44219 = n14136 & ~n44218 ;
  assign n44220 = n6084 | n8563 ;
  assign n44221 = n40974 ^ n31926 ^ 1'b0 ;
  assign n44222 = n10518 & n18531 ;
  assign n44223 = ( n6507 & n19192 ) | ( n6507 & ~n44222 ) | ( n19192 & ~n44222 ) ;
  assign n44224 = n44223 ^ n29132 ^ n5899 ;
  assign n44225 = n11020 & n41169 ;
  assign n44226 = n9101 | n44225 ;
  assign n44227 = ( n8865 & ~n39339 ) | ( n8865 & n44226 ) | ( ~n39339 & n44226 ) ;
  assign n44228 = n10247 | n18256 ;
  assign n44229 = n44228 ^ n33044 ^ 1'b0 ;
  assign n44230 = n13502 | n13721 ;
  assign n44231 = n23055 | n44230 ;
  assign n44236 = n39303 ^ n12378 ^ n1288 ;
  assign n44237 = n9918 & ~n44236 ;
  assign n44238 = n44237 ^ n37864 ^ 1'b0 ;
  assign n44235 = n4797 & ~n7887 ;
  assign n44232 = n33252 ^ n13068 ^ 1'b0 ;
  assign n44233 = n37439 & n44232 ;
  assign n44234 = n44233 ^ n37148 ^ n6008 ;
  assign n44239 = n44238 ^ n44235 ^ n44234 ;
  assign n44240 = n4449 & n33313 ;
  assign n44241 = n27485 & n44240 ;
  assign n44242 = ( n3020 & n20544 ) | ( n3020 & n44241 ) | ( n20544 & n44241 ) ;
  assign n44243 = n25005 ^ n21146 ^ n12239 ;
  assign n44244 = n37882 ^ n27981 ^ 1'b0 ;
  assign n44245 = n44243 | n44244 ;
  assign n44247 = n21538 ^ n10932 ^ 1'b0 ;
  assign n44248 = n44247 ^ n39020 ^ n19260 ;
  assign n44246 = ~n15171 & n36927 ;
  assign n44249 = n44248 ^ n44246 ^ 1'b0 ;
  assign n44250 = ~n7522 & n17961 ;
  assign n44251 = n39478 ^ n30531 ^ 1'b0 ;
  assign n44252 = n15430 & ~n44251 ;
  assign n44253 = n29957 ^ n7087 ^ n3296 ;
  assign n44254 = n5662 & ~n22357 ;
  assign n44255 = ( n21753 & n44253 ) | ( n21753 & n44254 ) | ( n44253 & n44254 ) ;
  assign n44256 = n25937 ^ n22306 ^ n440 ;
  assign n44257 = ( n21063 & ~n22349 ) | ( n21063 & n38050 ) | ( ~n22349 & n38050 ) ;
  assign n44258 = n17313 & n36441 ;
  assign n44259 = n32751 & ~n44258 ;
  assign n44260 = n32994 & n44259 ;
  assign n44261 = n16284 ^ n11424 ^ 1'b0 ;
  assign n44262 = n10601 ^ n6737 ^ 1'b0 ;
  assign n44263 = ~n5466 & n44262 ;
  assign n44264 = ~n3093 & n44263 ;
  assign n44265 = n44264 ^ n32898 ^ 1'b0 ;
  assign n44266 = n2140 | n42658 ;
  assign n44267 = n44265 | n44266 ;
  assign n44269 = ~n5484 & n10573 ;
  assign n44270 = n44269 ^ n21661 ^ 1'b0 ;
  assign n44271 = n22608 & n44270 ;
  assign n44268 = n10052 & ~n20319 ;
  assign n44272 = n44271 ^ n44268 ^ 1'b0 ;
  assign n44275 = n3389 | n5686 ;
  assign n44273 = n37553 ^ n14050 ^ 1'b0 ;
  assign n44274 = n23666 & n44273 ;
  assign n44276 = n44275 ^ n44274 ^ n18182 ;
  assign n44277 = n24186 & n29888 ;
  assign n44278 = n21340 & ~n32111 ;
  assign n44279 = n2608 & ~n33637 ;
  assign n44280 = n23742 & n44279 ;
  assign n44281 = n1185 & n44280 ;
  assign n44282 = n44281 ^ n30367 ^ 1'b0 ;
  assign n44283 = ~n22821 & n44282 ;
  assign n44284 = n2266 & n3233 ;
  assign n44285 = n44284 ^ n25656 ^ 1'b0 ;
  assign n44286 = ~n6338 & n44285 ;
  assign n44287 = ~n6051 & n44286 ;
  assign n44288 = ~n1318 & n7184 ;
  assign n44289 = ~n4889 & n18197 ;
  assign n44290 = n10801 & ~n44289 ;
  assign n44291 = x53 & n5825 ;
  assign n44292 = n44290 & n44291 ;
  assign n44293 = n2735 | n4752 ;
  assign n44294 = n4752 & ~n44293 ;
  assign n44295 = ~n1034 & n3864 ;
  assign n44296 = n1034 & n44295 ;
  assign n44297 = n44296 ^ n16738 ^ 1'b0 ;
  assign n44298 = ~n44294 & n44297 ;
  assign n44299 = n32009 ^ n3740 ^ 1'b0 ;
  assign n44300 = n20924 & ~n44299 ;
  assign n44301 = n44298 & n44300 ;
  assign n44302 = n11099 ^ n10663 ^ 1'b0 ;
  assign n44303 = ( n6605 & ~n26049 ) | ( n6605 & n44302 ) | ( ~n26049 & n44302 ) ;
  assign n44304 = ( n4743 & n23631 ) | ( n4743 & ~n33209 ) | ( n23631 & ~n33209 ) ;
  assign n44305 = n29448 ^ n668 ^ 1'b0 ;
  assign n44306 = ( n15610 & ~n33173 ) | ( n15610 & n44305 ) | ( ~n33173 & n44305 ) ;
  assign n44307 = n37274 ^ n17963 ^ 1'b0 ;
  assign n44308 = n11536 & ~n44307 ;
  assign n44309 = n774 & n9222 ;
  assign n44310 = ~n44308 & n44309 ;
  assign n44311 = n33060 ^ n18924 ^ n11283 ;
  assign n44312 = n44311 ^ n33198 ^ 1'b0 ;
  assign n44313 = ~n1422 & n37790 ;
  assign n44314 = n12342 & ~n44313 ;
  assign n44315 = n1236 | n10543 ;
  assign n44316 = n44315 ^ n15169 ^ 1'b0 ;
  assign n44317 = n3100 | n4587 ;
  assign n44318 = n44317 ^ n17603 ^ 1'b0 ;
  assign n44319 = n9447 & ~n44318 ;
  assign n44320 = n44319 ^ n16264 ^ 1'b0 ;
  assign n44321 = ~n7639 & n13281 ;
  assign n44322 = n44321 ^ n10056 ^ 1'b0 ;
  assign n44323 = n44322 ^ n21029 ^ 1'b0 ;
  assign n44324 = ~n11837 & n42616 ;
  assign n44325 = n44324 ^ n17279 ^ 1'b0 ;
  assign n44326 = ( ~n6515 & n13604 ) | ( ~n6515 & n44325 ) | ( n13604 & n44325 ) ;
  assign n44327 = n40369 ^ n11322 ^ 1'b0 ;
  assign n44328 = n10220 ^ n1795 ^ 1'b0 ;
  assign n44329 = n41429 ^ n9185 ^ 1'b0 ;
  assign n44330 = n18825 ^ n15180 ^ n5863 ;
  assign n44331 = ~n21361 & n44330 ;
  assign n44332 = n44331 ^ n19129 ^ 1'b0 ;
  assign n44333 = n27840 & n44332 ;
  assign n44334 = n24681 ^ n3614 ^ 1'b0 ;
  assign n44335 = n35951 & n44334 ;
  assign n44336 = n36725 ^ n23754 ^ 1'b0 ;
  assign n44337 = n44335 & n44336 ;
  assign n44339 = n16908 & n18560 ;
  assign n44340 = ( n4080 & n4381 ) | ( n4080 & ~n44339 ) | ( n4381 & ~n44339 ) ;
  assign n44338 = n6821 ^ n4001 ^ 1'b0 ;
  assign n44341 = n44340 ^ n44338 ^ n2885 ;
  assign n44342 = n22216 ^ n3302 ^ 1'b0 ;
  assign n44343 = n5103 | n44342 ;
  assign n44344 = n44343 ^ n17587 ^ 1'b0 ;
  assign n44347 = n10358 | n21570 ;
  assign n44345 = n20127 ^ n18575 ^ 1'b0 ;
  assign n44346 = n5044 & ~n44345 ;
  assign n44348 = n44347 ^ n44346 ^ 1'b0 ;
  assign n44349 = n44348 ^ n43455 ^ n9447 ;
  assign n44350 = n27921 ^ n18143 ^ 1'b0 ;
  assign n44351 = n25180 & ~n44350 ;
  assign n44352 = n44351 ^ n10370 ^ n3130 ;
  assign n44353 = n3052 | n30546 ;
  assign n44354 = n35385 | n44353 ;
  assign n44355 = n12842 & ~n44354 ;
  assign n44356 = n8919 | n21761 ;
  assign n44357 = n5929 | n19216 ;
  assign n44358 = n24092 & ~n31772 ;
  assign n44359 = n4404 | n44358 ;
  assign n44360 = n44359 ^ n16221 ^ 1'b0 ;
  assign n44361 = ~n26352 & n38457 ;
  assign n44362 = n20142 & ~n34330 ;
  assign n44363 = n18797 & n44362 ;
  assign n44366 = n10963 | n17001 ;
  assign n44364 = n30641 ^ n3991 ^ 1'b0 ;
  assign n44365 = n44364 ^ n30958 ^ 1'b0 ;
  assign n44367 = n44366 ^ n44365 ^ n26203 ;
  assign n44368 = n42057 ^ n23367 ^ n1781 ;
  assign n44369 = n42333 ^ n21331 ^ 1'b0 ;
  assign n44370 = n6296 & ~n32674 ;
  assign n44371 = ( n11414 & n21204 ) | ( n11414 & n33934 ) | ( n21204 & n33934 ) ;
  assign n44372 = ( n44281 & n44370 ) | ( n44281 & n44371 ) | ( n44370 & n44371 ) ;
  assign n44373 = ( n2299 & n36840 ) | ( n2299 & ~n44372 ) | ( n36840 & ~n44372 ) ;
  assign n44374 = n27732 & n43567 ;
  assign n44375 = n44374 ^ n26711 ^ 1'b0 ;
  assign n44376 = ~n1486 & n11861 ;
  assign n44377 = n11880 ^ n11861 ^ n6822 ;
  assign n44378 = ~n3591 & n44377 ;
  assign n44379 = n2204 & ~n35107 ;
  assign n44380 = n44378 & n44379 ;
  assign n44381 = n9382 | n20119 ;
  assign n44382 = n620 | n44381 ;
  assign n44383 = n40369 & ~n44382 ;
  assign n44384 = n15955 ^ n13893 ^ 1'b0 ;
  assign n44385 = ~n22832 & n44384 ;
  assign n44386 = ~n15214 & n44385 ;
  assign n44387 = n6284 & n44386 ;
  assign n44388 = n21543 ^ n9011 ^ 1'b0 ;
  assign n44389 = n22355 & n44388 ;
  assign n44390 = ( n35522 & n40087 ) | ( n35522 & ~n44389 ) | ( n40087 & ~n44389 ) ;
  assign n44391 = ( ~n3820 & n15714 ) | ( ~n3820 & n36923 ) | ( n15714 & n36923 ) ;
  assign n44392 = ( ~n17592 & n18963 ) | ( ~n17592 & n23950 ) | ( n18963 & n23950 ) ;
  assign n44393 = n44392 ^ n42847 ^ 1'b0 ;
  assign n44394 = n11113 & ~n25975 ;
  assign n44395 = ~n16034 & n34397 ;
  assign n44396 = n16580 & n34295 ;
  assign n44397 = n44396 ^ n16510 ^ 1'b0 ;
  assign n44398 = n43019 & ~n44397 ;
  assign n44399 = n22951 ^ n10016 ^ 1'b0 ;
  assign n44400 = n23265 ^ n15132 ^ 1'b0 ;
  assign n44401 = ~n44399 & n44400 ;
  assign n44402 = x234 & ~n22150 ;
  assign n44403 = n44402 ^ n675 ^ 1'b0 ;
  assign n44404 = n1035 & n13506 ;
  assign n44405 = n38195 ^ n35582 ^ n7055 ;
  assign n44406 = n19264 | n25855 ;
  assign n44407 = n44405 | n44406 ;
  assign n44408 = n37761 ^ n24568 ^ 1'b0 ;
  assign n44409 = ( ~n1830 & n2682 ) | ( ~n1830 & n19321 ) | ( n2682 & n19321 ) ;
  assign n44410 = n44409 ^ n15953 ^ n6459 ;
  assign n44411 = n17394 & ~n30134 ;
  assign n44412 = n32084 ^ n14721 ^ 1'b0 ;
  assign n44413 = ~n14370 & n44412 ;
  assign n44414 = n37916 ^ n15123 ^ 1'b0 ;
  assign n44415 = n3583 ^ x25 ^ 1'b0 ;
  assign n44416 = ( ~n11279 & n21166 ) | ( ~n11279 & n44415 ) | ( n21166 & n44415 ) ;
  assign n44417 = n44416 ^ n21574 ^ 1'b0 ;
  assign n44418 = ( n14743 & ~n27906 ) | ( n14743 & n35852 ) | ( ~n27906 & n35852 ) ;
  assign n44419 = n44418 ^ n6571 ^ 1'b0 ;
  assign n44420 = n36414 & ~n44419 ;
  assign n44421 = n12210 & n12614 ;
  assign n44422 = n44421 ^ n24239 ^ 1'b0 ;
  assign n44423 = n10342 & ~n18359 ;
  assign n44424 = n806 & n14703 ;
  assign n44425 = n9408 ^ n8781 ^ n516 ;
  assign n44426 = ( n2293 & n44424 ) | ( n2293 & n44425 ) | ( n44424 & n44425 ) ;
  assign n44427 = n7027 & ~n44426 ;
  assign n44428 = ~n40566 & n44427 ;
  assign n44429 = ~n5377 & n35392 ;
  assign n44430 = n20831 ^ n11391 ^ 1'b0 ;
  assign n44431 = n44429 & ~n44430 ;
  assign n44432 = n39459 ^ n18522 ^ n9545 ;
  assign n44433 = n3724 & ~n14107 ;
  assign n44434 = n21316 & n44433 ;
  assign n44435 = n10375 & ~n44434 ;
  assign n44436 = ( ~n24438 & n32032 ) | ( ~n24438 & n44435 ) | ( n32032 & n44435 ) ;
  assign n44437 = n2984 & ~n5076 ;
  assign n44438 = n44437 ^ n13306 ^ 1'b0 ;
  assign n44439 = n22053 & n44438 ;
  assign n44440 = n44439 ^ n29135 ^ 1'b0 ;
  assign n44441 = n44440 ^ n13538 ^ 1'b0 ;
  assign n44443 = n25498 ^ n12885 ^ 1'b0 ;
  assign n44444 = n13327 | n44443 ;
  assign n44442 = n30275 | n42319 ;
  assign n44445 = n44444 ^ n44442 ^ 1'b0 ;
  assign n44446 = x141 & ~n23517 ;
  assign n44447 = ~n15423 & n44446 ;
  assign n44448 = ~n6143 & n44447 ;
  assign n44449 = n14619 ^ n14295 ^ 1'b0 ;
  assign n44450 = n16625 ^ n7782 ^ 1'b0 ;
  assign n44451 = n44449 & n44450 ;
  assign n44452 = n7832 ^ n5453 ^ 1'b0 ;
  assign n44453 = ( n557 & n6976 ) | ( n557 & ~n33915 ) | ( n6976 & ~n33915 ) ;
  assign n44454 = n2767 ^ n1922 ^ 1'b0 ;
  assign n44455 = n27772 | n44454 ;
  assign n44456 = ( ~n2804 & n42488 ) | ( ~n2804 & n44455 ) | ( n42488 & n44455 ) ;
  assign n44457 = n4405 & n33104 ;
  assign n44458 = ~n4756 & n44457 ;
  assign n44459 = n22449 & ~n44458 ;
  assign n44460 = n11242 & n44459 ;
  assign n44461 = n3444 | n10794 ;
  assign n44462 = n44461 ^ n30327 ^ 1'b0 ;
  assign n44465 = n38879 ^ n14785 ^ 1'b0 ;
  assign n44463 = ( n2875 & n15329 ) | ( n2875 & ~n20634 ) | ( n15329 & ~n20634 ) ;
  assign n44464 = n19955 & ~n44463 ;
  assign n44466 = n44465 ^ n44464 ^ 1'b0 ;
  assign n44467 = n1332 | n17372 ;
  assign n44468 = n5781 & ~n44467 ;
  assign n44469 = n7435 & ~n12471 ;
  assign n44470 = ( ~n2238 & n10193 ) | ( ~n2238 & n12359 ) | ( n10193 & n12359 ) ;
  assign n44471 = ( n35222 & ~n44469 ) | ( n35222 & n44470 ) | ( ~n44469 & n44470 ) ;
  assign n44472 = n3353 & n18121 ;
  assign n44473 = n44472 ^ n17542 ^ n16653 ;
  assign n44474 = n43814 ^ n29894 ^ 1'b0 ;
  assign n44475 = ~n16844 & n41290 ;
  assign n44476 = n44475 ^ n15104 ^ 1'b0 ;
  assign n44477 = n32080 ^ n1347 ^ 1'b0 ;
  assign n44478 = n19874 & ~n44477 ;
  assign n44479 = n33967 ^ n13007 ^ 1'b0 ;
  assign n44480 = n44478 & n44479 ;
  assign n44481 = n15650 ^ n12410 ^ 1'b0 ;
  assign n44482 = n12959 & n20410 ;
  assign n44483 = n8584 | n44482 ;
  assign n44484 = n44483 ^ n43565 ^ n35097 ;
  assign n44485 = ( n6342 & n12700 ) | ( n6342 & n38485 ) | ( n12700 & n38485 ) ;
  assign n44486 = n35860 ^ n34891 ^ 1'b0 ;
  assign n44487 = n8755 & n25373 ;
  assign n44488 = ( n2908 & n44486 ) | ( n2908 & ~n44487 ) | ( n44486 & ~n44487 ) ;
  assign n44489 = n690 & ~n13353 ;
  assign n44490 = ~n9359 & n44489 ;
  assign n44491 = ~n13629 & n44490 ;
  assign n44492 = n30140 ^ n12841 ^ 1'b0 ;
  assign n44493 = n10777 | n44138 ;
  assign n44494 = n8197 & ~n32006 ;
  assign n44495 = n31382 ^ n13583 ^ 1'b0 ;
  assign n44496 = n30882 & ~n44495 ;
  assign n44497 = n15195 ^ n7915 ^ 1'b0 ;
  assign n44498 = n2951 & n4523 ;
  assign n44499 = n44498 ^ n17621 ^ 1'b0 ;
  assign n44500 = ( n11181 & ~n38906 ) | ( n11181 & n44458 ) | ( ~n38906 & n44458 ) ;
  assign n44502 = n26452 ^ n6221 ^ 1'b0 ;
  assign n44501 = n5602 & ~n33361 ;
  assign n44503 = n44502 ^ n44501 ^ 1'b0 ;
  assign n44504 = n15001 | n18268 ;
  assign n44505 = n44503 | n44504 ;
  assign n44506 = n1285 & ~n28899 ;
  assign n44507 = n3170 ^ x62 ^ 1'b0 ;
  assign n44508 = n30789 & n44507 ;
  assign n44509 = n5173 | n26635 ;
  assign n44510 = ( n12817 & ~n33541 ) | ( n12817 & n37565 ) | ( ~n33541 & n37565 ) ;
  assign n44511 = n38259 ^ n13515 ^ 1'b0 ;
  assign n44512 = n4912 & n21249 ;
  assign n44513 = n15359 | n44512 ;
  assign n44514 = n44513 ^ n42072 ^ n19874 ;
  assign n44515 = n29516 ^ n6048 ^ 1'b0 ;
  assign n44516 = ( ~n11875 & n13135 ) | ( ~n11875 & n44515 ) | ( n13135 & n44515 ) ;
  assign n44517 = n24934 ^ n8502 ^ 1'b0 ;
  assign n44518 = n4963 | n31811 ;
  assign n44519 = n4854 | n13407 ;
  assign n44520 = n43343 ^ n42459 ^ 1'b0 ;
  assign n44521 = n23077 | n42886 ;
  assign n44523 = n5377 | n23694 ;
  assign n44522 = n2577 | n13981 ;
  assign n44524 = n44523 ^ n44522 ^ 1'b0 ;
  assign n44525 = n3426 | n8422 ;
  assign n44535 = n16241 | n43807 ;
  assign n44527 = n5803 & ~n13252 ;
  assign n44528 = n13252 & n44527 ;
  assign n44529 = n9831 | n44528 ;
  assign n44530 = n44529 ^ n27689 ^ 1'b0 ;
  assign n44531 = n31769 | n44530 ;
  assign n44532 = n44531 ^ n2260 ^ 1'b0 ;
  assign n44533 = n44532 ^ n2297 ^ 1'b0 ;
  assign n44526 = ( n1661 & n18234 ) | ( n1661 & ~n28997 ) | ( n18234 & ~n28997 ) ;
  assign n44534 = n44533 ^ n44526 ^ 1'b0 ;
  assign n44536 = n44535 ^ n44534 ^ n4395 ;
  assign n44537 = n39880 ^ n28142 ^ 1'b0 ;
  assign n44538 = n12153 & ~n44537 ;
  assign n44539 = n12842 ^ n4405 ^ 1'b0 ;
  assign n44540 = n40908 ^ n19964 ^ n5550 ;
  assign n44541 = n43978 ^ n15096 ^ 1'b0 ;
  assign n44542 = n44541 ^ n36413 ^ n16012 ;
  assign n44543 = n44542 ^ n18968 ^ 1'b0 ;
  assign n44544 = ~n44540 & n44543 ;
  assign n44545 = n44544 ^ n5763 ^ 1'b0 ;
  assign n44546 = n41987 ^ n7135 ^ 1'b0 ;
  assign n44547 = n44545 & ~n44546 ;
  assign n44548 = ( x96 & ~n9428 ) | ( x96 & n29319 ) | ( ~n9428 & n29319 ) ;
  assign n44549 = n5833 ^ n3027 ^ 1'b0 ;
  assign n44550 = n44548 & ~n44549 ;
  assign n44551 = n43209 ^ n16605 ^ 1'b0 ;
  assign n44552 = ( ~n12865 & n13523 ) | ( ~n12865 & n16431 ) | ( n13523 & n16431 ) ;
  assign n44553 = n44552 ^ n7215 ^ 1'b0 ;
  assign n44554 = n10368 & n27655 ;
  assign n44555 = n44554 ^ n23236 ^ 1'b0 ;
  assign n44556 = n37325 ^ n7990 ^ 1'b0 ;
  assign n44557 = n9683 | n44556 ;
  assign n44558 = n44557 ^ n20857 ^ n4154 ;
  assign n44559 = n44558 ^ n27643 ^ 1'b0 ;
  assign n44560 = n15098 | n21892 ;
  assign n44561 = ( ~n14827 & n37237 ) | ( ~n14827 & n44560 ) | ( n37237 & n44560 ) ;
  assign n44562 = ( n3261 & n16751 ) | ( n3261 & ~n19379 ) | ( n16751 & ~n19379 ) ;
  assign n44563 = n44562 ^ n19632 ^ 1'b0 ;
  assign n44564 = ~n44561 & n44563 ;
  assign n44565 = ~n4273 & n34398 ;
  assign n44566 = ~n44564 & n44565 ;
  assign n44567 = n13786 ^ n264 ^ 1'b0 ;
  assign n44568 = n7535 & n10275 ;
  assign n44569 = n44568 ^ n5813 ^ n2642 ;
  assign n44570 = n5827 ^ n2991 ^ 1'b0 ;
  assign n44571 = n1736 | n44570 ;
  assign n44572 = n44571 ^ n17610 ^ n5165 ;
  assign n44573 = n7689 ^ n6558 ^ 1'b0 ;
  assign n44574 = n9694 & ~n44573 ;
  assign n44575 = ( n3173 & ~n12929 ) | ( n3173 & n44574 ) | ( ~n12929 & n44574 ) ;
  assign n44576 = ~n16378 & n44575 ;
  assign n44577 = ( n438 & n44572 ) | ( n438 & n44576 ) | ( n44572 & n44576 ) ;
  assign n44578 = ( n13102 & n30384 ) | ( n13102 & n34735 ) | ( n30384 & n34735 ) ;
  assign n44579 = n17481 ^ n6924 ^ n5947 ;
  assign n44580 = n30243 ^ n20883 ^ 1'b0 ;
  assign n44581 = n44579 & n44580 ;
  assign n44582 = ~n33025 & n44581 ;
  assign n44583 = ~n31402 & n44582 ;
  assign n44584 = n44583 ^ n40756 ^ n38187 ;
  assign n44585 = n417 & ~n9386 ;
  assign n44586 = ~n2110 & n44585 ;
  assign n44587 = n16311 & ~n27127 ;
  assign n44588 = ~n4958 & n44587 ;
  assign n44589 = n22953 | n25049 ;
  assign n44590 = n44589 ^ n3029 ^ 1'b0 ;
  assign n44591 = n9032 ^ n8806 ^ n1481 ;
  assign n44592 = n23367 & n44591 ;
  assign n44593 = n11064 ^ x22 ^ 1'b0 ;
  assign n44594 = n3775 & n44593 ;
  assign n44595 = n17598 | n25209 ;
  assign n44596 = n44594 | n44595 ;
  assign n44597 = ~n5349 & n44596 ;
  assign n44598 = n44597 ^ n7900 ^ 1'b0 ;
  assign n44599 = n7260 ^ n4572 ^ 1'b0 ;
  assign n44600 = n4084 & n44599 ;
  assign n44601 = n44600 ^ n1769 ^ 1'b0 ;
  assign n44602 = n5259 & ~n24837 ;
  assign n44605 = n19627 ^ n13104 ^ 1'b0 ;
  assign n44606 = n3710 | n44605 ;
  assign n44603 = n1527 & n22355 ;
  assign n44604 = n44603 ^ n35960 ^ 1'b0 ;
  assign n44607 = n44606 ^ n44604 ^ n11449 ;
  assign n44608 = n16209 & n21181 ;
  assign n44609 = ~n5942 & n44608 ;
  assign n44610 = n11921 & n43153 ;
  assign n44611 = n43338 ^ n17840 ^ 1'b0 ;
  assign n44612 = n28955 | n44611 ;
  assign n44613 = n38507 ^ n34832 ^ 1'b0 ;
  assign n44615 = n12029 & n21723 ;
  assign n44614 = ( ~n6310 & n25732 ) | ( ~n6310 & n27841 ) | ( n25732 & n27841 ) ;
  assign n44616 = n44615 ^ n44614 ^ n3745 ;
  assign n44617 = n21274 | n25762 ;
  assign n44618 = n1552 & ~n14055 ;
  assign n44619 = n44618 ^ n16104 ^ 1'b0 ;
  assign n44620 = n23706 ^ n9165 ^ n8655 ;
  assign n44621 = ( n41924 & n44619 ) | ( n41924 & n44620 ) | ( n44619 & n44620 ) ;
  assign n44622 = n12072 & n17826 ;
  assign n44623 = n16317 | n44622 ;
  assign n44624 = n15246 ^ n5055 ^ 1'b0 ;
  assign n44625 = n3315 & ~n44624 ;
  assign n44626 = n27876 ^ n6053 ^ 1'b0 ;
  assign n44627 = n4537 & ~n31716 ;
  assign n44628 = n26403 ^ n12859 ^ 1'b0 ;
  assign n44629 = n10894 | n44628 ;
  assign n44630 = ~n11972 & n34364 ;
  assign n44631 = ( n944 & n994 ) | ( n944 & n44630 ) | ( n994 & n44630 ) ;
  assign n44632 = ( n5589 & ~n38777 ) | ( n5589 & n44631 ) | ( ~n38777 & n44631 ) ;
  assign n44633 = n23755 ^ n19614 ^ n12231 ;
  assign n44634 = n21357 & ~n44633 ;
  assign n44635 = n34613 & n44634 ;
  assign n44636 = n44635 ^ n8851 ^ 1'b0 ;
  assign n44637 = ( n2724 & n24013 ) | ( n2724 & n44636 ) | ( n24013 & n44636 ) ;
  assign n44641 = ( n6728 & ~n6750 ) | ( n6728 & n44067 ) | ( ~n6750 & n44067 ) ;
  assign n44642 = n40842 & n44641 ;
  assign n44640 = n10959 & n29027 ;
  assign n44638 = n20416 ^ n5675 ^ 1'b0 ;
  assign n44639 = ~n14785 & n44638 ;
  assign n44643 = n44642 ^ n44640 ^ n44639 ;
  assign n44644 = n10318 & n12356 ;
  assign n44645 = n44644 ^ n15686 ^ 1'b0 ;
  assign n44646 = n25392 ^ n5039 ^ 1'b0 ;
  assign n44647 = n3389 & n5781 ;
  assign n44648 = n5376 ^ x235 ^ 1'b0 ;
  assign n44654 = n2750 | n5020 ;
  assign n44653 = n24518 ^ n6272 ^ n1829 ;
  assign n44649 = n23301 ^ n9344 ^ 1'b0 ;
  assign n44650 = n15629 & ~n44649 ;
  assign n44651 = ( n10927 & n26916 ) | ( n10927 & n44650 ) | ( n26916 & n44650 ) ;
  assign n44652 = n44651 ^ n27101 ^ n26376 ;
  assign n44655 = n44654 ^ n44653 ^ n44652 ;
  assign n44656 = ~n12818 & n22168 ;
  assign n44657 = n35559 ^ n15108 ^ n6776 ;
  assign n44658 = n7843 ^ n2523 ^ 1'b0 ;
  assign n44659 = n4795 & n44658 ;
  assign n44660 = n1383 & n44659 ;
  assign n44661 = n13587 & n15893 ;
  assign n44662 = n14677 & n44661 ;
  assign n44663 = n36430 | n44662 ;
  assign n44664 = n31843 | n44663 ;
  assign n44665 = n23581 | n29380 ;
  assign n44666 = n44665 ^ n23427 ^ 1'b0 ;
  assign n44667 = n40304 ^ n4550 ^ 1'b0 ;
  assign n44668 = ( n3029 & n41879 ) | ( n3029 & ~n42209 ) | ( n41879 & ~n42209 ) ;
  assign n44669 = ~n6176 & n8900 ;
  assign n44670 = n14422 | n16867 ;
  assign n44671 = n19875 & ~n44670 ;
  assign n44672 = n12850 & ~n44671 ;
  assign n44673 = n12133 & ~n14370 ;
  assign n44674 = n44673 ^ n29507 ^ 1'b0 ;
  assign n44675 = n3620 | n44674 ;
  assign n44676 = n44675 ^ n29206 ^ 1'b0 ;
  assign n44677 = n22265 ^ n7066 ^ 1'b0 ;
  assign n44678 = n18138 & ~n44677 ;
  assign n44679 = n31733 & ~n37526 ;
  assign n44680 = n11066 & n44679 ;
  assign n44681 = n7199 & ~n33134 ;
  assign n44682 = n41569 ^ n12863 ^ 1'b0 ;
  assign n44683 = n44681 & n44682 ;
  assign n44684 = n952 & ~n1938 ;
  assign n44685 = n633 ^ n632 ^ 1'b0 ;
  assign n44686 = n34967 ^ n10634 ^ n3233 ;
  assign n44687 = n30633 & ~n44686 ;
  assign n44689 = n12520 ^ n8678 ^ n6509 ;
  assign n44688 = n8228 | n20449 ;
  assign n44690 = n44689 ^ n44688 ^ 1'b0 ;
  assign n44691 = n1667 & n3674 ;
  assign n44692 = ~n22916 & n44691 ;
  assign n44693 = n44692 ^ n8491 ^ 1'b0 ;
  assign n44694 = ~n32336 & n44693 ;
  assign n44695 = n29112 ^ n14288 ^ 1'b0 ;
  assign n44696 = ~n27749 & n44695 ;
  assign n44697 = n14559 ^ n12938 ^ 1'b0 ;
  assign n44698 = n29252 | n42090 ;
  assign n44699 = n16521 | n44698 ;
  assign n44700 = n3960 & n31462 ;
  assign n44701 = n44700 ^ n31262 ^ 1'b0 ;
  assign n44702 = n28795 ^ n23431 ^ 1'b0 ;
  assign n44703 = ~n13494 & n17381 ;
  assign n44704 = n2701 & n44703 ;
  assign n44705 = ( x196 & ~n29666 ) | ( x196 & n44633 ) | ( ~n29666 & n44633 ) ;
  assign n44706 = ~n44704 & n44705 ;
  assign n44707 = ~n4543 & n35310 ;
  assign n44708 = n27711 ^ n10173 ^ 1'b0 ;
  assign n44709 = n44707 & n44708 ;
  assign n44710 = n44709 ^ n12392 ^ 1'b0 ;
  assign n44711 = n16898 & ~n44710 ;
  assign n44712 = n2245 & n34610 ;
  assign n44713 = n3613 & n44712 ;
  assign n44714 = ( n4274 & ~n12203 ) | ( n4274 & n13363 ) | ( ~n12203 & n13363 ) ;
  assign n44715 = ~n21531 & n44714 ;
  assign n44716 = n41767 ^ n22199 ^ n19529 ;
  assign n44717 = ( ~n27690 & n30836 ) | ( ~n27690 & n44716 ) | ( n30836 & n44716 ) ;
  assign n44718 = n6620 | n12799 ;
  assign n44719 = n44718 ^ n40173 ^ 1'b0 ;
  assign n44720 = n12916 & ~n44719 ;
  assign n44721 = n44717 & n44720 ;
  assign n44722 = ~n28370 & n44721 ;
  assign n44723 = n10174 | n22256 ;
  assign n44724 = ( ~x17 & n28033 ) | ( ~x17 & n44723 ) | ( n28033 & n44723 ) ;
  assign n44727 = n3568 ^ x92 ^ 1'b0 ;
  assign n44726 = n5631 | n12617 ;
  assign n44728 = n44727 ^ n44726 ^ 1'b0 ;
  assign n44725 = n595 & ~n15022 ;
  assign n44729 = n44728 ^ n44725 ^ 1'b0 ;
  assign n44730 = ( n2779 & n22152 ) | ( n2779 & n39653 ) | ( n22152 & n39653 ) ;
  assign n44731 = ( n24501 & n44729 ) | ( n24501 & ~n44730 ) | ( n44729 & ~n44730 ) ;
  assign n44732 = n35040 ^ n1250 ^ 1'b0 ;
  assign n44733 = ( n3160 & ~n11020 ) | ( n3160 & n12354 ) | ( ~n11020 & n12354 ) ;
  assign n44734 = n44733 ^ n34632 ^ n23191 ;
  assign n44735 = n25599 & ~n28531 ;
  assign n44736 = n512 & ~n19897 ;
  assign n44737 = n18034 ^ n1895 ^ 1'b0 ;
  assign n44738 = n36606 & n44737 ;
  assign n44739 = x147 & n37518 ;
  assign n44740 = ~n11634 & n13648 ;
  assign n44741 = n44740 ^ n2613 ^ n1690 ;
  assign n44742 = n44741 ^ n31161 ^ 1'b0 ;
  assign n44743 = n42581 ^ n19015 ^ n17428 ;
  assign n44744 = n17071 ^ n3351 ^ n563 ;
  assign n44745 = n15652 & ~n15767 ;
  assign n44746 = n31103 & n44745 ;
  assign n44750 = n14827 | n15070 ;
  assign n44751 = n44750 ^ n44372 ^ 1'b0 ;
  assign n44752 = ~n5880 & n44751 ;
  assign n44747 = n1944 & ~n30501 ;
  assign n44748 = ~n3317 & n44747 ;
  assign n44749 = n38765 & ~n44748 ;
  assign n44753 = n44752 ^ n44749 ^ 1'b0 ;
  assign n44754 = n24013 ^ n11670 ^ 1'b0 ;
  assign n44755 = n4669 & n44754 ;
  assign n44756 = n22817 ^ n9572 ^ n2481 ;
  assign n44757 = n24487 & n44756 ;
  assign n44758 = n44757 ^ n9864 ^ 1'b0 ;
  assign n44759 = ~n20991 & n34576 ;
  assign n44760 = n44759 ^ n43352 ^ 1'b0 ;
  assign n44762 = n33411 & ~n42744 ;
  assign n44763 = n44762 ^ n10334 ^ 1'b0 ;
  assign n44764 = ~n5524 & n38325 ;
  assign n44765 = n44764 ^ n5337 ^ 1'b0 ;
  assign n44766 = n44765 ^ n6123 ^ 1'b0 ;
  assign n44767 = n44763 & ~n44766 ;
  assign n44761 = ~n2445 & n14576 ;
  assign n44768 = n44767 ^ n44761 ^ 1'b0 ;
  assign n44769 = n27199 & ~n37305 ;
  assign n44770 = ~n1326 & n44769 ;
  assign n44771 = n44770 ^ n13120 ^ 1'b0 ;
  assign n44772 = n44771 ^ n5464 ^ 1'b0 ;
  assign n44773 = ( n6345 & n32671 ) | ( n6345 & n44772 ) | ( n32671 & n44772 ) ;
  assign n44774 = n39420 ^ n18295 ^ 1'b0 ;
  assign n44775 = n17570 & ~n18735 ;
  assign n44776 = n30601 ^ n5077 ^ 1'b0 ;
  assign n44777 = n40727 ^ n31478 ^ 1'b0 ;
  assign n44779 = n9698 | n29550 ;
  assign n44778 = n28211 & n41100 ;
  assign n44780 = n44779 ^ n44778 ^ 1'b0 ;
  assign n44781 = n37701 ^ n33231 ^ n21816 ;
  assign n44784 = n14980 & n20005 ;
  assign n44785 = n6413 & n44784 ;
  assign n44782 = n4970 ^ n3654 ^ n1262 ;
  assign n44783 = ~n9379 & n44782 ;
  assign n44786 = n44785 ^ n44783 ^ n23055 ;
  assign n44787 = n40549 & ~n42801 ;
  assign n44788 = n17710 & n44787 ;
  assign n44789 = ( n3466 & ~n29568 ) | ( n3466 & n44788 ) | ( ~n29568 & n44788 ) ;
  assign n44791 = n27912 ^ n19574 ^ n4538 ;
  assign n44790 = n44727 ^ n21793 ^ 1'b0 ;
  assign n44792 = n44791 ^ n44790 ^ n38898 ;
  assign n44793 = n44792 ^ n7678 ^ n4367 ;
  assign n44794 = n371 & n32946 ;
  assign n44795 = ( n10160 & n23914 ) | ( n10160 & n24518 ) | ( n23914 & n24518 ) ;
  assign n44796 = ~n22496 & n32339 ;
  assign n44797 = n44795 & n44796 ;
  assign n44798 = n3487 | n18717 ;
  assign n44799 = n44798 ^ n1206 ^ 1'b0 ;
  assign n44800 = ~n24461 & n44799 ;
  assign n44801 = n37590 & n44800 ;
  assign n44802 = n25439 ^ n17072 ^ n14612 ;
  assign n44803 = n27626 ^ n7326 ^ 1'b0 ;
  assign n44804 = n9189 & n43537 ;
  assign n44805 = n16252 & n27620 ;
  assign n44806 = n17735 & n44805 ;
  assign n44807 = n42052 | n44806 ;
  assign n44808 = n748 & n17572 ;
  assign n44809 = ~n748 & n44808 ;
  assign n44810 = ~n3254 & n44809 ;
  assign n44811 = n27798 & n44810 ;
  assign n44812 = n320 & ~n8689 ;
  assign n44813 = n8689 & n44812 ;
  assign n44814 = ( ~n6073 & n10468 ) | ( ~n6073 & n44813 ) | ( n10468 & n44813 ) ;
  assign n44815 = n44814 ^ n8684 ^ 1'b0 ;
  assign n44816 = ~n44811 & n44815 ;
  assign n44817 = n44816 ^ n23455 ^ 1'b0 ;
  assign n44818 = n43978 ^ n7368 ^ n2321 ;
  assign n44819 = ~n4103 & n5366 ;
  assign n44820 = ~n44818 & n44819 ;
  assign n44821 = n4496 | n14779 ;
  assign n44822 = n1118 & n22147 ;
  assign n44824 = n21365 ^ n6999 ^ n2088 ;
  assign n44823 = n16743 | n16795 ;
  assign n44825 = n44824 ^ n44823 ^ 1'b0 ;
  assign n44826 = n5786 & n26524 ;
  assign n44827 = n44826 ^ n3621 ^ 1'b0 ;
  assign n44828 = n20908 ^ n6681 ^ 1'b0 ;
  assign n44829 = ( n15035 & ~n41133 ) | ( n15035 & n44828 ) | ( ~n41133 & n44828 ) ;
  assign n44830 = n19572 ^ n14487 ^ n12360 ;
  assign n44831 = n44830 ^ n29929 ^ n14413 ;
  assign n44832 = n33672 | n38628 ;
  assign n44833 = n7674 | n44832 ;
  assign n44834 = n27130 ^ n2857 ^ 1'b0 ;
  assign n44835 = ~n9154 & n44834 ;
  assign n44836 = ( ~n2059 & n4966 ) | ( ~n2059 & n9953 ) | ( n4966 & n9953 ) ;
  assign n44837 = ( n25485 & n27968 ) | ( n25485 & ~n44836 ) | ( n27968 & ~n44836 ) ;
  assign n44838 = ( n10028 & n18367 ) | ( n10028 & n20685 ) | ( n18367 & n20685 ) ;
  assign n44839 = ( n4655 & n10875 ) | ( n4655 & ~n15590 ) | ( n10875 & ~n15590 ) ;
  assign n44840 = n1934 | n31185 ;
  assign n44841 = ( n2998 & ~n28651 ) | ( n2998 & n44840 ) | ( ~n28651 & n44840 ) ;
  assign n44842 = n44841 ^ n26733 ^ 1'b0 ;
  assign n44843 = n26944 & ~n44842 ;
  assign n44844 = n3389 & n44843 ;
  assign n44845 = n7613 | n44844 ;
  assign n44846 = n42339 ^ n29933 ^ 1'b0 ;
  assign n44847 = n27381 & n44846 ;
  assign n44848 = n14404 & n41327 ;
  assign n44849 = n44848 ^ n24597 ^ 1'b0 ;
  assign n44850 = n19018 ^ n3589 ^ 1'b0 ;
  assign n44851 = n44850 ^ n17011 ^ 1'b0 ;
  assign n44852 = n38930 ^ n14867 ^ 1'b0 ;
  assign n44853 = n36782 ^ n27802 ^ n4516 ;
  assign n44854 = n22003 ^ n19486 ^ 1'b0 ;
  assign n44855 = n44853 & ~n44854 ;
  assign n44856 = n39513 ^ n3689 ^ 1'b0 ;
  assign n44857 = n13920 & ~n34119 ;
  assign n44858 = n8453 & n44857 ;
  assign n44859 = n36522 ^ n9308 ^ 1'b0 ;
  assign n44860 = ~n44858 & n44859 ;
  assign n44861 = ( ~n2932 & n44856 ) | ( ~n2932 & n44860 ) | ( n44856 & n44860 ) ;
  assign n44862 = ~n7810 & n13357 ;
  assign n44863 = n1933 | n16858 ;
  assign n44864 = n2118 | n7647 ;
  assign n44865 = n44863 | n44864 ;
  assign n44866 = n29650 | n44865 ;
  assign n44867 = n31066 ^ n29816 ^ n5245 ;
  assign n44868 = ( n7791 & n7887 ) | ( n7791 & ~n44867 ) | ( n7887 & ~n44867 ) ;
  assign n44869 = n7526 ^ n2610 ^ n369 ;
  assign n44870 = n33064 | n44869 ;
  assign n44871 = n31216 & n44870 ;
  assign n44872 = n1337 | n6134 ;
  assign n44873 = n11372 | n44872 ;
  assign n44874 = ~n557 & n669 ;
  assign n44875 = ( ~n17467 & n26554 ) | ( ~n17467 & n44874 ) | ( n26554 & n44874 ) ;
  assign n44876 = n44875 ^ n19819 ^ 1'b0 ;
  assign n44877 = ( n5707 & n8302 ) | ( n5707 & ~n44876 ) | ( n8302 & ~n44876 ) ;
  assign n44878 = n7077 & n8760 ;
  assign n44879 = ( n2149 & n10851 ) | ( n2149 & ~n27185 ) | ( n10851 & ~n27185 ) ;
  assign n44880 = n44879 ^ n26571 ^ 1'b0 ;
  assign n44881 = n3568 & ~n14847 ;
  assign n44882 = n44881 ^ n1797 ^ 1'b0 ;
  assign n44883 = n14086 & ~n14717 ;
  assign n44884 = n38634 ^ n28727 ^ 1'b0 ;
  assign n44885 = ~n27327 & n44884 ;
  assign n44886 = ~n5502 & n15121 ;
  assign n44887 = ~n4895 & n44886 ;
  assign n44888 = n34187 | n44887 ;
  assign n44889 = n2962 & ~n26173 ;
  assign n44890 = ~n10371 & n44889 ;
  assign n44891 = n13503 & ~n44890 ;
  assign n44892 = n4554 ^ n4300 ^ 1'b0 ;
  assign n44893 = n4807 | n8742 ;
  assign n44894 = n44893 ^ n32243 ^ n8909 ;
  assign n44895 = n38901 ^ n19823 ^ n1604 ;
  assign n44896 = n23188 & n30808 ;
  assign n44897 = n27193 ^ n1048 ^ 1'b0 ;
  assign n44898 = n21227 | n23660 ;
  assign n44899 = n5754 ^ n1847 ^ 1'b0 ;
  assign n44900 = ~n44898 & n44899 ;
  assign n44901 = n44328 ^ n36752 ^ 1'b0 ;
  assign n44902 = ~n20219 & n44901 ;
  assign n44903 = n36818 | n38656 ;
  assign n44904 = n44903 ^ n17104 ^ 1'b0 ;
  assign n44905 = ~n9746 & n18094 ;
  assign n44906 = n27633 & ~n44905 ;
  assign n44907 = n17388 ^ n12102 ^ n9433 ;
  assign n44908 = n44907 ^ n28044 ^ n4705 ;
  assign n44913 = n7220 & ~n14663 ;
  assign n44909 = x145 & n485 ;
  assign n44910 = n44909 ^ n14548 ^ 1'b0 ;
  assign n44911 = n44910 ^ n1873 ^ 1'b0 ;
  assign n44912 = n44911 ^ n15394 ^ n13067 ;
  assign n44914 = n44913 ^ n44912 ^ n41014 ;
  assign n44915 = ~n10255 & n25323 ;
  assign n44916 = n44915 ^ n33510 ^ 1'b0 ;
  assign n44917 = ( n27816 & n37482 ) | ( n27816 & ~n44916 ) | ( n37482 & ~n44916 ) ;
  assign n44918 = n35279 ^ x148 ^ 1'b0 ;
  assign n44919 = n5075 & ~n38625 ;
  assign n44920 = ~n2680 & n6390 ;
  assign n44921 = ~n42405 & n44920 ;
  assign n44922 = n6533 & ~n40461 ;
  assign n44923 = n44922 ^ n3125 ^ 1'b0 ;
  assign n44924 = n27194 | n32867 ;
  assign n44925 = n42017 ^ n8247 ^ n5737 ;
  assign n44926 = n22888 ^ n3826 ^ 1'b0 ;
  assign n44927 = n21669 ^ n11152 ^ 1'b0 ;
  assign n44928 = n44927 ^ n15539 ^ 1'b0 ;
  assign n44929 = n10440 & n29725 ;
  assign n44930 = n44929 ^ n36580 ^ n13722 ;
  assign n44931 = ~n37746 & n44930 ;
  assign n44932 = n15051 | n25687 ;
  assign n44933 = n44932 ^ n14543 ^ 1'b0 ;
  assign n44934 = n20335 | n20780 ;
  assign n44935 = n44933 | n44934 ;
  assign n44936 = n18694 ^ n2670 ^ 1'b0 ;
  assign n44937 = n31249 & n44936 ;
  assign n44938 = n15273 | n43560 ;
  assign n44939 = n20829 | n44938 ;
  assign n44940 = x233 & ~n44939 ;
  assign n44941 = n30219 ^ n2879 ^ 1'b0 ;
  assign n44942 = n25447 | n44941 ;
  assign n44943 = ~n15102 & n44942 ;
  assign n44944 = n34760 ^ n3950 ^ x145 ;
  assign n44945 = ( n8534 & ~n10408 ) | ( n8534 & n17612 ) | ( ~n10408 & n17612 ) ;
  assign n44946 = ( n9966 & n18367 ) | ( n9966 & ~n44945 ) | ( n18367 & ~n44945 ) ;
  assign n44947 = n41177 ^ n2989 ^ 1'b0 ;
  assign n44950 = n262 | n17881 ;
  assign n44949 = n16489 & ~n33041 ;
  assign n44948 = n12753 | n15693 ;
  assign n44951 = n44950 ^ n44949 ^ n44948 ;
  assign n44952 = ~n2788 & n10285 ;
  assign n44953 = n44952 ^ n27096 ^ 1'b0 ;
  assign n44954 = n36405 ^ n31803 ^ 1'b0 ;
  assign n44955 = n2868 & n44954 ;
  assign n44958 = n15979 & n36668 ;
  assign n44959 = n8488 & n44958 ;
  assign n44956 = n7670 & ~n12895 ;
  assign n44957 = n44956 ^ n19871 ^ 1'b0 ;
  assign n44960 = n44959 ^ n44957 ^ n4271 ;
  assign n44961 = n14297 & n27875 ;
  assign n44962 = n44960 & n44961 ;
  assign n44963 = n19908 ^ n4546 ^ 1'b0 ;
  assign n44964 = n1629 & ~n44963 ;
  assign n44966 = n8954 | n21059 ;
  assign n44967 = n16236 & ~n44966 ;
  assign n44965 = n8909 ^ n1142 ^ 1'b0 ;
  assign n44968 = n44967 ^ n44965 ^ n39648 ;
  assign n44969 = n23159 & ~n42612 ;
  assign n44970 = n44969 ^ n38411 ^ n19178 ;
  assign n44971 = ~n44968 & n44970 ;
  assign n44972 = n18476 ^ n17699 ^ n12329 ;
  assign n44973 = ( n11883 & n23301 ) | ( n11883 & n44972 ) | ( n23301 & n44972 ) ;
  assign n44974 = n13067 & ~n35108 ;
  assign n44975 = n40621 ^ n24844 ^ 1'b0 ;
  assign n44976 = n44767 & n44975 ;
  assign n44977 = ~n29036 & n44976 ;
  assign n44978 = n2752 & n27131 ;
  assign n44979 = n2255 | n35179 ;
  assign n44980 = n8658 & n26747 ;
  assign n44981 = n44980 ^ n4623 ^ 1'b0 ;
  assign n44982 = x167 & n25250 ;
  assign n44983 = n44982 ^ n34056 ^ 1'b0 ;
  assign n44984 = n24094 | n44983 ;
  assign n44985 = n10036 ^ n6674 ^ 1'b0 ;
  assign n44986 = n25625 | n44985 ;
  assign n44987 = n8034 & ~n44986 ;
  assign n44988 = n44987 ^ n32049 ^ n13384 ;
  assign n44989 = n12392 | n13690 ;
  assign n44991 = ( n1475 & ~n10777 ) | ( n1475 & n16817 ) | ( ~n10777 & n16817 ) ;
  assign n44990 = n26350 ^ n25629 ^ n4243 ;
  assign n44992 = n44991 ^ n44990 ^ 1'b0 ;
  assign n44993 = n19256 ^ n6001 ^ 1'b0 ;
  assign n44994 = ~n4723 & n44993 ;
  assign n44995 = ~n15888 & n44994 ;
  assign n44996 = n16508 ^ n15738 ^ 1'b0 ;
  assign n44999 = n18904 ^ n9040 ^ n8375 ;
  assign n44997 = n43267 ^ n37324 ^ n35473 ;
  assign n44998 = n6618 & ~n44997 ;
  assign n45000 = n44999 ^ n44998 ^ 1'b0 ;
  assign n45001 = n10163 & ~n38128 ;
  assign n45002 = n16878 & n45001 ;
  assign n45003 = ~n39738 & n45002 ;
  assign n45004 = n37485 ^ n32997 ^ n4416 ;
  assign n45005 = ~n2179 & n25400 ;
  assign n45006 = ~n7818 & n45005 ;
  assign n45007 = ( n18840 & n35116 ) | ( n18840 & ~n45006 ) | ( n35116 & ~n45006 ) ;
  assign n45008 = n16992 & n45007 ;
  assign n45009 = ~n21837 & n30776 ;
  assign n45010 = n45009 ^ n16819 ^ 1'b0 ;
  assign n45013 = n12875 ^ n3624 ^ n952 ;
  assign n45011 = n15486 ^ n6063 ^ n3984 ;
  assign n45012 = n33885 & n45011 ;
  assign n45014 = n45013 ^ n45012 ^ 1'b0 ;
  assign n45015 = n14550 ^ n11934 ^ 1'b0 ;
  assign n45016 = ~n31846 & n45015 ;
  assign n45019 = ~n12281 & n31471 ;
  assign n45020 = n27596 & n45019 ;
  assign n45021 = n45020 ^ n28136 ^ n20671 ;
  assign n45017 = n38493 ^ n1873 ^ x116 ;
  assign n45018 = n8534 & ~n45017 ;
  assign n45022 = n45021 ^ n45018 ^ 1'b0 ;
  assign n45023 = ( n7551 & n14619 ) | ( n7551 & ~n38924 ) | ( n14619 & ~n38924 ) ;
  assign n45024 = n2548 & n12836 ;
  assign n45025 = n16687 & ~n45024 ;
  assign n45026 = n45023 & ~n45025 ;
  assign n45027 = ( ~n9538 & n9861 ) | ( ~n9538 & n26837 ) | ( n9861 & n26837 ) ;
  assign n45028 = n27668 | n35086 ;
  assign n45029 = n12050 & ~n43473 ;
  assign n45032 = ( n2045 & ~n2715 ) | ( n2045 & n18175 ) | ( ~n2715 & n18175 ) ;
  assign n45033 = n45032 ^ n35130 ^ n26181 ;
  assign n45030 = n26328 ^ n13393 ^ n7293 ;
  assign n45031 = n42216 & ~n45030 ;
  assign n45034 = n45033 ^ n45031 ^ 1'b0 ;
  assign n45035 = n18962 | n23917 ;
  assign n45036 = n31011 ^ n17607 ^ 1'b0 ;
  assign n45037 = ~n39612 & n45036 ;
  assign n45038 = ( n1959 & n10342 ) | ( n1959 & n28271 ) | ( n10342 & n28271 ) ;
  assign n45039 = n4111 & n37255 ;
  assign n45040 = n45039 ^ n19644 ^ 1'b0 ;
  assign n45041 = ( n23708 & ~n39291 ) | ( n23708 & n45040 ) | ( ~n39291 & n45040 ) ;
  assign n45042 = n45041 ^ n40304 ^ 1'b0 ;
  assign n45044 = n11383 | n22251 ;
  assign n45045 = n42666 | n45044 ;
  assign n45043 = n11933 ^ n10593 ^ n3368 ;
  assign n45046 = n45045 ^ n45043 ^ n24169 ;
  assign n45047 = n18267 | n19250 ;
  assign n45048 = n45047 ^ n6424 ^ 1'b0 ;
  assign n45049 = n12600 | n15793 ;
  assign n45050 = n19675 & ~n45049 ;
  assign n45051 = ( n885 & ~n3648 ) | ( n885 & n5446 ) | ( ~n3648 & n5446 ) ;
  assign n45052 = n45051 ^ n23274 ^ n10416 ;
  assign n45053 = n45052 ^ n30075 ^ n21905 ;
  assign n45054 = n23724 | n45053 ;
  assign n45055 = n33696 ^ n10084 ^ n9139 ;
  assign n45056 = n43573 ^ n8850 ^ 1'b0 ;
  assign n45057 = n11809 | n16559 ;
  assign n45058 = n45057 ^ n1298 ^ 1'b0 ;
  assign n45059 = n45058 ^ n31433 ^ n30849 ;
  assign n45060 = n6506 & ~n11439 ;
  assign n45061 = ~n5690 & n40436 ;
  assign n45062 = n27041 ^ n4587 ^ 1'b0 ;
  assign n45063 = n16105 | n22802 ;
  assign n45064 = n39739 & n45063 ;
  assign n45065 = n11936 ^ n6024 ^ 1'b0 ;
  assign n45066 = n42424 ^ n25407 ^ n24250 ;
  assign n45067 = n1913 & ~n21052 ;
  assign n45068 = n14714 & ~n45067 ;
  assign n45069 = ~n39280 & n45068 ;
  assign n45075 = n1023 & n14662 ;
  assign n45076 = ~n1023 & n45075 ;
  assign n45070 = n8975 & n22467 ;
  assign n45071 = ~n8975 & n45070 ;
  assign n45072 = n3329 & ~n14559 ;
  assign n45073 = n45072 ^ n1805 ^ 1'b0 ;
  assign n45074 = ~n45071 & n45073 ;
  assign n45077 = n45076 ^ n45074 ^ 1'b0 ;
  assign n45078 = n24270 & n45077 ;
  assign n45079 = n18519 | n38206 ;
  assign n45080 = n45079 ^ n10456 ^ 1'b0 ;
  assign n45081 = n45080 ^ n24641 ^ 1'b0 ;
  assign n45082 = n32996 ^ n25942 ^ n23074 ;
  assign n45083 = ( n23686 & n26877 ) | ( n23686 & ~n35939 ) | ( n26877 & ~n35939 ) ;
  assign n45084 = n36097 ^ n26503 ^ n9352 ;
  assign n45086 = n20458 | n34862 ;
  assign n45085 = ~n8418 & n16126 ;
  assign n45087 = n45086 ^ n45085 ^ 1'b0 ;
  assign n45088 = n3773 & ~n10643 ;
  assign n45089 = n45088 ^ n34186 ^ 1'b0 ;
  assign n45090 = n37259 ^ n14548 ^ 1'b0 ;
  assign n45091 = n45089 & n45090 ;
  assign n45092 = ( n6352 & n20900 ) | ( n6352 & n41625 ) | ( n20900 & n41625 ) ;
  assign n45093 = n22032 ^ n21045 ^ 1'b0 ;
  assign n45094 = n45092 & n45093 ;
  assign n45095 = n18963 | n26773 ;
  assign n45096 = n45095 ^ n32901 ^ n6916 ;
  assign n45097 = n6371 ^ n5528 ^ 1'b0 ;
  assign n45098 = n1043 | n45097 ;
  assign n45099 = ( n5798 & n11653 ) | ( n5798 & n45098 ) | ( n11653 & n45098 ) ;
  assign n45100 = n20220 & n45099 ;
  assign n45101 = n33691 ^ n1194 ^ 1'b0 ;
  assign n45102 = n11921 ^ n8552 ^ 1'b0 ;
  assign n45103 = n36639 & n45102 ;
  assign n45104 = n17140 & n44102 ;
  assign n45105 = n45103 & n45104 ;
  assign n45106 = n34559 ^ n8835 ^ n4891 ;
  assign n45107 = n12371 ^ n12144 ^ 1'b0 ;
  assign n45108 = n18306 | n45107 ;
  assign n45109 = n45108 ^ n27743 ^ 1'b0 ;
  assign n45110 = n30564 & n45109 ;
  assign n45111 = n14393 & ~n14430 ;
  assign n45112 = n45111 ^ n1689 ^ 1'b0 ;
  assign n45113 = n30012 ^ n10234 ^ 1'b0 ;
  assign n45114 = n28719 ^ n3349 ^ 1'b0 ;
  assign n45115 = n41635 ^ n17990 ^ 1'b0 ;
  assign n45116 = n7022 & ~n18428 ;
  assign n45117 = n12342 & n45116 ;
  assign n45118 = n45117 ^ n13538 ^ 1'b0 ;
  assign n45119 = n33568 & n45118 ;
  assign n45120 = n45119 ^ n6769 ^ 1'b0 ;
  assign n45122 = n19216 ^ n11920 ^ n3892 ;
  assign n45121 = n7376 | n30912 ;
  assign n45123 = n45122 ^ n45121 ^ 1'b0 ;
  assign n45124 = ~n5345 & n45123 ;
  assign n45125 = ~n21615 & n45124 ;
  assign n45127 = n3961 & ~n35251 ;
  assign n45126 = ~n4855 & n42804 ;
  assign n45128 = n45127 ^ n45126 ^ 1'b0 ;
  assign n45129 = n42097 & n42175 ;
  assign n45130 = n12236 & n45129 ;
  assign n45132 = ( ~n1204 & n4273 ) | ( ~n1204 & n22004 ) | ( n4273 & n22004 ) ;
  assign n45131 = n17629 | n36644 ;
  assign n45133 = n45132 ^ n45131 ^ 1'b0 ;
  assign n45134 = n44238 ^ n10723 ^ 1'b0 ;
  assign n45135 = ~n3943 & n45134 ;
  assign n45136 = n11926 & ~n31332 ;
  assign n45137 = n7326 & n45136 ;
  assign n45138 = n5603 & ~n45137 ;
  assign n45139 = n9492 | n20995 ;
  assign n45140 = n13146 & n18800 ;
  assign n45141 = n5817 & n43856 ;
  assign n45142 = n45141 ^ n20810 ^ 1'b0 ;
  assign n45143 = ( n25569 & ~n45140 ) | ( n25569 & n45142 ) | ( ~n45140 & n45142 ) ;
  assign n45144 = n23427 ^ n19819 ^ 1'b0 ;
  assign n45145 = n1102 & n45144 ;
  assign n45165 = n35256 ^ n32753 ^ n13389 ;
  assign n45146 = ~n692 & n952 ;
  assign n45147 = ~n952 & n45146 ;
  assign n45148 = n6266 | n45147 ;
  assign n45149 = n6266 & ~n45148 ;
  assign n45150 = n302 | n1106 ;
  assign n45151 = n1106 & ~n45150 ;
  assign n45152 = x55 & ~n45151 ;
  assign n45153 = n45151 & n45152 ;
  assign n45154 = n45149 | n45153 ;
  assign n45155 = n45149 & ~n45154 ;
  assign n45156 = n578 & n14108 ;
  assign n45157 = ~n578 & n45156 ;
  assign n45158 = n6249 | n6620 ;
  assign n45159 = n6620 & ~n45158 ;
  assign n45160 = n2507 | n45159 ;
  assign n45161 = n45160 ^ n6157 ^ 1'b0 ;
  assign n45162 = n3898 & ~n45161 ;
  assign n45163 = n45162 ^ n10105 ^ 1'b0 ;
  assign n45164 = ( ~n45155 & n45157 ) | ( ~n45155 & n45163 ) | ( n45157 & n45163 ) ;
  assign n45166 = n45165 ^ n45164 ^ n14575 ;
  assign n45167 = n16530 & n40264 ;
  assign n45168 = ~n27978 & n45167 ;
  assign n45169 = n36791 ^ n21345 ^ 1'b0 ;
  assign n45170 = n15634 | n45169 ;
  assign n45171 = n2047 | n8277 ;
  assign n45172 = n45171 ^ n28376 ^ 1'b0 ;
  assign n45173 = n10072 ^ n1309 ^ 1'b0 ;
  assign n45174 = x198 & ~n40258 ;
  assign n45175 = n26175 ^ n22381 ^ 1'b0 ;
  assign n45176 = n45175 ^ n32655 ^ n26944 ;
  assign n45177 = n4217 & n32292 ;
  assign n45178 = ~n32257 & n45177 ;
  assign n45179 = n17799 | n45178 ;
  assign n45180 = n6441 & n8164 ;
  assign n45181 = ( n14026 & n29707 ) | ( n14026 & n45180 ) | ( n29707 & n45180 ) ;
  assign n45183 = n12032 & n38015 ;
  assign n45184 = n21968 & n45183 ;
  assign n45182 = ~n1222 & n2672 ;
  assign n45185 = n45184 ^ n45182 ^ 1'b0 ;
  assign n45186 = n9626 & n24747 ;
  assign n45187 = n10176 ^ n2462 ^ 1'b0 ;
  assign n45188 = n23784 ^ n3564 ^ 1'b0 ;
  assign n45189 = n45187 & n45188 ;
  assign n45190 = ~n27309 & n41990 ;
  assign n45191 = n4421 & n8376 ;
  assign n45192 = n45191 ^ n13416 ^ 1'b0 ;
  assign n45193 = n29872 ^ n23600 ^ n19876 ;
  assign n45194 = n45192 & n45193 ;
  assign n45195 = n16003 ^ n4922 ^ 1'b0 ;
  assign n45196 = n2142 & ~n45195 ;
  assign n45197 = n13822 & n45196 ;
  assign n45198 = n45197 ^ n12269 ^ 1'b0 ;
  assign n45199 = n45198 ^ n5816 ^ 1'b0 ;
  assign n45200 = n17794 ^ n2314 ^ n2278 ;
  assign n45201 = n16202 & ~n18276 ;
  assign n45202 = n26156 & n37671 ;
  assign n45203 = ~n18667 & n45202 ;
  assign n45204 = n44654 & ~n45203 ;
  assign n45207 = ~n637 & n13032 ;
  assign n45208 = n45207 ^ n33090 ^ 1'b0 ;
  assign n45205 = n39121 ^ n31311 ^ n29880 ;
  assign n45206 = n18209 | n45205 ;
  assign n45209 = n45208 ^ n45206 ^ 1'b0 ;
  assign n45210 = ~n2577 & n43523 ;
  assign n45211 = ~n32406 & n45210 ;
  assign n45212 = n19533 ^ n15528 ^ 1'b0 ;
  assign n45213 = n33008 | n45212 ;
  assign n45214 = n17888 & n26112 ;
  assign n45215 = n45214 ^ n12572 ^ 1'b0 ;
  assign n45216 = ( n3051 & ~n5253 ) | ( n3051 & n15186 ) | ( ~n5253 & n15186 ) ;
  assign n45217 = ( n17959 & ~n33097 ) | ( n17959 & n45216 ) | ( ~n33097 & n45216 ) ;
  assign n45218 = n18528 ^ n7077 ^ 1'b0 ;
  assign n45219 = x98 & ~n45218 ;
  assign n45220 = n45219 ^ n17036 ^ 1'b0 ;
  assign n45221 = ~n27193 & n34508 ;
  assign n45222 = ~n26718 & n45221 ;
  assign n45223 = n45222 ^ n40833 ^ 1'b0 ;
  assign n45224 = n6980 | n13395 ;
  assign n45225 = n26485 & ~n45224 ;
  assign n45226 = ~n20491 & n38865 ;
  assign n45227 = ~n36506 & n45226 ;
  assign n45228 = n36776 | n44023 ;
  assign n45229 = n45228 ^ n29071 ^ 1'b0 ;
  assign n45230 = n16521 ^ n256 ^ 1'b0 ;
  assign n45231 = n25781 | n45230 ;
  assign n45232 = n25619 ^ n14355 ^ 1'b0 ;
  assign n45233 = n17816 | n45232 ;
  assign n45234 = ~n2628 & n32393 ;
  assign n45235 = n18865 & n45234 ;
  assign n45237 = n10941 & ~n13179 ;
  assign n45236 = n13708 ^ n925 ^ 1'b0 ;
  assign n45238 = n45237 ^ n45236 ^ n39020 ;
  assign n45239 = n20456 ^ n8246 ^ 1'b0 ;
  assign n45240 = n7497 | n15632 ;
  assign n45241 = n23798 | n45240 ;
  assign n45242 = n36112 ^ n14107 ^ 1'b0 ;
  assign n45243 = n31521 & ~n45242 ;
  assign n45244 = n31002 ^ n12624 ^ 1'b0 ;
  assign n45245 = n13167 & n24096 ;
  assign n45246 = n45244 & n45245 ;
  assign n45247 = n21062 ^ n1352 ^ 1'b0 ;
  assign n45248 = n28407 ^ n25582 ^ 1'b0 ;
  assign n45249 = n980 | n19399 ;
  assign n45250 = n5241 | n45249 ;
  assign n45251 = n11708 & ~n45250 ;
  assign n45252 = ~n45248 & n45251 ;
  assign n45253 = n10216 & n45092 ;
  assign n45254 = n31543 ^ n12828 ^ 1'b0 ;
  assign n45255 = n18864 ^ n7827 ^ x113 ;
  assign n45256 = n13453 ^ n12539 ^ 1'b0 ;
  assign n45257 = n2130 | n45256 ;
  assign n45258 = ~n45255 & n45257 ;
  assign n45259 = ~n2558 & n45258 ;
  assign n45260 = ( n11551 & ~n28327 ) | ( n11551 & n43483 ) | ( ~n28327 & n43483 ) ;
  assign n45261 = n18372 & n30719 ;
  assign n45262 = n45261 ^ n5744 ^ 1'b0 ;
  assign n45263 = n45262 ^ n33438 ^ 1'b0 ;
  assign n45264 = n13249 ^ n4767 ^ 1'b0 ;
  assign n45265 = n45263 | n45264 ;
  assign n45266 = n7195 ^ x42 ^ 1'b0 ;
  assign n45267 = n27122 & n45266 ;
  assign n45268 = n5818 & n36656 ;
  assign n45269 = ~n35661 & n45268 ;
  assign n45270 = n39114 ^ n33117 ^ n12190 ;
  assign n45271 = ( n28020 & ~n42430 ) | ( n28020 & n45270 ) | ( ~n42430 & n45270 ) ;
  assign n45272 = n34605 & n41322 ;
  assign n45273 = ~n34197 & n45272 ;
  assign n45274 = ~n5398 & n19382 ;
  assign n45275 = n45273 & n45274 ;
  assign n45276 = ( n4944 & n5991 ) | ( n4944 & n45275 ) | ( n5991 & n45275 ) ;
  assign n45277 = n28981 ^ n26674 ^ n15836 ;
  assign n45278 = n14437 ^ n7291 ^ n2562 ;
  assign n45279 = n22319 ^ n18848 ^ 1'b0 ;
  assign n45280 = n11510 & n45279 ;
  assign n45282 = ( n13837 & n14262 ) | ( n13837 & n27832 ) | ( n14262 & n27832 ) ;
  assign n45283 = n45282 ^ n24764 ^ 1'b0 ;
  assign n45284 = n20680 & ~n45283 ;
  assign n45281 = n10910 | n23587 ;
  assign n45285 = n45284 ^ n45281 ^ 1'b0 ;
  assign n45286 = n45095 ^ n35287 ^ 1'b0 ;
  assign n45287 = n18675 | n38668 ;
  assign n45288 = ~n3877 & n4355 ;
  assign n45289 = n18709 ^ n1688 ^ 1'b0 ;
  assign n45290 = n45289 ^ n4840 ^ 1'b0 ;
  assign n45291 = n35135 | n39464 ;
  assign n45292 = n45291 ^ n11511 ^ 1'b0 ;
  assign n45293 = n45292 ^ n6111 ^ 1'b0 ;
  assign n45302 = ( n4067 & n5226 ) | ( n4067 & ~n13114 ) | ( n5226 & ~n13114 ) ;
  assign n45294 = n10220 ^ n1294 ^ 1'b0 ;
  assign n45295 = ~n28486 & n45294 ;
  assign n45296 = ( n8808 & n12255 ) | ( n8808 & ~n30832 ) | ( n12255 & ~n30832 ) ;
  assign n45297 = n45296 ^ n4388 ^ 1'b0 ;
  assign n45298 = n25261 & n45297 ;
  assign n45299 = ( n11811 & ~n45295 ) | ( n11811 & n45298 ) | ( ~n45295 & n45298 ) ;
  assign n45300 = ( n24146 & n43598 ) | ( n24146 & n45299 ) | ( n43598 & n45299 ) ;
  assign n45301 = ~n2033 & n45300 ;
  assign n45303 = n45302 ^ n45301 ^ 1'b0 ;
  assign n45304 = n45173 ^ n8739 ^ 1'b0 ;
  assign n45305 = n13062 ^ n3053 ^ 1'b0 ;
  assign n45306 = ~n7254 & n14662 ;
  assign n45307 = n33690 ^ n30116 ^ 1'b0 ;
  assign n45309 = n9793 | n15890 ;
  assign n45308 = ~n9967 & n22373 ;
  assign n45310 = n45309 ^ n45308 ^ n22371 ;
  assign n45311 = ( n17678 & ~n45307 ) | ( n17678 & n45310 ) | ( ~n45307 & n45310 ) ;
  assign n45312 = n25970 ^ n12105 ^ n11293 ;
  assign n45317 = n11467 ^ n7542 ^ 1'b0 ;
  assign n45318 = n7672 | n45317 ;
  assign n45313 = n10847 & ~n14273 ;
  assign n45314 = ~n5937 & n45313 ;
  assign n45315 = n45314 ^ n2731 ^ 1'b0 ;
  assign n45316 = n17887 | n45315 ;
  assign n45319 = n45318 ^ n45316 ^ 1'b0 ;
  assign n45320 = ~n929 & n25354 ;
  assign n45321 = ~n7620 & n45320 ;
  assign n45322 = ~n18569 & n42097 ;
  assign n45323 = n45322 ^ n20436 ^ 1'b0 ;
  assign n45324 = ( n5114 & ~n24575 ) | ( n5114 & n45006 ) | ( ~n24575 & n45006 ) ;
  assign n45325 = n33912 ^ n29698 ^ n16221 ;
  assign n45326 = n4746 | n45325 ;
  assign n45327 = n31427 ^ n29192 ^ n21003 ;
  assign n45328 = n13561 ^ n13281 ^ 1'b0 ;
  assign n45329 = n45328 ^ n40614 ^ n27670 ;
  assign n45330 = n28924 & n45329 ;
  assign n45331 = n45327 & n45330 ;
  assign n45332 = n10422 & ~n25116 ;
  assign n45333 = ~n24060 & n45332 ;
  assign n45334 = n1126 | n2227 ;
  assign n45335 = ( n7451 & n17794 ) | ( n7451 & n45334 ) | ( n17794 & n45334 ) ;
  assign n45336 = n15430 & ~n45335 ;
  assign n45337 = ~n7692 & n23584 ;
  assign n45338 = n45337 ^ n44534 ^ 1'b0 ;
  assign n45339 = n35094 & ~n45338 ;
  assign n45340 = ~n45336 & n45339 ;
  assign n45341 = n15202 ^ n8655 ^ 1'b0 ;
  assign n45343 = n5824 & ~n8058 ;
  assign n45342 = ~n11501 & n12463 ;
  assign n45344 = n45343 ^ n45342 ^ 1'b0 ;
  assign n45345 = ( n932 & n5362 ) | ( n932 & n5521 ) | ( n5362 & n5521 ) ;
  assign n45347 = n4621 ^ x139 ^ 1'b0 ;
  assign n45348 = n2430 & n45347 ;
  assign n45346 = n8787 & n20530 ;
  assign n45349 = n45348 ^ n45346 ^ n19723 ;
  assign n45350 = n7262 & n15486 ;
  assign n45351 = ~n30506 & n45350 ;
  assign n45352 = ( n4215 & ~n5499 ) | ( n4215 & n26907 ) | ( ~n5499 & n26907 ) ;
  assign n45353 = ~n31779 & n43893 ;
  assign n45357 = ~n18895 & n24383 ;
  assign n45358 = ~n28362 & n45357 ;
  assign n45359 = n7822 ^ n2103 ^ 1'b0 ;
  assign n45360 = n45358 | n45359 ;
  assign n45354 = n20945 ^ n3305 ^ 1'b0 ;
  assign n45355 = n42160 | n45354 ;
  assign n45356 = n6581 & ~n45355 ;
  assign n45361 = n45360 ^ n45356 ^ 1'b0 ;
  assign n45365 = n5417 & ~n6886 ;
  assign n45366 = n14363 & n45365 ;
  assign n45367 = ( n5491 & n25444 ) | ( n5491 & ~n45366 ) | ( n25444 & ~n45366 ) ;
  assign n45362 = n22486 ^ n6865 ^ 1'b0 ;
  assign n45363 = n6082 | n45362 ;
  assign n45364 = n11706 | n45363 ;
  assign n45368 = n45367 ^ n45364 ^ n26298 ;
  assign n45369 = n17570 ^ n16467 ^ 1'b0 ;
  assign n45370 = ~n16728 & n25177 ;
  assign n45371 = n45370 ^ n23236 ^ n3250 ;
  assign n45372 = n23392 ^ n21555 ^ n9858 ;
  assign n45373 = n45372 ^ n34252 ^ n15648 ;
  assign n45374 = n35951 ^ n21185 ^ n10564 ;
  assign n45375 = n45374 ^ n9594 ^ 1'b0 ;
  assign n45377 = ~n9741 & n19065 ;
  assign n45378 = n45377 ^ n26638 ^ 1'b0 ;
  assign n45376 = n14820 ^ n11651 ^ n6154 ;
  assign n45379 = n45378 ^ n45376 ^ 1'b0 ;
  assign n45380 = n22710 & ~n45379 ;
  assign n45381 = ( n13396 & n19571 ) | ( n13396 & n25521 ) | ( n19571 & n25521 ) ;
  assign n45382 = n24191 ^ n5362 ^ 1'b0 ;
  assign n45383 = n45382 ^ n7440 ^ 1'b0 ;
  assign n45384 = n34766 | n45383 ;
  assign n45385 = ( ~n1094 & n12060 ) | ( ~n1094 & n20690 ) | ( n12060 & n20690 ) ;
  assign n45386 = n24423 & n45385 ;
  assign n45387 = n45386 ^ n2756 ^ 1'b0 ;
  assign n45388 = n32898 ^ n6164 ^ 1'b0 ;
  assign n45389 = n38991 & ~n45388 ;
  assign n45390 = n45389 ^ n39576 ^ 1'b0 ;
  assign n45391 = ~n567 & n44763 ;
  assign n45392 = n33227 | n45391 ;
  assign n45393 = n45390 & ~n45392 ;
  assign n45394 = n11795 ^ n6219 ^ 1'b0 ;
  assign n45395 = n1626 | n45394 ;
  assign n45396 = n45395 ^ n9221 ^ 1'b0 ;
  assign n45397 = ~n5439 & n45396 ;
  assign n45398 = n33785 ^ n11486 ^ 1'b0 ;
  assign n45399 = n3466 & n4474 ;
  assign n45400 = n13121 ^ n11330 ^ n2454 ;
  assign n45401 = ~n2950 & n10349 ;
  assign n45402 = n45401 ^ n5480 ^ 1'b0 ;
  assign n45403 = n45402 ^ n20466 ^ 1'b0 ;
  assign n45404 = ( n1778 & n5133 ) | ( n1778 & ~n10094 ) | ( n5133 & ~n10094 ) ;
  assign n45405 = n3439 & n7027 ;
  assign n45406 = ~n38716 & n45405 ;
  assign n45407 = n28486 | n45406 ;
  assign n45408 = n45407 ^ n40832 ^ 1'b0 ;
  assign n45409 = ( n9937 & n45404 ) | ( n9937 & ~n45408 ) | ( n45404 & ~n45408 ) ;
  assign n45410 = n23391 ^ x192 ^ 1'b0 ;
  assign n45411 = n3086 & n12380 ;
  assign n45412 = n45411 ^ n5619 ^ 1'b0 ;
  assign n45413 = ~n9868 & n45412 ;
  assign n45414 = n42160 ^ n30948 ^ 1'b0 ;
  assign n45415 = n36381 & ~n45414 ;
  assign n45416 = n37485 & ~n44976 ;
  assign n45417 = n9906 & ~n10076 ;
  assign n45418 = ~n14734 & n45417 ;
  assign n45419 = ( n4107 & ~n42896 ) | ( n4107 & n45418 ) | ( ~n42896 & n45418 ) ;
  assign n45420 = n29233 ^ n4498 ^ 1'b0 ;
  assign n45421 = n34341 ^ n17341 ^ 1'b0 ;
  assign n45422 = n4498 & ~n12663 ;
  assign n45423 = ~n7795 & n45422 ;
  assign n45424 = n3544 & n45423 ;
  assign n45425 = n45424 ^ n31179 ^ n10487 ;
  assign n45426 = n38641 ^ n24506 ^ 1'b0 ;
  assign n45427 = n45144 & n45426 ;
  assign n45428 = n30201 ^ n22372 ^ n11381 ;
  assign n45429 = n22371 & n45428 ;
  assign n45430 = n28236 ^ n14510 ^ 1'b0 ;
  assign n45431 = n45429 & n45430 ;
  assign n45432 = ( n14417 & n22610 ) | ( n14417 & ~n36303 ) | ( n22610 & ~n36303 ) ;
  assign n45433 = n24681 & ~n45432 ;
  assign n45434 = n9995 & ~n23840 ;
  assign n45435 = n45434 ^ n13353 ^ 1'b0 ;
  assign n45436 = n403 | n37411 ;
  assign n45437 = n45435 & ~n45436 ;
  assign n45438 = n2482 & ~n4185 ;
  assign n45439 = n45438 ^ n2823 ^ 1'b0 ;
  assign n45440 = n37389 & ~n45439 ;
  assign n45441 = n10034 & ~n21822 ;
  assign n45442 = n316 & ~n9933 ;
  assign n45443 = n45442 ^ n28272 ^ 1'b0 ;
  assign n45444 = ( n19993 & n45441 ) | ( n19993 & n45443 ) | ( n45441 & n45443 ) ;
  assign n45446 = n12886 ^ n8979 ^ 1'b0 ;
  assign n45447 = n13211 | n45446 ;
  assign n45445 = ~n1707 & n18892 ;
  assign n45448 = n45447 ^ n45445 ^ 1'b0 ;
  assign n45449 = n31817 & ~n45448 ;
  assign n45450 = n22682 & ~n26658 ;
  assign n45451 = n33240 ^ n16416 ^ 1'b0 ;
  assign n45452 = n13438 ^ n679 ^ 1'b0 ;
  assign n45453 = n15611 & ~n19113 ;
  assign n45454 = n45453 ^ n6075 ^ 1'b0 ;
  assign n45455 = n45454 ^ n42507 ^ n37511 ;
  assign n45456 = n5996 ^ n4966 ^ 1'b0 ;
  assign n45457 = n23253 | n30489 ;
  assign n45458 = ~n18248 & n21164 ;
  assign n45459 = n45458 ^ n2017 ^ 1'b0 ;
  assign n45460 = n31279 ^ n845 ^ 1'b0 ;
  assign n45461 = n1454 & n2594 ;
  assign n45462 = n45461 ^ n38323 ^ 1'b0 ;
  assign n45463 = ( n5071 & n9807 ) | ( n5071 & n30874 ) | ( n9807 & n30874 ) ;
  assign n45464 = n45463 ^ n13786 ^ 1'b0 ;
  assign n45465 = n6674 & ~n13116 ;
  assign n45466 = ~n45464 & n45465 ;
  assign n45467 = n45466 ^ n4159 ^ 1'b0 ;
  assign n45468 = ~x46 & n21978 ;
  assign n45469 = n45468 ^ n33057 ^ 1'b0 ;
  assign n45470 = n43109 & ~n45469 ;
  assign n45471 = ( n12585 & ~n12634 ) | ( n12585 & n45470 ) | ( ~n12634 & n45470 ) ;
  assign n45472 = n4369 | n12684 ;
  assign n45473 = ( n14023 & n17751 ) | ( n14023 & n45472 ) | ( n17751 & n45472 ) ;
  assign n45474 = n2818 & n14014 ;
  assign n45475 = n45474 ^ n10690 ^ 1'b0 ;
  assign n45476 = n4026 | n45475 ;
  assign n45477 = ( ~n38088 & n44343 ) | ( ~n38088 & n45476 ) | ( n44343 & n45476 ) ;
  assign n45478 = n5595 | n18774 ;
  assign n45479 = n30354 ^ n9958 ^ 1'b0 ;
  assign n45480 = ~n13947 & n45479 ;
  assign n45481 = n45480 ^ n4537 ^ 1'b0 ;
  assign n45482 = n14810 & n45481 ;
  assign n45483 = ~n45478 & n45482 ;
  assign n45484 = n10497 & ~n45483 ;
  assign n45485 = n45484 ^ n8346 ^ 1'b0 ;
  assign n45486 = n27381 ^ n17239 ^ 1'b0 ;
  assign n45487 = ~n44981 & n45486 ;
  assign n45488 = n22923 ^ n7294 ^ n2939 ;
  assign n45489 = n12026 & ~n13102 ;
  assign n45490 = n45488 & n45489 ;
  assign n45491 = n15039 & n28235 ;
  assign n45492 = n45491 ^ n23068 ^ n2200 ;
  assign n45493 = n45492 ^ n9834 ^ 1'b0 ;
  assign n45495 = n22928 & n22930 ;
  assign n45496 = n5004 & n45495 ;
  assign n45494 = n10994 & n35196 ;
  assign n45497 = n45496 ^ n45494 ^ 1'b0 ;
  assign n45498 = n1598 & n3688 ;
  assign n45499 = n45498 ^ n42250 ^ 1'b0 ;
  assign n45500 = ( n3273 & n22850 ) | ( n3273 & ~n23089 ) | ( n22850 & ~n23089 ) ;
  assign n45501 = ( n37757 & n45499 ) | ( n37757 & ~n45500 ) | ( n45499 & ~n45500 ) ;
  assign n45502 = n2945 & n8935 ;
  assign n45503 = n2847 & n45502 ;
  assign n45504 = n18877 & n45503 ;
  assign n45505 = n42143 ^ n14551 ^ n10031 ;
  assign n45506 = ( n17880 & ~n45504 ) | ( n17880 & n45505 ) | ( ~n45504 & n45505 ) ;
  assign n45507 = n28157 ^ n23218 ^ n11882 ;
  assign n45508 = ( n9480 & n17397 ) | ( n9480 & ~n32826 ) | ( n17397 & ~n32826 ) ;
  assign n45509 = n1962 & ~n6334 ;
  assign n45510 = n45509 ^ n1775 ^ 1'b0 ;
  assign n45511 = ~n13115 & n16301 ;
  assign n45512 = n30525 & n45511 ;
  assign n45513 = n34269 | n45512 ;
  assign n45514 = n20637 & ~n24664 ;
  assign n45515 = n13234 & n45514 ;
  assign n45516 = n24434 ^ n14322 ^ 1'b0 ;
  assign n45517 = ~n20785 & n45516 ;
  assign n45518 = n11907 | n40619 ;
  assign n45523 = n43751 ^ n43466 ^ n13151 ;
  assign n45519 = n10240 & n32319 ;
  assign n45520 = n45519 ^ n14641 ^ 1'b0 ;
  assign n45521 = n18641 | n45520 ;
  assign n45522 = n25278 & ~n45521 ;
  assign n45524 = n45523 ^ n45522 ^ 1'b0 ;
  assign n45525 = n34671 ^ n503 ^ 1'b0 ;
  assign n45526 = ( n13241 & ~n39506 ) | ( n13241 & n45525 ) | ( ~n39506 & n45525 ) ;
  assign n45527 = ~n814 & n4792 ;
  assign n45528 = n45527 ^ n9376 ^ 1'b0 ;
  assign n45531 = n23469 ^ n6310 ^ 1'b0 ;
  assign n45532 = x202 & ~n45531 ;
  assign n45529 = n24802 ^ n4590 ^ 1'b0 ;
  assign n45530 = n31501 & n45529 ;
  assign n45533 = n45532 ^ n45530 ^ 1'b0 ;
  assign n45534 = n6728 & ~n28159 ;
  assign n45535 = ~n1770 & n45534 ;
  assign n45536 = n23839 | n33785 ;
  assign n45537 = n45535 & ~n45536 ;
  assign n45538 = ( ~n378 & n24293 ) | ( ~n378 & n45537 ) | ( n24293 & n45537 ) ;
  assign n45539 = n1969 & ~n5296 ;
  assign n45540 = n6717 & n45539 ;
  assign n45541 = n27208 | n45540 ;
  assign n45542 = n41477 & ~n45541 ;
  assign n45543 = n10401 & n26064 ;
  assign n45544 = n45543 ^ n8894 ^ 1'b0 ;
  assign n45545 = n45544 ^ n43807 ^ 1'b0 ;
  assign n45546 = n9113 & ~n10333 ;
  assign n45547 = n24668 & n45546 ;
  assign n45548 = n1079 & n5800 ;
  assign n45549 = ( ~n10557 & n16993 ) | ( ~n10557 & n31155 ) | ( n16993 & n31155 ) ;
  assign n45550 = n3281 ^ n692 ^ 1'b0 ;
  assign n45551 = n45550 ^ n28266 ^ n9707 ;
  assign n45552 = n1009 & ~n6435 ;
  assign n45553 = n45552 ^ n12885 ^ 1'b0 ;
  assign n45554 = n28230 ^ n20661 ^ 1'b0 ;
  assign n45555 = ~n25112 & n45554 ;
  assign n45556 = n36348 & ~n37287 ;
  assign n45557 = n45556 ^ n10248 ^ 1'b0 ;
  assign n45558 = n45557 ^ n5475 ^ 1'b0 ;
  assign n45559 = n19004 | n45558 ;
  assign n45560 = n21580 ^ n3965 ^ 1'b0 ;
  assign n45561 = n15270 ^ n3840 ^ 1'b0 ;
  assign n45562 = n45560 & ~n45561 ;
  assign n45563 = n41998 ^ n21726 ^ 1'b0 ;
  assign n45564 = ( ~n3025 & n16430 ) | ( ~n3025 & n20116 ) | ( n16430 & n20116 ) ;
  assign n45565 = n18440 | n41980 ;
  assign n45566 = n8611 & ~n22315 ;
  assign n45567 = ~n25627 & n26217 ;
  assign n45568 = n40262 ^ n438 ^ 1'b0 ;
  assign n45569 = n12513 | n45568 ;
  assign n45571 = n23448 ^ n10165 ^ n3080 ;
  assign n45570 = ~n28122 & n32799 ;
  assign n45572 = n45571 ^ n45570 ^ 1'b0 ;
  assign n45573 = n35116 & n44578 ;
  assign n45574 = n38391 & n45573 ;
  assign n45575 = n25586 ^ n24474 ^ x75 ;
  assign n45576 = ( n8088 & n13576 ) | ( n8088 & n23753 ) | ( n13576 & n23753 ) ;
  assign n45577 = n20148 ^ n12118 ^ 1'b0 ;
  assign n45578 = ~n943 & n25247 ;
  assign n45579 = n45578 ^ n7536 ^ 1'b0 ;
  assign n45580 = n43124 ^ n16157 ^ 1'b0 ;
  assign n45581 = ~n20431 & n45580 ;
  assign n45582 = n9953 & n28669 ;
  assign n45583 = n45582 ^ n16702 ^ 1'b0 ;
  assign n45584 = n8569 ^ n3178 ^ 1'b0 ;
  assign n45585 = n45584 ^ n32602 ^ 1'b0 ;
  assign n45586 = n7715 & n45585 ;
  assign n45587 = ( n8000 & n41830 ) | ( n8000 & ~n43907 ) | ( n41830 & ~n43907 ) ;
  assign n45588 = n45587 ^ n1374 ^ 1'b0 ;
  assign n45589 = n20256 & ~n31304 ;
  assign n45594 = n3575 | n19109 ;
  assign n45595 = n1154 | n45594 ;
  assign n45590 = n19190 | n44377 ;
  assign n45591 = n45590 ^ n25630 ^ 1'b0 ;
  assign n45592 = n45591 ^ n17445 ^ 1'b0 ;
  assign n45593 = ~n32691 & n45592 ;
  assign n45596 = n45595 ^ n45593 ^ 1'b0 ;
  assign n45597 = n27612 ^ n8333 ^ 1'b0 ;
  assign n45598 = n13738 | n23788 ;
  assign n45599 = n45598 ^ n8300 ^ 1'b0 ;
  assign n45600 = x184 & ~n23096 ;
  assign n45601 = n22430 & n45600 ;
  assign n45602 = n8282 | n36267 ;
  assign n45603 = n45602 ^ n6005 ^ 1'b0 ;
  assign n45604 = n44654 ^ n29453 ^ n24908 ;
  assign n45605 = ( n21062 & n31782 ) | ( n21062 & ~n34067 ) | ( n31782 & ~n34067 ) ;
  assign n45606 = n45605 ^ n28767 ^ n13722 ;
  assign n45607 = n19350 | n33179 ;
  assign n45608 = n45607 ^ n31794 ^ 1'b0 ;
  assign n45609 = n34855 ^ n12004 ^ 1'b0 ;
  assign n45610 = n20983 ^ n20808 ^ 1'b0 ;
  assign n45611 = n45610 ^ n36793 ^ 1'b0 ;
  assign n45612 = n16600 | n18894 ;
  assign n45613 = n11109 & ~n45612 ;
  assign n45614 = n4243 & ~n19402 ;
  assign n45615 = n45614 ^ n17507 ^ 1'b0 ;
  assign n45616 = ( n30387 & n41389 ) | ( n30387 & ~n45615 ) | ( n41389 & ~n45615 ) ;
  assign n45617 = n32484 ^ n16497 ^ n5228 ;
  assign n45618 = ( n8798 & n16351 ) | ( n8798 & n17572 ) | ( n16351 & n17572 ) ;
  assign n45619 = ~n8911 & n45618 ;
  assign n45620 = n45619 ^ n21875 ^ n13984 ;
  assign n45621 = n17163 & n27467 ;
  assign n45622 = n13733 | n16757 ;
  assign n45623 = n29852 ^ n2613 ^ 1'b0 ;
  assign n45624 = n45622 & ~n45623 ;
  assign n45625 = n2331 & ~n37828 ;
  assign n45626 = n10373 & n45625 ;
  assign n45627 = n40099 ^ n37829 ^ 1'b0 ;
  assign n45628 = n4214 & n9388 ;
  assign n45630 = n4525 | n12041 ;
  assign n45631 = ~n1842 & n6229 ;
  assign n45632 = n1842 & n45631 ;
  assign n45633 = n2302 | n7560 ;
  assign n45634 = n7560 & ~n45633 ;
  assign n45635 = n8762 & ~n45634 ;
  assign n45636 = n45632 & n45635 ;
  assign n45637 = n10866 | n45636 ;
  assign n45638 = n45636 & ~n45637 ;
  assign n45639 = n12569 | n45638 ;
  assign n45640 = n12569 & ~n45639 ;
  assign n45641 = ( n21256 & n45630 ) | ( n21256 & ~n45640 ) | ( n45630 & ~n45640 ) ;
  assign n45629 = n37608 ^ n21431 ^ 1'b0 ;
  assign n45642 = n45641 ^ n45629 ^ n8254 ;
  assign n45643 = n29612 ^ n16344 ^ n3188 ;
  assign n45644 = n40221 ^ n30367 ^ n1347 ;
  assign n45645 = n45644 ^ n39244 ^ n23156 ;
  assign n45646 = ( n6596 & ~n18651 ) | ( n6596 & n20538 ) | ( ~n18651 & n20538 ) ;
  assign n45647 = n45646 ^ n43710 ^ n7460 ;
  assign n45648 = n7512 | n15006 ;
  assign n45649 = n24968 ^ n13126 ^ n2196 ;
  assign n45650 = ( n1082 & n23470 ) | ( n1082 & ~n45649 ) | ( n23470 & ~n45649 ) ;
  assign n45651 = n14027 & n22854 ;
  assign n45652 = n21429 & n45651 ;
  assign n45653 = n15701 | n45652 ;
  assign n45654 = n45650 & ~n45653 ;
  assign n45656 = ( n5318 & n6931 ) | ( n5318 & ~n8843 ) | ( n6931 & ~n8843 ) ;
  assign n45657 = n45656 ^ n31432 ^ n19711 ;
  assign n45658 = n32125 & n45657 ;
  assign n45655 = n7481 & n24096 ;
  assign n45659 = n45658 ^ n45655 ^ 1'b0 ;
  assign n45663 = ~n11366 & n13645 ;
  assign n45660 = ~n10429 & n11936 ;
  assign n45661 = n2423 & n45660 ;
  assign n45662 = n32172 | n45661 ;
  assign n45664 = n45663 ^ n45662 ^ 1'b0 ;
  assign n45665 = ~n3194 & n43696 ;
  assign n45666 = n41832 ^ n1320 ^ 1'b0 ;
  assign n45667 = n45666 ^ n24868 ^ 1'b0 ;
  assign n45668 = ( n12779 & ~n17292 ) | ( n12779 & n39161 ) | ( ~n17292 & n39161 ) ;
  assign n45669 = n3391 & ~n45668 ;
  assign n45670 = n20752 ^ n17068 ^ n16743 ;
  assign n45671 = x73 | n45670 ;
  assign n45672 = ( n7582 & ~n16254 ) | ( n7582 & n45671 ) | ( ~n16254 & n45671 ) ;
  assign n45673 = n17284 ^ n3125 ^ 1'b0 ;
  assign n45674 = n5441 & n45673 ;
  assign n45675 = n44415 ^ n29652 ^ 1'b0 ;
  assign n45676 = ~n15272 & n23672 ;
  assign n45677 = n45675 & n45676 ;
  assign n45678 = n31168 & ~n45677 ;
  assign n45679 = n10450 ^ n6003 ^ 1'b0 ;
  assign n45680 = n26049 & ~n45679 ;
  assign n45681 = ~n1482 & n37470 ;
  assign n45682 = ~n32006 & n45681 ;
  assign n45683 = n45682 ^ x44 ^ 1'b0 ;
  assign n45684 = n44652 | n45683 ;
  assign n45685 = n12297 | n18004 ;
  assign n45686 = n39041 | n45685 ;
  assign n45687 = ( n3581 & ~n21437 ) | ( n3581 & n45686 ) | ( ~n21437 & n45686 ) ;
  assign n45688 = ( n1190 & n17319 ) | ( n1190 & n22816 ) | ( n17319 & n22816 ) ;
  assign n45689 = n19996 & ~n45688 ;
  assign n45696 = ( ~n14014 & n15411 ) | ( ~n14014 & n16345 ) | ( n15411 & n16345 ) ;
  assign n45693 = n20626 ^ n8626 ^ 1'b0 ;
  assign n45694 = n8669 ^ x176 ^ 1'b0 ;
  assign n45695 = ~n45693 & n45694 ;
  assign n45690 = n31047 ^ n27707 ^ 1'b0 ;
  assign n45691 = ~n11875 & n13139 ;
  assign n45692 = n45690 & ~n45691 ;
  assign n45697 = n45696 ^ n45695 ^ n45692 ;
  assign n45698 = n28181 ^ n13041 ^ n11177 ;
  assign n45699 = n8047 ^ n1377 ^ x187 ;
  assign n45700 = n34570 & n45699 ;
  assign n45701 = n45700 ^ n4919 ^ 1'b0 ;
  assign n45702 = n31421 & n45701 ;
  assign n45706 = n29338 ^ n13402 ^ n9342 ;
  assign n45703 = ~n23785 & n36203 ;
  assign n45704 = n45703 ^ n19954 ^ 1'b0 ;
  assign n45705 = ( ~n6216 & n11368 ) | ( ~n6216 & n45704 ) | ( n11368 & n45704 ) ;
  assign n45707 = n45706 ^ n45705 ^ 1'b0 ;
  assign n45708 = ~n2039 & n44977 ;
  assign n45709 = n45708 ^ n4154 ^ 1'b0 ;
  assign n45710 = n16349 ^ n6781 ^ 1'b0 ;
  assign n45711 = n13453 & n45710 ;
  assign n45716 = n8621 & ~n9658 ;
  assign n45717 = n5298 & n45716 ;
  assign n45712 = n6302 & n16998 ;
  assign n45713 = n24173 & n45712 ;
  assign n45714 = n43719 | n45713 ;
  assign n45715 = n11152 | n45714 ;
  assign n45718 = n45717 ^ n45715 ^ n3305 ;
  assign n45724 = x161 & ~n3288 ;
  assign n45725 = ~x161 & n45724 ;
  assign n45720 = n15316 & n17887 ;
  assign n45721 = n45720 ^ n1369 ^ 1'b0 ;
  assign n45722 = ( ~x150 & n7800 ) | ( ~x150 & n45721 ) | ( n7800 & n45721 ) ;
  assign n45719 = ~n9729 & n36411 ;
  assign n45723 = n45722 ^ n45719 ^ 1'b0 ;
  assign n45726 = n45725 ^ n45723 ^ n4214 ;
  assign n45727 = n21789 ^ n14562 ^ n4542 ;
  assign n45728 = ~n10298 & n45727 ;
  assign n45736 = ( n9212 & ~n12764 ) | ( n9212 & n13505 ) | ( ~n12764 & n13505 ) ;
  assign n45737 = ~n35965 & n45736 ;
  assign n45729 = n26546 ^ n6313 ^ 1'b0 ;
  assign n45730 = n36687 & n45729 ;
  assign n45731 = n2516 & ~n26228 ;
  assign n45732 = ~n45730 & n45731 ;
  assign n45733 = ~n1071 & n7657 ;
  assign n45734 = n45732 & n45733 ;
  assign n45735 = n38605 | n45734 ;
  assign n45738 = n45737 ^ n45735 ^ 1'b0 ;
  assign n45739 = n22048 & ~n40366 ;
  assign n45740 = ~n322 & n38745 ;
  assign n45741 = n45740 ^ n4341 ^ 1'b0 ;
  assign n45742 = n45741 ^ n5257 ^ 1'b0 ;
  assign n45743 = n11387 | n45742 ;
  assign n45744 = n3690 | n45743 ;
  assign n45745 = n12408 & n12522 ;
  assign n45746 = n40639 & n45745 ;
  assign n45747 = n41500 ^ n28681 ^ n26920 ;
  assign n45748 = n39827 ^ n29876 ^ n4544 ;
  assign n45749 = ~n2910 & n12343 ;
  assign n45750 = n45749 ^ n29802 ^ n9102 ;
  assign n45751 = n19079 & n27377 ;
  assign n45752 = n45751 ^ n18757 ^ 1'b0 ;
  assign n45753 = n5637 | n45752 ;
  assign n45754 = n10121 ^ n6742 ^ 1'b0 ;
  assign n45755 = n25618 & n45754 ;
  assign n45756 = n45755 ^ n12872 ^ 1'b0 ;
  assign n45757 = n2727 ^ n2411 ^ n1386 ;
  assign n45758 = ~n45756 & n45757 ;
  assign n45759 = ( ~n12415 & n14138 ) | ( ~n12415 & n36863 ) | ( n14138 & n36863 ) ;
  assign n45760 = n6644 & n28768 ;
  assign n45761 = ( n4901 & n10620 ) | ( n4901 & n27269 ) | ( n10620 & n27269 ) ;
  assign n45762 = n887 | n28437 ;
  assign n45763 = n45762 ^ n33742 ^ n20750 ;
  assign n45764 = n39759 & n45763 ;
  assign n45766 = n10894 | n11897 ;
  assign n45765 = n10654 | n42412 ;
  assign n45767 = n45766 ^ n45765 ^ n3516 ;
  assign n45768 = n45349 ^ n35076 ^ 1'b0 ;
  assign n45769 = n45767 | n45768 ;
  assign n45770 = n12041 & n36737 ;
  assign n45771 = n45770 ^ n24400 ^ 1'b0 ;
  assign n45772 = ~n6988 & n40500 ;
  assign n45773 = ~n16342 & n45772 ;
  assign n45774 = n12836 & ~n21983 ;
  assign n45775 = n45774 ^ n2173 ^ 1'b0 ;
  assign n45776 = n45775 ^ n10211 ^ n5868 ;
  assign n45777 = n8218 ^ n1680 ^ 1'b0 ;
  assign n45778 = ~n12255 & n45777 ;
  assign n45779 = n45778 ^ n23069 ^ n5681 ;
  assign n45780 = n23224 ^ n8171 ^ n7586 ;
  assign n45781 = ( ~n17537 & n39538 ) | ( ~n17537 & n45089 ) | ( n39538 & n45089 ) ;
  assign n45782 = n9799 & ~n16402 ;
  assign n45783 = n44917 | n45782 ;
  assign n45784 = n25184 & ~n45783 ;
  assign n45785 = n259 & ~n23351 ;
  assign n45786 = n6950 & ~n21380 ;
  assign n45787 = ~n23907 & n45786 ;
  assign n45788 = n45787 ^ n15130 ^ 1'b0 ;
  assign n45789 = n28719 ^ n27537 ^ 1'b0 ;
  assign n45790 = n43955 ^ n8431 ^ 1'b0 ;
  assign n45791 = n45789 & n45790 ;
  assign n45792 = n2791 & n26783 ;
  assign n45793 = n1232 & n22854 ;
  assign n45794 = ~n39432 & n45793 ;
  assign n45795 = n27655 ^ n5039 ^ 1'b0 ;
  assign n45796 = ( n3312 & ~n25080 ) | ( n3312 & n45795 ) | ( ~n25080 & n45795 ) ;
  assign n45797 = n21354 ^ n6656 ^ 1'b0 ;
  assign n45798 = ~n30196 & n45797 ;
  assign n45799 = ~n39530 & n45798 ;
  assign n45800 = n4128 | n7850 ;
  assign n45801 = n40649 & n45800 ;
  assign n45802 = n7691 ^ n3361 ^ n1893 ;
  assign n45803 = n26268 & n45802 ;
  assign n45804 = n45803 ^ n2088 ^ 1'b0 ;
  assign n45805 = n11315 | n45804 ;
  assign n45806 = n5544 & ~n5928 ;
  assign n45807 = n45806 ^ n10535 ^ 1'b0 ;
  assign n45808 = n2164 | n22030 ;
  assign n45809 = n37608 | n45808 ;
  assign n45810 = n26780 ^ n6627 ^ 1'b0 ;
  assign n45815 = ~n12190 & n43362 ;
  assign n45816 = ~n23223 & n45815 ;
  assign n45811 = n28118 ^ n15537 ^ n3932 ;
  assign n45812 = ( x24 & n949 ) | ( x24 & ~n3702 ) | ( n949 & ~n3702 ) ;
  assign n45813 = ( n37729 & n45811 ) | ( n37729 & n45812 ) | ( n45811 & n45812 ) ;
  assign n45814 = n15614 | n45813 ;
  assign n45817 = n45816 ^ n45814 ^ 1'b0 ;
  assign n45818 = n7302 & ~n9927 ;
  assign n45819 = n24651 & n45818 ;
  assign n45820 = ( n31044 & n33339 ) | ( n31044 & ~n45819 ) | ( n33339 & ~n45819 ) ;
  assign n45821 = n17619 ^ n11601 ^ 1'b0 ;
  assign n45822 = n15873 & n45821 ;
  assign n45823 = n13202 | n39740 ;
  assign n45824 = n25666 & ~n45823 ;
  assign n45825 = ( n15528 & n17837 ) | ( n15528 & n21111 ) | ( n17837 & n21111 ) ;
  assign n45826 = n45825 ^ n23148 ^ 1'b0 ;
  assign n45827 = ( n7070 & n9161 ) | ( n7070 & ~n11518 ) | ( n9161 & ~n11518 ) ;
  assign n45828 = n36380 ^ n7331 ^ 1'b0 ;
  assign n45829 = n24611 & ~n45828 ;
  assign n45830 = n16653 & n45488 ;
  assign n45831 = n45829 | n45830 ;
  assign n45832 = n19004 ^ n6738 ^ n3609 ;
  assign n45833 = n8094 ^ n1369 ^ 1'b0 ;
  assign n45834 = n8005 | n45833 ;
  assign n45835 = n27754 | n38922 ;
  assign n45836 = n18380 & ~n22367 ;
  assign n45837 = n28750 ^ n21866 ^ 1'b0 ;
  assign n45838 = ( ~n6908 & n16080 ) | ( ~n6908 & n16366 ) | ( n16080 & n16366 ) ;
  assign n45839 = n45838 ^ n5454 ^ 1'b0 ;
  assign n45840 = ~n45837 & n45839 ;
  assign n45841 = n41329 ^ n26747 ^ 1'b0 ;
  assign n45844 = ~n1885 & n13278 ;
  assign n45842 = n21020 | n34559 ;
  assign n45843 = n35014 & ~n45842 ;
  assign n45845 = n45844 ^ n45843 ^ 1'b0 ;
  assign n45846 = n16847 ^ n5377 ^ 1'b0 ;
  assign n45847 = n33287 & n45846 ;
  assign n45848 = n9287 ^ n1285 ^ 1'b0 ;
  assign n45849 = n45847 & ~n45848 ;
  assign n45850 = n45849 ^ n25098 ^ 1'b0 ;
  assign n45851 = n10970 & n29136 ;
  assign n45852 = ~n23279 & n31507 ;
  assign n45853 = n5609 ^ n4361 ^ 1'b0 ;
  assign n45854 = n13498 | n45853 ;
  assign n45855 = n2192 & ~n41254 ;
  assign n45856 = n12624 & ~n39162 ;
  assign n45857 = n5030 & n41554 ;
  assign n45858 = ~n10804 & n45857 ;
  assign n45859 = n27050 ^ n17202 ^ x90 ;
  assign n45860 = ( n6250 & n9187 ) | ( n6250 & ~n30960 ) | ( n9187 & ~n30960 ) ;
  assign n45863 = ~n3981 & n22023 ;
  assign n45864 = n45863 ^ n9344 ^ 1'b0 ;
  assign n45861 = n5394 & n9063 ;
  assign n45862 = n45861 ^ n31749 ^ 1'b0 ;
  assign n45865 = n45864 ^ n45862 ^ n34543 ;
  assign n45867 = n4118 & n13361 ;
  assign n45868 = ~n16846 & n45867 ;
  assign n45866 = n1144 | n4067 ;
  assign n45869 = n45868 ^ n45866 ^ 1'b0 ;
  assign n45870 = n3687 & ~n8116 ;
  assign n45871 = ( n14618 & n32572 ) | ( n14618 & ~n45870 ) | ( n32572 & ~n45870 ) ;
  assign n45872 = ( n9068 & n15075 ) | ( n9068 & n45871 ) | ( n15075 & n45871 ) ;
  assign n45873 = n4237 & ~n45872 ;
  assign n45874 = n39001 ^ n2643 ^ 1'b0 ;
  assign n45875 = ( n6341 & ~n18992 ) | ( n6341 & n45874 ) | ( ~n18992 & n45874 ) ;
  assign n45876 = n24754 & ~n38869 ;
  assign n45877 = n6537 & n45876 ;
  assign n45878 = n45437 | n45877 ;
  assign n45879 = n45875 & ~n45878 ;
  assign n45880 = n8563 ^ n7807 ^ 1'b0 ;
  assign n45881 = ~n16187 & n45880 ;
  assign n45882 = n33519 ^ n20075 ^ n8454 ;
  assign n45883 = ( n13082 & ~n29878 ) | ( n13082 & n45500 ) | ( ~n29878 & n45500 ) ;
  assign n45884 = ( ~n10902 & n13968 ) | ( ~n10902 & n21768 ) | ( n13968 & n21768 ) ;
  assign n45885 = ( ~n4529 & n6088 ) | ( ~n4529 & n8966 ) | ( n6088 & n8966 ) ;
  assign n45886 = n23207 | n45668 ;
  assign n45887 = n45886 ^ n2600 ^ 1'b0 ;
  assign n45888 = n28863 & n34057 ;
  assign n45889 = n38515 & n45888 ;
  assign n45890 = ~n21743 & n28790 ;
  assign n45891 = n45890 ^ n20979 ^ 1'b0 ;
  assign n45892 = n4930 | n5151 ;
  assign n45893 = n14127 ^ n7584 ^ 1'b0 ;
  assign n45894 = n45892 & ~n45893 ;
  assign n45895 = n10774 & ~n45894 ;
  assign n45896 = ( ~n325 & n3592 ) | ( ~n325 & n20327 ) | ( n3592 & n20327 ) ;
  assign n45897 = n2573 & n13821 ;
  assign n45900 = n11852 & n35769 ;
  assign n45898 = n19267 ^ n3564 ^ 1'b0 ;
  assign n45899 = n45898 ^ n19801 ^ n18884 ;
  assign n45901 = n45900 ^ n45899 ^ 1'b0 ;
  assign n45902 = ( n27923 & n34910 ) | ( n27923 & n45901 ) | ( n34910 & n45901 ) ;
  assign n45903 = n8328 | n13877 ;
  assign n45904 = ~n2690 & n40810 ;
  assign n45905 = n15130 | n45904 ;
  assign n45906 = n45903 | n45905 ;
  assign n45907 = n1963 & n5311 ;
  assign n45908 = n15392 & n45907 ;
  assign n45909 = n4827 | n10645 ;
  assign n45910 = n1981 & ~n45909 ;
  assign n45911 = n5334 & ~n25100 ;
  assign n45912 = n32253 ^ n21098 ^ 1'b0 ;
  assign n45913 = n6645 & n35951 ;
  assign n45914 = n16286 & n45913 ;
  assign n45915 = n19994 | n33327 ;
  assign n45916 = n20342 ^ n4411 ^ 1'b0 ;
  assign n45917 = n11934 & ~n45916 ;
  assign n45918 = ( n40740 & ~n44487 ) | ( n40740 & n45917 ) | ( ~n44487 & n45917 ) ;
  assign n45919 = ( n13566 & ~n28214 ) | ( n13566 & n28982 ) | ( ~n28214 & n28982 ) ;
  assign n45920 = ( n5261 & n12667 ) | ( n5261 & ~n36895 ) | ( n12667 & ~n36895 ) ;
  assign n45921 = n14598 ^ n12241 ^ n12164 ;
  assign n45922 = n45921 ^ n29443 ^ n11405 ;
  assign n45923 = n45922 ^ n10984 ^ 1'b0 ;
  assign n45924 = n35411 ^ n3991 ^ 1'b0 ;
  assign n45925 = n14510 | n45924 ;
  assign n45926 = n23831 | n34153 ;
  assign n45927 = n6703 ^ n5413 ^ 1'b0 ;
  assign n45928 = ~n45926 & n45927 ;
  assign n45929 = n15841 & ~n28441 ;
  assign n45930 = n13877 & ~n21303 ;
  assign n45931 = n8160 & n45930 ;
  assign n45932 = n7051 & ~n39290 ;
  assign n45933 = n34230 | n45932 ;
  assign n45934 = n45933 ^ n26141 ^ 1'b0 ;
  assign n45935 = n45806 ^ n7327 ^ 1'b0 ;
  assign n45936 = n13848 & n44385 ;
  assign n45937 = n45936 ^ n13607 ^ 1'b0 ;
  assign n45938 = n26945 & n45937 ;
  assign n45939 = n20219 & n45938 ;
  assign n45940 = n8278 ^ n4130 ^ 1'b0 ;
  assign n45941 = ~n10894 & n45940 ;
  assign n45942 = n11223 | n45941 ;
  assign n45943 = ( n5992 & n11370 ) | ( n5992 & ~n31630 ) | ( n11370 & ~n31630 ) ;
  assign n45944 = n27886 & n45943 ;
  assign n45945 = ( n15037 & n45942 ) | ( n15037 & ~n45944 ) | ( n45942 & ~n45944 ) ;
  assign n45946 = n20597 ^ n11330 ^ 1'b0 ;
  assign n45947 = n45946 ^ n30367 ^ n6472 ;
  assign n45948 = n31888 & ~n33891 ;
  assign n45949 = ( n9685 & n9860 ) | ( n9685 & n35453 ) | ( n9860 & n35453 ) ;
  assign n45950 = n3096 & ~n17321 ;
  assign n45951 = ~n22092 & n45950 ;
  assign n45952 = n45951 ^ n44476 ^ 1'b0 ;
  assign n45953 = ~n34722 & n45952 ;
  assign n45954 = n12616 | n13658 ;
  assign n45955 = n45954 ^ n31121 ^ 1'b0 ;
  assign n45956 = n11571 & ~n12704 ;
  assign n45957 = ~n16452 & n45956 ;
  assign n45958 = n16346 ^ n343 ^ 1'b0 ;
  assign n45959 = n13597 & ~n45958 ;
  assign n45960 = ~n25861 & n36752 ;
  assign n45961 = n45959 & n45960 ;
  assign n45962 = n12260 ^ n1733 ^ 1'b0 ;
  assign n45963 = ~n39209 & n45962 ;
  assign n45964 = ~n4793 & n45963 ;
  assign n45965 = n7664 & ~n16083 ;
  assign n45966 = n30686 ^ n21421 ^ n17673 ;
  assign n45967 = ( n31370 & n45965 ) | ( n31370 & ~n45966 ) | ( n45965 & ~n45966 ) ;
  assign n45968 = n1989 | n17340 ;
  assign n45969 = n45968 ^ n16706 ^ 1'b0 ;
  assign n45970 = ~n5056 & n5467 ;
  assign n45971 = ~n23123 & n45970 ;
  assign n45972 = ~n5839 & n45971 ;
  assign n45973 = n45969 & ~n45972 ;
  assign n45974 = n18731 & ~n19627 ;
  assign n45975 = n8685 & n45974 ;
  assign n45976 = n8792 & ~n34219 ;
  assign n45977 = n24002 & n45976 ;
  assign n45978 = ( n7142 & n45975 ) | ( n7142 & ~n45977 ) | ( n45975 & ~n45977 ) ;
  assign n45979 = ( ~n1182 & n12476 ) | ( ~n1182 & n45978 ) | ( n12476 & n45978 ) ;
  assign n45980 = n13085 ^ n11749 ^ 1'b0 ;
  assign n45981 = n40564 | n45980 ;
  assign n45982 = n15892 ^ n4055 ^ 1'b0 ;
  assign n45983 = n6084 & ~n45982 ;
  assign n45984 = n19753 ^ n13104 ^ 1'b0 ;
  assign n45985 = n2445 & n43178 ;
  assign n45986 = n34568 & ~n45985 ;
  assign n45987 = n24664 ^ n8085 ^ n1476 ;
  assign n45988 = n45986 & ~n45987 ;
  assign n45989 = n36883 ^ n18349 ^ 1'b0 ;
  assign n45990 = ~n28262 & n45989 ;
  assign n45991 = n36990 ^ n21769 ^ n9282 ;
  assign n45992 = n19839 ^ n7079 ^ n1492 ;
  assign n45993 = n45992 ^ n39109 ^ 1'b0 ;
  assign n45994 = ~n6990 & n45993 ;
  assign n45995 = n5520 & n45994 ;
  assign n45996 = n23450 & ~n45995 ;
  assign n45997 = ( n8387 & n42134 ) | ( n8387 & ~n45996 ) | ( n42134 & ~n45996 ) ;
  assign n45998 = n40040 ^ n23710 ^ 1'b0 ;
  assign n45999 = n1674 | n45998 ;
  assign n46000 = n39653 | n45999 ;
  assign n46001 = n44526 ^ n4132 ^ n2849 ;
  assign n46002 = n46001 ^ n45171 ^ n40210 ;
  assign n46003 = n36642 & ~n39935 ;
  assign n46004 = n40197 ^ n11870 ^ 1'b0 ;
  assign n46005 = ~x102 & n15327 ;
  assign n46006 = x226 & ~n46005 ;
  assign n46007 = n46006 ^ n41990 ^ 1'b0 ;
  assign n46008 = n3739 & ~n8042 ;
  assign n46009 = n17263 & n46008 ;
  assign n46010 = n46009 ^ n3386 ^ 1'b0 ;
  assign n46011 = n28225 | n46010 ;
  assign n46012 = n25124 ^ n7986 ^ 1'b0 ;
  assign n46013 = n30882 & n46012 ;
  assign n46014 = n10926 & n46013 ;
  assign n46015 = ~n4428 & n46014 ;
  assign n46016 = n354 | n46015 ;
  assign n46017 = n20570 & ~n46016 ;
  assign n46018 = n1327 & ~n31108 ;
  assign n46019 = ~n41942 & n46018 ;
  assign n46020 = ( n11056 & n37053 ) | ( n11056 & n39023 ) | ( n37053 & n39023 ) ;
  assign n46021 = n43549 ^ n32673 ^ n7035 ;
  assign n46022 = n35513 & ~n36677 ;
  assign n46023 = ( n1877 & ~n18032 ) | ( n1877 & n46022 ) | ( ~n18032 & n46022 ) ;
  assign n46024 = n11673 | n21073 ;
  assign n46025 = n16564 | n46024 ;
  assign n46026 = ~n19762 & n20950 ;
  assign n46027 = n16213 & n46026 ;
  assign n46028 = n8313 & ~n19065 ;
  assign n46029 = n21985 & ~n39102 ;
  assign n46030 = ~n24542 & n46029 ;
  assign n46031 = ( n5872 & n9534 ) | ( n5872 & ~n18853 ) | ( n9534 & ~n18853 ) ;
  assign n46032 = n46031 ^ n8254 ^ 1'b0 ;
  assign n46033 = n46030 & ~n46032 ;
  assign n46034 = ( ~n5246 & n7044 ) | ( ~n5246 & n34443 ) | ( n7044 & n34443 ) ;
  assign n46035 = n46034 ^ n11715 ^ n8129 ;
  assign n46036 = n19734 | n27047 ;
  assign n46037 = n46036 ^ n22907 ^ 1'b0 ;
  assign n46038 = ~n9861 & n21080 ;
  assign n46039 = n8026 & n46038 ;
  assign n46040 = n42834 | n46039 ;
  assign n46041 = n8306 & n18176 ;
  assign n46042 = n10524 & n46041 ;
  assign n46043 = n1107 & ~n3430 ;
  assign n46044 = n21561 & n36116 ;
  assign n46045 = n24160 ^ n18333 ^ 1'b0 ;
  assign n46046 = n14444 | n46045 ;
  assign n46047 = n46046 ^ n31952 ^ 1'b0 ;
  assign n46048 = ~n46044 & n46047 ;
  assign n46050 = ( n1050 & n12761 ) | ( n1050 & ~n24375 ) | ( n12761 & ~n24375 ) ;
  assign n46049 = ( n22090 & n35526 ) | ( n22090 & ~n40887 ) | ( n35526 & ~n40887 ) ;
  assign n46051 = n46050 ^ n46049 ^ n30398 ;
  assign n46052 = n41852 ^ n34916 ^ 1'b0 ;
  assign n46053 = ~n5598 & n46052 ;
  assign n46054 = n46053 ^ n34525 ^ n4458 ;
  assign n46055 = ~n3851 & n6517 ;
  assign n46056 = ( n29961 & n31014 ) | ( n29961 & ~n46055 ) | ( n31014 & ~n46055 ) ;
  assign n46057 = ( n6821 & n8517 ) | ( n6821 & ~n26179 ) | ( n8517 & ~n26179 ) ;
  assign n46058 = n15914 ^ n11531 ^ 1'b0 ;
  assign n46059 = n46058 ^ n13543 ^ 1'b0 ;
  assign n46060 = ~n46057 & n46059 ;
  assign n46061 = n37178 ^ x123 ^ 1'b0 ;
  assign n46062 = n28717 ^ n28482 ^ 1'b0 ;
  assign n46063 = n9615 | n38270 ;
  assign n46064 = n46063 ^ n25320 ^ 1'b0 ;
  assign n46065 = n3247 & n15877 ;
  assign n46066 = n46065 ^ n1716 ^ 1'b0 ;
  assign n46067 = n46066 ^ n28681 ^ n12834 ;
  assign n46068 = n46067 ^ n44765 ^ n35451 ;
  assign n46069 = n21583 | n30740 ;
  assign n46070 = n38115 ^ n24911 ^ 1'b0 ;
  assign n46071 = n3256 & ~n36304 ;
  assign n46072 = n4890 & n46071 ;
  assign n46073 = n19519 | n45603 ;
  assign n46074 = n11559 | n46073 ;
  assign n46078 = ~n3044 & n7649 ;
  assign n46075 = ( n6310 & n8453 ) | ( n6310 & n18850 ) | ( n8453 & n18850 ) ;
  assign n46076 = ( n4469 & n34271 ) | ( n4469 & ~n46075 ) | ( n34271 & ~n46075 ) ;
  assign n46077 = n8275 | n46076 ;
  assign n46079 = n46078 ^ n46077 ^ 1'b0 ;
  assign n46080 = n6699 ^ n6556 ^ n637 ;
  assign n46081 = ~n24150 & n46080 ;
  assign n46082 = n36960 ^ n15590 ^ 1'b0 ;
  assign n46083 = ~n24784 & n46082 ;
  assign n46084 = n19476 & ~n29578 ;
  assign n46085 = n46084 ^ n30655 ^ 1'b0 ;
  assign n46086 = n5022 & n9099 ;
  assign n46087 = n9872 & n46086 ;
  assign n46088 = n46085 & n46087 ;
  assign n46089 = ( n31806 & n36781 ) | ( n31806 & ~n46088 ) | ( n36781 & ~n46088 ) ;
  assign n46090 = n33315 & ~n41420 ;
  assign n46091 = n10919 | n46090 ;
  assign n46092 = n46091 ^ n42803 ^ 1'b0 ;
  assign n46093 = ~n9899 & n24902 ;
  assign n46094 = ~n21181 & n46093 ;
  assign n46099 = ~n1299 & n40588 ;
  assign n46095 = n4569 & ~n24319 ;
  assign n46096 = n13863 & n46095 ;
  assign n46097 = n9299 & ~n24991 ;
  assign n46098 = ( n6218 & n46096 ) | ( n6218 & ~n46097 ) | ( n46096 & ~n46097 ) ;
  assign n46100 = n46099 ^ n46098 ^ n493 ;
  assign n46101 = n14430 | n27024 ;
  assign n46102 = n46101 ^ n34489 ^ 1'b0 ;
  assign n46103 = n5389 | n46102 ;
  assign n46104 = ~n4314 & n7794 ;
  assign n46105 = n46104 ^ n44313 ^ n14999 ;
  assign n46106 = ( n654 & n1030 ) | ( n654 & n36154 ) | ( n1030 & n36154 ) ;
  assign n46107 = n33752 ^ n27737 ^ 1'b0 ;
  assign n46108 = n14151 & n46107 ;
  assign n46109 = n4227 | n27393 ;
  assign n46110 = n39664 ^ n6190 ^ n2209 ;
  assign n46111 = ~n18732 & n39571 ;
  assign n46112 = n11766 & n35805 ;
  assign n46113 = n46111 & n46112 ;
  assign n46114 = n27712 ^ n10543 ^ 1'b0 ;
  assign n46115 = n14796 & ~n46114 ;
  assign n46116 = n40146 ^ n15964 ^ 1'b0 ;
  assign n46117 = n14721 | n46116 ;
  assign n46118 = n21857 ^ n19480 ^ 1'b0 ;
  assign n46119 = n46118 ^ n44405 ^ n3900 ;
  assign n46122 = n2449 | n7135 ;
  assign n46120 = n18825 & ~n19507 ;
  assign n46121 = n9261 | n46120 ;
  assign n46123 = n46122 ^ n46121 ^ 1'b0 ;
  assign n46124 = n41552 ^ n1844 ^ 1'b0 ;
  assign n46126 = n27912 | n31058 ;
  assign n46127 = n46126 ^ n31209 ^ 1'b0 ;
  assign n46125 = n2394 & n3300 ;
  assign n46128 = n46127 ^ n46125 ^ 1'b0 ;
  assign n46129 = n7965 & ~n30245 ;
  assign n46133 = ( ~n8651 & n12906 ) | ( ~n8651 & n16882 ) | ( n12906 & n16882 ) ;
  assign n46130 = n483 & n39789 ;
  assign n46131 = ~n33653 & n46130 ;
  assign n46132 = n5360 | n46131 ;
  assign n46134 = n46133 ^ n46132 ^ 1'b0 ;
  assign n46135 = n12194 ^ n6172 ^ n1367 ;
  assign n46136 = n46135 ^ n11400 ^ 1'b0 ;
  assign n46137 = n16152 | n36966 ;
  assign n46138 = ( n14529 & n19731 ) | ( n14529 & n46137 ) | ( n19731 & n46137 ) ;
  assign n46139 = n1817 | n10696 ;
  assign n46140 = n46139 ^ n5976 ^ n4561 ;
  assign n46141 = n46140 ^ n10787 ^ 1'b0 ;
  assign n46142 = ~x198 & n46141 ;
  assign n46143 = n18463 & n34149 ;
  assign n46144 = n18488 & n46143 ;
  assign n46145 = n17821 ^ n1050 ^ 1'b0 ;
  assign n46146 = n11363 & n46145 ;
  assign n46147 = n41667 ^ n19176 ^ 1'b0 ;
  assign n46148 = n4322 & ~n46147 ;
  assign n46149 = n23391 & n46148 ;
  assign n46150 = ( n9816 & ~n18487 ) | ( n9816 & n46149 ) | ( ~n18487 & n46149 ) ;
  assign n46151 = n46150 ^ n8996 ^ 1'b0 ;
  assign n46152 = ( ~n4214 & n37933 ) | ( ~n4214 & n38391 ) | ( n37933 & n38391 ) ;
  assign n46153 = n17068 ^ n16649 ^ 1'b0 ;
  assign n46154 = n2529 | n46153 ;
  assign n46155 = n2827 & n39329 ;
  assign n46156 = n46155 ^ n21238 ^ 1'b0 ;
  assign n46158 = n20323 & ~n42851 ;
  assign n46159 = ~n46127 & n46158 ;
  assign n46157 = n17022 & ~n38709 ;
  assign n46160 = n46159 ^ n46157 ^ 1'b0 ;
  assign n46161 = n18202 ^ n4522 ^ 1'b0 ;
  assign n46162 = n15211 & ~n46161 ;
  assign n46163 = ~n37511 & n44707 ;
  assign n46164 = ( x110 & n12630 ) | ( x110 & ~n24553 ) | ( n12630 & ~n24553 ) ;
  assign n46165 = ~n1176 & n1760 ;
  assign n46166 = n46165 ^ n7732 ^ 1'b0 ;
  assign n46167 = n20752 ^ n14648 ^ 1'b0 ;
  assign n46168 = ~n46166 & n46167 ;
  assign n46169 = n46168 ^ n25993 ^ n6422 ;
  assign n46170 = n36593 ^ n8278 ^ 1'b0 ;
  assign n46171 = ~n16624 & n46170 ;
  assign n46172 = n46171 ^ n38413 ^ n20166 ;
  assign n46173 = n42964 ^ n11933 ^ 1'b0 ;
  assign n46174 = n15681 & ~n24909 ;
  assign n46175 = n5330 & ~n46174 ;
  assign n46178 = n40151 ^ n17758 ^ 1'b0 ;
  assign n46176 = n13437 ^ n2005 ^ n1985 ;
  assign n46177 = n36999 & n46176 ;
  assign n46179 = n46178 ^ n46177 ^ 1'b0 ;
  assign n46180 = n3766 & n28185 ;
  assign n46182 = n7753 ^ n1489 ^ 1'b0 ;
  assign n46181 = n2414 & n22131 ;
  assign n46183 = n46182 ^ n46181 ^ 1'b0 ;
  assign n46184 = n46183 ^ n19364 ^ 1'b0 ;
  assign n46185 = n45374 | n46184 ;
  assign n46186 = n22021 & ~n42650 ;
  assign n46187 = n17930 & n46186 ;
  assign n46188 = n15884 ^ n5056 ^ 1'b0 ;
  assign n46189 = n11667 & n46188 ;
  assign n46190 = n34911 ^ n3624 ^ 1'b0 ;
  assign n46191 = n1669 & n38965 ;
  assign n46192 = n46191 ^ n36299 ^ 1'b0 ;
  assign n46193 = ( n23563 & n26788 ) | ( n23563 & ~n37959 ) | ( n26788 & ~n37959 ) ;
  assign n46194 = ( n13497 & n46192 ) | ( n13497 & n46193 ) | ( n46192 & n46193 ) ;
  assign n46195 = n15568 | n21421 ;
  assign n46196 = n40561 ^ n11104 ^ n7998 ;
  assign n46197 = n37249 ^ n1256 ^ 1'b0 ;
  assign n46198 = ( n1715 & n33508 ) | ( n1715 & ~n40164 ) | ( n33508 & ~n40164 ) ;
  assign n46199 = n19317 & ~n46198 ;
  assign n46200 = n46199 ^ n18623 ^ 1'b0 ;
  assign n46201 = n22404 ^ n14679 ^ 1'b0 ;
  assign n46202 = n32437 & n46201 ;
  assign n46203 = n9637 ^ n660 ^ 1'b0 ;
  assign n46204 = n586 & ~n46203 ;
  assign n46205 = ~n4711 & n6839 ;
  assign n46206 = n46205 ^ n1025 ^ 1'b0 ;
  assign n46207 = n10509 & ~n18335 ;
  assign n46208 = n14116 & ~n46207 ;
  assign n46209 = n46208 ^ n2086 ^ 1'b0 ;
  assign n46210 = n2253 | n46209 ;
  assign n46211 = n46206 | n46210 ;
  assign n46212 = n8001 & n46211 ;
  assign n46213 = n46212 ^ n30350 ^ 1'b0 ;
  assign n46214 = ( n15699 & n15745 ) | ( n15699 & n40533 ) | ( n15745 & n40533 ) ;
  assign n46215 = n7528 & n9916 ;
  assign n46216 = n46215 ^ n8676 ^ 1'b0 ;
  assign n46217 = ( n16603 & n25166 ) | ( n16603 & n46216 ) | ( n25166 & n46216 ) ;
  assign n46218 = n29255 ^ n8690 ^ 1'b0 ;
  assign n46219 = n22413 & ~n34345 ;
  assign n46220 = ~n1580 & n46219 ;
  assign n46221 = n35648 ^ n5988 ^ n4659 ;
  assign n46222 = n21595 ^ n12703 ^ 1'b0 ;
  assign n46223 = n46221 & ~n46222 ;
  assign n46224 = n46220 | n46223 ;
  assign n46226 = n10806 ^ n2319 ^ 1'b0 ;
  assign n46227 = n40258 | n46226 ;
  assign n46225 = n21327 & ~n39443 ;
  assign n46228 = n46227 ^ n46225 ^ 1'b0 ;
  assign n46229 = ( n1024 & n1460 ) | ( n1024 & n1831 ) | ( n1460 & n1831 ) ;
  assign n46230 = n4982 ^ n4460 ^ n1961 ;
  assign n46231 = n46230 ^ n13741 ^ n12860 ;
  assign n46232 = n7721 ^ n7051 ^ 1'b0 ;
  assign n46233 = n46231 & ~n46232 ;
  assign n46234 = n46233 ^ n15875 ^ 1'b0 ;
  assign n46235 = n46229 | n46234 ;
  assign n46236 = n31715 ^ n3358 ^ n2326 ;
  assign n46237 = n2774 ^ x50 ^ 1'b0 ;
  assign n46238 = n797 & n46237 ;
  assign n46239 = n6822 | n20170 ;
  assign n46241 = n15579 | n34853 ;
  assign n46242 = n15579 & ~n46241 ;
  assign n46243 = n1969 & ~n18752 ;
  assign n46244 = n46242 & n46243 ;
  assign n46240 = n6052 | n30130 ;
  assign n46245 = n46244 ^ n46240 ^ 1'b0 ;
  assign n46246 = n46245 ^ n29684 ^ n28086 ;
  assign n46249 = n32004 ^ n20065 ^ 1'b0 ;
  assign n46250 = ( n13678 & n37729 ) | ( n13678 & n46249 ) | ( n37729 & n46249 ) ;
  assign n46247 = n12930 & n27462 ;
  assign n46248 = n41412 | n46247 ;
  assign n46251 = n46250 ^ n46248 ^ 1'b0 ;
  assign n46252 = n907 & ~n16144 ;
  assign n46253 = n41573 ^ n17167 ^ n2028 ;
  assign n46254 = n10232 | n22485 ;
  assign n46255 = n46254 ^ n24707 ^ 1'b0 ;
  assign n46256 = x176 & ~n7869 ;
  assign n46257 = ~n18374 & n46256 ;
  assign n46258 = ~n976 & n35074 ;
  assign n46259 = n46258 ^ n2936 ^ 1'b0 ;
  assign n46262 = n26478 & ~n34730 ;
  assign n46263 = n966 & n46262 ;
  assign n46260 = n1203 & ~n2083 ;
  assign n46261 = n34583 | n46260 ;
  assign n46264 = n46263 ^ n46261 ^ 1'b0 ;
  assign n46265 = n32386 ^ n9136 ^ 1'b0 ;
  assign n46266 = n21430 & ~n46265 ;
  assign n46267 = ~n2067 & n15506 ;
  assign n46268 = n46267 ^ x81 ^ 1'b0 ;
  assign n46269 = n35339 | n46268 ;
  assign n46270 = n46269 ^ n19874 ^ 1'b0 ;
  assign n46271 = n34199 & n46270 ;
  assign n46272 = ~n28780 & n46271 ;
  assign n46273 = n19293 ^ n8858 ^ 1'b0 ;
  assign n46274 = n38050 ^ n21225 ^ n444 ;
  assign n46275 = ~n36031 & n46274 ;
  assign n46276 = ~x208 & n46275 ;
  assign n46277 = n3016 & n25162 ;
  assign n46278 = n46277 ^ n403 ^ 1'b0 ;
  assign n46279 = n1327 & ~n26628 ;
  assign n46280 = n46279 ^ n33856 ^ 1'b0 ;
  assign n46281 = n21928 | n37328 ;
  assign n46282 = ~n2506 & n4034 ;
  assign n46283 = n46282 ^ n13984 ^ n7586 ;
  assign n46284 = ( n854 & ~n3817 ) | ( n854 & n4498 ) | ( ~n3817 & n4498 ) ;
  assign n46285 = n10489 ^ n862 ^ 1'b0 ;
  assign n46286 = n24464 & n27243 ;
  assign n46287 = n12112 & n14619 ;
  assign n46288 = n14082 | n46287 ;
  assign n46289 = ( ~n12470 & n25671 ) | ( ~n12470 & n25993 ) | ( n25671 & n25993 ) ;
  assign n46290 = ( n19741 & n41499 ) | ( n19741 & n46289 ) | ( n41499 & n46289 ) ;
  assign n46291 = n46288 | n46290 ;
  assign n46292 = n46286 | n46291 ;
  assign n46293 = ~n15863 & n26090 ;
  assign n46294 = n6414 & ~n27403 ;
  assign n46295 = n14448 & n46294 ;
  assign n46296 = n46293 & ~n46295 ;
  assign n46297 = n31425 & n46296 ;
  assign n46298 = n29963 & ~n35939 ;
  assign n46299 = n46298 ^ n29922 ^ 1'b0 ;
  assign n46300 = n27656 & n40596 ;
  assign n46301 = n46300 ^ n26129 ^ 1'b0 ;
  assign n46302 = n15658 ^ n10925 ^ 1'b0 ;
  assign n46303 = n11984 & ~n46302 ;
  assign n46304 = n38599 ^ n36922 ^ 1'b0 ;
  assign n46305 = n46303 & n46304 ;
  assign n46306 = n46305 ^ n1372 ^ 1'b0 ;
  assign n46307 = n22842 & n46306 ;
  assign n46308 = ~n5433 & n27801 ;
  assign n46309 = ~n27610 & n46308 ;
  assign n46310 = n46309 ^ n12989 ^ n2738 ;
  assign n46311 = ( n629 & n17948 ) | ( n629 & n36863 ) | ( n17948 & n36863 ) ;
  assign n46312 = n46311 ^ n25467 ^ 1'b0 ;
  assign n46313 = ~n14227 & n36946 ;
  assign n46314 = n2769 | n24037 ;
  assign n46315 = ~n25523 & n46314 ;
  assign n46316 = n46315 ^ n4327 ^ 1'b0 ;
  assign n46317 = ~n1365 & n2331 ;
  assign n46318 = ~x221 & n46317 ;
  assign n46319 = n14517 | n34682 ;
  assign n46320 = n26012 | n46319 ;
  assign n46321 = ~n46318 & n46320 ;
  assign n46322 = n46321 ^ n9903 ^ 1'b0 ;
  assign n46323 = n14815 ^ n1638 ^ 1'b0 ;
  assign n46324 = ~n16199 & n26541 ;
  assign n46325 = n3064 & n46324 ;
  assign n46326 = ( n11285 & n23669 ) | ( n11285 & n29123 ) | ( n23669 & n29123 ) ;
  assign n46327 = ( n11070 & n33365 ) | ( n11070 & ~n46326 ) | ( n33365 & ~n46326 ) ;
  assign n46328 = n17285 & ~n28308 ;
  assign n46329 = n46328 ^ n16403 ^ 1'b0 ;
  assign n46330 = n29068 ^ n11676 ^ 1'b0 ;
  assign n46331 = n27936 | n46330 ;
  assign n46332 = ~n7240 & n17923 ;
  assign n46333 = n15520 & ~n46332 ;
  assign n46334 = n46333 ^ n11739 ^ 1'b0 ;
  assign n46335 = n26247 & ~n46334 ;
  assign n46336 = n33434 ^ n15957 ^ 1'b0 ;
  assign n46337 = n40877 & ~n46336 ;
  assign n46338 = n13032 & n22873 ;
  assign n46339 = n8777 & n27734 ;
  assign n46340 = n38413 ^ n23807 ^ 1'b0 ;
  assign n46341 = n22691 | n32852 ;
  assign n46342 = ( n11668 & n13148 ) | ( n11668 & n23012 ) | ( n13148 & n23012 ) ;
  assign n46343 = ( ~n22221 & n46341 ) | ( ~n22221 & n46342 ) | ( n46341 & n46342 ) ;
  assign n46344 = n46343 ^ n45917 ^ n38087 ;
  assign n46345 = n38366 ^ n665 ^ x65 ;
  assign n46346 = n2830 & ~n7431 ;
  assign n46347 = n46346 ^ n17952 ^ 1'b0 ;
  assign n46348 = ~n46345 & n46347 ;
  assign n46349 = ~n18602 & n46348 ;
  assign n46350 = n40154 ^ n39326 ^ 1'b0 ;
  assign n46351 = ~n30021 & n46350 ;
  assign n46352 = n1705 & ~n5766 ;
  assign n46353 = n46352 ^ n2875 ^ 1'b0 ;
  assign n46354 = n46353 ^ n15971 ^ n3358 ;
  assign n46355 = n24673 & ~n46354 ;
  assign n46356 = n12220 & n46355 ;
  assign n46357 = n19002 & ~n43241 ;
  assign n46358 = ~n25608 & n46357 ;
  assign n46359 = n9751 & ~n19017 ;
  assign n46360 = ~x136 & n46359 ;
  assign n46361 = n29481 ^ n12217 ^ 1'b0 ;
  assign n46362 = n46360 | n46361 ;
  assign n46363 = ( ~n6728 & n40097 ) | ( ~n6728 & n40482 ) | ( n40097 & n40482 ) ;
  assign n46364 = n46363 ^ n14992 ^ 1'b0 ;
  assign n46365 = ( n9711 & n18053 ) | ( n9711 & n21983 ) | ( n18053 & n21983 ) ;
  assign n46366 = n25170 ^ n14431 ^ n2594 ;
  assign n46367 = n9887 & ~n16524 ;
  assign n46368 = ~n46366 & n46367 ;
  assign n46369 = ~n24909 & n31430 ;
  assign n46370 = n46369 ^ n24195 ^ 1'b0 ;
  assign n46371 = n28094 & n46370 ;
  assign n46372 = n10124 & ~n21093 ;
  assign n46373 = n4292 & n46372 ;
  assign n46374 = n14696 | n46373 ;
  assign n46375 = n40843 ^ n14986 ^ 1'b0 ;
  assign n46376 = ~n20269 & n39825 ;
  assign n46377 = n46375 & n46376 ;
  assign n46378 = n18991 & n31122 ;
  assign n46379 = ~n1787 & n46378 ;
  assign n46380 = n7906 ^ x224 ^ 1'b0 ;
  assign n46381 = n10080 & ~n46380 ;
  assign n46382 = n46381 ^ n32881 ^ n9100 ;
  assign n46383 = n35012 ^ n23236 ^ n1858 ;
  assign n46384 = ( ~n1234 & n5741 ) | ( ~n1234 & n37537 ) | ( n5741 & n37537 ) ;
  assign n46385 = n2901 & ~n8238 ;
  assign n46386 = n26179 ^ n24550 ^ 1'b0 ;
  assign n46387 = ~n46385 & n46386 ;
  assign n46388 = n3085 | n6986 ;
  assign n46389 = n16185 ^ n5495 ^ 1'b0 ;
  assign n46390 = n14691 | n46389 ;
  assign n46391 = n31258 ^ n11223 ^ 1'b0 ;
  assign n46392 = ~n892 & n2355 ;
  assign n46393 = n46392 ^ n4776 ^ 1'b0 ;
  assign n46394 = n11418 ^ n8252 ^ 1'b0 ;
  assign n46395 = ~n42467 & n46394 ;
  assign n46398 = n12524 ^ n4067 ^ 1'b0 ;
  assign n46399 = ~n15278 & n46398 ;
  assign n46397 = ~n3986 & n25354 ;
  assign n46400 = n46399 ^ n46397 ^ 1'b0 ;
  assign n46396 = n17901 | n44916 ;
  assign n46401 = n46400 ^ n46396 ^ 1'b0 ;
  assign n46402 = n46401 ^ n19428 ^ 1'b0 ;
  assign n46403 = ( n2032 & ~n29975 ) | ( n2032 & n43640 ) | ( ~n29975 & n43640 ) ;
  assign n46404 = n20265 & ~n35772 ;
  assign n46405 = n28129 ^ n24608 ^ 1'b0 ;
  assign n46406 = n13393 | n44458 ;
  assign n46407 = n21832 | n43170 ;
  assign n46408 = n46407 ^ n42196 ^ 1'b0 ;
  assign n46409 = n8006 ^ n3651 ^ n3575 ;
  assign n46410 = ( n3629 & n17841 ) | ( n3629 & ~n21829 ) | ( n17841 & ~n21829 ) ;
  assign n46411 = n25349 & ~n35314 ;
  assign n46412 = n10201 & ~n15750 ;
  assign n46413 = n46411 & n46412 ;
  assign n46414 = n10506 & ~n15991 ;
  assign n46415 = ~n15987 & n46414 ;
  assign n46416 = n46415 ^ n41209 ^ n1030 ;
  assign n46417 = n11159 ^ n9897 ^ 1'b0 ;
  assign n46418 = n46416 | n46417 ;
  assign n46419 = n8521 & n44417 ;
  assign n46420 = n24273 & n46419 ;
  assign n46422 = n15800 ^ n7196 ^ 1'b0 ;
  assign n46423 = n479 & n46422 ;
  assign n46424 = ~n5475 & n46423 ;
  assign n46421 = ~n9182 & n32133 ;
  assign n46425 = n46424 ^ n46421 ^ 1'b0 ;
  assign n46426 = n19250 ^ n18139 ^ 1'b0 ;
  assign n46427 = n43252 ^ n27841 ^ 1'b0 ;
  assign n46428 = n46427 ^ n22615 ^ n13725 ;
  assign n46429 = n25328 ^ n20465 ^ n18280 ;
  assign n46430 = n42497 ^ n12352 ^ 1'b0 ;
  assign n46431 = ~n4556 & n46430 ;
  assign n46432 = n24638 ^ n1486 ^ n929 ;
  assign n46433 = n34416 ^ n12202 ^ 1'b0 ;
  assign n46434 = n46432 & n46433 ;
  assign n46435 = n1034 | n11486 ;
  assign n46436 = ( n6879 & n16581 ) | ( n6879 & n22365 ) | ( n16581 & n22365 ) ;
  assign n46437 = ~n11988 & n46436 ;
  assign n46438 = n46437 ^ x114 ^ 1'b0 ;
  assign n46439 = n19065 & ~n46438 ;
  assign n46440 = ( n1842 & ~n8927 ) | ( n1842 & n20096 ) | ( ~n8927 & n20096 ) ;
  assign n46441 = n22801 | n46440 ;
  assign n46442 = n5370 | n29335 ;
  assign n46443 = n43200 ^ n6642 ^ 1'b0 ;
  assign n46444 = n46442 | n46443 ;
  assign n46445 = n10998 ^ n3705 ^ 1'b0 ;
  assign n46446 = n8945 | n46445 ;
  assign n46447 = ( n2534 & n5667 ) | ( n2534 & n12227 ) | ( n5667 & n12227 ) ;
  assign n46448 = n46446 | n46447 ;
  assign n46449 = n29914 & ~n46448 ;
  assign n46450 = ~n24424 & n46449 ;
  assign n46451 = ( n13086 & n15126 ) | ( n13086 & n39102 ) | ( n15126 & n39102 ) ;
  assign n46452 = ( n16878 & n46450 ) | ( n16878 & n46451 ) | ( n46450 & n46451 ) ;
  assign n46453 = n46452 ^ n13614 ^ n12736 ;
  assign n46454 = ~n7132 & n13775 ;
  assign n46455 = n12543 | n46454 ;
  assign n46456 = ~n15841 & n20789 ;
  assign n46457 = ( n390 & ~n30421 ) | ( n390 & n46456 ) | ( ~n30421 & n46456 ) ;
  assign n46458 = ~n5049 & n46457 ;
  assign n46459 = n33094 & n46458 ;
  assign n46460 = n41640 ^ n28646 ^ 1'b0 ;
  assign n46461 = n17359 | n17765 ;
  assign n46462 = n571 | n46461 ;
  assign n46463 = n22960 & n46462 ;
  assign n46464 = n46460 & n46463 ;
  assign n46465 = n1350 ^ n292 ^ 1'b0 ;
  assign n46466 = n26443 ^ n18321 ^ 1'b0 ;
  assign n46467 = n22043 & ~n46466 ;
  assign n46468 = ~n9578 & n33177 ;
  assign n46469 = n332 & n24787 ;
  assign n46470 = n33424 & ~n43663 ;
  assign n46472 = n8816 & n16254 ;
  assign n46471 = n12030 | n32729 ;
  assign n46473 = n46472 ^ n46471 ^ n23359 ;
  assign n46474 = n15686 ^ n7090 ^ 1'b0 ;
  assign n46475 = n1250 & ~n46474 ;
  assign n46476 = n24008 ^ n19513 ^ 1'b0 ;
  assign n46477 = n46475 & ~n46476 ;
  assign n46478 = n923 | n36062 ;
  assign n46479 = n1441 & ~n46478 ;
  assign n46480 = ~n12703 & n25796 ;
  assign n46481 = n46480 ^ n4004 ^ 1'b0 ;
  assign n46482 = n15443 & ~n43587 ;
  assign n46483 = n35113 ^ n24039 ^ 1'b0 ;
  assign n46484 = n29963 ^ n13675 ^ 1'b0 ;
  assign n46485 = n14091 & n21030 ;
  assign n46486 = ~n10735 & n39938 ;
  assign n46487 = n46485 & n46486 ;
  assign n46488 = n46487 ^ n31083 ^ 1'b0 ;
  assign n46489 = n29603 ^ n20605 ^ n8266 ;
  assign n46490 = n42430 & n46489 ;
  assign n46491 = n6094 & n13019 ;
  assign n46492 = ~n37466 & n46491 ;
  assign n46493 = ~n6602 & n17821 ;
  assign n46494 = n46493 ^ n40183 ^ 1'b0 ;
  assign n46495 = n32792 ^ n15436 ^ n7115 ;
  assign n46496 = ( ~n2264 & n23069 ) | ( ~n2264 & n46495 ) | ( n23069 & n46495 ) ;
  assign n46497 = ( ~n11781 & n36194 ) | ( ~n11781 & n41533 ) | ( n36194 & n41533 ) ;
  assign n46498 = n6247 ^ n4585 ^ 1'b0 ;
  assign n46500 = n1444 & n15044 ;
  assign n46501 = ~n10708 & n46500 ;
  assign n46499 = n16067 & n23427 ;
  assign n46502 = n46501 ^ n46499 ^ n20461 ;
  assign n46503 = n23045 ^ n6983 ^ 1'b0 ;
  assign n46504 = n8375 & n46503 ;
  assign n46505 = ( x114 & ~n3267 ) | ( x114 & n16728 ) | ( ~n3267 & n16728 ) ;
  assign n46506 = n46505 ^ n12344 ^ 1'b0 ;
  assign n46507 = n15822 & ~n27585 ;
  assign n46508 = ~n763 & n46507 ;
  assign n46509 = ( n6407 & n24254 ) | ( n6407 & n31420 ) | ( n24254 & n31420 ) ;
  assign n46510 = ~n21593 & n39983 ;
  assign n46511 = n30516 & n35541 ;
  assign n46512 = n46511 ^ n9165 ^ 1'b0 ;
  assign n46513 = n33055 ^ n31780 ^ n3259 ;
  assign n46514 = n44548 | n46513 ;
  assign n46515 = n9106 ^ n5988 ^ n1916 ;
  assign n46516 = n8878 & ~n46515 ;
  assign n46517 = n25805 ^ n10116 ^ n6310 ;
  assign n46518 = n46517 ^ n5062 ^ 1'b0 ;
  assign n46519 = n39621 & n46518 ;
  assign n46520 = n4978 | n23448 ;
  assign n46521 = ( n5731 & ~n17525 ) | ( n5731 & n39352 ) | ( ~n17525 & n39352 ) ;
  assign n46522 = n29314 ^ n18492 ^ 1'b0 ;
  assign n46523 = n46522 ^ n42138 ^ n17823 ;
  assign n46524 = n17923 ^ n6839 ^ n1814 ;
  assign n46525 = n3229 & ~n7631 ;
  assign n46527 = ( n9682 & n10830 ) | ( n9682 & n37586 ) | ( n10830 & n37586 ) ;
  assign n46526 = n9390 & ~n35286 ;
  assign n46528 = n46527 ^ n46526 ^ 1'b0 ;
  assign n46529 = n39628 ^ n28842 ^ 1'b0 ;
  assign n46530 = ~n4431 & n12733 ;
  assign n46531 = n46530 ^ n30092 ^ 1'b0 ;
  assign n46532 = n12522 & ~n46531 ;
  assign n46533 = ( n5800 & n7111 ) | ( n5800 & n13082 ) | ( n7111 & n13082 ) ;
  assign n46534 = ( ~n4700 & n6209 ) | ( ~n4700 & n11135 ) | ( n6209 & n11135 ) ;
  assign n46535 = n8179 | n30455 ;
  assign n46539 = n10846 ^ n627 ^ 1'b0 ;
  assign n46540 = ~n25184 & n46539 ;
  assign n46536 = n25125 ^ n21676 ^ 1'b0 ;
  assign n46537 = ~n21213 & n46536 ;
  assign n46538 = n31615 & n46537 ;
  assign n46541 = n46540 ^ n46538 ^ 1'b0 ;
  assign n46542 = n18240 ^ n10767 ^ n3691 ;
  assign n46543 = n46542 ^ n2354 ^ 1'b0 ;
  assign n46544 = ~n46541 & n46543 ;
  assign n46545 = n35196 & n41409 ;
  assign n46546 = ~n31173 & n34747 ;
  assign n46547 = n22609 & ~n29217 ;
  assign n46548 = ~n10003 & n46547 ;
  assign n46549 = n15091 ^ n5389 ^ 1'b0 ;
  assign n46550 = ( n1755 & n17275 ) | ( n1755 & ~n18841 ) | ( n17275 & ~n18841 ) ;
  assign n46551 = ~n2868 & n44714 ;
  assign n46552 = n17596 ^ n11579 ^ 1'b0 ;
  assign n46553 = n8024 | n46552 ;
  assign n46554 = n4755 & ~n46553 ;
  assign n46555 = ~n14019 & n23176 ;
  assign n46556 = n46555 ^ n33296 ^ 1'b0 ;
  assign n46557 = n5073 & ~n21851 ;
  assign n46558 = n42544 ^ n15407 ^ 1'b0 ;
  assign n46559 = n46557 & n46558 ;
  assign n46563 = n1206 & n13196 ;
  assign n46560 = n43693 ^ n39337 ^ n15483 ;
  assign n46561 = n18934 ^ n530 ^ 1'b0 ;
  assign n46562 = n46560 | n46561 ;
  assign n46564 = n46563 ^ n46562 ^ n18972 ;
  assign n46565 = n46564 ^ n841 ^ 1'b0 ;
  assign n46566 = n46559 & n46565 ;
  assign n46567 = n26733 & n37929 ;
  assign n46568 = ~n1524 & n46567 ;
  assign n46569 = n46568 ^ n3551 ^ 1'b0 ;
  assign n46570 = ~n14627 & n19511 ;
  assign n46571 = ~n36463 & n46570 ;
  assign n46572 = n13711 | n27006 ;
  assign n46573 = n46572 ^ n1336 ^ 1'b0 ;
  assign n46574 = n8490 | n29983 ;
  assign n46575 = n31450 ^ n9257 ^ n362 ;
  assign n46576 = n13911 | n21598 ;
  assign n46577 = n46576 ^ n20726 ^ 1'b0 ;
  assign n46578 = n717 & n46577 ;
  assign n46579 = n10683 & n13153 ;
  assign n46580 = n46579 ^ n14224 ^ 1'b0 ;
  assign n46581 = n46580 ^ n12246 ^ 1'b0 ;
  assign n46582 = ~n8743 & n46581 ;
  assign n46583 = n46582 ^ n21822 ^ n15485 ;
  assign n46584 = ~n4480 & n19281 ;
  assign n46585 = n13098 & ~n24982 ;
  assign n46586 = ~x103 & n46585 ;
  assign n46587 = n39351 | n46586 ;
  assign n46588 = n46587 ^ n14881 ^ 1'b0 ;
  assign n46589 = n42851 ^ n11653 ^ 1'b0 ;
  assign n46590 = n42669 ^ n28148 ^ n14871 ;
  assign n46591 = n17379 ^ n1150 ^ 1'b0 ;
  assign n46592 = n44089 ^ n9203 ^ 1'b0 ;
  assign n46593 = ~n35499 & n37513 ;
  assign n46594 = n30154 ^ n4597 ^ n2582 ;
  assign n46595 = ( n10491 & n44182 ) | ( n10491 & ~n46594 ) | ( n44182 & ~n46594 ) ;
  assign n46596 = n8799 & n21827 ;
  assign n46597 = n46596 ^ n8435 ^ 1'b0 ;
  assign n46598 = n19692 | n46597 ;
  assign n46599 = n46598 ^ n1636 ^ 1'b0 ;
  assign n46600 = ( n11398 & n27085 ) | ( n11398 & n31802 ) | ( n27085 & n31802 ) ;
  assign n46601 = ( n19619 & n46599 ) | ( n19619 & ~n46600 ) | ( n46599 & ~n46600 ) ;
  assign n46602 = n46601 ^ n34665 ^ 1'b0 ;
  assign n46603 = n4207 ^ n2543 ^ 1'b0 ;
  assign n46604 = n23263 & ~n46603 ;
  assign n46605 = n15808 & n46604 ;
  assign n46606 = n14833 & ~n27439 ;
  assign n46607 = n18896 & n46606 ;
  assign n46608 = n20104 & ~n23361 ;
  assign n46609 = n46608 ^ n13067 ^ 1'b0 ;
  assign n46610 = ( n3928 & n14366 ) | ( n3928 & ~n46609 ) | ( n14366 & ~n46609 ) ;
  assign n46611 = n46610 ^ n31430 ^ n1463 ;
  assign n46612 = n10739 | n11612 ;
  assign n46613 = n46611 | n46612 ;
  assign n46614 = ~n518 & n15224 ;
  assign n46615 = n46614 ^ n6123 ^ 1'b0 ;
  assign n46616 = n22048 | n46615 ;
  assign n46617 = n1977 & ~n46616 ;
  assign n46618 = ~n16726 & n46617 ;
  assign n46619 = ~n1422 & n46618 ;
  assign n46620 = n41746 ^ n39077 ^ n3398 ;
  assign n46621 = n31995 ^ n26097 ^ n5181 ;
  assign n46624 = n10325 ^ n4761 ^ 1'b0 ;
  assign n46622 = n9152 & ~n16289 ;
  assign n46623 = n46622 ^ n33163 ^ 1'b0 ;
  assign n46625 = n46624 ^ n46623 ^ n6638 ;
  assign n46626 = n9176 & ~n16600 ;
  assign n46627 = n46626 ^ n45382 ^ n4946 ;
  assign n46628 = n5782 & ~n38766 ;
  assign n46629 = n46628 ^ n12570 ^ 1'b0 ;
  assign n46630 = ~n36002 & n45687 ;
  assign n46631 = n5337 | n46630 ;
  assign n46632 = n46629 & ~n46631 ;
  assign n46633 = n39986 ^ n38411 ^ n14279 ;
  assign n46634 = n21042 & ~n46633 ;
  assign n46635 = n42087 ^ n18866 ^ 1'b0 ;
  assign n46636 = n3310 & ~n12267 ;
  assign n46637 = n9634 & n46636 ;
  assign n46638 = n46637 ^ n37406 ^ 1'b0 ;
  assign n46639 = n5885 & ~n46638 ;
  assign n46640 = ( n3376 & n8942 ) | ( n3376 & n29876 ) | ( n8942 & n29876 ) ;
  assign n46641 = ~n1260 & n46640 ;
  assign n46642 = n46641 ^ n14798 ^ 1'b0 ;
  assign n46643 = n6497 & ~n40750 ;
  assign n46644 = ~n46642 & n46643 ;
  assign n46645 = ~n15976 & n32051 ;
  assign n46646 = n45652 | n46637 ;
  assign n46647 = n29747 | n44243 ;
  assign n46648 = n46647 ^ n31013 ^ 1'b0 ;
  assign n46649 = n30670 ^ n26323 ^ n14578 ;
  assign n46650 = n46648 & n46649 ;
  assign n46651 = n11870 & n46650 ;
  assign n46652 = n2998 & ~n41143 ;
  assign n46653 = n15417 | n46652 ;
  assign n46654 = ~n15836 & n46653 ;
  assign n46655 = ~n27099 & n46654 ;
  assign n46656 = n759 & ~n12473 ;
  assign n46657 = n33493 ^ n20097 ^ n4140 ;
  assign n46658 = n46657 ^ n19059 ^ 1'b0 ;
  assign n46659 = ( ~n6264 & n45302 ) | ( ~n6264 & n46658 ) | ( n45302 & n46658 ) ;
  assign n46660 = n24536 ^ n21856 ^ 1'b0 ;
  assign n46661 = n46659 | n46660 ;
  assign n46662 = ( ~n12259 & n37816 ) | ( ~n12259 & n38444 ) | ( n37816 & n38444 ) ;
  assign n46663 = n22337 | n23951 ;
  assign n46664 = n4439 | n46663 ;
  assign n46665 = ~n29248 & n46664 ;
  assign n46666 = n15121 & ~n22260 ;
  assign n46667 = ~n5637 & n17148 ;
  assign n46668 = ~n12196 & n25237 ;
  assign n46669 = n46668 ^ n36971 ^ 1'b0 ;
  assign n46670 = ~n12807 & n46669 ;
  assign n46671 = n33373 & ~n46670 ;
  assign n46672 = n27320 ^ n15816 ^ n4646 ;
  assign n46673 = n23672 ^ n22521 ^ 1'b0 ;
  assign n46674 = n4153 & ~n46673 ;
  assign n46675 = n33131 ^ n31211 ^ 1'b0 ;
  assign n46676 = n16959 | n33996 ;
  assign n46677 = n46675 | n46676 ;
  assign n46678 = n46677 ^ n29847 ^ 1'b0 ;
  assign n46679 = n4041 & ~n46678 ;
  assign n46680 = n6012 & n6325 ;
  assign n46681 = n15536 & n46680 ;
  assign n46682 = n30891 ^ n6882 ^ 1'b0 ;
  assign n46683 = ~n17507 & n46682 ;
  assign n46684 = ~n3358 & n46683 ;
  assign n46685 = n46681 & n46684 ;
  assign n46686 = ( ~n3552 & n32781 ) | ( ~n3552 & n46457 ) | ( n32781 & n46457 ) ;
  assign n46687 = n43933 ^ n32375 ^ n955 ;
  assign n46688 = n2907 & ~n44733 ;
  assign n46689 = n10660 & n24113 ;
  assign n46690 = n18566 ^ n10960 ^ 1'b0 ;
  assign n46691 = ~n36580 & n46690 ;
  assign n46692 = n13847 | n14064 ;
  assign n46693 = n25608 & ~n46692 ;
  assign n46694 = n6979 & n25908 ;
  assign n46695 = n15819 & n46694 ;
  assign n46696 = ( n8613 & ~n15121 ) | ( n8613 & n23264 ) | ( ~n15121 & n23264 ) ;
  assign n46697 = n41646 ^ n2954 ^ 1'b0 ;
  assign n46698 = n46696 & n46697 ;
  assign n46699 = n27458 ^ n4174 ^ 1'b0 ;
  assign n46700 = n46699 ^ n31136 ^ 1'b0 ;
  assign n46701 = ( n2912 & n13722 ) | ( n2912 & ~n46700 ) | ( n13722 & ~n46700 ) ;
  assign n46702 = n46701 ^ n3282 ^ 1'b0 ;
  assign n46705 = n1197 & n4948 ;
  assign n46706 = n46705 ^ n10269 ^ 1'b0 ;
  assign n46703 = n16656 | n34177 ;
  assign n46704 = n12622 & ~n46703 ;
  assign n46707 = n46706 ^ n46704 ^ 1'b0 ;
  assign n46708 = n11059 | n45686 ;
  assign n46709 = n9803 & n46624 ;
  assign n46710 = n3309 & ~n46709 ;
  assign n46711 = n25531 ^ n7454 ^ 1'b0 ;
  assign n46712 = n4641 | n46711 ;
  assign n46713 = ( n5592 & n27991 ) | ( n5592 & ~n46712 ) | ( n27991 & ~n46712 ) ;
  assign n46714 = n3389 | n11790 ;
  assign n46715 = n23892 | n27705 ;
  assign n46716 = n39003 ^ n11684 ^ 1'b0 ;
  assign n46717 = n5959 & ~n46716 ;
  assign n46718 = n28222 ^ n20634 ^ n12423 ;
  assign n46719 = n27971 ^ n26321 ^ 1'b0 ;
  assign n46721 = n6689 ^ n4994 ^ n4097 ;
  assign n46720 = n32681 ^ n17490 ^ 1'b0 ;
  assign n46722 = n46721 ^ n46720 ^ 1'b0 ;
  assign n46723 = n34207 ^ n23280 ^ n2680 ;
  assign n46724 = ~n5484 & n22361 ;
  assign n46725 = ~n4827 & n5786 ;
  assign n46726 = ~n9838 & n46725 ;
  assign n46727 = n5203 & n5833 ;
  assign n46728 = n46727 ^ n2017 ^ 1'b0 ;
  assign n46729 = n23870 ^ n11979 ^ n5689 ;
  assign n46730 = n23439 & ~n38009 ;
  assign n46731 = n14789 ^ n2476 ^ 1'b0 ;
  assign n46732 = ( n21769 & n25762 ) | ( n21769 & n46731 ) | ( n25762 & n46731 ) ;
  assign n46733 = n26200 | n46732 ;
  assign n46734 = n19278 & ~n24706 ;
  assign n46735 = n46734 ^ n12828 ^ 1'b0 ;
  assign n46736 = n13987 | n17562 ;
  assign n46737 = n32799 | n46736 ;
  assign n46739 = n12987 ^ n9512 ^ 1'b0 ;
  assign n46740 = n5580 & n46739 ;
  assign n46741 = n46740 ^ n7566 ^ 1'b0 ;
  assign n46738 = n7777 | n18059 ;
  assign n46742 = n46741 ^ n46738 ^ 1'b0 ;
  assign n46743 = n7794 & n36514 ;
  assign n46744 = ( ~n5263 & n12858 ) | ( ~n5263 & n19854 ) | ( n12858 & n19854 ) ;
  assign n46745 = n3898 & n46744 ;
  assign n46746 = n41157 ^ n10026 ^ 1'b0 ;
  assign n46747 = ~n22150 & n46746 ;
  assign n46748 = n6012 & ~n46747 ;
  assign n46749 = ~n1536 & n46748 ;
  assign n46750 = n2030 | n12967 ;
  assign n46751 = n27647 ^ n20821 ^ 1'b0 ;
  assign n46752 = n13531 | n46751 ;
  assign n46753 = n46750 | n46752 ;
  assign n46754 = ( ~n6018 & n10127 ) | ( ~n6018 & n29537 ) | ( n10127 & n29537 ) ;
  assign n46755 = n14575 | n23196 ;
  assign n46756 = ~n9408 & n46755 ;
  assign n46757 = n45358 | n46756 ;
  assign n46758 = ( ~n4292 & n18008 ) | ( ~n4292 & n23676 ) | ( n18008 & n23676 ) ;
  assign n46759 = n30327 ^ n23484 ^ n12098 ;
  assign n46760 = n46759 ^ n37701 ^ 1'b0 ;
  assign n46761 = n46758 & ~n46760 ;
  assign n46762 = n22720 ^ n1536 ^ 1'b0 ;
  assign n46765 = n25959 | n35769 ;
  assign n46763 = n15204 & n15291 ;
  assign n46764 = ~n17935 & n46763 ;
  assign n46766 = n46765 ^ n46764 ^ n32950 ;
  assign n46767 = ~n11552 & n16512 ;
  assign n46768 = n46766 & n46767 ;
  assign n46769 = n7237 | n18602 ;
  assign n46770 = n18004 & ~n46769 ;
  assign n46771 = n26432 | n46770 ;
  assign n46772 = ~n23956 & n37903 ;
  assign n46773 = n40894 ^ n3432 ^ 1'b0 ;
  assign n46774 = ~n18604 & n46773 ;
  assign n46775 = n28490 & ~n34053 ;
  assign n46776 = n14228 & n26696 ;
  assign n46777 = ~n46775 & n46776 ;
  assign n46781 = ( n4001 & n13512 ) | ( n4001 & n18746 ) | ( n13512 & n18746 ) ;
  assign n46780 = ~n12682 & n16619 ;
  assign n46778 = n1658 | n4292 ;
  assign n46779 = n46778 ^ n19666 ^ 1'b0 ;
  assign n46782 = n46781 ^ n46780 ^ n46779 ;
  assign n46783 = n46777 & n46782 ;
  assign n46784 = n40953 ^ n25817 ^ n13680 ;
  assign n46785 = ( x142 & n12592 ) | ( x142 & n46784 ) | ( n12592 & n46784 ) ;
  assign n46786 = n46785 ^ n10531 ^ 1'b0 ;
  assign n46787 = n12954 & n46786 ;
  assign n46788 = ~n7956 & n16321 ;
  assign n46789 = n35327 & ~n46788 ;
  assign n46790 = ( n6074 & n46787 ) | ( n6074 & ~n46789 ) | ( n46787 & ~n46789 ) ;
  assign n46791 = ~n6074 & n28851 ;
  assign n46792 = ( n3755 & n13668 ) | ( n3755 & n20412 ) | ( n13668 & n20412 ) ;
  assign n46793 = n13905 & ~n46792 ;
  assign n46794 = ~n18649 & n23782 ;
  assign n46795 = ~n34061 & n45290 ;
  assign n46796 = n23298 & n46795 ;
  assign n46797 = ~n2425 & n44668 ;
  assign n46798 = n46797 ^ n545 ^ 1'b0 ;
  assign n46799 = n23032 ^ n5628 ^ 1'b0 ;
  assign n46800 = ~n41574 & n46799 ;
  assign n46801 = n17957 & ~n46800 ;
  assign n46802 = n29243 ^ n2500 ^ 1'b0 ;
  assign n46803 = n28352 | n46802 ;
  assign n46804 = n46803 ^ n36994 ^ n10129 ;
  assign n46807 = n1447 | n6399 ;
  assign n46808 = n46807 ^ n23952 ^ 1'b0 ;
  assign n46809 = n19995 | n46808 ;
  assign n46805 = ~n18360 & n25307 ;
  assign n46806 = n46805 ^ n28767 ^ n704 ;
  assign n46810 = n46809 ^ n46806 ^ 1'b0 ;
  assign n46811 = n302 & ~n1106 ;
  assign n46812 = ( n9012 & n32594 ) | ( n9012 & n46811 ) | ( n32594 & n46811 ) ;
  assign n46813 = n42897 ^ n490 ^ 1'b0 ;
  assign n46814 = n24769 ^ n9035 ^ 1'b0 ;
  assign n46815 = n44170 ^ n20328 ^ 1'b0 ;
  assign n46816 = n7339 ^ n4784 ^ 1'b0 ;
  assign n46817 = n23840 | n46816 ;
  assign n46818 = n26736 & ~n45922 ;
  assign n46819 = ( n18208 & n29069 ) | ( n18208 & ~n46818 ) | ( n29069 & ~n46818 ) ;
  assign n46820 = n16581 | n30903 ;
  assign n46821 = n10259 ^ n9567 ^ 1'b0 ;
  assign n46822 = n46820 & ~n46821 ;
  assign n46823 = ( ~n9408 & n16411 ) | ( ~n9408 & n46822 ) | ( n16411 & n46822 ) ;
  assign n46824 = n9418 ^ n6054 ^ n5155 ;
  assign n46825 = n26483 & n41999 ;
  assign n46826 = n4961 & ~n18702 ;
  assign n46827 = n46826 ^ n21057 ^ n18617 ;
  assign n46828 = n3770 & n4304 ;
  assign n46830 = n6453 & ~n10255 ;
  assign n46829 = n10740 & ~n16964 ;
  assign n46831 = n46830 ^ n46829 ^ 1'b0 ;
  assign n46832 = n15382 & ~n32741 ;
  assign n46833 = ~n43364 & n46832 ;
  assign n46834 = n46833 ^ n12677 ^ 1'b0 ;
  assign n46835 = ( ~n23812 & n31733 ) | ( ~n23812 & n40154 ) | ( n31733 & n40154 ) ;
  assign n46836 = n34269 ^ n32642 ^ 1'b0 ;
  assign n46837 = n21689 ^ n4875 ^ 1'b0 ;
  assign n46838 = n46837 ^ n45587 ^ n839 ;
  assign n46839 = n5234 & ~n32686 ;
  assign n46840 = n46839 ^ n8477 ^ 1'b0 ;
  assign n46841 = n7037 & n26686 ;
  assign n46842 = n5009 & n34164 ;
  assign n46843 = n46842 ^ n44850 ^ 1'b0 ;
  assign n46844 = n4929 & ~n27362 ;
  assign n46845 = n46844 ^ n45978 ^ 1'b0 ;
  assign n46846 = n37925 ^ n21316 ^ 1'b0 ;
  assign n46847 = n42282 ^ n21477 ^ n6912 ;
  assign n46848 = ( ~n2560 & n7231 ) | ( ~n2560 & n44912 ) | ( n7231 & n44912 ) ;
  assign n46849 = n5834 & n15617 ;
  assign n46850 = n46849 ^ n15966 ^ 1'b0 ;
  assign n46851 = ( n25439 & n26531 ) | ( n25439 & ~n46850 ) | ( n26531 & ~n46850 ) ;
  assign n46852 = n14470 ^ n13214 ^ n7145 ;
  assign n46853 = n46852 ^ n574 ^ 1'b0 ;
  assign n46854 = n12454 | n33666 ;
  assign n46855 = n30722 & ~n46854 ;
  assign n46856 = n29890 ^ n7854 ^ 1'b0 ;
  assign n46857 = ~n46855 & n46856 ;
  assign n46858 = n16325 | n43678 ;
  assign n46859 = n10429 & ~n46858 ;
  assign n46860 = ~n21179 & n46859 ;
  assign n46861 = n14225 | n15927 ;
  assign n46862 = n46861 ^ n10364 ^ 1'b0 ;
  assign n46863 = n11531 ^ n4961 ^ 1'b0 ;
  assign n46864 = ~n16940 & n46863 ;
  assign n46865 = n46864 ^ n38748 ^ n3085 ;
  assign n46867 = n28125 ^ n20634 ^ n17544 ;
  assign n46866 = n6016 & n14689 ;
  assign n46868 = n46867 ^ n46866 ^ n9803 ;
  assign n46869 = n12241 ^ n11308 ^ n5259 ;
  assign n46870 = n33406 ^ n22695 ^ 1'b0 ;
  assign n46871 = n15774 & n17978 ;
  assign n46872 = n46870 & n46871 ;
  assign n46874 = n2092 ^ n266 ^ 1'b0 ;
  assign n46875 = ~n23659 & n46874 ;
  assign n46873 = n19669 | n21203 ;
  assign n46876 = n46875 ^ n46873 ^ 1'b0 ;
  assign n46877 = n21146 ^ n17414 ^ n6393 ;
  assign n46878 = n46877 ^ n13847 ^ 1'b0 ;
  assign n46879 = n2669 | n11625 ;
  assign n46880 = n46879 ^ n14679 ^ 1'b0 ;
  assign n46881 = ( n6193 & ~n7006 ) | ( n6193 & n22297 ) | ( ~n7006 & n22297 ) ;
  assign n46882 = ( n21056 & n26462 ) | ( n21056 & n36470 ) | ( n26462 & n36470 ) ;
  assign n46883 = n32790 ^ n27845 ^ 1'b0 ;
  assign n46884 = n33328 ^ n20796 ^ 1'b0 ;
  assign n46885 = n513 & n45295 ;
  assign n46886 = n16722 | n46885 ;
  assign n46887 = n46886 ^ n2943 ^ 1'b0 ;
  assign n46888 = n14403 | n46887 ;
  assign n46889 = n46888 ^ n21344 ^ 1'b0 ;
  assign n46890 = ( ~n34378 & n35987 ) | ( ~n34378 & n38985 ) | ( n35987 & n38985 ) ;
  assign n46891 = n46890 ^ n18849 ^ 1'b0 ;
  assign n46892 = n24438 & ~n46891 ;
  assign n46893 = ( n4763 & ~n7991 ) | ( n4763 & n20725 ) | ( ~n7991 & n20725 ) ;
  assign n46895 = n41177 ^ n3470 ^ 1'b0 ;
  assign n46894 = ~n15415 & n35875 ;
  assign n46896 = n46895 ^ n46894 ^ n1780 ;
  assign n46897 = ( ~n25380 & n46893 ) | ( ~n25380 & n46896 ) | ( n46893 & n46896 ) ;
  assign n46898 = n23217 ^ n13244 ^ n7569 ;
  assign n46899 = n12036 ^ n8012 ^ n447 ;
  assign n46900 = ( x39 & n20168 ) | ( x39 & ~n46899 ) | ( n20168 & ~n46899 ) ;
  assign n46901 = ~n785 & n15264 ;
  assign n46902 = n10250 & ~n24430 ;
  assign n46903 = ~n32545 & n46902 ;
  assign n46904 = ( ~n1324 & n13734 ) | ( ~n1324 & n46903 ) | ( n13734 & n46903 ) ;
  assign n46905 = n13625 ^ n1879 ^ 1'b0 ;
  assign n46906 = n21951 | n46905 ;
  assign n46907 = n46906 ^ x234 ^ 1'b0 ;
  assign n46908 = n46904 | n46907 ;
  assign n46909 = n46287 ^ n37967 ^ 1'b0 ;
  assign n46910 = n17579 | n46909 ;
  assign n46911 = ~n21214 & n30318 ;
  assign n46912 = n18610 ^ n15540 ^ 1'b0 ;
  assign n46913 = n1025 | n1387 ;
  assign n46914 = n5054 | n42886 ;
  assign n46915 = n46913 | n46914 ;
  assign n46916 = n22459 & ~n46915 ;
  assign n46917 = ( x204 & n7390 ) | ( x204 & ~n8085 ) | ( n7390 & ~n8085 ) ;
  assign n46918 = n1239 & ~n20794 ;
  assign n46919 = n46918 ^ n31789 ^ 1'b0 ;
  assign n46920 = n46917 & ~n46919 ;
  assign n46921 = ( ~x229 & n21363 ) | ( ~x229 & n28511 ) | ( n21363 & n28511 ) ;
  assign n46922 = n15132 & n46921 ;
  assign n46926 = n24143 | n33433 ;
  assign n46927 = n32304 & ~n46926 ;
  assign n46923 = ( ~n1541 & n6831 ) | ( ~n1541 & n23807 ) | ( n6831 & n23807 ) ;
  assign n46924 = n30865 ^ n2013 ^ 1'b0 ;
  assign n46925 = ( n25377 & n46923 ) | ( n25377 & n46924 ) | ( n46923 & n46924 ) ;
  assign n46928 = n46927 ^ n46925 ^ n8172 ;
  assign n46929 = ( n36031 & ~n46922 ) | ( n36031 & n46928 ) | ( ~n46922 & n46928 ) ;
  assign n46930 = n35661 ^ n16890 ^ 1'b0 ;
  assign n46931 = n15057 & n46930 ;
  assign n46932 = n46931 ^ n43796 ^ n16371 ;
  assign n46933 = n28222 ^ n9757 ^ n4776 ;
  assign n46934 = ~n3369 & n40074 ;
  assign n46935 = ~n46933 & n46934 ;
  assign n46936 = n46935 ^ n39979 ^ 1'b0 ;
  assign n46937 = n6952 | n41465 ;
  assign n46938 = n11895 & ~n18864 ;
  assign n46939 = n41558 & ~n46938 ;
  assign n46940 = n34050 ^ n27361 ^ 1'b0 ;
  assign n46941 = n654 & n46940 ;
  assign n46942 = ( n763 & n11076 ) | ( n763 & ~n32959 ) | ( n11076 & ~n32959 ) ;
  assign n46943 = n22346 ^ n6270 ^ 1'b0 ;
  assign n46944 = n46943 ^ n26948 ^ n2678 ;
  assign n46945 = n7878 & ~n10848 ;
  assign n46946 = ( ~n13982 & n40436 ) | ( ~n13982 & n46945 ) | ( n40436 & n46945 ) ;
  assign n46947 = n15574 ^ n6673 ^ n947 ;
  assign n46948 = n46947 ^ n30716 ^ 1'b0 ;
  assign n46949 = ~n23260 & n43199 ;
  assign n46950 = n46949 ^ n22174 ^ n17870 ;
  assign n46951 = n18259 ^ n1816 ^ 1'b0 ;
  assign n46952 = n46951 ^ n23853 ^ n6156 ;
  assign n46953 = n39032 ^ n31909 ^ n10837 ;
  assign n46954 = x174 & n46953 ;
  assign n46955 = n38984 ^ n9606 ^ 1'b0 ;
  assign n46956 = n6020 | n46955 ;
  assign n46957 = n44365 & ~n46956 ;
  assign n46958 = n28786 & ~n46957 ;
  assign n46959 = n20518 & ~n30868 ;
  assign n46960 = ( n8238 & ~n19485 ) | ( n8238 & n46959 ) | ( ~n19485 & n46959 ) ;
  assign n46961 = ( n28224 & n40491 ) | ( n28224 & n46960 ) | ( n40491 & n46960 ) ;
  assign n46962 = n34854 ^ n11299 ^ 1'b0 ;
  assign n46963 = n2920 & ~n22788 ;
  assign n46964 = n46963 ^ n32872 ^ 1'b0 ;
  assign n46965 = n46964 ^ n28582 ^ n3905 ;
  assign n46966 = n8591 ^ n2282 ^ 1'b0 ;
  assign n46967 = n8718 & ~n46966 ;
  assign n46968 = n46965 & ~n46967 ;
  assign n46969 = n1145 | n36853 ;
  assign n46970 = n16334 ^ n10228 ^ 1'b0 ;
  assign n46971 = ~n38763 & n46970 ;
  assign n46973 = n40154 ^ n23771 ^ 1'b0 ;
  assign n46974 = n10426 & ~n46973 ;
  assign n46972 = n23052 | n28319 ;
  assign n46975 = n46974 ^ n46972 ^ 1'b0 ;
  assign n46976 = n46287 ^ n18963 ^ n8169 ;
  assign n46977 = ~n8754 & n46976 ;
  assign n46978 = n46977 ^ n15335 ^ 1'b0 ;
  assign n46979 = n582 & n46978 ;
  assign n46980 = ~n46975 & n46979 ;
  assign n46981 = n41173 ^ n18696 ^ 1'b0 ;
  assign n46982 = n13227 & ~n46981 ;
  assign n46983 = n27186 | n37830 ;
  assign n46984 = n46983 ^ n37589 ^ 1'b0 ;
  assign n46985 = n6218 | n46984 ;
  assign n46986 = n25003 & ~n46985 ;
  assign n46987 = n4521 & n6568 ;
  assign n46988 = ~x146 & n46987 ;
  assign n46989 = ( n2058 & n39248 ) | ( n2058 & ~n46988 ) | ( n39248 & ~n46988 ) ;
  assign n46990 = n16850 ^ n9853 ^ n4355 ;
  assign n46991 = ( ~n21188 & n36598 ) | ( ~n21188 & n46990 ) | ( n36598 & n46990 ) ;
  assign n46992 = ~n7750 & n46991 ;
  assign n46993 = n7739 & n26557 ;
  assign n46994 = n46993 ^ n12015 ^ 1'b0 ;
  assign n46995 = ( n20731 & n22425 ) | ( n20731 & n46994 ) | ( n22425 & n46994 ) ;
  assign n46996 = n25904 ^ n12147 ^ n7573 ;
  assign n46997 = ( n2174 & ~n41524 ) | ( n2174 & n46996 ) | ( ~n41524 & n46996 ) ;
  assign n46998 = n1105 | n9028 ;
  assign n46999 = n46998 ^ n8870 ^ 1'b0 ;
  assign n47000 = n46999 ^ n15638 ^ 1'b0 ;
  assign n47001 = n35669 ^ n14519 ^ 1'b0 ;
  assign n47002 = n32386 | n47001 ;
  assign n47003 = n29914 ^ n1532 ^ 1'b0 ;
  assign n47004 = n6272 & ~n47003 ;
  assign n47005 = n12930 ^ n6663 ^ x8 ;
  assign n47006 = n19046 ^ n10333 ^ n2247 ;
  assign n47007 = n16337 & n40396 ;
  assign n47008 = n22724 & n47007 ;
  assign n47009 = n47008 ^ n29231 ^ n8927 ;
  assign n47010 = n42647 ^ n9957 ^ n4945 ;
  assign n47011 = ~n913 & n47010 ;
  assign n47012 = n39667 & n47011 ;
  assign n47013 = n1116 & ~n18905 ;
  assign n47014 = ~n7302 & n47013 ;
  assign n47015 = n40740 | n47014 ;
  assign n47016 = n39363 ^ n13177 ^ 1'b0 ;
  assign n47017 = n13171 & n47016 ;
  assign n47018 = n23674 ^ n22574 ^ n16172 ;
  assign n47019 = ( n6047 & n47017 ) | ( n6047 & n47018 ) | ( n47017 & n47018 ) ;
  assign n47020 = n30830 ^ n29398 ^ n9061 ;
  assign n47022 = n15967 ^ n12066 ^ 1'b0 ;
  assign n47021 = n2566 & n19775 ;
  assign n47023 = n47022 ^ n47021 ^ n41120 ;
  assign n47024 = n30055 ^ n1858 ^ 1'b0 ;
  assign n47025 = ~n2107 & n27164 ;
  assign n47026 = ~n35147 & n47025 ;
  assign n47027 = n29556 ^ n9887 ^ 1'b0 ;
  assign n47028 = ~n13148 & n47027 ;
  assign n47029 = n26585 | n45207 ;
  assign n47030 = n47029 ^ n20107 ^ 1'b0 ;
  assign n47031 = n33996 ^ n24076 ^ 1'b0 ;
  assign n47033 = n5389 ^ n2562 ^ 1'b0 ;
  assign n47034 = n6551 & ~n47033 ;
  assign n47035 = n47034 ^ n24446 ^ n15645 ;
  assign n47032 = n10873 ^ n4371 ^ 1'b0 ;
  assign n47036 = n47035 ^ n47032 ^ n12060 ;
  assign n47037 = n25287 ^ n16366 ^ 1'b0 ;
  assign n47038 = n11501 ^ n10195 ^ n4243 ;
  assign n47039 = n36737 ^ n994 ^ 1'b0 ;
  assign n47040 = ~n369 & n47039 ;
  assign n47041 = n47040 ^ n37522 ^ n7416 ;
  assign n47042 = x229 & ~n20341 ;
  assign n47044 = n10970 | n18504 ;
  assign n47043 = n11418 & n41763 ;
  assign n47045 = n47044 ^ n47043 ^ n10171 ;
  assign n47046 = n31433 ^ n16982 ^ 1'b0 ;
  assign n47047 = n3545 & ~n9779 ;
  assign n47048 = n6028 & n47047 ;
  assign n47050 = n981 | n32570 ;
  assign n47049 = n4426 & ~n16703 ;
  assign n47051 = n47050 ^ n47049 ^ 1'b0 ;
  assign n47052 = n30597 | n42028 ;
  assign n47053 = n47052 ^ n7208 ^ 1'b0 ;
  assign n47054 = ~n4827 & n27887 ;
  assign n47055 = n47054 ^ n30615 ^ 1'b0 ;
  assign n47056 = ~n14079 & n47055 ;
  assign n47057 = n10517 & ~n11197 ;
  assign n47058 = n47057 ^ n9118 ^ 1'b0 ;
  assign n47059 = n47058 ^ n45117 ^ n16417 ;
  assign n47060 = n5007 & ~n11112 ;
  assign n47061 = ( n7689 & n17789 ) | ( n7689 & n35429 ) | ( n17789 & n35429 ) ;
  assign n47062 = ( n676 & n19700 ) | ( n676 & ~n47061 ) | ( n19700 & ~n47061 ) ;
  assign n47063 = ( ~n40839 & n47060 ) | ( ~n40839 & n47062 ) | ( n47060 & n47062 ) ;
  assign n47064 = n32832 ^ n4341 ^ 1'b0 ;
  assign n47065 = ~n8114 & n10886 ;
  assign n47066 = n47065 ^ n12157 ^ 1'b0 ;
  assign n47067 = n1185 & n29271 ;
  assign n47068 = n13916 ^ n1360 ^ 1'b0 ;
  assign n47069 = n1569 & n34332 ;
  assign n47070 = n47069 ^ n37764 ^ 1'b0 ;
  assign n47071 = n36087 ^ n35341 ^ n2639 ;
  assign n47072 = n37027 ^ n8576 ^ 1'b0 ;
  assign n47074 = n9170 & ~n20062 ;
  assign n47075 = ~n9069 & n47074 ;
  assign n47073 = n9765 ^ n8800 ^ 1'b0 ;
  assign n47076 = n47075 ^ n47073 ^ n2993 ;
  assign n47077 = ( n2772 & n34519 ) | ( n2772 & n39471 ) | ( n34519 & n39471 ) ;
  assign n47078 = ( n13403 & n20669 ) | ( n13403 & ~n25319 ) | ( n20669 & ~n25319 ) ;
  assign n47079 = n11277 | n15913 ;
  assign n47080 = n47078 & ~n47079 ;
  assign n47081 = n3891 & ~n15939 ;
  assign n47082 = n47080 & n47081 ;
  assign n47083 = n47082 ^ n4446 ^ 1'b0 ;
  assign n47084 = n9295 | n47083 ;
  assign n47085 = n30128 ^ n6605 ^ 1'b0 ;
  assign n47086 = n28292 & ~n47085 ;
  assign n47087 = n37712 ^ n6474 ^ 1'b0 ;
  assign n47088 = n4097 & ~n47087 ;
  assign n47089 = n46947 ^ n39108 ^ 1'b0 ;
  assign n47090 = n47088 & ~n47089 ;
  assign n47091 = n3624 & n3691 ;
  assign n47092 = ~n25783 & n47091 ;
  assign n47093 = n24927 | n47092 ;
  assign n47094 = n13452 & ~n47093 ;
  assign n47095 = n33078 & ~n47094 ;
  assign n47096 = n18275 ^ n4958 ^ 1'b0 ;
  assign n47097 = n38552 ^ n33806 ^ 1'b0 ;
  assign n47098 = n35772 ^ n33843 ^ n2489 ;
  assign n47099 = n25864 & ~n43204 ;
  assign n47100 = n17795 & ~n23113 ;
  assign n47101 = n47100 ^ n14022 ^ 1'b0 ;
  assign n47102 = n6267 & n17957 ;
  assign n47103 = n11534 & n47102 ;
  assign n47104 = n10636 & ~n47103 ;
  assign n47105 = n28554 ^ n7058 ^ 1'b0 ;
  assign n47106 = n9390 & ~n47105 ;
  assign n47108 = ( ~n14446 & n17530 ) | ( ~n14446 & n35459 ) | ( n17530 & n35459 ) ;
  assign n47107 = n38699 & ~n45200 ;
  assign n47109 = n47108 ^ n47107 ^ 1'b0 ;
  assign n47110 = n26142 & ~n37284 ;
  assign n47111 = ( n12529 & n22897 ) | ( n12529 & n35260 ) | ( n22897 & n35260 ) ;
  assign n47112 = n13150 & ~n28304 ;
  assign n47113 = n19540 & n20334 ;
  assign n47114 = n47113 ^ n953 ^ 1'b0 ;
  assign n47115 = n18087 | n47114 ;
  assign n47116 = n20263 | n23142 ;
  assign n47117 = n47115 & ~n47116 ;
  assign n47118 = n35909 ^ n12222 ^ 1'b0 ;
  assign n47119 = n25170 ^ n7134 ^ 1'b0 ;
  assign n47120 = n9173 | n47119 ;
  assign n47121 = n7141 | n8218 ;
  assign n47122 = n47121 ^ n26915 ^ n11913 ;
  assign n47123 = n4503 & n9820 ;
  assign n47124 = ( n7331 & ~n16627 ) | ( n7331 & n47123 ) | ( ~n16627 & n47123 ) ;
  assign n47125 = ( n17130 & n47122 ) | ( n17130 & n47124 ) | ( n47122 & n47124 ) ;
  assign n47126 = n20556 ^ n8049 ^ 1'b0 ;
  assign n47127 = ( ~n4471 & n30778 ) | ( ~n4471 & n47126 ) | ( n30778 & n47126 ) ;
  assign n47128 = n6652 | n13951 ;
  assign n47129 = n7983 & ~n13475 ;
  assign n47130 = n24723 & ~n28787 ;
  assign n47131 = ~n12102 & n47130 ;
  assign n47132 = n3331 & ~n4290 ;
  assign n47133 = n8104 & n47132 ;
  assign n47134 = n19656 ^ n1494 ^ 1'b0 ;
  assign n47135 = n1971 | n47134 ;
  assign n47136 = n8409 ^ n4547 ^ 1'b0 ;
  assign n47137 = n20405 ^ n19018 ^ 1'b0 ;
  assign n47138 = ~n901 & n13693 ;
  assign n47139 = ~n26134 & n47138 ;
  assign n47140 = n31359 & ~n47139 ;
  assign n47141 = n29925 ^ n22873 ^ n2567 ;
  assign n47142 = n38456 ^ n26402 ^ 1'b0 ;
  assign n47143 = ~n5706 & n11364 ;
  assign n47144 = n23213 | n43511 ;
  assign n47145 = n1713 & ~n40173 ;
  assign n47146 = n26279 & n47145 ;
  assign n47147 = ~n4303 & n47146 ;
  assign n47148 = n33702 | n47147 ;
  assign n47149 = n38559 & ~n47148 ;
  assign n47150 = n35823 ^ n20055 ^ n13944 ;
  assign n47151 = n46260 & n47150 ;
  assign n47152 = n16430 | n47151 ;
  assign n47153 = n30830 | n47152 ;
  assign n47154 = n22269 ^ n1734 ^ 1'b0 ;
  assign n47155 = ~n763 & n47154 ;
  assign n47156 = ~n3707 & n47155 ;
  assign n47157 = ( ~n4623 & n40482 ) | ( ~n4623 & n44455 ) | ( n40482 & n44455 ) ;
  assign n47159 = n16696 & n17236 ;
  assign n47158 = n13690 & n28390 ;
  assign n47160 = n47159 ^ n47158 ^ 1'b0 ;
  assign n47161 = n47160 ^ n34037 ^ 1'b0 ;
  assign n47162 = n44454 ^ n4695 ^ 1'b0 ;
  assign n47163 = n4968 ^ n1836 ^ 1'b0 ;
  assign n47164 = n37410 ^ n17006 ^ 1'b0 ;
  assign n47165 = n22257 & n47164 ;
  assign n47166 = n35690 ^ n18589 ^ 1'b0 ;
  assign n47167 = n47165 & ~n47166 ;
  assign n47168 = n27240 ^ n11398 ^ 1'b0 ;
  assign n47169 = n6414 & ~n12418 ;
  assign n47170 = n47169 ^ n28614 ^ 1'b0 ;
  assign n47171 = n8343 & ~n11749 ;
  assign n47172 = n47170 & n47171 ;
  assign n47173 = n18151 | n47172 ;
  assign n47174 = n8580 | n47173 ;
  assign n47175 = n16357 ^ n15005 ^ n2202 ;
  assign n47176 = n32584 ^ n21371 ^ 1'b0 ;
  assign n47177 = ~n17841 & n33993 ;
  assign n47178 = n42701 ^ n29758 ^ 1'b0 ;
  assign n47179 = ~n32166 & n47178 ;
  assign n47180 = n47179 ^ n13648 ^ 1'b0 ;
  assign n47181 = ( ~n23881 & n43926 ) | ( ~n23881 & n47180 ) | ( n43926 & n47180 ) ;
  assign n47182 = ~n6719 & n13141 ;
  assign n47183 = n29242 & ~n47182 ;
  assign n47184 = n11289 & n47183 ;
  assign n47185 = n27794 ^ n6674 ^ 1'b0 ;
  assign n47186 = ~n25270 & n47185 ;
  assign n47187 = n20408 ^ n10258 ^ 1'b0 ;
  assign n47188 = n16233 & ~n28305 ;
  assign n47189 = ~n47187 & n47188 ;
  assign n47190 = n15000 & ~n45675 ;
  assign n47191 = n47190 ^ n2077 ^ 1'b0 ;
  assign n47192 = n42284 ^ n14770 ^ 1'b0 ;
  assign n47193 = n47191 & n47192 ;
  assign n47194 = ~n292 & n47193 ;
  assign n47197 = n9534 ^ n1778 ^ 1'b0 ;
  assign n47195 = n22035 ^ n4848 ^ n720 ;
  assign n47196 = n47195 ^ n10065 ^ 1'b0 ;
  assign n47198 = n47197 ^ n47196 ^ n38276 ;
  assign n47199 = ( ~n22689 & n32508 ) | ( ~n22689 & n47198 ) | ( n32508 & n47198 ) ;
  assign n47200 = ( n5106 & ~n24522 ) | ( n5106 & n32292 ) | ( ~n24522 & n32292 ) ;
  assign n47201 = ~n20739 & n32529 ;
  assign n47202 = ~n12604 & n47201 ;
  assign n47203 = n26809 & n47202 ;
  assign n47204 = n43299 ^ n20716 ^ n9263 ;
  assign n47205 = n3742 | n13556 ;
  assign n47206 = n47205 ^ n4193 ^ 1'b0 ;
  assign n47207 = n11025 ^ x141 ^ 1'b0 ;
  assign n47208 = n7696 & n47207 ;
  assign n47209 = ~n12113 & n47208 ;
  assign n47210 = n1132 & ~n10346 ;
  assign n47211 = n47210 ^ n12520 ^ 1'b0 ;
  assign n47212 = n33461 & ~n42720 ;
  assign n47213 = ~n47211 & n47212 ;
  assign n47214 = n16882 & ~n47213 ;
  assign n47215 = ~n41124 & n47214 ;
  assign n47216 = n13111 & ~n13944 ;
  assign n47217 = n43437 ^ n33099 ^ 1'b0 ;
  assign n47218 = n7701 & ~n47217 ;
  assign n47219 = n47216 & ~n47218 ;
  assign n47220 = n30003 ^ n25270 ^ n10720 ;
  assign n47221 = n45943 ^ n43728 ^ 1'b0 ;
  assign n47222 = n22432 ^ n7975 ^ n4842 ;
  assign n47223 = n10525 | n44913 ;
  assign n47224 = n39853 & ~n47223 ;
  assign n47225 = ~n2677 & n7475 ;
  assign n47226 = ~n23335 & n47225 ;
  assign n47227 = n6858 | n14997 ;
  assign n47228 = n1906 & ~n47227 ;
  assign n47229 = ( n2296 & ~n16004 ) | ( n2296 & n40239 ) | ( ~n16004 & n40239 ) ;
  assign n47230 = n7757 & ~n47229 ;
  assign n47231 = n42553 ^ n8829 ^ 1'b0 ;
  assign n47232 = ( n7512 & n16671 ) | ( n7512 & n42339 ) | ( n16671 & n42339 ) ;
  assign n47233 = ( ~n10953 & n16640 ) | ( ~n10953 & n47232 ) | ( n16640 & n47232 ) ;
  assign n47234 = n8116 ^ n4904 ^ 1'b0 ;
  assign n47235 = ( n13704 & n29468 ) | ( n13704 & ~n47234 ) | ( n29468 & ~n47234 ) ;
  assign n47236 = n47235 ^ n43979 ^ n14978 ;
  assign n47237 = n8858 ^ n7810 ^ 1'b0 ;
  assign n47238 = n6832 & ~n47237 ;
  assign n47239 = n4150 & n22288 ;
  assign n47240 = ~n36070 & n47239 ;
  assign n47241 = ( n16386 & n47238 ) | ( n16386 & n47240 ) | ( n47238 & n47240 ) ;
  assign n47242 = n26004 ^ n7385 ^ n1069 ;
  assign n47243 = n43095 & n47242 ;
  assign n47244 = n22146 ^ n11983 ^ n10573 ;
  assign n47245 = ~n11248 & n46432 ;
  assign n47246 = n47245 ^ n18201 ^ 1'b0 ;
  assign n47247 = n31593 & n47246 ;
  assign n47248 = n29314 & n47247 ;
  assign n47251 = n44222 ^ n1261 ^ 1'b0 ;
  assign n47250 = n6048 ^ n5645 ^ 1'b0 ;
  assign n47249 = ( n8926 & ~n12792 ) | ( n8926 & n36848 ) | ( ~n12792 & n36848 ) ;
  assign n47252 = n47251 ^ n47250 ^ n47249 ;
  assign n47253 = ( n10289 & n21154 ) | ( n10289 & n31107 ) | ( n21154 & n31107 ) ;
  assign n47254 = n16926 | n30733 ;
  assign n47255 = n31707 | n47254 ;
  assign n47256 = ( n12410 & n27733 ) | ( n12410 & n47255 ) | ( n27733 & n47255 ) ;
  assign n47257 = n47253 & n47256 ;
  assign n47258 = n19503 & ~n44651 ;
  assign n47259 = n375 & ~n3970 ;
  assign n47260 = n47259 ^ n25838 ^ 1'b0 ;
  assign n47261 = ~n41686 & n47260 ;
  assign n47262 = n24890 & n47261 ;
  assign n47263 = ~n2082 & n41680 ;
  assign n47264 = n47263 ^ n469 ^ 1'b0 ;
  assign n47265 = n1329 & n20433 ;
  assign n47268 = ( ~n8236 & n36805 ) | ( ~n8236 & n45406 ) | ( n36805 & n45406 ) ;
  assign n47266 = n2715 | n10020 ;
  assign n47267 = n12408 | n47266 ;
  assign n47269 = n47268 ^ n47267 ^ 1'b0 ;
  assign n47270 = ( n1103 & n10075 ) | ( n1103 & n15707 ) | ( n10075 & n15707 ) ;
  assign n47271 = n8776 | n47270 ;
  assign n47272 = ~n729 & n1294 ;
  assign n47273 = n38215 & n47272 ;
  assign n47274 = n10188 | n43229 ;
  assign n47275 = n23790 ^ n11852 ^ n3387 ;
  assign n47276 = n47275 ^ n23224 ^ 1'b0 ;
  assign n47277 = ~n5516 & n33004 ;
  assign n47278 = n47277 ^ n25037 ^ 1'b0 ;
  assign n47279 = n37659 | n42090 ;
  assign n47280 = n729 & ~n47279 ;
  assign n47281 = n30156 ^ n28276 ^ 1'b0 ;
  assign n47282 = n2083 & ~n47281 ;
  assign n47283 = ~n40810 & n47282 ;
  assign n47284 = n2802 | n9438 ;
  assign n47285 = n47284 ^ n38089 ^ x97 ;
  assign n47286 = n11140 & ~n28190 ;
  assign n47287 = ~n17541 & n23630 ;
  assign n47290 = n27801 ^ n16012 ^ 1'b0 ;
  assign n47291 = n10480 & ~n47290 ;
  assign n47288 = n21209 ^ n18503 ^ 1'b0 ;
  assign n47289 = n43236 & n47288 ;
  assign n47292 = n47291 ^ n47289 ^ n45512 ;
  assign n47293 = n26686 ^ n10793 ^ n329 ;
  assign n47294 = n24566 | n47293 ;
  assign n47295 = n13743 | n47294 ;
  assign n47296 = n16370 & n29589 ;
  assign n47297 = n30859 | n32709 ;
  assign n47298 = n18204 | n41197 ;
  assign n47299 = n23342 & ~n47298 ;
  assign n47300 = ( ~n862 & n8965 ) | ( ~n862 & n25730 ) | ( n8965 & n25730 ) ;
  assign n47301 = ( n1110 & ~n8433 ) | ( n1110 & n47300 ) | ( ~n8433 & n47300 ) ;
  assign n47303 = n2638 & ~n12382 ;
  assign n47302 = n3621 & ~n11202 ;
  assign n47304 = n47303 ^ n47302 ^ 1'b0 ;
  assign n47305 = ( n3695 & n28575 ) | ( n3695 & n47304 ) | ( n28575 & n47304 ) ;
  assign n47306 = n15487 | n47305 ;
  assign n47307 = n21035 & ~n47306 ;
  assign n47308 = ~n47301 & n47307 ;
  assign n47309 = n47308 ^ n9731 ^ 1'b0 ;
  assign n47310 = n31089 ^ n13555 ^ n9075 ;
  assign n47311 = n33177 ^ n12634 ^ 1'b0 ;
  assign n47312 = ~n16911 & n27751 ;
  assign n47313 = n18292 & ~n18486 ;
  assign n47314 = n4490 | n38419 ;
  assign n47315 = n2035 & n26400 ;
  assign n47316 = n47315 ^ n11596 ^ 1'b0 ;
  assign n47317 = n36659 ^ n10537 ^ 1'b0 ;
  assign n47318 = n5374 & ~n32605 ;
  assign n47319 = ~n29975 & n47318 ;
  assign n47320 = n6948 ^ n5705 ^ 1'b0 ;
  assign n47323 = n15704 ^ n2307 ^ 1'b0 ;
  assign n47324 = ~n15142 & n47323 ;
  assign n47325 = n47324 ^ n12993 ^ 1'b0 ;
  assign n47326 = n24448 | n47325 ;
  assign n47321 = n27885 ^ n6127 ^ 1'b0 ;
  assign n47322 = ~n34748 & n47321 ;
  assign n47327 = n47326 ^ n47322 ^ 1'b0 ;
  assign n47328 = ( n26381 & n47320 ) | ( n26381 & n47327 ) | ( n47320 & n47327 ) ;
  assign n47329 = n19156 ^ n14714 ^ 1'b0 ;
  assign n47330 = n47329 ^ n16073 ^ n604 ;
  assign n47331 = x148 & ~n26646 ;
  assign n47332 = n47331 ^ n17051 ^ 1'b0 ;
  assign n47333 = ( ~n15737 & n22924 ) | ( ~n15737 & n47332 ) | ( n22924 & n47332 ) ;
  assign n47334 = n10552 & n42276 ;
  assign n47335 = ~n23230 & n28238 ;
  assign n47336 = ~n15126 & n20448 ;
  assign n47337 = n47336 ^ n520 ^ 1'b0 ;
  assign n47338 = ~n22076 & n47337 ;
  assign n47339 = n21304 ^ n17932 ^ n7851 ;
  assign n47340 = ~n817 & n2832 ;
  assign n47341 = n47339 & n47340 ;
  assign n47342 = ( n9181 & n9783 ) | ( n9181 & n39149 ) | ( n9783 & n39149 ) ;
  assign n47343 = n44446 & n47342 ;
  assign n47344 = ( n7172 & ~n11221 ) | ( n7172 & n47343 ) | ( ~n11221 & n47343 ) ;
  assign n47345 = ( n2227 & n9596 ) | ( n2227 & n47344 ) | ( n9596 & n47344 ) ;
  assign n47346 = n7707 & n23972 ;
  assign n47347 = ( n1168 & n10165 ) | ( n1168 & ~n47346 ) | ( n10165 & ~n47346 ) ;
  assign n47349 = ~n1626 & n22065 ;
  assign n47350 = n47349 ^ n574 ^ 1'b0 ;
  assign n47351 = n47350 ^ n5991 ^ 1'b0 ;
  assign n47352 = ~n33977 & n47351 ;
  assign n47348 = ( ~n2403 & n17985 ) | ( ~n2403 & n26658 ) | ( n17985 & n26658 ) ;
  assign n47353 = n47352 ^ n47348 ^ 1'b0 ;
  assign n47354 = n39283 ^ n5775 ^ n1595 ;
  assign n47355 = ~n42890 & n47354 ;
  assign n47356 = n47355 ^ n4024 ^ n2394 ;
  assign n47357 = n3605 & ~n41871 ;
  assign n47358 = n29932 ^ n620 ^ 1'b0 ;
  assign n47359 = n7029 & ~n47358 ;
  assign n47360 = n5975 & n25765 ;
  assign n47361 = n47360 ^ n33036 ^ 1'b0 ;
  assign n47362 = n47361 ^ n43224 ^ 1'b0 ;
  assign n47363 = n47359 & n47362 ;
  assign n47364 = n35118 ^ n7125 ^ 1'b0 ;
  assign n47365 = ~n19669 & n47364 ;
  assign n47366 = n6815 | n27707 ;
  assign n47367 = n14054 | n47366 ;
  assign n47368 = ( n4970 & n8124 ) | ( n4970 & ~n43959 ) | ( n8124 & ~n43959 ) ;
  assign n47369 = n36033 | n37072 ;
  assign n47370 = n35713 ^ n21100 ^ n11957 ;
  assign n47371 = n6958 ^ n4402 ^ 1'b0 ;
  assign n47372 = n23294 ^ n18635 ^ n3335 ;
  assign n47373 = n47372 ^ n14509 ^ 1'b0 ;
  assign n47374 = ~n47371 & n47373 ;
  assign n47375 = ~n4986 & n27475 ;
  assign n47376 = n47375 ^ n24501 ^ 1'b0 ;
  assign n47377 = ~n33032 & n43973 ;
  assign n47378 = n4937 | n8893 ;
  assign n47379 = n47378 ^ n23457 ^ 1'b0 ;
  assign n47380 = n39313 & n47379 ;
  assign n47381 = n39178 ^ n25867 ^ 1'b0 ;
  assign n47382 = ~n20596 & n47381 ;
  assign n47383 = n22747 ^ n3698 ^ 1'b0 ;
  assign n47384 = n47382 & ~n47383 ;
  assign n47385 = n36598 ^ n29302 ^ 1'b0 ;
  assign n47386 = ( ~n15832 & n36249 ) | ( ~n15832 & n38806 ) | ( n36249 & n38806 ) ;
  assign n47389 = n23531 ^ n12215 ^ 1'b0 ;
  assign n47390 = n3660 & ~n47389 ;
  assign n47387 = n21018 ^ n9231 ^ 1'b0 ;
  assign n47388 = x226 | n47387 ;
  assign n47391 = n47390 ^ n47388 ^ n20664 ;
  assign n47392 = ~n30508 & n41198 ;
  assign n47393 = n47392 ^ n4792 ^ 1'b0 ;
  assign n47394 = ( n10203 & ~n41082 ) | ( n10203 & n47393 ) | ( ~n41082 & n47393 ) ;
  assign n47395 = n47394 ^ n26646 ^ n14739 ;
  assign n47396 = n27256 ^ n2572 ^ 1'b0 ;
  assign n47397 = n1542 & ~n47396 ;
  assign n47398 = n47397 ^ n26900 ^ 1'b0 ;
  assign n47399 = n33235 & ~n33939 ;
  assign n47400 = n21576 ^ n2189 ^ 1'b0 ;
  assign n47401 = ~n4567 & n11064 ;
  assign n47402 = ~n47400 & n47401 ;
  assign n47403 = n1053 | n40925 ;
  assign n47404 = n32736 & ~n47403 ;
  assign n47405 = ( n5011 & n17161 ) | ( n5011 & n18914 ) | ( n17161 & n18914 ) ;
  assign n47406 = n47405 ^ n42697 ^ 1'b0 ;
  assign n47412 = n17748 | n42784 ;
  assign n47413 = n12043 | n47412 ;
  assign n47407 = n9515 ^ n5381 ^ 1'b0 ;
  assign n47408 = ~n21550 & n47407 ;
  assign n47409 = ~n10516 & n47408 ;
  assign n47410 = n47409 ^ n44605 ^ n5690 ;
  assign n47411 = n25090 & n47410 ;
  assign n47414 = n47413 ^ n47411 ^ 1'b0 ;
  assign n47415 = ~n10636 & n41831 ;
  assign n47416 = ~n13588 & n47415 ;
  assign n47417 = n47416 ^ n20205 ^ 1'b0 ;
  assign n47418 = n42189 & n47417 ;
  assign n47419 = n14725 & ~n18435 ;
  assign n47420 = n47419 ^ n29825 ^ 1'b0 ;
  assign n47421 = n28861 & ~n30573 ;
  assign n47422 = n24578 ^ n22845 ^ n17033 ;
  assign n47423 = n28823 ^ n22777 ^ n7339 ;
  assign n47424 = n2437 ^ n2209 ^ 1'b0 ;
  assign n47425 = n47424 ^ n41220 ^ n12232 ;
  assign n47426 = n45030 ^ n5609 ^ 1'b0 ;
  assign n47427 = n44498 ^ n25278 ^ 1'b0 ;
  assign n47428 = n5961 & n7621 ;
  assign n47429 = ~n15275 & n38595 ;
  assign n47430 = n47428 & n47429 ;
  assign n47431 = ~n9382 & n11217 ;
  assign n47432 = ~n33178 & n47431 ;
  assign n47433 = ( n9618 & n13066 ) | ( n9618 & n23374 ) | ( n13066 & n23374 ) ;
  assign n47434 = n47433 ^ n40949 ^ 1'b0 ;
  assign n47435 = ~n34255 & n47434 ;
  assign n47437 = n25726 ^ n20821 ^ 1'b0 ;
  assign n47436 = ( n498 & n22797 ) | ( n498 & n31410 ) | ( n22797 & n31410 ) ;
  assign n47438 = n47437 ^ n47436 ^ n41051 ;
  assign n47439 = n7766 | n26293 ;
  assign n47440 = n36098 & ~n47439 ;
  assign n47441 = ( n2833 & n24324 ) | ( n2833 & ~n47440 ) | ( n24324 & ~n47440 ) ;
  assign n47442 = n15575 ^ n12950 ^ 1'b0 ;
  assign n47443 = n47442 ^ n42790 ^ n24796 ;
  assign n47444 = n43978 ^ n17489 ^ 1'b0 ;
  assign n47445 = n13226 | n47444 ;
  assign n47446 = n20772 ^ n14454 ^ 1'b0 ;
  assign n47447 = n42322 | n47446 ;
  assign n47448 = n1387 & n41406 ;
  assign n47449 = n47448 ^ n22649 ^ 1'b0 ;
  assign n47450 = ~n15037 & n16749 ;
  assign n47451 = n1530 & n47450 ;
  assign n47452 = n27600 ^ n18472 ^ n4286 ;
  assign n47453 = n19655 ^ n3865 ^ n1294 ;
  assign n47454 = ~n31781 & n33085 ;
  assign n47455 = n47453 & n47454 ;
  assign n47456 = ~n19278 & n47455 ;
  assign n47457 = ( ~n2986 & n36834 ) | ( ~n2986 & n47456 ) | ( n36834 & n47456 ) ;
  assign n47458 = n19903 ^ n11372 ^ 1'b0 ;
  assign n47459 = ( n16227 & n41471 ) | ( n16227 & ~n47458 ) | ( n41471 & ~n47458 ) ;
  assign n47460 = n30013 & ~n32145 ;
  assign n47461 = n47460 ^ n18757 ^ 1'b0 ;
  assign n47462 = ( ~n24293 & n43643 ) | ( ~n24293 & n47461 ) | ( n43643 & n47461 ) ;
  assign n47463 = n14942 ^ n2618 ^ 1'b0 ;
  assign n47464 = ~n2677 & n47463 ;
  assign n47465 = ~n16008 & n47464 ;
  assign n47466 = ~n5432 & n47465 ;
  assign n47467 = n775 | n9885 ;
  assign n47468 = n9885 & ~n47467 ;
  assign n47469 = n31547 | n47468 ;
  assign n47470 = n17488 & n21026 ;
  assign n47471 = ~n21026 & n47470 ;
  assign n47472 = n14936 & ~n22691 ;
  assign n47473 = ~n2529 & n47472 ;
  assign n47474 = n3887 | n47473 ;
  assign n47475 = n47473 & ~n47474 ;
  assign n47476 = n47471 | n47475 ;
  assign n47477 = n47469 & ~n47476 ;
  assign n47478 = n47477 ^ n4668 ^ 1'b0 ;
  assign n47479 = ~n1527 & n20691 ;
  assign n47480 = n3260 & n35578 ;
  assign n47481 = n1635 & n47480 ;
  assign n47482 = ~n19712 & n24019 ;
  assign n47483 = n39105 & n47482 ;
  assign n47484 = ~n31700 & n47483 ;
  assign n47485 = ( n24065 & n29945 ) | ( n24065 & n40742 ) | ( n29945 & n40742 ) ;
  assign n47486 = ( n1258 & n2278 ) | ( n1258 & ~n12049 ) | ( n2278 & ~n12049 ) ;
  assign n47487 = ( n25960 & n40046 ) | ( n25960 & ~n47486 ) | ( n40046 & ~n47486 ) ;
  assign n47488 = x10 & ~n9234 ;
  assign n47489 = ~n403 & n27176 ;
  assign n47490 = n47489 ^ n38358 ^ 1'b0 ;
  assign n47491 = n41451 ^ n31700 ^ n17994 ;
  assign n47492 = n17820 & ~n47491 ;
  assign n47493 = n47492 ^ n45706 ^ 1'b0 ;
  assign n47494 = n35211 ^ n22120 ^ 1'b0 ;
  assign n47495 = n37607 ^ n27507 ^ n21850 ;
  assign n47496 = n15909 ^ n3071 ^ 1'b0 ;
  assign n47497 = n15134 | n30045 ;
  assign n47498 = n20747 | n47497 ;
  assign n47499 = n30623 ^ n30114 ^ n4955 ;
  assign n47500 = n6103 | n47499 ;
  assign n47501 = n38190 ^ n34933 ^ 1'b0 ;
  assign n47502 = n36737 ^ n24397 ^ 1'b0 ;
  assign n47503 = n34559 ^ n2389 ^ 1'b0 ;
  assign n47504 = n33864 ^ n14221 ^ n3629 ;
  assign n47505 = n8908 & n47504 ;
  assign n47506 = n702 ^ x188 ^ 1'b0 ;
  assign n47507 = n22004 ^ n5680 ^ 1'b0 ;
  assign n47508 = n6276 & n47507 ;
  assign n47509 = ( n27295 & n47506 ) | ( n27295 & n47508 ) | ( n47506 & n47508 ) ;
  assign n47510 = x106 & ~n22335 ;
  assign n47511 = n16954 & n47510 ;
  assign n47512 = n7838 & ~n16992 ;
  assign n47513 = n1769 & n11270 ;
  assign n47514 = ~n19459 & n29408 ;
  assign n47515 = n47514 ^ n12749 ^ 1'b0 ;
  assign n47516 = n9617 ^ n7848 ^ 1'b0 ;
  assign n47517 = n39725 | n47516 ;
  assign n47518 = n8138 ^ n2774 ^ 1'b0 ;
  assign n47519 = ( n4039 & n25901 ) | ( n4039 & ~n47518 ) | ( n25901 & ~n47518 ) ;
  assign n47520 = n47519 ^ n42525 ^ n19604 ;
  assign n47521 = n7151 & n34654 ;
  assign n47522 = n39134 ^ n34649 ^ n17553 ;
  assign n47524 = ( ~n7490 & n12174 ) | ( ~n7490 & n13497 ) | ( n12174 & n13497 ) ;
  assign n47523 = n35470 ^ n30230 ^ n23509 ;
  assign n47525 = n47524 ^ n47523 ^ n20501 ;
  assign n47526 = n23128 ^ n21623 ^ n2334 ;
  assign n47527 = n13275 | n47526 ;
  assign n47528 = n47527 ^ n23873 ^ 1'b0 ;
  assign n47529 = ( n16714 & n35506 ) | ( n16714 & n47528 ) | ( n35506 & n47528 ) ;
  assign n47530 = n47529 ^ n38593 ^ 1'b0 ;
  assign n47531 = n20493 & n47530 ;
  assign n47532 = n19874 ^ n9488 ^ 1'b0 ;
  assign n47533 = n30923 | n47532 ;
  assign n47534 = n2046 & n21525 ;
  assign n47535 = ~n14621 & n16519 ;
  assign n47536 = n47534 & n47535 ;
  assign n47537 = ~n28989 & n46962 ;
  assign n47538 = n47536 & n47537 ;
  assign n47539 = n47454 ^ n11207 ^ n5688 ;
  assign n47540 = ( n6484 & ~n9627 ) | ( n6484 & n17545 ) | ( ~n9627 & n17545 ) ;
  assign n47541 = ( n1104 & n38906 ) | ( n1104 & n47540 ) | ( n38906 & n47540 ) ;
  assign n47542 = n7665 ^ n1011 ^ 1'b0 ;
  assign n47543 = ~n30222 & n37518 ;
  assign n47544 = n22304 ^ n3542 ^ 1'b0 ;
  assign n47545 = n29186 ^ n14929 ^ n13863 ;
  assign n47546 = ( ~n22311 & n30129 ) | ( ~n22311 & n47545 ) | ( n30129 & n47545 ) ;
  assign n47547 = n15302 ^ n6448 ^ 1'b0 ;
  assign n47548 = n24522 ^ n5534 ^ 1'b0 ;
  assign n47549 = ~n47547 & n47548 ;
  assign n47550 = ~n47546 & n47549 ;
  assign n47551 = n13734 & ~n29042 ;
  assign n47552 = n5094 ^ n2231 ^ 1'b0 ;
  assign n47553 = n47551 & ~n47552 ;
  assign n47554 = n15933 ^ n13250 ^ n2149 ;
  assign n47555 = n43654 ^ n1069 ^ 1'b0 ;
  assign n47556 = n47554 & n47555 ;
  assign n47557 = n44949 ^ n35181 ^ n5030 ;
  assign n47558 = n27980 ^ n17175 ^ 1'b0 ;
  assign n47559 = n47558 ^ n32381 ^ n18780 ;
  assign n47560 = n47559 ^ n33433 ^ 1'b0 ;
  assign n47562 = n2662 & ~n5032 ;
  assign n47563 = n10938 & n47562 ;
  assign n47561 = n11895 ^ n5102 ^ 1'b0 ;
  assign n47564 = n47563 ^ n47561 ^ n29469 ;
  assign n47565 = n47564 ^ n4538 ^ 1'b0 ;
  assign n47566 = n2831 & n47565 ;
  assign n47567 = n27249 & n46913 ;
  assign n47568 = ~n5434 & n28109 ;
  assign n47569 = n13678 & n47568 ;
  assign n47570 = ( n4311 & n14957 ) | ( n4311 & ~n17676 ) | ( n14957 & ~n17676 ) ;
  assign n47571 = n14265 | n15546 ;
  assign n47572 = n47571 ^ n17976 ^ 1'b0 ;
  assign n47573 = ~n4448 & n47572 ;
  assign n47574 = n4816 & ~n46287 ;
  assign n47575 = ( ~n2082 & n39862 ) | ( ~n2082 & n47574 ) | ( n39862 & n47574 ) ;
  assign n47576 = n47575 ^ n19049 ^ 1'b0 ;
  assign n47577 = n20338 ^ n8927 ^ 1'b0 ;
  assign n47578 = n44167 ^ n4243 ^ 1'b0 ;
  assign n47579 = n37502 & ~n47578 ;
  assign n47580 = n24899 & n47579 ;
  assign n47581 = ( n3728 & n23557 ) | ( n3728 & n47580 ) | ( n23557 & n47580 ) ;
  assign n47582 = ( n3364 & ~n7075 ) | ( n3364 & n13009 ) | ( ~n7075 & n13009 ) ;
  assign n47583 = ~n8263 & n13593 ;
  assign n47584 = ~n7504 & n47583 ;
  assign n47585 = n47584 ^ n5599 ^ 1'b0 ;
  assign n47586 = n20647 ^ n18365 ^ 1'b0 ;
  assign n47587 = n36859 | n47586 ;
  assign n47590 = n6517 ^ n4724 ^ 1'b0 ;
  assign n47591 = ~n34547 & n47590 ;
  assign n47588 = ( x196 & ~n15229 ) | ( x196 & n40515 ) | ( ~n15229 & n40515 ) ;
  assign n47589 = ~n11949 & n47588 ;
  assign n47592 = n47591 ^ n47589 ^ 1'b0 ;
  assign n47593 = ~n7966 & n37536 ;
  assign n47594 = n25601 ^ n18112 ^ 1'b0 ;
  assign n47595 = ~n8739 & n47594 ;
  assign n47596 = n13555 | n33339 ;
  assign n47597 = ( n24231 & n26894 ) | ( n24231 & n36007 ) | ( n26894 & n36007 ) ;
  assign n47598 = n12124 & n47597 ;
  assign n47599 = ( n8810 & n11593 ) | ( n8810 & n37101 ) | ( n11593 & n37101 ) ;
  assign n47600 = n19126 | n39191 ;
  assign n47601 = n33676 ^ n8124 ^ 1'b0 ;
  assign n47602 = n19244 | n47601 ;
  assign n47603 = n47602 ^ n18746 ^ n15086 ;
  assign n47604 = n29652 ^ n3900 ^ 1'b0 ;
  assign n47605 = n284 & ~n3812 ;
  assign n47606 = n44163 & ~n47605 ;
  assign n47607 = n21272 & n36750 ;
  assign n47609 = n38313 ^ n13887 ^ n8039 ;
  assign n47608 = n16765 ^ n2927 ^ 1'b0 ;
  assign n47610 = n47609 ^ n47608 ^ 1'b0 ;
  assign n47611 = ( n12214 & n24642 ) | ( n12214 & ~n41612 ) | ( n24642 & ~n41612 ) ;
  assign n47612 = n18806 | n47611 ;
  assign n47613 = n47612 ^ n6422 ^ 1'b0 ;
  assign n47614 = n29473 ^ n27107 ^ n20283 ;
  assign n47615 = n23651 ^ n16937 ^ 1'b0 ;
  assign n47616 = n20433 & ~n47615 ;
  assign n47617 = n47616 ^ n30106 ^ n16373 ;
  assign n47618 = ( n12129 & n15660 ) | ( n12129 & n47617 ) | ( n15660 & n47617 ) ;
  assign n47619 = ~n25819 & n47618 ;
  assign n47625 = n4609 ^ n4243 ^ 1'b0 ;
  assign n47620 = n3471 & n22407 ;
  assign n47621 = ~n13527 & n47620 ;
  assign n47622 = ( ~n17841 & n33676 ) | ( ~n17841 & n47621 ) | ( n33676 & n47621 ) ;
  assign n47623 = n31918 ^ n21831 ^ 1'b0 ;
  assign n47624 = n47622 | n47623 ;
  assign n47626 = n47625 ^ n47624 ^ n10220 ;
  assign n47633 = n12646 | n31652 ;
  assign n47634 = n12267 & ~n47633 ;
  assign n47628 = n2804 | n30877 ;
  assign n47629 = n17626 | n47628 ;
  assign n47627 = n7439 | n14600 ;
  assign n47630 = n47629 ^ n47627 ^ n17810 ;
  assign n47631 = n47630 ^ n7280 ^ 1'b0 ;
  assign n47632 = ~n24195 & n47631 ;
  assign n47635 = n47634 ^ n47632 ^ n23202 ;
  assign n47636 = n8375 & n28986 ;
  assign n47637 = n34623 ^ n21963 ^ n17753 ;
  assign n47638 = n18153 & ~n47637 ;
  assign n47639 = n28924 ^ n22850 ^ 1'b0 ;
  assign n47640 = n47638 | n47639 ;
  assign n47641 = ( n3425 & ~n6141 ) | ( n3425 & n19388 ) | ( ~n6141 & n19388 ) ;
  assign n47642 = n14328 ^ n5747 ^ 1'b0 ;
  assign n47643 = n47641 & ~n47642 ;
  assign n47644 = n24466 ^ n22420 ^ 1'b0 ;
  assign n47645 = n10014 & ~n12115 ;
  assign n47646 = ( n7761 & n26633 ) | ( n7761 & ~n31657 ) | ( n26633 & ~n31657 ) ;
  assign n47647 = ( n21058 & ~n22782 ) | ( n21058 & n47646 ) | ( ~n22782 & n47646 ) ;
  assign n47648 = n41976 ^ n17551 ^ 1'b0 ;
  assign n47649 = ~n6332 & n12065 ;
  assign n47650 = n5081 ^ n679 ^ 1'b0 ;
  assign n47651 = n6827 | n47650 ;
  assign n47652 = n9966 & ~n27485 ;
  assign n47653 = n47652 ^ n30147 ^ 1'b0 ;
  assign n47654 = n33780 & ~n47653 ;
  assign n47655 = n33620 ^ n2406 ^ 1'b0 ;
  assign n47656 = n28832 ^ n14855 ^ 1'b0 ;
  assign n47657 = ~n47655 & n47656 ;
  assign n47658 = n2566 & ~n3732 ;
  assign n47659 = n26274 ^ n21781 ^ 1'b0 ;
  assign n47660 = ~n12478 & n47659 ;
  assign n47661 = ( ~n3212 & n3989 ) | ( ~n3212 & n6228 ) | ( n3989 & n6228 ) ;
  assign n47662 = ( n34662 & n47660 ) | ( n34662 & n47661 ) | ( n47660 & n47661 ) ;
  assign n47663 = n19728 ^ n5610 ^ 1'b0 ;
  assign n47664 = ( ~n13235 & n46788 ) | ( ~n13235 & n47663 ) | ( n46788 & n47663 ) ;
  assign n47667 = ~n2172 & n38015 ;
  assign n47668 = n47667 ^ n27835 ^ 1'b0 ;
  assign n47669 = n44465 ^ n7590 ^ 1'b0 ;
  assign n47670 = n47668 & n47669 ;
  assign n47666 = n14196 ^ n5538 ^ 1'b0 ;
  assign n47665 = n26049 ^ n20966 ^ n10758 ;
  assign n47671 = n47670 ^ n47666 ^ n47665 ;
  assign n47672 = n35298 ^ n9492 ^ 1'b0 ;
  assign n47673 = n6660 & ~n47672 ;
  assign n47674 = n38809 ^ n738 ^ 1'b0 ;
  assign n47675 = n12779 | n17212 ;
  assign n47676 = n15239 & ~n47675 ;
  assign n47677 = n8545 | n12285 ;
  assign n47678 = n47677 ^ n461 ^ 1'b0 ;
  assign n47679 = n17581 ^ n13182 ^ n3943 ;
  assign n47680 = n47679 ^ n27775 ^ n13878 ;
  assign n47681 = ( ~n17086 & n32260 ) | ( ~n17086 & n45532 ) | ( n32260 & n45532 ) ;
  assign n47682 = n26067 ^ n19367 ^ 1'b0 ;
  assign n47683 = n22430 & n32319 ;
  assign n47684 = n994 & n8695 ;
  assign n47685 = ( ~n18748 & n47683 ) | ( ~n18748 & n47684 ) | ( n47683 & n47684 ) ;
  assign n47686 = n43429 & n47685 ;
  assign n47687 = n7770 & n36170 ;
  assign n47688 = n41081 & n47687 ;
  assign n47689 = ( ~n47682 & n47686 ) | ( ~n47682 & n47688 ) | ( n47686 & n47688 ) ;
  assign n47690 = n26008 ^ n21898 ^ 1'b0 ;
  assign n47691 = n8074 | n24639 ;
  assign n47692 = n47691 ^ n11367 ^ 1'b0 ;
  assign n47693 = n47690 & n47692 ;
  assign n47694 = ~n18995 & n34107 ;
  assign n47695 = n47694 ^ n14427 ^ 1'b0 ;
  assign n47696 = n46696 ^ n6032 ^ 1'b0 ;
  assign n47697 = n13452 & ~n18872 ;
  assign n47698 = n36686 ^ n4827 ^ 1'b0 ;
  assign n47699 = n47698 ^ n33537 ^ 1'b0 ;
  assign n47700 = ~n24335 & n47699 ;
  assign n47701 = n4621 & n46842 ;
  assign n47702 = n496 & ~n10894 ;
  assign n47703 = n47702 ^ n34829 ^ 1'b0 ;
  assign n47704 = ( n20034 & n22227 ) | ( n20034 & ~n38487 ) | ( n22227 & ~n38487 ) ;
  assign n47705 = ( ~n715 & n3956 ) | ( ~n715 & n40900 ) | ( n3956 & n40900 ) ;
  assign n47706 = n15027 ^ n1209 ^ 1'b0 ;
  assign n47707 = n47706 ^ n26458 ^ n24955 ;
  assign n47708 = n35229 | n46805 ;
  assign n47709 = n33850 ^ n4592 ^ 1'b0 ;
  assign n47710 = n39523 ^ n1376 ^ 1'b0 ;
  assign n47711 = n47709 & n47710 ;
  assign n47712 = n4666 ^ n4158 ^ 1'b0 ;
  assign n47713 = n23741 ^ n23092 ^ n789 ;
  assign n47714 = n5124 | n47713 ;
  assign n47715 = n47712 | n47714 ;
  assign n47716 = ~n537 & n2769 ;
  assign n47717 = n17999 & n21872 ;
  assign n47722 = n5062 & ~n13424 ;
  assign n47723 = ~n5062 & n47722 ;
  assign n47724 = x52 & ~n554 ;
  assign n47725 = ~x52 & n47724 ;
  assign n47726 = n7376 | n14965 ;
  assign n47727 = n47725 & ~n47726 ;
  assign n47728 = n47723 | n47727 ;
  assign n47729 = n47723 & ~n47728 ;
  assign n47730 = n4487 & n16375 ;
  assign n47731 = n47729 & n47730 ;
  assign n47732 = n47731 ^ n12636 ^ n1327 ;
  assign n47718 = x72 & n673 ;
  assign n47719 = n47718 ^ n16640 ^ 1'b0 ;
  assign n47720 = ( n9019 & ~n11582 ) | ( n9019 & n33097 ) | ( ~n11582 & n33097 ) ;
  assign n47721 = ( n36056 & ~n47719 ) | ( n36056 & n47720 ) | ( ~n47719 & n47720 ) ;
  assign n47733 = n47732 ^ n47721 ^ 1'b0 ;
  assign n47734 = n36562 ^ n4697 ^ 1'b0 ;
  assign n47735 = n25351 & n47734 ;
  assign n47736 = ( n32025 & n42136 ) | ( n32025 & ~n47735 ) | ( n42136 & ~n47735 ) ;
  assign n47737 = ( ~n12703 & n32614 ) | ( ~n12703 & n43461 ) | ( n32614 & n43461 ) ;
  assign n47738 = n47737 ^ n21623 ^ 1'b0 ;
  assign n47739 = ( n6153 & n14257 ) | ( n6153 & ~n32207 ) | ( n14257 & ~n32207 ) ;
  assign n47740 = ( ~n4973 & n15418 ) | ( ~n4973 & n47739 ) | ( n15418 & n47739 ) ;
  assign n47741 = n6534 & ~n26219 ;
  assign n47742 = ( n3052 & n43562 ) | ( n3052 & ~n47741 ) | ( n43562 & ~n47741 ) ;
  assign n47743 = n27789 ^ n23815 ^ n4928 ;
  assign n47744 = ~n7536 & n47743 ;
  assign n47745 = n13942 | n15634 ;
  assign n47746 = n47745 ^ n29647 ^ 1'b0 ;
  assign n47747 = n9026 ^ n1028 ^ 1'b0 ;
  assign n47748 = n23764 & n47747 ;
  assign n47749 = n37051 ^ n9654 ^ 1'b0 ;
  assign n47750 = n19875 & n23743 ;
  assign n47751 = n43685 ^ n1154 ^ n1088 ;
  assign n47752 = x88 & n47751 ;
  assign n47753 = n39016 | n47752 ;
  assign n47754 = n3782 | n44409 ;
  assign n47755 = n47754 ^ n26236 ^ 1'b0 ;
  assign n47756 = n4928 & n47755 ;
  assign n47757 = n47756 ^ n7827 ^ n2875 ;
  assign n47758 = n12440 | n14663 ;
  assign n47759 = n22656 & ~n47758 ;
  assign n47760 = n47759 ^ n32779 ^ 1'b0 ;
  assign n47761 = n2331 & ~n16638 ;
  assign n47762 = n47761 ^ n21235 ^ n11791 ;
  assign n47763 = n47762 ^ n25135 ^ 1'b0 ;
  assign n47764 = ( n18557 & n27880 ) | ( n18557 & n47763 ) | ( n27880 & n47763 ) ;
  assign n47765 = n4579 & n22227 ;
  assign n47766 = n33842 ^ n2680 ^ 1'b0 ;
  assign n47767 = ~n27393 & n47766 ;
  assign n47768 = n23822 & ~n30973 ;
  assign n47769 = n47768 ^ n13102 ^ 1'b0 ;
  assign n47770 = n4785 ^ n4243 ^ 1'b0 ;
  assign n47771 = n9882 | n43915 ;
  assign n47772 = n20634 ^ n20185 ^ n5246 ;
  assign n47780 = n20040 ^ n13009 ^ n4254 ;
  assign n47777 = n2262 & ~n14023 ;
  assign n47775 = n15546 & n21658 ;
  assign n47776 = ~n43358 & n47775 ;
  assign n47778 = n47777 ^ n47776 ^ n42535 ;
  assign n47774 = n25646 ^ n13097 ^ 1'b0 ;
  assign n47779 = n47778 ^ n47774 ^ 1'b0 ;
  assign n47773 = n30101 ^ n7812 ^ 1'b0 ;
  assign n47781 = n47780 ^ n47779 ^ n47773 ;
  assign n47782 = n42333 ^ n28384 ^ 1'b0 ;
  assign n47783 = n12576 ^ n9803 ^ 1'b0 ;
  assign n47784 = ~n46947 & n47783 ;
  assign n47785 = n39833 ^ n28877 ^ 1'b0 ;
  assign n47786 = n2452 & n47785 ;
  assign n47787 = n6618 & n41374 ;
  assign n47788 = n16006 & n47787 ;
  assign n47789 = ~n10517 & n47788 ;
  assign n47790 = n6362 & ~n25851 ;
  assign n47791 = n7810 & n47790 ;
  assign n47792 = ( n10201 & ~n13967 ) | ( n10201 & n18742 ) | ( ~n13967 & n18742 ) ;
  assign n47793 = ~n7918 & n27509 ;
  assign n47794 = n7739 | n28577 ;
  assign n47795 = n4581 & n25319 ;
  assign n47796 = ~n40294 & n47795 ;
  assign n47797 = ~n9699 & n26160 ;
  assign n47798 = n9906 & n47797 ;
  assign n47799 = ( n10758 & n11125 ) | ( n10758 & n24862 ) | ( n11125 & n24862 ) ;
  assign n47800 = n47799 ^ x103 ^ 1'b0 ;
  assign n47801 = n310 & n47800 ;
  assign n47802 = n33573 ^ n9422 ^ n8523 ;
  assign n47803 = n47802 ^ n13569 ^ 1'b0 ;
  assign n47806 = n20722 ^ n1026 ^ 1'b0 ;
  assign n47804 = n2551 ^ x159 ^ 1'b0 ;
  assign n47805 = ~n17301 & n47804 ;
  assign n47807 = n47806 ^ n47805 ^ n37283 ;
  assign n47808 = n29020 ^ n7008 ^ 1'b0 ;
  assign n47809 = n30731 & n47808 ;
  assign n47810 = n11659 ^ n602 ^ 1'b0 ;
  assign n47811 = n47810 ^ n29653 ^ n7325 ;
  assign n47812 = ( n3351 & n6453 ) | ( n3351 & n44568 ) | ( n6453 & n44568 ) ;
  assign n47815 = ( ~n7142 & n9084 ) | ( ~n7142 & n10825 ) | ( n9084 & n10825 ) ;
  assign n47813 = n4623 ^ n1324 ^ 1'b0 ;
  assign n47814 = ~n44654 & n47813 ;
  assign n47816 = n47815 ^ n47814 ^ 1'b0 ;
  assign n47817 = n9650 & ~n23301 ;
  assign n47818 = n47817 ^ n19696 ^ 1'b0 ;
  assign n47819 = n18440 & ~n47818 ;
  assign n47822 = n654 & n9659 ;
  assign n47823 = ~n13888 & n47822 ;
  assign n47824 = n2993 & n47823 ;
  assign n47820 = n9890 ^ n2771 ^ x210 ;
  assign n47821 = n22492 | n47820 ;
  assign n47825 = n47824 ^ n47821 ^ 1'b0 ;
  assign n47826 = n13888 ^ n10185 ^ n888 ;
  assign n47827 = n47826 ^ n39038 ^ 1'b0 ;
  assign n47828 = n25813 & n47827 ;
  assign n47829 = n922 & ~n21736 ;
  assign n47830 = n20353 ^ n1775 ^ 1'b0 ;
  assign n47831 = n9676 ^ n9332 ^ n2888 ;
  assign n47832 = ( ~n31591 & n42618 ) | ( ~n31591 & n47831 ) | ( n42618 & n47831 ) ;
  assign n47833 = n47832 ^ n37748 ^ n23059 ;
  assign n47835 = n11970 ^ n297 ^ 1'b0 ;
  assign n47834 = ~n11454 & n21180 ;
  assign n47836 = n47835 ^ n47834 ^ 1'b0 ;
  assign n47837 = n22408 | n47836 ;
  assign n47841 = ( n5497 & n19212 ) | ( n5497 & ~n44057 ) | ( n19212 & ~n44057 ) ;
  assign n47840 = n7210 ^ n1327 ^ 1'b0 ;
  assign n47838 = n7326 & ~n15518 ;
  assign n47839 = ( n11945 & ~n29797 ) | ( n11945 & n47838 ) | ( ~n29797 & n47838 ) ;
  assign n47842 = n47841 ^ n47840 ^ n47839 ;
  assign n47843 = n31331 ^ n9949 ^ 1'b0 ;
  assign n47844 = n16031 | n47843 ;
  assign n47845 = n18493 ^ n2821 ^ 1'b0 ;
  assign n47846 = n5123 & n47845 ;
  assign n47847 = n47846 ^ n15776 ^ 1'b0 ;
  assign n47848 = ~n47844 & n47847 ;
  assign n47849 = ( n22716 & n26557 ) | ( n22716 & n47848 ) | ( n26557 & n47848 ) ;
  assign n47850 = n34508 ^ n5756 ^ 1'b0 ;
  assign n47851 = n15896 ^ n11941 ^ n4628 ;
  assign n47852 = n2809 | n4890 ;
  assign n47853 = n47852 ^ n20843 ^ n3310 ;
  assign n47854 = ( n29653 & ~n47851 ) | ( n29653 & n47853 ) | ( ~n47851 & n47853 ) ;
  assign n47855 = n47854 ^ n30730 ^ 1'b0 ;
  assign n47856 = n8142 & n47855 ;
  assign n47857 = ~n26791 & n47856 ;
  assign n47858 = n7693 & n33002 ;
  assign n47859 = n10712 & n47858 ;
  assign n47861 = n31696 ^ n931 ^ 1'b0 ;
  assign n47860 = ~n23664 & n26431 ;
  assign n47862 = n47861 ^ n47860 ^ 1'b0 ;
  assign n47863 = n33041 ^ n30926 ^ 1'b0 ;
  assign n47864 = ( n3354 & n8839 ) | ( n3354 & n47863 ) | ( n8839 & n47863 ) ;
  assign n47865 = n47864 ^ n19795 ^ 1'b0 ;
  assign n47866 = n20776 & ~n47865 ;
  assign n47867 = n3977 & n47866 ;
  assign n47868 = n25678 & ~n35309 ;
  assign n47869 = n13895 & n47868 ;
  assign n47870 = n47869 ^ n41404 ^ n10606 ;
  assign n47871 = n14422 | n33239 ;
  assign n47872 = n6538 & n25254 ;
  assign n47873 = n47872 ^ n25927 ^ n22916 ;
  assign n47874 = n41741 ^ n6693 ^ n4471 ;
  assign n47875 = n12789 ^ n5546 ^ 1'b0 ;
  assign n47876 = n27324 | n35323 ;
  assign n47877 = n47875 & ~n47876 ;
  assign n47878 = ~n10753 & n22114 ;
  assign n47879 = n47878 ^ n20215 ^ 1'b0 ;
  assign n47880 = n47879 ^ n6350 ^ 1'b0 ;
  assign n47881 = n14446 | n22190 ;
  assign n47882 = n18880 & ~n29192 ;
  assign n47883 = n47882 ^ n38769 ^ 1'b0 ;
  assign n47884 = n31331 ^ n19633 ^ 1'b0 ;
  assign n47885 = ( n9835 & n19424 ) | ( n9835 & n24157 ) | ( n19424 & n24157 ) ;
  assign n47886 = n7110 | n40239 ;
  assign n47887 = n10120 ^ x87 ^ 1'b0 ;
  assign n47888 = n14586 | n47887 ;
  assign n47889 = n24991 | n40545 ;
  assign n47890 = n47888 & ~n47889 ;
  assign n47891 = n47890 ^ n43359 ^ n32529 ;
  assign n47892 = n13905 | n35582 ;
  assign n47893 = n17898 & ~n47892 ;
  assign n47894 = n23685 ^ n20347 ^ n16022 ;
  assign n47895 = ~n37481 & n47894 ;
  assign n47896 = n47895 ^ n7379 ^ 1'b0 ;
  assign n47897 = n43604 ^ n3050 ^ 1'b0 ;
  assign n47898 = n30660 & ~n47897 ;
  assign n47899 = n500 & n6363 ;
  assign n47900 = ~n12880 & n47899 ;
  assign n47901 = n47900 ^ n32573 ^ n32141 ;
  assign n47902 = n47901 ^ n9132 ^ 1'b0 ;
  assign n47903 = n7561 & ~n47902 ;
  assign n47904 = n4536 & n47903 ;
  assign n47905 = ( n2611 & n7468 ) | ( n2611 & n17685 ) | ( n7468 & n17685 ) ;
  assign n47906 = n47905 ^ n1476 ^ 1'b0 ;
  assign n47907 = n47904 & ~n47906 ;
  assign n47908 = n34647 ^ n2809 ^ 1'b0 ;
  assign n47909 = ~n21439 & n47908 ;
  assign n47910 = n3263 | n13372 ;
  assign n47911 = n1635 & ~n8114 ;
  assign n47912 = n47911 ^ n17108 ^ n3857 ;
  assign n47913 = ( n4709 & n9206 ) | ( n4709 & n28070 ) | ( n9206 & n28070 ) ;
  assign n47914 = n47913 ^ n29649 ^ n8459 ;
  assign n47915 = n33590 ^ n25455 ^ x181 ;
  assign n47916 = n24545 ^ n8363 ^ n1512 ;
  assign n47917 = n38847 ^ n32471 ^ n22346 ;
  assign n47918 = ~n6221 & n47917 ;
  assign n47919 = ~n7747 & n43765 ;
  assign n47920 = n6382 ^ n4985 ^ 1'b0 ;
  assign n47921 = n15873 & ~n21654 ;
  assign n47922 = ~n47920 & n47921 ;
  assign n47923 = n14366 ^ n921 ^ 1'b0 ;
  assign n47924 = n47923 ^ n15991 ^ 1'b0 ;
  assign n47925 = n1403 & n6606 ;
  assign n47926 = ~n16171 & n47925 ;
  assign n47927 = ~n2910 & n31119 ;
  assign n47928 = ~n30880 & n47927 ;
  assign n47929 = n22513 | n47928 ;
  assign n47930 = ( n13512 & n34332 ) | ( n13512 & ~n47929 ) | ( n34332 & ~n47929 ) ;
  assign n47931 = n46657 & n47930 ;
  assign n47932 = n12748 ^ n3470 ^ 1'b0 ;
  assign n47933 = ( n7805 & ~n35309 ) | ( n7805 & n47932 ) | ( ~n35309 & n47932 ) ;
  assign n47934 = n47933 ^ n6992 ^ 1'b0 ;
  assign n47935 = n47934 ^ n13267 ^ 1'b0 ;
  assign n47936 = n22469 ^ n10061 ^ 1'b0 ;
  assign n47937 = n33530 ^ n5729 ^ 1'b0 ;
  assign n47938 = ~n11163 & n47937 ;
  assign n47939 = n47938 ^ n1644 ^ 1'b0 ;
  assign n47941 = ~n7064 & n7160 ;
  assign n47940 = ~n24824 & n29326 ;
  assign n47942 = n47941 ^ n47940 ^ 1'b0 ;
  assign n47943 = n405 & ~n32357 ;
  assign n47944 = n47943 ^ n22575 ^ 1'b0 ;
  assign n47945 = n46649 ^ n8507 ^ 1'b0 ;
  assign n47946 = ~n39935 & n47945 ;
  assign n47947 = n6041 | n16038 ;
  assign n47948 = n28508 & ~n47947 ;
  assign n47949 = n14333 | n32089 ;
  assign n47950 = n47949 ^ n26311 ^ n22127 ;
  assign n47951 = n47327 ^ n24968 ^ n6023 ;
  assign n47952 = n17333 ^ n13262 ^ 1'b0 ;
  assign n47953 = n41010 ^ n35392 ^ n18015 ;
  assign n47954 = n44203 & n47953 ;
  assign n47955 = n13863 | n18138 ;
  assign n47956 = ~n18971 & n47955 ;
  assign n47957 = ~n12524 & n47956 ;
  assign n47958 = n6459 ^ n4592 ^ 1'b0 ;
  assign n47959 = n35164 ^ n10140 ^ n870 ;
  assign n47960 = ~n25303 & n47959 ;
  assign n47961 = n47960 ^ n22515 ^ 1'b0 ;
  assign n47962 = n1104 & n47961 ;
  assign n47963 = ~n46475 & n47962 ;
  assign n47964 = n47963 ^ n24422 ^ 1'b0 ;
  assign n47965 = n25645 ^ n2929 ^ 1'b0 ;
  assign n47966 = n47965 ^ n41633 ^ n1828 ;
  assign n47967 = n8539 | n13678 ;
  assign n47968 = n47967 ^ n30066 ^ n4209 ;
  assign n47969 = n47968 ^ n33453 ^ 1'b0 ;
  assign n47970 = n42076 ^ n11579 ^ 1'b0 ;
  assign n47971 = n45207 & n47970 ;
  assign n47972 = n19097 & n29677 ;
  assign n47973 = n1927 & n47972 ;
  assign n47974 = n6147 ^ n578 ^ 1'b0 ;
  assign n47975 = ~n47973 & n47974 ;
  assign n47976 = ~n14266 & n32763 ;
  assign n47977 = n44416 & n47976 ;
  assign n47978 = n38375 ^ n32649 ^ n14711 ;
  assign n47979 = n47978 ^ n14714 ^ 1'b0 ;
  assign n47983 = n32514 ^ n2983 ^ 1'b0 ;
  assign n47984 = n33779 | n47983 ;
  assign n47980 = n46009 ^ n33330 ^ n21471 ;
  assign n47981 = n25207 & n29453 ;
  assign n47982 = ~n47980 & n47981 ;
  assign n47985 = n47984 ^ n47982 ^ 1'b0 ;
  assign n47986 = ( ~n7004 & n15473 ) | ( ~n7004 & n16735 ) | ( n15473 & n16735 ) ;
  assign n47987 = n35294 ^ n25079 ^ n997 ;
  assign n47988 = n35106 ^ n9115 ^ 1'b0 ;
  assign n47989 = n19688 & n47988 ;
  assign n47990 = n42847 ^ n30258 ^ 1'b0 ;
  assign n47991 = ( n4398 & n11739 ) | ( n4398 & n23455 ) | ( n11739 & n23455 ) ;
  assign n47992 = n10799 & ~n14965 ;
  assign n47993 = n47992 ^ n16333 ^ 1'b0 ;
  assign n47994 = n47993 ^ n19239 ^ n10325 ;
  assign n47995 = n44742 ^ n43742 ^ 1'b0 ;
  assign n47996 = n8222 & ~n47995 ;
  assign n47997 = ( n7433 & n32213 ) | ( n7433 & n47996 ) | ( n32213 & n47996 ) ;
  assign n47998 = n26783 ^ n25213 ^ 1'b0 ;
  assign n47999 = n318 & ~n36686 ;
  assign n48000 = ~n25144 & n47999 ;
  assign n48001 = n37094 & ~n48000 ;
  assign n48002 = n48001 ^ n13679 ^ 1'b0 ;
  assign n48003 = n41809 ^ n12488 ^ 1'b0 ;
  assign n48004 = ~n48002 & n48003 ;
  assign n48005 = ( n12167 & ~n13356 ) | ( n12167 & n18722 ) | ( ~n13356 & n18722 ) ;
  assign n48006 = n48005 ^ n11766 ^ 1'b0 ;
  assign n48007 = n31258 ^ n14741 ^ 1'b0 ;
  assign n48008 = n1061 | n13689 ;
  assign n48009 = n17690 | n48008 ;
  assign n48010 = n30878 ^ n3500 ^ 1'b0 ;
  assign n48011 = n29090 & n38552 ;
  assign n48012 = ~n15149 & n48011 ;
  assign n48013 = n47268 ^ n11140 ^ 1'b0 ;
  assign n48014 = ( ~n11379 & n19659 ) | ( ~n11379 & n35933 ) | ( n19659 & n35933 ) ;
  assign n48015 = n48014 ^ n3817 ^ 1'b0 ;
  assign n48016 = n23242 & ~n40219 ;
  assign n48017 = ~n41680 & n48016 ;
  assign n48018 = n37633 ^ n34783 ^ 1'b0 ;
  assign n48019 = n5674 ^ n4701 ^ 1'b0 ;
  assign n48020 = ~n14101 & n48019 ;
  assign n48021 = n48020 ^ n10727 ^ 1'b0 ;
  assign n48022 = n37621 | n48021 ;
  assign n48023 = n18524 & ~n48022 ;
  assign n48024 = n27026 ^ n12450 ^ n11000 ;
  assign n48025 = n39283 & n48024 ;
  assign n48029 = n43065 ^ n11554 ^ n304 ;
  assign n48028 = n5235 | n31330 ;
  assign n48030 = n48029 ^ n48028 ^ 1'b0 ;
  assign n48026 = n29488 ^ n10024 ^ 1'b0 ;
  assign n48027 = n1000 | n48026 ;
  assign n48031 = n48030 ^ n48027 ^ n35548 ;
  assign n48032 = n16390 ^ n12607 ^ 1'b0 ;
  assign n48033 = n48031 | n48032 ;
  assign n48034 = n8573 ^ n5611 ^ 1'b0 ;
  assign n48035 = ~n24035 & n48034 ;
  assign n48036 = n18138 ^ n7897 ^ 1'b0 ;
  assign n48037 = n48036 ^ n27005 ^ n4694 ;
  assign n48038 = n26312 ^ n15886 ^ n938 ;
  assign n48039 = ( n30037 & n46286 ) | ( n30037 & ~n48038 ) | ( n46286 & ~n48038 ) ;
  assign n48040 = n28613 ^ n5965 ^ n3589 ;
  assign n48041 = n24304 & ~n33784 ;
  assign n48045 = n7068 ^ n5712 ^ 1'b0 ;
  assign n48046 = n966 & n48045 ;
  assign n48047 = n48046 ^ n3541 ^ n945 ;
  assign n48048 = n30525 & ~n48047 ;
  assign n48042 = n9566 ^ n3512 ^ 1'b0 ;
  assign n48043 = n2219 & ~n48042 ;
  assign n48044 = n5798 & n48043 ;
  assign n48049 = n48048 ^ n48044 ^ n35771 ;
  assign n48050 = n20299 ^ n4164 ^ 1'b0 ;
  assign n48051 = n48049 | n48050 ;
  assign n48052 = x211 ^ x114 ^ 1'b0 ;
  assign n48053 = n2118 | n9996 ;
  assign n48054 = n48053 ^ n14395 ^ 1'b0 ;
  assign n48055 = n12539 | n48054 ;
  assign n48056 = n48052 | n48055 ;
  assign n48057 = n25757 & n27238 ;
  assign n48058 = n48057 ^ n1512 ^ 1'b0 ;
  assign n48059 = n48058 ^ n8668 ^ 1'b0 ;
  assign n48060 = n14829 | n33879 ;
  assign n48061 = n48060 ^ n25630 ^ 1'b0 ;
  assign n48062 = n48061 ^ n8352 ^ 1'b0 ;
  assign n48063 = n23140 & n39339 ;
  assign n48064 = n48063 ^ n40499 ^ 1'b0 ;
  assign n48065 = ( n4367 & ~n43691 ) | ( n4367 & n48064 ) | ( ~n43691 & n48064 ) ;
  assign n48066 = n19624 ^ n1536 ^ 1'b0 ;
  assign n48067 = n12944 & ~n48066 ;
  assign n48068 = ( ~n7848 & n36220 ) | ( ~n7848 & n48067 ) | ( n36220 & n48067 ) ;
  assign n48069 = ( n3045 & n23619 ) | ( n3045 & ~n29020 ) | ( n23619 & ~n29020 ) ;
  assign n48070 = n12359 ^ n7097 ^ 1'b0 ;
  assign n48072 = ( ~n3798 & n13879 ) | ( ~n3798 & n19737 ) | ( n13879 & n19737 ) ;
  assign n48071 = n12742 & n24293 ;
  assign n48073 = n48072 ^ n48071 ^ 1'b0 ;
  assign n48074 = n1766 | n32914 ;
  assign n48075 = n18941 ^ n843 ^ 1'b0 ;
  assign n48076 = ~n12219 & n48075 ;
  assign n48077 = n48076 ^ n9594 ^ 1'b0 ;
  assign n48078 = n48074 & ~n48077 ;
  assign n48079 = n38023 ^ n6272 ^ 1'b0 ;
  assign n48080 = n44449 & n48079 ;
  assign n48081 = n8970 & n42868 ;
  assign n48082 = n4357 & n48081 ;
  assign n48083 = n7694 | n33541 ;
  assign n48084 = n46228 ^ n31045 ^ 1'b0 ;
  assign n48085 = n37757 | n48084 ;
  assign n48086 = n3869 | n24129 ;
  assign n48087 = n48086 ^ n35689 ^ 1'b0 ;
  assign n48088 = n9807 | n48087 ;
  assign n48089 = ( ~n13554 & n20512 ) | ( ~n13554 & n32629 ) | ( n20512 & n32629 ) ;
  assign n48090 = n28281 ^ n27537 ^ n19572 ;
  assign n48093 = n16715 ^ n16613 ^ n1318 ;
  assign n48091 = n7701 | n31696 ;
  assign n48092 = n48091 ^ n32972 ^ 1'b0 ;
  assign n48094 = n48093 ^ n48092 ^ n15078 ;
  assign n48095 = n30629 ^ n10174 ^ 1'b0 ;
  assign n48096 = n8463 ^ n4407 ^ 1'b0 ;
  assign n48097 = n15081 & ~n48096 ;
  assign n48098 = ~n2440 & n48097 ;
  assign n48099 = n11603 | n13061 ;
  assign n48100 = n21658 | n48099 ;
  assign n48101 = n48100 ^ n39776 ^ n23448 ;
  assign n48102 = n4928 | n48101 ;
  assign n48103 = n23732 & ~n26809 ;
  assign n48104 = n43639 ^ n29224 ^ 1'b0 ;
  assign n48105 = n7808 ^ n5011 ^ 1'b0 ;
  assign n48106 = n873 & n27495 ;
  assign n48107 = n48106 ^ n629 ^ 1'b0 ;
  assign n48108 = n40397 & ~n48107 ;
  assign n48109 = ( ~n48104 & n48105 ) | ( ~n48104 & n48108 ) | ( n48105 & n48108 ) ;
  assign n48110 = ( n6745 & n11489 ) | ( n6745 & ~n22701 ) | ( n11489 & ~n22701 ) ;
  assign n48111 = ~n18209 & n48110 ;
  assign n48112 = n48111 ^ n22896 ^ 1'b0 ;
  assign n48113 = ( ~n12711 & n35196 ) | ( ~n12711 & n48112 ) | ( n35196 & n48112 ) ;
  assign n48114 = ( ~n8507 & n26606 ) | ( ~n8507 & n35892 ) | ( n26606 & n35892 ) ;
  assign n48115 = n48114 ^ n12657 ^ 1'b0 ;
  assign n48116 = ~n10704 & n37680 ;
  assign n48117 = n6287 & ~n16086 ;
  assign n48118 = ~n22918 & n48117 ;
  assign n48119 = n48118 ^ n25101 ^ 1'b0 ;
  assign n48120 = n11733 & n17921 ;
  assign n48121 = n15989 & n48120 ;
  assign n48122 = n23593 ^ n1980 ^ 1'b0 ;
  assign n48123 = ~n32570 & n48122 ;
  assign n48124 = n48123 ^ n33143 ^ n14549 ;
  assign n48125 = n48124 ^ n37963 ^ 1'b0 ;
  assign n48126 = ( ~n3521 & n12291 ) | ( ~n3521 & n48125 ) | ( n12291 & n48125 ) ;
  assign n48131 = n22162 | n23745 ;
  assign n48127 = n30474 & n40347 ;
  assign n48128 = n34199 & n38644 ;
  assign n48129 = n34023 & n48128 ;
  assign n48130 = n48127 & n48129 ;
  assign n48132 = n48131 ^ n48130 ^ 1'b0 ;
  assign n48133 = n38335 ^ n36644 ^ n9907 ;
  assign n48139 = ~n16870 & n33177 ;
  assign n48140 = n16815 & n48139 ;
  assign n48134 = n15192 ^ n8660 ^ 1'b0 ;
  assign n48135 = n10611 & ~n48134 ;
  assign n48136 = n48135 ^ n15769 ^ 1'b0 ;
  assign n48137 = n11393 | n48136 ;
  assign n48138 = n48137 ^ n9468 ^ 1'b0 ;
  assign n48141 = n48140 ^ n48138 ^ n31374 ;
  assign n48142 = n40842 ^ n39813 ^ 1'b0 ;
  assign n48143 = ~n20327 & n48142 ;
  assign n48144 = ~n3726 & n40589 ;
  assign n48145 = n13762 & n17415 ;
  assign n48146 = n48145 ^ n8305 ^ 1'b0 ;
  assign n48147 = ~n5897 & n48146 ;
  assign n48148 = n2676 | n12151 ;
  assign n48149 = n14159 & ~n14628 ;
  assign n48150 = n17751 ^ n10172 ^ 1'b0 ;
  assign n48151 = n18297 & n48150 ;
  assign n48152 = n18967 & ~n48151 ;
  assign n48153 = n11416 & n27840 ;
  assign n48154 = n48153 ^ n13365 ^ 1'b0 ;
  assign n48155 = ( n32569 & ~n32574 ) | ( n32569 & n48154 ) | ( ~n32574 & n48154 ) ;
  assign n48156 = ( ~n6287 & n7961 ) | ( ~n6287 & n20299 ) | ( n7961 & n20299 ) ;
  assign n48157 = n48156 ^ n9739 ^ n2584 ;
  assign n48158 = n7267 & ~n40701 ;
  assign n48159 = n6060 & ~n20597 ;
  assign n48160 = n38360 & n48159 ;
  assign n48161 = n18087 | n32950 ;
  assign n48162 = n2099 & ~n15435 ;
  assign n48163 = n48162 ^ n1499 ^ 1'b0 ;
  assign n48164 = n48163 ^ n32337 ^ 1'b0 ;
  assign n48165 = n33903 ^ n26673 ^ 1'b0 ;
  assign n48166 = n14737 & ~n48165 ;
  assign n48167 = ( n9008 & n14300 ) | ( n9008 & n39523 ) | ( n14300 & n39523 ) ;
  assign n48168 = n1455 & n12356 ;
  assign n48169 = n35369 ^ n25303 ^ n18238 ;
  assign n48170 = n16191 ^ n1641 ^ 1'b0 ;
  assign n48171 = ~n7446 & n41783 ;
  assign n48172 = ~n36442 & n48171 ;
  assign n48173 = ~n19411 & n21382 ;
  assign n48174 = n48173 ^ n18646 ^ 1'b0 ;
  assign n48175 = n3546 | n6589 ;
  assign n48176 = n48175 ^ n8900 ^ 1'b0 ;
  assign n48177 = ( n4163 & ~n9221 ) | ( n4163 & n37761 ) | ( ~n9221 & n37761 ) ;
  assign n48178 = n5159 | n45868 ;
  assign n48179 = n48177 & ~n48178 ;
  assign n48180 = n31205 | n48179 ;
  assign n48181 = n33116 & ~n48180 ;
  assign n48182 = ~n39861 & n47937 ;
  assign n48183 = ~n5591 & n21591 ;
  assign n48184 = n48183 ^ n26203 ^ n19775 ;
  assign n48185 = n47698 ^ n44472 ^ 1'b0 ;
  assign n48186 = n22827 ^ n1760 ^ 1'b0 ;
  assign n48187 = n48186 ^ n18516 ^ 1'b0 ;
  assign n48188 = n41105 ^ n38818 ^ 1'b0 ;
  assign n48189 = ~n27523 & n35019 ;
  assign n48191 = n17756 ^ n5875 ^ 1'b0 ;
  assign n48190 = n2499 & n21855 ;
  assign n48192 = n48191 ^ n48190 ^ 1'b0 ;
  assign n48193 = n3408 & ~n25974 ;
  assign n48194 = x192 & n10332 ;
  assign n48195 = ~n48193 & n48194 ;
  assign n48196 = n12275 ^ n3999 ^ 1'b0 ;
  assign n48197 = n4955 | n48196 ;
  assign n48198 = n43374 | n48197 ;
  assign n48199 = n19324 ^ n12600 ^ n5616 ;
  assign n48200 = n6905 & n16678 ;
  assign n48201 = n48200 ^ n11623 ^ 1'b0 ;
  assign n48202 = x117 & n5814 ;
  assign n48203 = n48104 ^ n27172 ^ n19482 ;
  assign n48204 = ( ~n2313 & n48202 ) | ( ~n2313 & n48203 ) | ( n48202 & n48203 ) ;
  assign n48205 = n11285 ^ n5938 ^ 1'b0 ;
  assign n48206 = n11871 | n48205 ;
  assign n48207 = n48206 ^ n30746 ^ n24400 ;
  assign n48208 = ( ~n9138 & n13374 ) | ( ~n9138 & n25410 ) | ( n13374 & n25410 ) ;
  assign n48209 = ( ~n23559 & n42647 ) | ( ~n23559 & n45307 ) | ( n42647 & n45307 ) ;
  assign n48210 = ~n9373 & n46306 ;
  assign n48211 = n48210 ^ n3642 ^ 1'b0 ;
  assign n48212 = n38338 ^ n12378 ^ 1'b0 ;
  assign n48213 = n22497 | n48212 ;
  assign n48214 = n12713 & n41554 ;
  assign n48215 = n48213 & n48214 ;
  assign n48216 = ( n25893 & n26913 ) | ( n25893 & n32795 ) | ( n26913 & n32795 ) ;
  assign n48217 = n12378 & n48216 ;
  assign n48218 = ( n10162 & n18713 ) | ( n10162 & n34149 ) | ( n18713 & n34149 ) ;
  assign n48219 = ( ~n1351 & n25354 ) | ( ~n1351 & n48218 ) | ( n25354 & n48218 ) ;
  assign n48220 = n29364 ^ n8838 ^ 1'b0 ;
  assign n48221 = n24370 | n48220 ;
  assign n48222 = n46782 ^ n6502 ^ 1'b0 ;
  assign n48223 = n34860 & ~n40919 ;
  assign n48224 = n4548 | n22070 ;
  assign n48225 = n48224 ^ n3080 ^ 1'b0 ;
  assign n48226 = n30109 | n39246 ;
  assign n48227 = n14600 | n18365 ;
  assign n48228 = n11288 ^ n10705 ^ n9845 ;
  assign n48229 = n9529 | n37979 ;
  assign n48230 = n37607 ^ n3954 ^ 1'b0 ;
  assign n48231 = n39313 ^ n18364 ^ 1'b0 ;
  assign n48232 = n803 & n7359 ;
  assign n48233 = x32 & n36657 ;
  assign n48234 = ( ~n8116 & n23845 ) | ( ~n8116 & n36275 ) | ( n23845 & n36275 ) ;
  assign n48235 = n18765 ^ n5274 ^ 1'b0 ;
  assign n48236 = n30994 ^ n27466 ^ n6436 ;
  assign n48237 = n5211 ^ n5114 ^ n729 ;
  assign n48238 = n48237 ^ n17098 ^ 1'b0 ;
  assign n48239 = n48238 ^ n26849 ^ n12288 ;
  assign n48240 = n42759 ^ n18997 ^ 1'b0 ;
  assign n48241 = n35972 ^ n30046 ^ 1'b0 ;
  assign n48242 = n24780 ^ n23099 ^ 1'b0 ;
  assign n48243 = n19764 & n48242 ;
  assign n48244 = n48243 ^ n12498 ^ n12314 ;
  assign n48245 = n48244 ^ n4769 ^ 1'b0 ;
  assign n48246 = n30636 ^ n3308 ^ 1'b0 ;
  assign n48247 = n15886 & ~n48246 ;
  assign n48248 = n40474 ^ n24058 ^ n5107 ;
  assign n48249 = n48248 ^ n5657 ^ 1'b0 ;
  assign n48250 = x2 & ~n7881 ;
  assign n48251 = n48250 ^ n7791 ^ n5031 ;
  assign n48252 = ( n22001 & ~n25306 ) | ( n22001 & n48251 ) | ( ~n25306 & n48251 ) ;
  assign n48253 = n6904 ^ n3657 ^ n3568 ;
  assign n48254 = ( x186 & ~n3385 ) | ( x186 & n41072 ) | ( ~n3385 & n41072 ) ;
  assign n48255 = n14971 | n34070 ;
  assign n48256 = n48255 ^ n4756 ^ 1'b0 ;
  assign n48257 = ~n2914 & n19541 ;
  assign n48258 = n48257 ^ n1285 ^ 1'b0 ;
  assign n48259 = n48258 ^ n38713 ^ 1'b0 ;
  assign n48260 = ~n21608 & n48259 ;
  assign n48261 = ~n48256 & n48260 ;
  assign n48262 = n33938 | n48261 ;
  assign n48263 = n48262 ^ n15686 ^ 1'b0 ;
  assign n48264 = n25180 & ~n43698 ;
  assign n48265 = n42844 ^ n23347 ^ n6051 ;
  assign n48266 = n27547 | n36417 ;
  assign n48267 = n35511 & n48266 ;
  assign n48268 = ~n48265 & n48267 ;
  assign n48269 = n48216 ^ n29193 ^ n16413 ;
  assign n48270 = n3640 & ~n48269 ;
  assign n48271 = n33063 & ~n42512 ;
  assign n48272 = n14878 & ~n22435 ;
  assign n48273 = ~n48271 & n48272 ;
  assign n48274 = n18576 ^ n10129 ^ 1'b0 ;
  assign n48275 = n21669 & n48274 ;
  assign n48276 = ( n8623 & n36056 ) | ( n8623 & ~n48275 ) | ( n36056 & ~n48275 ) ;
  assign n48277 = n28919 ^ n12164 ^ n7435 ;
  assign n48278 = n9099 & n48277 ;
  assign n48279 = ( n15546 & n17106 ) | ( n15546 & n35796 ) | ( n17106 & n35796 ) ;
  assign n48280 = ( n8966 & ~n28283 ) | ( n8966 & n29687 ) | ( ~n28283 & n29687 ) ;
  assign n48281 = ~n19585 & n35173 ;
  assign n48282 = n46664 ^ n13362 ^ 1'b0 ;
  assign n48283 = n10436 | n48282 ;
  assign n48284 = n3770 | n40879 ;
  assign n48285 = n48284 ^ n37534 ^ 1'b0 ;
  assign n48286 = ~n26893 & n31122 ;
  assign n48287 = n48286 ^ n27279 ^ 1'b0 ;
  assign n48288 = n42471 ^ n17471 ^ 1'b0 ;
  assign n48289 = n30078 | n41980 ;
  assign n48290 = n48289 ^ n8039 ^ n6047 ;
  assign n48291 = n42769 ^ n24237 ^ n11539 ;
  assign n48292 = n28528 | n48291 ;
  assign n48293 = n27024 & n31354 ;
  assign n48294 = n5807 | n48293 ;
  assign n48295 = n32239 ^ n4744 ^ 1'b0 ;
  assign n48296 = n24437 & ~n48295 ;
  assign n48297 = n5689 ^ n4685 ^ 1'b0 ;
  assign n48298 = n14416 & n48297 ;
  assign n48299 = n13694 & n28112 ;
  assign n48300 = n10533 | n29749 ;
  assign n48301 = n26571 | n48300 ;
  assign n48302 = n18737 & n48301 ;
  assign n48303 = ~n44247 & n48302 ;
  assign n48304 = ~n19874 & n47840 ;
  assign n48305 = n48304 ^ n32079 ^ 1'b0 ;
  assign n48306 = n41866 ^ n13241 ^ 1'b0 ;
  assign n48307 = n30104 | n48306 ;
  assign n48308 = n9266 & ~n10896 ;
  assign n48311 = ( ~n6182 & n7824 ) | ( ~n6182 & n30385 ) | ( n7824 & n30385 ) ;
  assign n48309 = ( ~x111 & n7530 ) | ( ~x111 & n18004 ) | ( n7530 & n18004 ) ;
  assign n48310 = n48309 ^ x40 ^ 1'b0 ;
  assign n48312 = n48311 ^ n48310 ^ n44719 ;
  assign n48313 = n28608 ^ x90 ^ 1'b0 ;
  assign n48314 = n44326 ^ n11762 ^ 1'b0 ;
  assign n48315 = n48313 & n48314 ;
  assign n48316 = n16761 & n31278 ;
  assign n48317 = n32978 ^ n17838 ^ 1'b0 ;
  assign n48318 = n18960 ^ n4334 ^ 1'b0 ;
  assign n48319 = ~n36327 & n48318 ;
  assign n48322 = n18345 ^ n13291 ^ n3956 ;
  assign n48321 = n13045 & n34528 ;
  assign n48323 = n48322 ^ n48321 ^ 1'b0 ;
  assign n48320 = n3629 & ~n30936 ;
  assign n48324 = n48323 ^ n48320 ^ 1'b0 ;
  assign n48325 = n44654 ^ n19610 ^ 1'b0 ;
  assign n48326 = n3109 & n48325 ;
  assign n48327 = n48326 ^ n14094 ^ n1817 ;
  assign n48328 = n3970 | n6377 ;
  assign n48329 = n25252 ^ n4736 ^ 1'b0 ;
  assign n48330 = n48329 ^ n46178 ^ n1275 ;
  assign n48331 = n23735 ^ n19077 ^ n5655 ;
  assign n48332 = n48331 ^ n46712 ^ n5653 ;
  assign n48333 = ( n6165 & ~n43710 ) | ( n6165 & n48332 ) | ( ~n43710 & n48332 ) ;
  assign n48334 = ~n28975 & n35212 ;
  assign n48335 = n4266 & ~n16354 ;
  assign n48336 = n3814 & ~n16546 ;
  assign n48337 = ~n44558 & n48336 ;
  assign n48338 = n4695 & n10909 ;
  assign n48339 = n48338 ^ n32755 ^ 1'b0 ;
  assign n48340 = n41613 ^ n7403 ^ 1'b0 ;
  assign n48341 = n48339 | n48340 ;
  assign n48342 = n18656 & n24281 ;
  assign n48343 = ~n28658 & n48342 ;
  assign n48344 = ( n6901 & n11361 ) | ( n6901 & ~n20959 ) | ( n11361 & ~n20959 ) ;
  assign n48345 = ( n22299 & n23718 ) | ( n22299 & ~n48344 ) | ( n23718 & ~n48344 ) ;
  assign n48346 = n16927 ^ n6152 ^ 1'b0 ;
  assign n48347 = ~n48345 & n48346 ;
  assign n48348 = n44842 ^ n37476 ^ n23994 ;
  assign n48349 = ( n13977 & n25476 ) | ( n13977 & ~n41728 ) | ( n25476 & ~n41728 ) ;
  assign n48350 = n37807 ^ n20315 ^ n19068 ;
  assign n48351 = n38419 & n42611 ;
  assign n48352 = n952 & ~n19884 ;
  assign n48353 = n48352 ^ n12289 ^ 1'b0 ;
  assign n48354 = ~n13876 & n37920 ;
  assign n48355 = n12803 ^ n11262 ^ 1'b0 ;
  assign n48356 = n23925 & ~n48355 ;
  assign n48357 = n32865 ^ n32145 ^ 1'b0 ;
  assign n48358 = n48357 ^ n15180 ^ n2297 ;
  assign n48359 = ( n1124 & n11930 ) | ( n1124 & n34218 ) | ( n11930 & n34218 ) ;
  assign n48360 = n48359 ^ n2387 ^ 1'b0 ;
  assign n48361 = n21082 & n36018 ;
  assign n48362 = n21829 ^ n976 ^ 1'b0 ;
  assign n48363 = n18944 | n48362 ;
  assign n48364 = n48361 & ~n48363 ;
  assign n48365 = n45112 & ~n46318 ;
  assign n48366 = n28487 & n48365 ;
  assign n48367 = n32282 ^ n24403 ^ 1'b0 ;
  assign n48368 = ~n6377 & n48367 ;
  assign n48369 = ~n31802 & n45702 ;
  assign n48370 = ~n48368 & n48369 ;
  assign n48371 = n7179 & ~n8776 ;
  assign n48372 = n8685 | n29602 ;
  assign n48373 = n36630 & n48372 ;
  assign n48374 = n33813 & n48373 ;
  assign n48375 = ~n10568 & n17988 ;
  assign n48376 = ~n14539 & n22798 ;
  assign n48377 = n48376 ^ n2118 ^ 1'b0 ;
  assign n48378 = ~n15092 & n20104 ;
  assign n48379 = n48378 ^ n8507 ^ 1'b0 ;
  assign n48380 = ( n21762 & ~n34525 ) | ( n21762 & n48379 ) | ( ~n34525 & n48379 ) ;
  assign n48381 = ( n8318 & n13284 ) | ( n8318 & n14466 ) | ( n13284 & n14466 ) ;
  assign n48382 = n1928 | n48381 ;
  assign n48383 = n9049 & ~n39948 ;
  assign n48384 = ( ~n48380 & n48382 ) | ( ~n48380 & n48383 ) | ( n48382 & n48383 ) ;
  assign n48385 = ( n1312 & n6195 ) | ( n1312 & n11886 ) | ( n6195 & n11886 ) ;
  assign n48386 = n48385 ^ n28558 ^ 1'b0 ;
  assign n48387 = ~n1321 & n48386 ;
  assign n48388 = n48387 ^ n37608 ^ 1'b0 ;
  assign n48389 = ( n729 & n9115 ) | ( n729 & ~n33643 ) | ( n9115 & ~n33643 ) ;
  assign n48390 = n827 & ~n12907 ;
  assign n48391 = n48390 ^ x230 ^ 1'b0 ;
  assign n48392 = n32629 ^ n5834 ^ 1'b0 ;
  assign n48393 = ~n18109 & n48392 ;
  assign n48394 = ~n9085 & n48393 ;
  assign n48395 = n13081 ^ n5245 ^ 1'b0 ;
  assign n48396 = ~n4783 & n48395 ;
  assign n48397 = n48394 & n48396 ;
  assign n48398 = n6967 & n44686 ;
  assign n48399 = n43300 ^ n20664 ^ 1'b0 ;
  assign n48400 = ~n17832 & n48399 ;
  assign n48401 = n4645 | n37243 ;
  assign n48402 = n14591 & ~n48401 ;
  assign n48403 = n28528 | n48402 ;
  assign n48404 = n34893 ^ n12868 ^ 1'b0 ;
  assign n48405 = n17174 ^ n2216 ^ 1'b0 ;
  assign n48406 = n39095 ^ n6457 ^ n5365 ;
  assign n48407 = n10546 ^ n268 ^ 1'b0 ;
  assign n48408 = ( n5219 & n9112 ) | ( n5219 & n48407 ) | ( n9112 & n48407 ) ;
  assign n48409 = ( n2230 & n11883 ) | ( n2230 & ~n48408 ) | ( n11883 & ~n48408 ) ;
  assign n48410 = n48409 ^ n7991 ^ 1'b0 ;
  assign n48411 = n42512 | n48410 ;
  assign n48412 = ( n13279 & n36779 ) | ( n13279 & ~n48411 ) | ( n36779 & ~n48411 ) ;
  assign n48413 = n9640 & ~n27727 ;
  assign n48414 = n48413 ^ n3979 ^ 1'b0 ;
  assign n48415 = ~n2906 & n48414 ;
  assign n48416 = n44875 ^ n8364 ^ 1'b0 ;
  assign n48417 = ~n44318 & n48416 ;
  assign n48419 = n23923 ^ n12440 ^ 1'b0 ;
  assign n48420 = n14712 & n48419 ;
  assign n48418 = n2336 & ~n30777 ;
  assign n48421 = n48420 ^ n48418 ^ 1'b0 ;
  assign n48422 = n23264 ^ n11855 ^ 1'b0 ;
  assign n48423 = n41422 & ~n48422 ;
  assign n48424 = ~n13545 & n39291 ;
  assign n48425 = n2667 & ~n17230 ;
  assign n48426 = n48425 ^ n33104 ^ 1'b0 ;
  assign n48427 = n20719 | n22553 ;
  assign n48428 = ( n5662 & n14246 ) | ( n5662 & ~n44594 ) | ( n14246 & ~n44594 ) ;
  assign n48430 = n36089 ^ n12859 ^ n2782 ;
  assign n48429 = n24685 | n26402 ;
  assign n48431 = n48430 ^ n48429 ^ 1'b0 ;
  assign n48432 = ( ~n20426 & n21804 ) | ( ~n20426 & n28028 ) | ( n21804 & n28028 ) ;
  assign n48433 = ( ~n2940 & n48431 ) | ( ~n2940 & n48432 ) | ( n48431 & n48432 ) ;
  assign n48434 = n18936 ^ n5374 ^ 1'b0 ;
  assign n48435 = ( ~n13284 & n15010 ) | ( ~n13284 & n48434 ) | ( n15010 & n48434 ) ;
  assign n48436 = ~n15403 & n48435 ;
  assign n48437 = n8640 ^ n3678 ^ 1'b0 ;
  assign n48438 = n31516 & ~n48437 ;
  assign n48439 = ~n15273 & n48438 ;
  assign n48440 = n30251 | n48439 ;
  assign n48441 = n1152 & ~n18569 ;
  assign n48442 = n29859 ^ n11719 ^ 1'b0 ;
  assign n48443 = n48441 & n48442 ;
  assign n48444 = n14576 & ~n22442 ;
  assign n48445 = n6773 ^ n4079 ^ 1'b0 ;
  assign n48446 = n48445 ^ n16195 ^ 1'b0 ;
  assign n48452 = ( n14675 & n17989 ) | ( n14675 & ~n26287 ) | ( n17989 & ~n26287 ) ;
  assign n48453 = n48452 ^ n27200 ^ 1'b0 ;
  assign n48454 = ~n13100 & n48453 ;
  assign n48447 = ~n4945 & n48250 ;
  assign n48448 = n48447 ^ n30808 ^ n26129 ;
  assign n48449 = n8624 ^ n6514 ^ 1'b0 ;
  assign n48450 = n31806 & ~n48449 ;
  assign n48451 = ~n48448 & n48450 ;
  assign n48455 = n48454 ^ n48451 ^ n15145 ;
  assign n48456 = n13405 & ~n23116 ;
  assign n48457 = n48456 ^ n1012 ^ 1'b0 ;
  assign n48458 = ( n8411 & n29204 ) | ( n8411 & n48457 ) | ( n29204 & n48457 ) ;
  assign n48459 = ~n1433 & n3767 ;
  assign n48460 = n48459 ^ n31083 ^ n11719 ;
  assign n48461 = ~n25096 & n48460 ;
  assign n48462 = n25313 ^ n6756 ^ n4345 ;
  assign n48463 = n48462 ^ n17107 ^ 1'b0 ;
  assign n48464 = n44828 ^ n44548 ^ 1'b0 ;
  assign n48465 = ( n5511 & n8211 ) | ( n5511 & ~n23099 ) | ( n8211 & ~n23099 ) ;
  assign n48466 = n10503 ^ n1129 ^ 1'b0 ;
  assign n48467 = n44415 ^ n30719 ^ 1'b0 ;
  assign n48468 = n31001 ^ n28517 ^ n17581 ;
  assign n48469 = n37135 & ~n38475 ;
  assign n48470 = n12084 & ~n40773 ;
  assign n48472 = n11191 ^ n8432 ^ 1'b0 ;
  assign n48471 = n2959 & n20213 ;
  assign n48473 = n48472 ^ n48471 ^ 1'b0 ;
  assign n48474 = ( n4670 & ~n5319 ) | ( n4670 & n16484 ) | ( ~n5319 & n16484 ) ;
  assign n48475 = ( n5327 & ~n12672 ) | ( n5327 & n48474 ) | ( ~n12672 & n48474 ) ;
  assign n48476 = ( n5706 & n45006 ) | ( n5706 & ~n48475 ) | ( n45006 & ~n48475 ) ;
  assign n48477 = n12385 & n48476 ;
  assign n48478 = n16952 & ~n39340 ;
  assign n48479 = n15607 ^ n11692 ^ 1'b0 ;
  assign n48480 = n48478 | n48479 ;
  assign n48481 = n19646 ^ n17335 ^ 1'b0 ;
  assign n48482 = n22351 & n46086 ;
  assign n48483 = n23126 & ~n38791 ;
  assign n48484 = n48483 ^ n12956 ^ 1'b0 ;
  assign n48485 = ~n17655 & n48484 ;
  assign n48486 = n24483 ^ n14832 ^ n4789 ;
  assign n48488 = ( n3152 & n4974 ) | ( n3152 & ~n7125 ) | ( n4974 & ~n7125 ) ;
  assign n48487 = ~n9834 & n15121 ;
  assign n48489 = n48488 ^ n48487 ^ 1'b0 ;
  assign n48490 = n34145 ^ n9242 ^ 1'b0 ;
  assign n48491 = n46791 & n48490 ;
  assign n48492 = ~n7376 & n40206 ;
  assign n48493 = n43659 & n48492 ;
  assign n48494 = n20714 ^ n11109 ^ 1'b0 ;
  assign n48495 = n6318 & ~n11407 ;
  assign n48496 = n48495 ^ n41696 ^ 1'b0 ;
  assign n48497 = ~n5480 & n38787 ;
  assign n48498 = n48497 ^ n14257 ^ 1'b0 ;
  assign n48500 = n7646 | n20040 ;
  assign n48499 = n3744 | n10211 ;
  assign n48501 = n48500 ^ n48499 ^ 1'b0 ;
  assign n48502 = n48501 ^ x233 ^ 1'b0 ;
  assign n48503 = n26606 ^ n12301 ^ n3151 ;
  assign n48504 = n12973 & ~n20992 ;
  assign n48505 = n19674 & n34649 ;
  assign n48506 = n48505 ^ n19556 ^ n6463 ;
  assign n48507 = n5471 | n18705 ;
  assign n48508 = n4616 | n48507 ;
  assign n48509 = n12306 ^ n12272 ^ 1'b0 ;
  assign n48510 = n9887 & ~n12407 ;
  assign n48511 = n48510 ^ n18845 ^ n5062 ;
  assign n48512 = n48511 ^ n22031 ^ 1'b0 ;
  assign n48513 = n4840 & ~n48512 ;
  assign n48514 = n23131 & ~n43000 ;
  assign n48515 = ~n48513 & n48514 ;
  assign n48516 = n17498 | n43880 ;
  assign n48517 = n14942 & ~n48516 ;
  assign n48518 = ~n46560 & n48517 ;
  assign n48519 = ( n26353 & n41540 ) | ( n26353 & ~n48518 ) | ( n41540 & ~n48518 ) ;
  assign n48520 = n47547 ^ n26602 ^ n11790 ;
  assign n48521 = n24681 ^ n22819 ^ 1'b0 ;
  assign n48522 = n8192 & ~n48521 ;
  assign n48523 = ~n18755 & n48522 ;
  assign n48524 = n38563 ^ n7998 ^ 1'b0 ;
  assign n48525 = ~n2124 & n12758 ;
  assign n48526 = n48524 & n48525 ;
  assign n48527 = n8335 & n34143 ;
  assign n48528 = n48527 ^ n26258 ^ 1'b0 ;
  assign n48529 = n13070 | n48528 ;
  assign n48530 = n33235 ^ n16073 ^ n10409 ;
  assign n48531 = n15484 & n48530 ;
  assign n48532 = n48531 ^ n32972 ^ 1'b0 ;
  assign n48533 = n3660 & ~n28791 ;
  assign n48534 = n4317 | n17642 ;
  assign n48535 = n48534 ^ n6725 ^ 1'b0 ;
  assign n48536 = n2042 & n29970 ;
  assign n48537 = ( n30078 & ~n43193 ) | ( n30078 & n44844 ) | ( ~n43193 & n44844 ) ;
  assign n48541 = n30010 ^ n16121 ^ 1'b0 ;
  assign n48539 = n10093 & ~n15965 ;
  assign n48540 = n48539 ^ n24863 ^ 1'b0 ;
  assign n48538 = n5337 & n47904 ;
  assign n48542 = n48541 ^ n48540 ^ n48538 ;
  assign n48543 = ~n28307 & n46703 ;
  assign n48544 = n20702 & ~n25946 ;
  assign n48545 = n1454 & n48544 ;
  assign n48546 = n41400 ^ n40018 ^ 1'b0 ;
  assign n48547 = n1434 | n48546 ;
  assign n48548 = n36049 ^ n6982 ^ 1'b0 ;
  assign n48549 = n45447 ^ n5907 ^ 1'b0 ;
  assign n48550 = n19369 & ~n30559 ;
  assign n48551 = ( n545 & n7302 ) | ( n545 & ~n48550 ) | ( n7302 & ~n48550 ) ;
  assign n48552 = n19766 & ~n24035 ;
  assign n48553 = n48552 ^ n2050 ^ 1'b0 ;
  assign n48554 = n5874 & n24501 ;
  assign n48555 = n48554 ^ n5936 ^ 1'b0 ;
  assign n48556 = ( n4232 & n42895 ) | ( n4232 & n48555 ) | ( n42895 & n48555 ) ;
  assign n48557 = n34160 ^ n17585 ^ 1'b0 ;
  assign n48558 = n1831 & ~n27057 ;
  assign n48559 = n11886 & ~n48558 ;
  assign n48560 = n48559 ^ n8679 ^ 1'b0 ;
  assign n48561 = n5721 | n48560 ;
  assign n48562 = n20205 & ~n48561 ;
  assign n48563 = n13291 & n40871 ;
  assign n48564 = n48562 & n48563 ;
  assign n48565 = n11905 ^ n8558 ^ 1'b0 ;
  assign n48566 = n39268 | n48565 ;
  assign n48567 = n21638 | n48566 ;
  assign n48568 = ( n3680 & n5203 ) | ( n3680 & n7676 ) | ( n5203 & n7676 ) ;
  assign n48569 = n18474 ^ n850 ^ 1'b0 ;
  assign n48570 = n48569 ^ n43241 ^ n29242 ;
  assign n48571 = n48570 ^ n25529 ^ n3106 ;
  assign n48572 = n30216 ^ n6427 ^ 1'b0 ;
  assign n48573 = n2750 | n16798 ;
  assign n48575 = n945 & ~n7298 ;
  assign n48574 = ~n3685 & n37960 ;
  assign n48576 = n48575 ^ n48574 ^ 1'b0 ;
  assign n48577 = n40299 | n48576 ;
  assign n48578 = n48573 & ~n48577 ;
  assign n48579 = n46452 ^ n26518 ^ 1'b0 ;
  assign n48580 = n2202 | n3060 ;
  assign n48581 = n48580 ^ n21087 ^ 1'b0 ;
  assign n48582 = n14189 ^ n6002 ^ 1'b0 ;
  assign n48583 = n4836 | n48582 ;
  assign n48584 = n13086 ^ n9807 ^ 1'b0 ;
  assign n48585 = n9209 ^ n5105 ^ 1'b0 ;
  assign n48586 = n23245 & ~n48585 ;
  assign n48587 = n31909 ^ n11045 ^ 1'b0 ;
  assign n48588 = n48587 ^ n38577 ^ 1'b0 ;
  assign n48589 = n36779 ^ n10493 ^ n1517 ;
  assign n48590 = n19261 ^ n1938 ^ 1'b0 ;
  assign n48591 = ~n4105 & n45591 ;
  assign n48592 = n15915 & ~n29052 ;
  assign n48594 = ( n3034 & ~n13248 ) | ( n3034 & n20379 ) | ( ~n13248 & n20379 ) ;
  assign n48593 = n1935 | n22923 ;
  assign n48595 = n48594 ^ n48593 ^ 1'b0 ;
  assign n48596 = n5292 & ~n12321 ;
  assign n48597 = n6990 & n48596 ;
  assign n48598 = n9044 & ~n11033 ;
  assign n48599 = ~n45023 & n48598 ;
  assign n48600 = n48599 ^ n25629 ^ 1'b0 ;
  assign n48605 = n12136 & n38411 ;
  assign n48602 = ( n11551 & n19752 ) | ( n11551 & ~n39694 ) | ( n19752 & ~n39694 ) ;
  assign n48601 = n9872 & n12653 ;
  assign n48603 = n48602 ^ n48601 ^ 1'b0 ;
  assign n48604 = n32796 & ~n48603 ;
  assign n48606 = n48605 ^ n48604 ^ 1'b0 ;
  assign n48607 = n17690 & n28554 ;
  assign n48608 = n47293 ^ n33781 ^ 1'b0 ;
  assign n48609 = n15704 ^ n10378 ^ 1'b0 ;
  assign n48610 = n1935 ^ n1369 ^ 1'b0 ;
  assign n48611 = ~n48609 & n48610 ;
  assign n48612 = n48611 ^ n44959 ^ 1'b0 ;
  assign n48613 = n36785 ^ n1727 ^ x254 ;
  assign n48614 = ~n31716 & n45782 ;
  assign n48615 = n4261 & n7739 ;
  assign n48616 = n48615 ^ n44158 ^ n28658 ;
  assign n48617 = ~n1028 & n48616 ;
  assign n48618 = ~n1150 & n48617 ;
  assign n48619 = n48618 ^ n12938 ^ 1'b0 ;
  assign n48620 = ~n9514 & n48619 ;
  assign n48621 = x18 & ~n32098 ;
  assign n48622 = n30124 & n48621 ;
  assign n48623 = n38415 ^ n16711 ^ 1'b0 ;
  assign n48624 = n43006 | n48623 ;
  assign n48625 = n12340 | n48624 ;
  assign n48626 = ( n10053 & ~n21769 ) | ( n10053 & n28393 ) | ( ~n21769 & n28393 ) ;
  assign n48627 = n33415 ^ n24148 ^ n2080 ;
  assign n48628 = n31451 ^ n12021 ^ n6510 ;
  assign n48629 = n317 | n3700 ;
  assign n48630 = n35100 & n40368 ;
  assign n48631 = n48630 ^ n21898 ^ 1'b0 ;
  assign n48633 = ( ~n9385 & n19052 ) | ( ~n9385 & n34955 ) | ( n19052 & n34955 ) ;
  assign n48632 = ~n13607 & n25400 ;
  assign n48634 = n48633 ^ n48632 ^ 1'b0 ;
  assign n48635 = n19920 ^ n9986 ^ 1'b0 ;
  assign n48636 = n5106 | n48635 ;
  assign n48637 = ~n17901 & n34715 ;
  assign n48638 = n48637 ^ n27948 ^ 1'b0 ;
  assign n48639 = n26638 ^ n21366 ^ 1'b0 ;
  assign n48640 = n4681 & n48639 ;
  assign n48641 = ~n34816 & n48640 ;
  assign n48642 = n47839 & n48641 ;
  assign n48643 = ( n13116 & n14125 ) | ( n13116 & ~n39883 ) | ( n14125 & ~n39883 ) ;
  assign n48644 = ( n1840 & n28239 ) | ( n1840 & ~n46366 ) | ( n28239 & ~n46366 ) ;
  assign n48645 = ( n14353 & n37870 ) | ( n14353 & ~n48644 ) | ( n37870 & ~n48644 ) ;
  assign n48646 = ~n13813 & n20714 ;
  assign n48647 = n48646 ^ n12648 ^ 1'b0 ;
  assign n48648 = n36738 & ~n48647 ;
  assign n48649 = n48648 ^ n17678 ^ 1'b0 ;
  assign n48650 = n2484 | n40421 ;
  assign n48651 = n48650 ^ n9925 ^ 1'b0 ;
  assign n48652 = ~n3277 & n43211 ;
  assign n48653 = n14460 | n17575 ;
  assign n48654 = n13644 & ~n48653 ;
  assign n48655 = n11636 | n48654 ;
  assign n48656 = ~n7155 & n30053 ;
  assign n48657 = n15539 & ~n48656 ;
  assign n48658 = ~n25292 & n48657 ;
  assign n48659 = n7540 ^ n3813 ^ n2106 ;
  assign n48661 = n10757 ^ n8375 ^ 1'b0 ;
  assign n48660 = n2633 | n14095 ;
  assign n48662 = n48661 ^ n48660 ^ n44910 ;
  assign n48663 = n14372 ^ n10492 ^ 1'b0 ;
  assign n48664 = n44898 ^ n15368 ^ 1'b0 ;
  assign n48665 = n29454 | n48664 ;
  assign n48666 = n47835 ^ n40270 ^ n40016 ;
  assign n48667 = ( n48663 & ~n48665 ) | ( n48663 & n48666 ) | ( ~n48665 & n48666 ) ;
  assign n48669 = n2734 & n4724 ;
  assign n48668 = n18746 & ~n33229 ;
  assign n48670 = n48669 ^ n48668 ^ 1'b0 ;
  assign n48671 = n48670 ^ n20382 ^ n15128 ;
  assign n48672 = n15461 & ~n45391 ;
  assign n48673 = n48672 ^ n5362 ^ 1'b0 ;
  assign n48674 = n5541 | n10712 ;
  assign n48675 = n2951 ^ n1980 ^ 1'b0 ;
  assign n48676 = ~n1761 & n48675 ;
  assign n48677 = n26638 ^ n10751 ^ n2228 ;
  assign n48678 = ( n575 & n3813 ) | ( n575 & n30619 ) | ( n3813 & n30619 ) ;
  assign n48679 = n27315 & n48678 ;
  assign n48680 = ~n36524 & n47073 ;
  assign n48681 = ~n11936 & n16443 ;
  assign n48682 = n3991 & n48681 ;
  assign n48683 = n15717 ^ n8850 ^ 1'b0 ;
  assign n48684 = n46683 & ~n48683 ;
  assign n48685 = n44705 ^ n1742 ^ 1'b0 ;
  assign n48686 = n48684 & n48685 ;
  assign n48687 = n9247 & n15420 ;
  assign n48688 = n48687 ^ n22747 ^ 1'b0 ;
  assign n48689 = n953 ^ n917 ^ 1'b0 ;
  assign n48690 = n16682 & ~n48689 ;
  assign n48691 = n42293 | n48690 ;
  assign n48692 = x126 & ~n18285 ;
  assign n48693 = n48692 ^ n39199 ^ 1'b0 ;
  assign n48698 = ( ~n4542 & n12956 ) | ( ~n4542 & n32257 ) | ( n12956 & n32257 ) ;
  assign n48696 = n10581 & n10621 ;
  assign n48697 = ~n14138 & n48696 ;
  assign n48694 = n35065 & ~n48345 ;
  assign n48695 = ~n44210 & n48694 ;
  assign n48699 = n48698 ^ n48697 ^ n48695 ;
  assign n48700 = ( n1399 & ~n15949 ) | ( n1399 & n36729 ) | ( ~n15949 & n36729 ) ;
  assign n48701 = n32679 ^ n14427 ^ n4193 ;
  assign n48702 = n12975 & n38112 ;
  assign n48703 = n48702 ^ n9726 ^ 1'b0 ;
  assign n48704 = n41787 & n48703 ;
  assign n48705 = n21496 ^ n6922 ^ 1'b0 ;
  assign n48706 = ~n27225 & n48705 ;
  assign n48707 = n48706 ^ n18716 ^ 1'b0 ;
  assign n48708 = n7506 & ~n48707 ;
  assign n48709 = n22332 & ~n48708 ;
  assign n48712 = ~n8062 & n12853 ;
  assign n48713 = ~n9628 & n48712 ;
  assign n48714 = n11458 & n48713 ;
  assign n48715 = n17909 | n48714 ;
  assign n48710 = n31475 ^ n22019 ^ n15384 ;
  assign n48711 = n15074 & ~n48710 ;
  assign n48716 = n48715 ^ n48711 ^ 1'b0 ;
  assign n48717 = n9463 & ~n48618 ;
  assign n48718 = ~n37809 & n48717 ;
  assign n48719 = ~n1912 & n4495 ;
  assign n48720 = n953 & ~n17454 ;
  assign n48721 = n48720 ^ n20234 ^ 1'b0 ;
  assign n48722 = n17914 & ~n19868 ;
  assign n48723 = n48722 ^ n16930 ^ 1'b0 ;
  assign n48724 = ( ~n21487 & n21951 ) | ( ~n21487 & n22423 ) | ( n21951 & n22423 ) ;
  assign n48725 = ~n15279 & n26648 ;
  assign n48726 = n358 & n48725 ;
  assign n48727 = ( ~n11076 & n43303 ) | ( ~n11076 & n48726 ) | ( n43303 & n48726 ) ;
  assign n48728 = n29762 ^ n20278 ^ n8067 ;
  assign n48729 = n25546 | n48728 ;
  assign n48730 = n48729 ^ n46964 ^ n27829 ;
  assign n48731 = n27435 ^ n12926 ^ n3532 ;
  assign n48732 = n4236 | n29465 ;
  assign n48733 = n46810 ^ n46295 ^ 1'b0 ;
  assign n48734 = n48732 & ~n48733 ;
  assign n48735 = n37234 ^ n32497 ^ 1'b0 ;
  assign n48736 = n38263 ^ n26394 ^ 1'b0 ;
  assign n48737 = n5188 | n48736 ;
  assign n48738 = n11598 & n20963 ;
  assign n48739 = ~n47464 & n48738 ;
  assign n48740 = n15533 ^ n14281 ^ 1'b0 ;
  assign n48741 = ~n17612 & n48740 ;
  assign n48742 = n2025 & ~n4854 ;
  assign n48743 = ~n48741 & n48742 ;
  assign n48744 = n18238 & n47249 ;
  assign n48745 = ~n18476 & n30836 ;
  assign n48746 = n9714 ^ n7604 ^ 1'b0 ;
  assign n48747 = n16412 ^ n13246 ^ 1'b0 ;
  assign n48748 = ~n1142 & n48747 ;
  assign n48749 = ~n10342 & n48748 ;
  assign n48750 = n43028 ^ n29533 ^ 1'b0 ;
  assign n48751 = ~n6237 & n15610 ;
  assign n48752 = n39515 | n48751 ;
  assign n48753 = ~n12346 & n27464 ;
  assign n48754 = n20840 & n41646 ;
  assign n48755 = n20691 & n48754 ;
  assign n48756 = n21057 & ~n48755 ;
  assign n48757 = n48756 ^ n45289 ^ 1'b0 ;
  assign n48758 = n10201 & ~n33855 ;
  assign n48759 = n6219 & ~n48758 ;
  assign n48760 = n15780 | n41480 ;
  assign n48761 = n6219 & n22648 ;
  assign n48762 = ~n26256 & n48761 ;
  assign n48763 = ( ~n4592 & n48760 ) | ( ~n4592 & n48762 ) | ( n48760 & n48762 ) ;
  assign n48764 = n2064 & ~n11599 ;
  assign n48765 = n2721 & n48764 ;
  assign n48766 = x104 & n3555 ;
  assign n48767 = ( n39491 & ~n48765 ) | ( n39491 & n48766 ) | ( ~n48765 & n48766 ) ;
  assign n48769 = ( n7686 & n26446 ) | ( n7686 & ~n34477 ) | ( n26446 & ~n34477 ) ;
  assign n48770 = ~n14168 & n19297 ;
  assign n48771 = ~n48769 & n48770 ;
  assign n48772 = n5699 & ~n48771 ;
  assign n48773 = n10416 & n48772 ;
  assign n48768 = ~n2836 & n34688 ;
  assign n48774 = n48773 ^ n48768 ^ 1'b0 ;
  assign n48775 = n37919 ^ n26485 ^ 1'b0 ;
  assign n48776 = n5935 | n48775 ;
  assign n48777 = ~n3160 & n43458 ;
  assign n48778 = n31353 & n36248 ;
  assign n48779 = n48778 ^ n18276 ^ 1'b0 ;
  assign n48780 = n4068 & ~n48779 ;
  assign n48782 = ( ~n8709 & n39382 ) | ( ~n8709 & n42858 ) | ( n39382 & n42858 ) ;
  assign n48781 = ~n8584 & n38031 ;
  assign n48783 = n48782 ^ n48781 ^ n19421 ;
  assign n48784 = n12267 ^ n2699 ^ 1'b0 ;
  assign n48785 = ~n41197 & n48784 ;
  assign n48786 = n48785 ^ n43814 ^ n28717 ;
  assign n48791 = n7159 | n8030 ;
  assign n48792 = n36371 | n48791 ;
  assign n48787 = n25625 ^ n2427 ^ 1'b0 ;
  assign n48788 = n16599 & ~n21423 ;
  assign n48789 = n10564 & ~n48788 ;
  assign n48790 = n48787 & n48789 ;
  assign n48793 = n48792 ^ n48790 ^ n47629 ;
  assign n48794 = n8922 & n13545 ;
  assign n48795 = ~n7299 & n14725 ;
  assign n48796 = n48795 ^ n31193 ^ 1'b0 ;
  assign n48797 = n26669 & n48796 ;
  assign n48798 = n48794 & n48797 ;
  assign n48799 = n10419 & ~n43944 ;
  assign n48800 = n7186 & ~n24298 ;
  assign n48801 = n2705 | n8426 ;
  assign n48802 = n48801 ^ n11484 ^ n8202 ;
  assign n48803 = n47283 | n48802 ;
  assign n48804 = n48800 | n48803 ;
  assign n48805 = n7913 ^ n1326 ^ 1'b0 ;
  assign n48806 = n5840 | n48805 ;
  assign n48807 = n48806 ^ n9215 ^ 1'b0 ;
  assign n48808 = n44825 ^ n38595 ^ 1'b0 ;
  assign n48809 = ~n48807 & n48808 ;
  assign n48810 = n1265 & ~n36927 ;
  assign n48811 = n16232 | n48810 ;
  assign n48812 = n11809 & ~n48811 ;
  assign n48813 = x33 & ~n41476 ;
  assign n48814 = n48813 ^ n9815 ^ 1'b0 ;
  assign n48815 = n33211 & n42369 ;
  assign n48816 = n33891 ^ n31524 ^ n16725 ;
  assign n48817 = n37740 ^ n13452 ^ 1'b0 ;
  assign n48818 = n13605 ^ n5083 ^ 1'b0 ;
  assign n48819 = n48818 ^ n17002 ^ n478 ;
  assign n48820 = n48819 ^ n4546 ^ 1'b0 ;
  assign n48821 = n10056 ^ n6795 ^ n3831 ;
  assign n48822 = n48821 ^ n26146 ^ 1'b0 ;
  assign n48823 = n12736 & ~n17619 ;
  assign n48824 = n20056 ^ n5628 ^ 1'b0 ;
  assign n48825 = n18441 | n40304 ;
  assign n48826 = n48825 ^ n39744 ^ 1'b0 ;
  assign n48829 = n19381 ^ n12860 ^ 1'b0 ;
  assign n48827 = n27754 ^ n26127 ^ 1'b0 ;
  assign n48828 = n8269 & n48827 ;
  assign n48830 = n48829 ^ n48828 ^ n22510 ;
  assign n48831 = n8271 & n25908 ;
  assign n48832 = n48831 ^ n36218 ^ 1'b0 ;
  assign n48833 = ( n11653 & n14355 ) | ( n11653 & ~n18293 ) | ( n14355 & ~n18293 ) ;
  assign n48834 = n43903 | n48833 ;
  assign n48836 = ( n4611 & ~n9075 ) | ( n4611 & n33811 ) | ( ~n9075 & n33811 ) ;
  assign n48837 = n48836 ^ n7630 ^ n6448 ;
  assign n48835 = ~n1609 & n3991 ;
  assign n48838 = n48837 ^ n48835 ^ 1'b0 ;
  assign n48839 = n48311 ^ n42016 ^ 1'b0 ;
  assign n48840 = n29956 ^ n10748 ^ 1'b0 ;
  assign n48841 = ~n29377 & n48840 ;
  assign n48842 = n48841 ^ n33259 ^ n17504 ;
  assign n48843 = n48842 ^ n24051 ^ n729 ;
  assign n48844 = n14304 ^ n10781 ^ n5885 ;
  assign n48845 = ~n28062 & n48844 ;
  assign n48846 = ~n14906 & n20849 ;
  assign n48847 = n20548 & ~n48846 ;
  assign n48848 = ~n2106 & n48847 ;
  assign n48849 = n48848 ^ n41979 ^ n23030 ;
  assign n48850 = n36897 ^ n19380 ^ n14071 ;
  assign n48851 = n46440 ^ n5170 ^ 1'b0 ;
  assign n48852 = n14025 ^ n5429 ^ 1'b0 ;
  assign n48853 = ~n8729 & n19968 ;
  assign n48854 = n41787 ^ n24270 ^ 1'b0 ;
  assign n48855 = n48853 | n48854 ;
  assign n48856 = n19088 ^ n831 ^ 1'b0 ;
  assign n48857 = n10826 | n48856 ;
  assign n48858 = ~n5851 & n8927 ;
  assign n48859 = n15542 ^ n10195 ^ 1'b0 ;
  assign n48860 = ( n1307 & ~n7883 ) | ( n1307 & n31583 ) | ( ~n7883 & n31583 ) ;
  assign n48861 = n48860 ^ n39420 ^ n15346 ;
  assign n48862 = n5836 & n18234 ;
  assign n48863 = n48862 ^ n44542 ^ 1'b0 ;
  assign n48864 = n10261 & ~n43520 ;
  assign n48866 = n14881 ^ n4781 ^ 1'b0 ;
  assign n48867 = n48866 ^ n15763 ^ 1'b0 ;
  assign n48868 = n21050 & ~n48867 ;
  assign n48865 = ~n8940 & n16749 ;
  assign n48869 = n48868 ^ n48865 ^ 1'b0 ;
  assign n48870 = n28373 ^ n18924 ^ 1'b0 ;
  assign n48871 = n9801 | n48870 ;
  assign n48872 = ~n4600 & n21729 ;
  assign n48873 = n17177 ^ n1795 ^ 1'b0 ;
  assign n48874 = n26303 | n48873 ;
  assign n48875 = ( n2099 & n8168 ) | ( n2099 & ~n30325 ) | ( n8168 & ~n30325 ) ;
  assign n48876 = ( n8980 & n36689 ) | ( n8980 & ~n48875 ) | ( n36689 & ~n48875 ) ;
  assign n48877 = n7273 & ~n48876 ;
  assign n48878 = n21274 ^ n8454 ^ 1'b0 ;
  assign n48879 = ~n1030 & n48878 ;
  assign n48880 = n48879 ^ n5057 ^ n382 ;
  assign n48881 = ~n868 & n5745 ;
  assign n48882 = n26497 ^ n7790 ^ 1'b0 ;
  assign n48883 = ~n1061 & n48882 ;
  assign n48884 = n22969 ^ n16022 ^ 1'b0 ;
  assign n48885 = n48884 ^ n45420 ^ 1'b0 ;
  assign n48886 = n47982 ^ n14274 ^ 1'b0 ;
  assign n48887 = ( n39117 & n43443 ) | ( n39117 & n43848 ) | ( n43443 & n43848 ) ;
  assign n48888 = n30365 ^ n10971 ^ 1'b0 ;
  assign n48889 = ~n38050 & n48888 ;
  assign n48890 = n48889 ^ n48020 ^ n18729 ;
  assign n48891 = n38499 ^ n35734 ^ n16668 ;
  assign n48892 = ~n7936 & n17694 ;
  assign n48893 = n48892 ^ n8370 ^ 1'b0 ;
  assign n48894 = n9222 & ~n33060 ;
  assign n48895 = n48894 ^ n29913 ^ 1'b0 ;
  assign n48896 = ( n35466 & ~n48893 ) | ( n35466 & n48895 ) | ( ~n48893 & n48895 ) ;
  assign n48897 = n6162 & ~n36342 ;
  assign n48898 = n48897 ^ n46029 ^ 1'b0 ;
  assign n48899 = n32795 | n39806 ;
  assign n48900 = n48899 ^ n27999 ^ 1'b0 ;
  assign n48901 = n48900 ^ n2590 ^ 1'b0 ;
  assign n48902 = n19600 & n48901 ;
  assign n48903 = n16293 ^ n1975 ^ 1'b0 ;
  assign n48904 = n2915 & ~n48903 ;
  assign n48905 = n29602 ^ n8755 ^ 1'b0 ;
  assign n48906 = n2832 & ~n48905 ;
  assign n48907 = ~n48904 & n48906 ;
  assign n48908 = n516 & ~n10994 ;
  assign n48909 = n48908 ^ n33585 ^ n32729 ;
  assign n48910 = ( n1076 & n9634 ) | ( n1076 & n10165 ) | ( n9634 & n10165 ) ;
  assign n48911 = n48910 ^ n42666 ^ 1'b0 ;
  assign n48912 = n5242 & ~n48911 ;
  assign n48913 = ~n48909 & n48912 ;
  assign n48914 = n16872 | n48913 ;
  assign n48915 = n30211 & ~n36734 ;
  assign n48916 = n32024 & n48915 ;
  assign n48917 = n48916 ^ n4862 ^ n3624 ;
  assign n48918 = x223 | n48917 ;
  assign n48919 = n42553 ^ n15766 ^ 1'b0 ;
  assign n48923 = n12473 ^ n5199 ^ 1'b0 ;
  assign n48920 = ( ~n5792 & n9400 ) | ( ~n5792 & n11068 ) | ( n9400 & n11068 ) ;
  assign n48921 = n6807 & n48920 ;
  assign n48922 = ~n32004 & n48921 ;
  assign n48924 = n48923 ^ n48922 ^ n5103 ;
  assign n48925 = n28409 | n34001 ;
  assign n48926 = n27137 & ~n48925 ;
  assign n48927 = n48926 ^ x61 ^ 1'b0 ;
  assign n48928 = n25555 ^ n8639 ^ 1'b0 ;
  assign n48929 = n15774 & n48928 ;
  assign n48930 = n31094 & n48929 ;
  assign n48931 = x53 & ~n20593 ;
  assign n48932 = n29418 ^ n26379 ^ 1'b0 ;
  assign n48933 = n7110 & ~n48932 ;
  assign n48934 = n22795 & ~n31352 ;
  assign n48935 = ~n25927 & n48934 ;
  assign n48936 = n48935 ^ n46356 ^ 1'b0 ;
  assign n48937 = n48933 & ~n48936 ;
  assign n48938 = ( n3492 & n30891 ) | ( n3492 & ~n38442 ) | ( n30891 & ~n38442 ) ;
  assign n48939 = ~n654 & n15213 ;
  assign n48940 = n4690 & ~n15996 ;
  assign n48941 = n32080 & ~n48940 ;
  assign n48942 = x138 & ~n2598 ;
  assign n48943 = n48941 & n48942 ;
  assign n48944 = n31926 & ~n48943 ;
  assign n48945 = n44335 ^ n12723 ^ n5458 ;
  assign n48946 = ( ~n12648 & n18279 ) | ( ~n12648 & n24211 ) | ( n18279 & n24211 ) ;
  assign n48947 = n46510 ^ n26551 ^ 1'b0 ;
  assign n48948 = n48946 & n48947 ;
  assign n48949 = n39178 ^ n30854 ^ 1'b0 ;
  assign n48950 = n3012 | n48949 ;
  assign n48951 = n19411 ^ n16470 ^ 1'b0 ;
  assign n48952 = n15417 | n16883 ;
  assign n48953 = n29782 & ~n48952 ;
  assign n48954 = n9430 & n46759 ;
  assign n48955 = n35394 ^ n15080 ^ 1'b0 ;
  assign n48956 = n13380 ^ n8374 ^ 1'b0 ;
  assign n48957 = n9217 | n48956 ;
  assign n48958 = n48957 ^ n45478 ^ n4719 ;
  assign n48959 = n17041 & ~n36000 ;
  assign n48960 = n48959 ^ n13395 ^ 1'b0 ;
  assign n48961 = ( ~n32049 & n38450 ) | ( ~n32049 & n48960 ) | ( n38450 & n48960 ) ;
  assign n48962 = n26260 ^ n26127 ^ 1'b0 ;
  assign n48963 = n44305 & n48962 ;
  assign n48964 = ~n13140 & n48963 ;
  assign n48965 = n3763 | n24658 ;
  assign n48966 = n45917 | n48965 ;
  assign n48967 = ( ~n3568 & n4151 ) | ( ~n3568 & n4241 ) | ( n4151 & n4241 ) ;
  assign n48968 = n48967 ^ n10522 ^ 1'b0 ;
  assign n48969 = n9555 ^ n3345 ^ 1'b0 ;
  assign n48970 = n48969 ^ n29577 ^ 1'b0 ;
  assign n48971 = n48968 & ~n48970 ;
  assign n48975 = n36303 ^ n32690 ^ n26323 ;
  assign n48973 = n12759 | n22040 ;
  assign n48972 = n8927 & ~n16068 ;
  assign n48974 = n48973 ^ n48972 ^ 1'b0 ;
  assign n48976 = n48975 ^ n48974 ^ 1'b0 ;
  assign n48977 = ( n6194 & ~n8026 ) | ( n6194 & n44972 ) | ( ~n8026 & n44972 ) ;
  assign n48978 = ( n5580 & ~n9375 ) | ( n5580 & n28239 ) | ( ~n9375 & n28239 ) ;
  assign n48979 = ( ~n2517 & n5088 ) | ( ~n2517 & n17932 ) | ( n5088 & n17932 ) ;
  assign n48980 = ( n2167 & n14035 ) | ( n2167 & n46075 ) | ( n14035 & n46075 ) ;
  assign n48981 = n48980 ^ n43829 ^ 1'b0 ;
  assign n48982 = n44364 & ~n48981 ;
  assign n48984 = n966 & n11043 ;
  assign n48985 = n48984 ^ n366 ^ 1'b0 ;
  assign n48983 = ~n7902 & n8348 ;
  assign n48986 = n48985 ^ n48983 ^ 1'b0 ;
  assign n48987 = n11227 & n16005 ;
  assign n48988 = n48987 ^ n7067 ^ 1'b0 ;
  assign n48989 = ~n1879 & n14661 ;
  assign n48990 = n48989 ^ n34068 ^ 1'b0 ;
  assign n48991 = ( ~n5665 & n6713 ) | ( ~n5665 & n28602 ) | ( n6713 & n28602 ) ;
  assign n48992 = ~n4890 & n48991 ;
  assign n48993 = n48992 ^ n11746 ^ 1'b0 ;
  assign n48994 = n45610 ^ n10581 ^ 1'b0 ;
  assign n48995 = n42763 ^ n1774 ^ 1'b0 ;
  assign n48996 = n37505 ^ n15933 ^ n2868 ;
  assign n48997 = n20798 & ~n30062 ;
  assign n48998 = x120 | n37322 ;
  assign n48999 = n8633 & ~n48998 ;
  assign n49000 = ~n14281 & n16811 ;
  assign n49001 = ~n11119 & n49000 ;
  assign n49002 = n8923 ^ n955 ^ 1'b0 ;
  assign n49003 = n43565 ^ n17519 ^ n12597 ;
  assign n49004 = n10816 ^ n3100 ^ 1'b0 ;
  assign n49005 = n41752 ^ n30982 ^ n21101 ;
  assign n49006 = ( x234 & ~n10041 ) | ( x234 & n49005 ) | ( ~n10041 & n49005 ) ;
  assign n49007 = n23854 | n27975 ;
  assign n49008 = n39581 ^ n14393 ^ n4529 ;
  assign n49009 = n8008 & n12946 ;
  assign n49010 = n21784 ^ n4340 ^ n1425 ;
  assign n49011 = n49010 ^ n38065 ^ 1'b0 ;
  assign n49012 = ~n3910 & n49011 ;
  assign n49013 = n25000 ^ n6930 ^ 1'b0 ;
  assign n49014 = n775 | n49013 ;
  assign n49015 = n3222 & ~n31852 ;
  assign n49016 = n49015 ^ n16977 ^ 1'b0 ;
  assign n49017 = n12188 | n27465 ;
  assign n49018 = n12127 | n49017 ;
  assign n49019 = n49018 ^ n37233 ^ n9422 ;
  assign n49020 = n32022 ^ n28196 ^ n6242 ;
  assign n49021 = n49020 ^ n42797 ^ 1'b0 ;
  assign n49022 = n37174 ^ n16581 ^ 1'b0 ;
  assign n49023 = ( n2505 & n5604 ) | ( n2505 & ~n12455 ) | ( n5604 & ~n12455 ) ;
  assign n49024 = n49023 ^ n24568 ^ n16063 ;
  assign n49025 = ( n6924 & ~n10296 ) | ( n6924 & n49024 ) | ( ~n10296 & n49024 ) ;
  assign n49026 = ( n8973 & n10533 ) | ( n8973 & n47017 ) | ( n10533 & n47017 ) ;
  assign n49027 = ~n33867 & n49026 ;
  assign n49028 = n49027 ^ n904 ^ 1'b0 ;
  assign n49029 = n2452 & ~n46514 ;
  assign n49030 = n49029 ^ n25996 ^ 1'b0 ;
  assign n49031 = ( n1403 & ~n4775 ) | ( n1403 & n11903 ) | ( ~n4775 & n11903 ) ;
  assign n49032 = n8885 & n49031 ;
  assign n49033 = n10917 & ~n45439 ;
  assign n49034 = x13 & ~n18430 ;
  assign n49035 = ( n3962 & n12973 ) | ( n3962 & n13875 ) | ( n12973 & n13875 ) ;
  assign n49036 = n7210 & n49035 ;
  assign n49037 = ~n49034 & n49036 ;
  assign n49038 = ( n3255 & n4654 ) | ( n3255 & ~n49037 ) | ( n4654 & ~n49037 ) ;
  assign n49039 = n16696 | n38840 ;
  assign n49040 = n49039 ^ n22910 ^ n19369 ;
  assign n49041 = n39504 ^ n27394 ^ n14742 ;
  assign n49043 = n22572 ^ n4715 ^ 1'b0 ;
  assign n49042 = n702 & ~n2348 ;
  assign n49044 = n49043 ^ n49042 ^ n41517 ;
  assign n49045 = n26349 ^ n8853 ^ 1'b0 ;
  assign n49046 = n5612 & n23765 ;
  assign n49047 = n49046 ^ n16845 ^ 1'b0 ;
  assign n49048 = n33875 ^ n9566 ^ 1'b0 ;
  assign n49049 = n13398 ^ n6251 ^ n6027 ;
  assign n49050 = ~n18224 & n49049 ;
  assign n49051 = n12546 & n49050 ;
  assign n49052 = n10089 & n49051 ;
  assign n49053 = ~n1750 & n5838 ;
  assign n49054 = n49053 ^ n7794 ^ 1'b0 ;
  assign n49055 = n14787 | n22342 ;
  assign n49056 = n49055 ^ n19540 ^ 1'b0 ;
  assign n49057 = n49054 | n49056 ;
  assign n49059 = ~n22203 & n46864 ;
  assign n49060 = n264 & n49059 ;
  assign n49058 = n18590 & ~n41656 ;
  assign n49061 = n49060 ^ n49058 ^ 1'b0 ;
  assign n49062 = ( n7632 & ~n28317 ) | ( n7632 & n29968 ) | ( ~n28317 & n29968 ) ;
  assign n49063 = n4869 & n49062 ;
  assign n49064 = n14482 ^ n5071 ^ 1'b0 ;
  assign n49065 = n17277 & ~n42055 ;
  assign n49066 = n22886 ^ n3020 ^ 1'b0 ;
  assign n49067 = n22593 ^ n6832 ^ 1'b0 ;
  assign n49068 = ( n13102 & ~n13377 ) | ( n13102 & n49067 ) | ( ~n13377 & n49067 ) ;
  assign n49069 = n32978 ^ n22345 ^ 1'b0 ;
  assign n49070 = n49068 & n49069 ;
  assign n49071 = n36545 | n38867 ;
  assign n49072 = n49071 ^ n29832 ^ 1'b0 ;
  assign n49073 = n37515 ^ n8553 ^ n663 ;
  assign n49074 = n4958 | n49073 ;
  assign n49075 = n19947 | n22699 ;
  assign n49076 = n25451 & ~n49075 ;
  assign n49077 = n5850 ^ n4498 ^ 1'b0 ;
  assign n49078 = ( n8466 & n16864 ) | ( n8466 & n24855 ) | ( n16864 & n24855 ) ;
  assign n49079 = ( n7447 & n49077 ) | ( n7447 & n49078 ) | ( n49077 & n49078 ) ;
  assign n49080 = ( n38129 & n49076 ) | ( n38129 & ~n49079 ) | ( n49076 & ~n49079 ) ;
  assign n49081 = n37379 ^ n28521 ^ n13231 ;
  assign n49082 = ~n9563 & n15756 ;
  assign n49083 = n49082 ^ n35272 ^ 1'b0 ;
  assign n49087 = ( n5567 & ~n9653 ) | ( n5567 & n17219 ) | ( ~n9653 & n17219 ) ;
  assign n49088 = n49087 ^ n18908 ^ n7528 ;
  assign n49084 = n12614 ^ n11058 ^ 1'b0 ;
  assign n49085 = n42355 & n49084 ;
  assign n49086 = ~n23395 & n49085 ;
  assign n49089 = n49088 ^ n49086 ^ n1412 ;
  assign n49090 = n40357 ^ n13356 ^ 1'b0 ;
  assign n49091 = n13134 & n49090 ;
  assign n49092 = n21651 | n30771 ;
  assign n49093 = n36303 | n49092 ;
  assign n49094 = ~n12980 & n49093 ;
  assign n49095 = n994 & ~n19921 ;
  assign n49096 = ~n43523 & n49095 ;
  assign n49097 = n25316 ^ n10767 ^ 1'b0 ;
  assign n49098 = n9712 & n49097 ;
  assign n49100 = n14248 ^ n5797 ^ 1'b0 ;
  assign n49101 = n26357 & ~n49100 ;
  assign n49102 = n21788 & n49101 ;
  assign n49103 = n49102 ^ n7865 ^ 1'b0 ;
  assign n49099 = n16064 & ~n36386 ;
  assign n49104 = n49103 ^ n49099 ^ 1'b0 ;
  assign n49105 = n31789 ^ n4695 ^ n2838 ;
  assign n49107 = ( ~n10081 & n20596 ) | ( ~n10081 & n27264 ) | ( n20596 & n27264 ) ;
  assign n49106 = n6048 | n36393 ;
  assign n49108 = n49107 ^ n49106 ^ 1'b0 ;
  assign n49109 = n49108 ^ n15195 ^ n11470 ;
  assign n49112 = ~n19876 & n26495 ;
  assign n49110 = ( n7354 & ~n17892 ) | ( n7354 & n29590 ) | ( ~n17892 & n29590 ) ;
  assign n49111 = ~n1593 & n49110 ;
  assign n49113 = n49112 ^ n49111 ^ n27476 ;
  assign n49114 = n20512 & n40368 ;
  assign n49115 = n49114 ^ n30903 ^ 1'b0 ;
  assign n49116 = n2155 & n49115 ;
  assign n49117 = n1998 | n36393 ;
  assign n49118 = n49117 ^ n10826 ^ 1'b0 ;
  assign n49119 = n19006 ^ n702 ^ 1'b0 ;
  assign n49120 = n1152 | n44721 ;
  assign n49121 = n13151 & n21374 ;
  assign n49122 = n7110 & n26099 ;
  assign n49123 = n49122 ^ n32679 ^ 1'b0 ;
  assign n49124 = n49123 ^ n47211 ^ n1187 ;
  assign n49125 = n36925 ^ n29896 ^ n3746 ;
  assign n49126 = ~n21941 & n30122 ;
  assign n49127 = ( ~n26903 & n31103 ) | ( ~n26903 & n49126 ) | ( n31103 & n49126 ) ;
  assign n49128 = n23255 ^ n15539 ^ 1'b0 ;
  assign n49129 = n20471 & ~n49128 ;
  assign n49130 = ( ~n6841 & n44534 ) | ( ~n6841 & n48269 ) | ( n44534 & n48269 ) ;
  assign n49131 = n40881 & n49130 ;
  assign n49132 = n49131 ^ n31221 ^ 1'b0 ;
  assign n49133 = n16350 & ~n19868 ;
  assign n49134 = n7692 | n49133 ;
  assign n49135 = n37701 & ~n49134 ;
  assign n49136 = n31199 ^ n18443 ^ 1'b0 ;
  assign n49137 = n34442 ^ n19946 ^ 1'b0 ;
  assign n49138 = n49136 & ~n49137 ;
  assign n49139 = n5069 & n18533 ;
  assign n49141 = n19844 ^ n13857 ^ 1'b0 ;
  assign n49140 = n1727 ^ x46 ^ 1'b0 ;
  assign n49142 = n49141 ^ n49140 ^ n48648 ;
  assign n49143 = n39578 ^ n24241 ^ n10842 ;
  assign n49144 = n36474 ^ n682 ^ 1'b0 ;
  assign n49145 = n30494 ^ n21413 ^ 1'b0 ;
  assign n49146 = n30547 & n49145 ;
  assign n49147 = n11037 & ~n34545 ;
  assign n49148 = n19440 ^ n13209 ^ 1'b0 ;
  assign n49149 = n16665 & ~n49148 ;
  assign n49150 = n47965 ^ n11032 ^ 1'b0 ;
  assign n49151 = ( n10151 & n16965 ) | ( n10151 & ~n49150 ) | ( n16965 & ~n49150 ) ;
  assign n49152 = n6395 | n16939 ;
  assign n49153 = n49151 & ~n49152 ;
  assign n49154 = n49153 ^ n37444 ^ n2657 ;
  assign n49155 = n49154 ^ n2118 ^ 1'b0 ;
  assign n49156 = n17778 ^ n6403 ^ 1'b0 ;
  assign n49157 = ( n18649 & n34310 ) | ( n18649 & ~n49156 ) | ( n34310 & ~n49156 ) ;
  assign n49158 = n49157 ^ n2794 ^ 1'b0 ;
  assign n49159 = n23968 & ~n49158 ;
  assign n49160 = ( n26321 & n30751 ) | ( n26321 & n34907 ) | ( n30751 & n34907 ) ;
  assign n49161 = n9530 | n32741 ;
  assign n49162 = ( n37931 & n49076 ) | ( n37931 & ~n49161 ) | ( n49076 & ~n49161 ) ;
  assign n49163 = n12733 & ~n14037 ;
  assign n49164 = n11703 | n11884 ;
  assign n49165 = n32176 & ~n49164 ;
  assign n49166 = n22221 | n49165 ;
  assign n49167 = n49163 | n49166 ;
  assign n49168 = ~n2695 & n4078 ;
  assign n49169 = ~n49167 & n49168 ;
  assign n49170 = n19132 ^ n7196 ^ 1'b0 ;
  assign n49171 = n42030 & ~n49170 ;
  assign n49172 = n23417 ^ n18827 ^ 1'b0 ;
  assign n49173 = n27366 & ~n40571 ;
  assign n49174 = ~n10720 & n23325 ;
  assign n49175 = ~n19342 & n49174 ;
  assign n49176 = n8186 & ~n49175 ;
  assign n49177 = n15921 ^ n14502 ^ 1'b0 ;
  assign n49178 = ( n7066 & ~n8112 ) | ( n7066 & n39709 ) | ( ~n8112 & n39709 ) ;
  assign n49179 = n47172 ^ n19490 ^ n11767 ;
  assign n49180 = ~n15127 & n16761 ;
  assign n49181 = n49180 ^ n14943 ^ 1'b0 ;
  assign n49182 = n809 & ~n48182 ;
  assign n49183 = n4269 & ~n7334 ;
  assign n49184 = ~n46787 & n49183 ;
  assign n49185 = n38211 ^ n28580 ^ 1'b0 ;
  assign n49186 = n35801 & ~n49185 ;
  assign n49188 = n25770 ^ n18910 ^ 1'b0 ;
  assign n49189 = ~n34270 & n49188 ;
  assign n49187 = n16350 | n21999 ;
  assign n49190 = n49189 ^ n49187 ^ 1'b0 ;
  assign n49191 = n37600 ^ n906 ^ 1'b0 ;
  assign n49192 = n20170 & ~n30824 ;
  assign n49193 = n43941 ^ n17112 ^ n8689 ;
  assign n49194 = n49193 ^ n31239 ^ 1'b0 ;
  assign n49195 = n46122 ^ n15931 ^ 1'b0 ;
  assign n49196 = n7983 & ~n49195 ;
  assign n49197 = n49196 ^ n22182 ^ n1004 ;
  assign n49198 = n20669 ^ n17411 ^ n10711 ;
  assign n49199 = n49198 ^ n49112 ^ n32263 ;
  assign n49200 = n12735 & ~n49199 ;
  assign n49201 = n49200 ^ n13798 ^ 1'b0 ;
  assign n49202 = n30832 ^ n15665 ^ n8015 ;
  assign n49203 = n49202 ^ n39197 ^ 1'b0 ;
  assign n49204 = n9894 & n36983 ;
  assign n49205 = ~n26781 & n49204 ;
  assign n49206 = n5402 & n49205 ;
  assign n49207 = ~n28053 & n48517 ;
  assign n49208 = n12162 | n49207 ;
  assign n49209 = n49208 ^ n2607 ^ 1'b0 ;
  assign n49210 = n29020 ^ n13992 ^ 1'b0 ;
  assign n49211 = n42216 & n49210 ;
  assign n49212 = n38904 ^ n280 ^ 1'b0 ;
  assign n49213 = n22121 ^ n1918 ^ 1'b0 ;
  assign n49214 = n18877 ^ x159 ^ 1'b0 ;
  assign n49215 = n3628 & n49214 ;
  assign n49220 = n22451 ^ n17828 ^ 1'b0 ;
  assign n49221 = n7804 & n49220 ;
  assign n49219 = ( n21520 & n23708 ) | ( n21520 & n34364 ) | ( n23708 & n34364 ) ;
  assign n49216 = ( n1847 & n3866 ) | ( n1847 & n19519 ) | ( n3866 & n19519 ) ;
  assign n49217 = n8305 | n32730 ;
  assign n49218 = n49216 & ~n49217 ;
  assign n49222 = n49221 ^ n49219 ^ n49218 ;
  assign n49223 = n49023 ^ n8182 ^ n7157 ;
  assign n49224 = n41050 ^ n37122 ^ 1'b0 ;
  assign n49225 = n32075 ^ n4823 ^ 1'b0 ;
  assign n49226 = n308 & n35933 ;
  assign n49227 = n49226 ^ n14765 ^ 1'b0 ;
  assign n49228 = n49227 ^ n33279 ^ n14962 ;
  assign n49229 = n4350 & ~n8310 ;
  assign n49230 = ( ~n26755 & n49228 ) | ( ~n26755 & n49229 ) | ( n49228 & n49229 ) ;
  assign n49231 = ~n15024 & n49230 ;
  assign n49232 = n956 | n29919 ;
  assign n49233 = n5624 & ~n49232 ;
  assign n49234 = n44043 ^ n20650 ^ 1'b0 ;
  assign n49235 = ( n10054 & ~n20556 ) | ( n10054 & n32769 ) | ( ~n20556 & n32769 ) ;
  assign n49239 = ~n16099 & n23764 ;
  assign n49240 = n49239 ^ n18325 ^ 1'b0 ;
  assign n49236 = n25674 | n41109 ;
  assign n49237 = n49236 ^ n11707 ^ 1'b0 ;
  assign n49238 = n49237 ^ n2013 ^ 1'b0 ;
  assign n49241 = n49240 ^ n49238 ^ n36348 ;
  assign n49242 = n32254 ^ n6294 ^ n3678 ;
  assign n49243 = n46030 | n49242 ;
  assign n49244 = n10619 & n36926 ;
  assign n49245 = n28668 | n46815 ;
  assign n49246 = n11737 | n49245 ;
  assign n49247 = n40973 ^ n4296 ^ 1'b0 ;
  assign n49248 = ( n5052 & n6428 ) | ( n5052 & ~n13973 ) | ( n6428 & ~n13973 ) ;
  assign n49249 = n17325 | n49248 ;
  assign n49250 = n49249 ^ n9557 ^ n2022 ;
  assign n49251 = n13100 ^ n4528 ^ 1'b0 ;
  assign n49252 = n27884 & n49251 ;
  assign n49253 = n24088 & ~n37841 ;
  assign n49254 = ~n6330 & n44659 ;
  assign n49255 = n2465 | n45257 ;
  assign n49256 = n49255 ^ n14943 ^ 1'b0 ;
  assign n49257 = n23655 | n49256 ;
  assign n49258 = n2088 | n49257 ;
  assign n49259 = n17597 ^ n4835 ^ 1'b0 ;
  assign n49260 = n22689 & ~n49259 ;
  assign n49261 = n49260 ^ n10637 ^ 1'b0 ;
  assign n49262 = n23343 ^ n9106 ^ 1'b0 ;
  assign n49263 = n29469 | n49262 ;
  assign n49264 = n4598 & n32810 ;
  assign n49265 = n1606 & ~n23484 ;
  assign n49266 = n17594 & n49265 ;
  assign n49267 = n5604 & ~n14997 ;
  assign n49268 = n32714 ^ n6357 ^ 1'b0 ;
  assign n49269 = ~n8836 & n49268 ;
  assign n49270 = ( n2092 & n49267 ) | ( n2092 & n49269 ) | ( n49267 & n49269 ) ;
  assign n49271 = n49266 & ~n49270 ;
  assign n49272 = n25652 | n44571 ;
  assign n49273 = n13848 ^ n9523 ^ 1'b0 ;
  assign n49274 = n12513 | n39642 ;
  assign n49275 = n49274 ^ n27057 ^ 1'b0 ;
  assign n49276 = n49275 ^ n5253 ^ 1'b0 ;
  assign n49277 = ( n49272 & n49273 ) | ( n49272 & ~n49276 ) | ( n49273 & ~n49276 ) ;
  assign n49278 = n20047 ^ n4963 ^ n300 ;
  assign n49280 = n7618 ^ n2435 ^ 1'b0 ;
  assign n49281 = n16572 & n49280 ;
  assign n49279 = n28248 ^ n14157 ^ n5288 ;
  assign n49282 = n49281 ^ n49279 ^ n8201 ;
  assign n49283 = n38439 ^ n29047 ^ n1294 ;
  assign n49284 = n2236 & n49283 ;
  assign n49285 = ~n22729 & n49284 ;
  assign n49286 = n49285 ^ n44226 ^ 1'b0 ;
  assign n49287 = n2229 & ~n4398 ;
  assign n49288 = n6117 ^ n1723 ^ 1'b0 ;
  assign n49289 = ~n17340 & n49288 ;
  assign n49290 = ( n15112 & n39418 ) | ( n15112 & ~n49289 ) | ( n39418 & ~n49289 ) ;
  assign n49291 = n7240 & n9464 ;
  assign n49292 = n49290 & n49291 ;
  assign n49293 = n40953 ^ n3381 ^ 1'b0 ;
  assign n49294 = ~n49292 & n49293 ;
  assign n49295 = ~n6001 & n11401 ;
  assign n49296 = n49295 ^ n5674 ^ 1'b0 ;
  assign n49297 = n49296 ^ n16149 ^ 1'b0 ;
  assign n49298 = n40542 ^ n11355 ^ 1'b0 ;
  assign n49299 = n49297 | n49298 ;
  assign n49300 = n17771 ^ n3631 ^ 1'b0 ;
  assign n49301 = ~n5009 & n11550 ;
  assign n49302 = n49300 & n49301 ;
  assign n49303 = n43200 ^ n25937 ^ 1'b0 ;
  assign n49304 = ~n5653 & n49303 ;
  assign n49305 = n16673 & n49304 ;
  assign n49306 = n49305 ^ n1969 ^ 1'b0 ;
  assign n49307 = n46952 & n49306 ;
  assign n49308 = n20335 ^ n6294 ^ 1'b0 ;
  assign n49309 = n49307 & n49308 ;
  assign n49310 = n39923 ^ n14183 ^ 1'b0 ;
  assign n49311 = n49309 & n49310 ;
  assign n49312 = ( x130 & n12922 ) | ( x130 & ~n24719 ) | ( n12922 & ~n24719 ) ;
  assign n49313 = ~n11152 & n21371 ;
  assign n49314 = n49313 ^ n7016 ^ 1'b0 ;
  assign n49315 = n49314 ^ n33289 ^ 1'b0 ;
  assign n49316 = ~n36659 & n49315 ;
  assign n49318 = n32934 ^ n18295 ^ 1'b0 ;
  assign n49317 = n9518 & n13342 ;
  assign n49319 = n49318 ^ n49317 ^ 1'b0 ;
  assign n49320 = n31258 & n49319 ;
  assign n49321 = n44463 ^ n36309 ^ n16403 ;
  assign n49322 = n10936 & ~n49321 ;
  assign n49323 = ~n12450 & n49322 ;
  assign n49324 = n35804 ^ n14397 ^ 1'b0 ;
  assign n49325 = n25875 | n49324 ;
  assign n49326 = n1881 | n2035 ;
  assign n49327 = ~n25633 & n46770 ;
  assign n49328 = ( n4780 & n25403 ) | ( n4780 & ~n49327 ) | ( n25403 & ~n49327 ) ;
  assign n49329 = n11957 & n49328 ;
  assign n49330 = ~n49326 & n49329 ;
  assign n49332 = n4121 & n19124 ;
  assign n49333 = n49332 ^ n21486 ^ 1'b0 ;
  assign n49331 = n2406 | n2790 ;
  assign n49334 = n49333 ^ n49331 ^ 1'b0 ;
  assign n49335 = ~n24860 & n45106 ;
  assign n49336 = n7442 & ~n49335 ;
  assign n49337 = n1806 | n5747 ;
  assign n49338 = n12212 & ~n49337 ;
  assign n49339 = ~n1227 & n24622 ;
  assign n49340 = n30743 ^ n23663 ^ n20751 ;
  assign n49341 = ( n1048 & n49339 ) | ( n1048 & n49340 ) | ( n49339 & n49340 ) ;
  assign n49342 = ~n49338 & n49341 ;
  assign n49343 = n49342 ^ n40555 ^ n24769 ;
  assign n49344 = n34662 ^ n26773 ^ n3604 ;
  assign n49345 = n31946 | n49344 ;
  assign n49346 = n49345 ^ n27585 ^ 1'b0 ;
  assign n49347 = n24986 ^ n15196 ^ 1'b0 ;
  assign n49348 = ~n12754 & n16689 ;
  assign n49349 = n48690 & n49348 ;
  assign n49350 = n45199 ^ n951 ^ 1'b0 ;
  assign n49351 = ~n34856 & n49350 ;
  assign n49352 = n26915 ^ n26348 ^ 1'b0 ;
  assign n49353 = n49352 ^ n40697 ^ n24817 ;
  assign n49354 = n49353 ^ n12852 ^ 1'b0 ;
  assign n49355 = n8838 | n49354 ;
  assign n49356 = n33811 ^ n33772 ^ 1'b0 ;
  assign n49357 = n29521 & n49356 ;
  assign n49358 = n8924 | n12883 ;
  assign n49359 = n49358 ^ x24 ^ 1'b0 ;
  assign n49360 = n4209 & n9869 ;
  assign n49361 = n49360 ^ n22152 ^ 1'b0 ;
  assign n49362 = n3658 | n7580 ;
  assign n49363 = n49362 ^ n18980 ^ 1'b0 ;
  assign n49364 = ~n8052 & n12418 ;
  assign n49365 = n17286 & ~n27411 ;
  assign n49366 = n13990 ^ n6528 ^ 1'b0 ;
  assign n49367 = n1869 & n49366 ;
  assign n49368 = n26595 ^ n17562 ^ 1'b0 ;
  assign n49369 = n19248 & ~n49368 ;
  assign n49370 = n2070 | n46309 ;
  assign n49371 = n49370 ^ n7850 ^ 1'b0 ;
  assign n49372 = n21421 | n49371 ;
  assign n49373 = n49372 ^ n11902 ^ 1'b0 ;
  assign n49374 = n9012 | n25640 ;
  assign n49375 = n49373 | n49374 ;
  assign n49376 = n30330 & n45055 ;
  assign n49377 = n18194 ^ n11379 ^ 1'b0 ;
  assign n49378 = n13423 & ~n24083 ;
  assign n49379 = n9391 & n49378 ;
  assign n49380 = ( n4111 & n6183 ) | ( n4111 & ~n11485 ) | ( n6183 & ~n11485 ) ;
  assign n49381 = n22546 | n25922 ;
  assign n49382 = n49380 | n49381 ;
  assign n49383 = n26403 ^ n9820 ^ 1'b0 ;
  assign n49384 = n42055 & ~n46744 ;
  assign n49385 = n10102 ^ n5881 ^ 1'b0 ;
  assign n49386 = n27965 ^ x21 ^ 1'b0 ;
  assign n49387 = n13708 ^ x164 ^ 1'b0 ;
  assign n49388 = ~n6020 & n49387 ;
  assign n49389 = ( n7578 & n15125 ) | ( n7578 & ~n49388 ) | ( n15125 & ~n49388 ) ;
  assign n49390 = n49389 ^ n45781 ^ 1'b0 ;
  assign n49391 = n2147 & ~n49390 ;
  assign n49393 = n18236 & ~n47851 ;
  assign n49394 = n49393 ^ n11322 ^ 1'b0 ;
  assign n49395 = n49394 ^ n11712 ^ 1'b0 ;
  assign n49396 = ~n489 & n49395 ;
  assign n49392 = n15213 & ~n16206 ;
  assign n49397 = n49396 ^ n49392 ^ 1'b0 ;
  assign n49398 = n27062 ^ n4449 ^ 1'b0 ;
  assign n49399 = n46211 ^ n14986 ^ 1'b0 ;
  assign n49400 = n43789 | n49399 ;
  assign n49401 = n10121 ^ n3475 ^ n2028 ;
  assign n49402 = n18303 ^ n2278 ^ n1067 ;
  assign n49403 = n49402 ^ n31782 ^ 1'b0 ;
  assign n49404 = ( ~n2575 & n49401 ) | ( ~n2575 & n49403 ) | ( n49401 & n49403 ) ;
  assign n49405 = ( ~n5694 & n15590 ) | ( ~n5694 & n49404 ) | ( n15590 & n49404 ) ;
  assign n49407 = ( n1727 & ~n15719 ) | ( n1727 & n44574 ) | ( ~n15719 & n44574 ) ;
  assign n49408 = ~n29983 & n49407 ;
  assign n49409 = ~n8368 & n49408 ;
  assign n49406 = n4158 | n34575 ;
  assign n49410 = n49409 ^ n49406 ^ 1'b0 ;
  assign n49411 = n5963 ^ n771 ^ 1'b0 ;
  assign n49412 = n49410 | n49411 ;
  assign n49413 = n49412 ^ n2106 ^ 1'b0 ;
  assign n49414 = ( n623 & n13880 ) | ( n623 & ~n20330 ) | ( n13880 & ~n20330 ) ;
  assign n49415 = n36138 | n49414 ;
  assign n49416 = ~n24319 & n49415 ;
  assign n49417 = n11798 & ~n42810 ;
  assign n49418 = n47371 ^ n27850 ^ 1'b0 ;
  assign n49419 = n10299 ^ n2849 ^ 1'b0 ;
  assign n49420 = n24078 | n49419 ;
  assign n49421 = n41822 ^ n30629 ^ 1'b0 ;
  assign n49422 = n49420 | n49421 ;
  assign n49424 = n347 | n12202 ;
  assign n49425 = n49424 ^ n19364 ^ 1'b0 ;
  assign n49423 = n8179 & n8214 ;
  assign n49426 = n49425 ^ n49423 ^ n684 ;
  assign n49427 = n49426 ^ n32442 ^ 1'b0 ;
  assign n49428 = n2714 & n37994 ;
  assign n49429 = ~n4226 & n49428 ;
  assign n49430 = ( n12471 & ~n17519 ) | ( n12471 & n18305 ) | ( ~n17519 & n18305 ) ;
  assign n49431 = ( ~n5519 & n23577 ) | ( ~n5519 & n49430 ) | ( n23577 & n49430 ) ;
  assign n49432 = n16779 ^ n3934 ^ n2039 ;
  assign n49433 = n27214 | n42604 ;
  assign n49434 = n41334 ^ n1695 ^ 1'b0 ;
  assign n49435 = n10791 & ~n49434 ;
  assign n49436 = ( ~n4719 & n7404 ) | ( ~n4719 & n44241 ) | ( n7404 & n44241 ) ;
  assign n49437 = ~n1123 & n49436 ;
  assign n49438 = n49437 ^ n3312 ^ 1'b0 ;
  assign n49439 = n18347 & ~n43704 ;
  assign n49440 = n49430 & n49439 ;
  assign n49441 = n32249 & ~n45173 ;
  assign n49442 = ~n17843 & n49441 ;
  assign n49443 = n13319 & ~n34295 ;
  assign n49444 = n8483 & n49443 ;
  assign n49445 = n4367 & n33045 ;
  assign n49446 = n49445 ^ n33640 ^ 1'b0 ;
  assign n49447 = n4650 | n14947 ;
  assign n49448 = n49447 ^ n36015 ^ n31240 ;
  assign n49449 = n11279 | n21641 ;
  assign n49450 = n49449 ^ n42548 ^ 1'b0 ;
  assign n49451 = ~n17228 & n49450 ;
  assign n49452 = ~n20669 & n30315 ;
  assign n49453 = ( n15130 & n49451 ) | ( n15130 & ~n49452 ) | ( n49451 & ~n49452 ) ;
  assign n49454 = n30106 & n33555 ;
  assign n49455 = n49454 ^ n17018 ^ 1'b0 ;
  assign n49456 = n49455 ^ n2306 ^ 1'b0 ;
  assign n49457 = ( n6652 & n6820 ) | ( n6652 & ~n39936 ) | ( n6820 & ~n39936 ) ;
  assign n49458 = ~n6522 & n13459 ;
  assign n49459 = n34345 ^ n24214 ^ 1'b0 ;
  assign n49460 = n11728 & ~n49459 ;
  assign n49461 = n49460 ^ n39829 ^ 1'b0 ;
  assign n49462 = n49458 & ~n49461 ;
  assign n49464 = n14046 ^ n10370 ^ 1'b0 ;
  assign n49463 = ~n38562 & n42651 ;
  assign n49465 = n49464 ^ n49463 ^ 1'b0 ;
  assign n49466 = n41490 ^ n27176 ^ 1'b0 ;
  assign n49467 = n19159 & ~n49466 ;
  assign n49468 = n16773 | n47257 ;
  assign n49469 = n31075 | n49468 ;
  assign n49470 = n2331 & ~n29192 ;
  assign n49471 = ~n43032 & n49470 ;
  assign n49472 = n13284 & n24419 ;
  assign n49473 = ~n45290 & n49472 ;
  assign n49475 = ( n341 & ~n30376 ) | ( n341 & n43672 ) | ( ~n30376 & n43672 ) ;
  assign n49474 = n1671 & ~n15681 ;
  assign n49476 = n49475 ^ n49474 ^ 1'b0 ;
  assign n49477 = n33009 ^ n6102 ^ 1'b0 ;
  assign n49478 = n42967 ^ n8077 ^ 1'b0 ;
  assign n49479 = n22175 & ~n49478 ;
  assign n49480 = ( ~n16662 & n49477 ) | ( ~n16662 & n49479 ) | ( n49477 & n49479 ) ;
  assign n49481 = n49314 ^ n27610 ^ n20780 ;
  assign n49482 = ~n609 & n19915 ;
  assign n49483 = n26049 ^ n24261 ^ 1'b0 ;
  assign n49484 = n5043 ^ n4670 ^ 1'b0 ;
  assign n49485 = ~n20332 & n49484 ;
  assign n49486 = n49485 ^ n31345 ^ 1'b0 ;
  assign n49487 = n13643 | n49486 ;
  assign n49488 = n25426 ^ n25048 ^ 1'b0 ;
  assign n49491 = n17271 & n31417 ;
  assign n49489 = n16532 ^ n12457 ^ 1'b0 ;
  assign n49490 = n42777 & n49489 ;
  assign n49492 = n49491 ^ n49490 ^ 1'b0 ;
  assign n49493 = n22218 ^ n16880 ^ 1'b0 ;
  assign n49494 = ( n12407 & n12923 ) | ( n12407 & ~n14779 ) | ( n12923 & ~n14779 ) ;
  assign n49495 = ~n1106 & n49494 ;
  assign n49496 = ~n3212 & n22017 ;
  assign n49497 = n49496 ^ n18783 ^ n2538 ;
  assign n49498 = n1368 & ~n20197 ;
  assign n49499 = n23376 & n49498 ;
  assign n49500 = n49499 ^ n9193 ^ 1'b0 ;
  assign n49501 = n13962 & n40896 ;
  assign n49502 = n12577 ^ n3848 ^ 1'b0 ;
  assign n49503 = n20971 | n49502 ;
  assign n49504 = n16631 & n19634 ;
  assign n49506 = ( n2637 & ~n2832 ) | ( n2637 & n18705 ) | ( ~n2832 & n18705 ) ;
  assign n49505 = n1154 & ~n16427 ;
  assign n49507 = n49506 ^ n49505 ^ 1'b0 ;
  assign n49508 = n9746 ^ n1503 ^ 1'b0 ;
  assign n49509 = n25546 & n49508 ;
  assign n49510 = n49509 ^ n27026 ^ n25494 ;
  assign n49511 = n7066 & n31394 ;
  assign n49512 = n12206 & ~n13215 ;
  assign n49513 = ( ~n26499 & n49511 ) | ( ~n26499 & n49512 ) | ( n49511 & n49512 ) ;
  assign n49514 = ~n9424 & n31556 ;
  assign n49515 = n31818 ^ n19174 ^ n1603 ;
  assign n49516 = ( n14238 & ~n14675 ) | ( n14238 & n21289 ) | ( ~n14675 & n21289 ) ;
  assign n49517 = n5895 & ~n49516 ;
  assign n49518 = n49517 ^ n3774 ^ 1'b0 ;
  assign n49519 = n41726 | n49518 ;
  assign n49520 = n49519 ^ n28401 ^ 1'b0 ;
  assign n49521 = n24899 & n33984 ;
  assign n49522 = ~n46303 & n49521 ;
  assign n49523 = ~n35596 & n43882 ;
  assign n49524 = n40547 ^ n4059 ^ 1'b0 ;
  assign n49525 = n5749 & n49524 ;
  assign n49526 = n49525 ^ n2169 ^ 1'b0 ;
  assign n49527 = n15680 & ~n49526 ;
  assign n49528 = n36961 ^ n7270 ^ 1'b0 ;
  assign n49529 = n49527 & n49528 ;
  assign y0 = x7 ;
  assign y1 = x14 ;
  assign y2 = x44 ;
  assign y3 = x47 ;
  assign y4 = x51 ;
  assign y5 = x57 ;
  assign y6 = x61 ;
  assign y7 = x67 ;
  assign y8 = x69 ;
  assign y9 = x72 ;
  assign y10 = x81 ;
  assign y11 = x85 ;
  assign y12 = x91 ;
  assign y13 = x93 ;
  assign y14 = x95 ;
  assign y15 = x99 ;
  assign y16 = x103 ;
  assign y17 = x112 ;
  assign y18 = x113 ;
  assign y19 = x114 ;
  assign y20 = x119 ;
  assign y21 = x125 ;
  assign y22 = x126 ;
  assign y23 = x128 ;
  assign y24 = x143 ;
  assign y25 = x146 ;
  assign y26 = x149 ;
  assign y27 = x151 ;
  assign y28 = x165 ;
  assign y29 = x169 ;
  assign y30 = x173 ;
  assign y31 = x174 ;
  assign y32 = x176 ;
  assign y33 = x184 ;
  assign y34 = x190 ;
  assign y35 = x197 ;
  assign y36 = x201 ;
  assign y37 = x203 ;
  assign y38 = x205 ;
  assign y39 = x207 ;
  assign y40 = x209 ;
  assign y41 = x210 ;
  assign y42 = x216 ;
  assign y43 = x217 ;
  assign y44 = x222 ;
  assign y45 = x226 ;
  assign y46 = x227 ;
  assign y47 = x229 ;
  assign y48 = x231 ;
  assign y49 = x235 ;
  assign y50 = x246 ;
  assign y51 = x248 ;
  assign y52 = x249 ;
  assign y53 = x250 ;
  assign y54 = x252 ;
  assign y55 = x253 ;
  assign y56 = ~n256 ;
  assign y57 = ~n257 ;
  assign y58 = ~n259 ;
  assign y59 = ~n260 ;
  assign y60 = ~n262 ;
  assign y61 = ~1'b0 ;
  assign y62 = ~1'b0 ;
  assign y63 = n263 ;
  assign y64 = ~n264 ;
  assign y65 = n266 ;
  assign y66 = ~n268 ;
  assign y67 = ~n270 ;
  assign y68 = n271 ;
  assign y69 = ~1'b0 ;
  assign y70 = ~n275 ;
  assign y71 = ~1'b0 ;
  assign y72 = ~1'b0 ;
  assign y73 = ~n277 ;
  assign y74 = ~1'b0 ;
  assign y75 = ~n280 ;
  assign y76 = ~n282 ;
  assign y77 = ~n284 ;
  assign y78 = ~n287 ;
  assign y79 = n290 ;
  assign y80 = n292 ;
  assign y81 = ~n293 ;
  assign y82 = n294 ;
  assign y83 = ~1'b0 ;
  assign y84 = ~1'b0 ;
  assign y85 = n295 ;
  assign y86 = n298 ;
  assign y87 = x146 ;
  assign y88 = n300 ;
  assign y89 = ~n303 ;
  assign y90 = ~1'b0 ;
  assign y91 = n308 ;
  assign y92 = ~1'b0 ;
  assign y93 = ~n310 ;
  assign y94 = ~n314 ;
  assign y95 = ~1'b0 ;
  assign y96 = ~n317 ;
  assign y97 = n318 ;
  assign y98 = ~n322 ;
  assign y99 = n327 ;
  assign y100 = ~n330 ;
  assign y101 = ~n334 ;
  assign y102 = ~1'b0 ;
  assign y103 = ~1'b0 ;
  assign y104 = ~n335 ;
  assign y105 = ~1'b0 ;
  assign y106 = n347 ;
  assign y107 = n350 ;
  assign y108 = ~n351 ;
  assign y109 = ~n354 ;
  assign y110 = ~1'b0 ;
  assign y111 = n363 ;
  assign y112 = n365 ;
  assign y113 = ~1'b0 ;
  assign y114 = ~1'b0 ;
  assign y115 = n366 ;
  assign y116 = ~n375 ;
  assign y117 = ~1'b0 ;
  assign y118 = ~1'b0 ;
  assign y119 = n385 ;
  assign y120 = ~n389 ;
  assign y121 = ~n390 ;
  assign y122 = ~1'b0 ;
  assign y123 = ~n391 ;
  assign y124 = n393 ;
  assign y125 = ~n396 ;
  assign y126 = ~n398 ;
  assign y127 = ~1'b0 ;
  assign y128 = ~1'b0 ;
  assign y129 = ~n401 ;
  assign y130 = n402 ;
  assign y131 = ~n403 ;
  assign y132 = ~1'b0 ;
  assign y133 = n407 ;
  assign y134 = n412 ;
  assign y135 = ~n413 ;
  assign y136 = n417 ;
  assign y137 = n430 ;
  assign y138 = n434 ;
  assign y139 = n442 ;
  assign y140 = ~n450 ;
  assign y141 = ~n453 ;
  assign y142 = ~1'b0 ;
  assign y143 = n454 ;
  assign y144 = ~1'b0 ;
  assign y145 = n457 ;
  assign y146 = n462 ;
  assign y147 = ~1'b0 ;
  assign y148 = ~n464 ;
  assign y149 = n475 ;
  assign y150 = n479 ;
  assign y151 = n483 ;
  assign y152 = n485 ;
  assign y153 = n500 ;
  assign y154 = ~n501 ;
  assign y155 = ~1'b0 ;
  assign y156 = ~1'b0 ;
  assign y157 = ~n503 ;
  assign y158 = n505 ;
  assign y159 = n512 ;
  assign y160 = n514 ;
  assign y161 = ~n515 ;
  assign y162 = ~1'b0 ;
  assign y163 = n516 ;
  assign y164 = ~n518 ;
  assign y165 = ~n530 ;
  assign y166 = ~n533 ;
  assign y167 = n536 ;
  assign y168 = ~n542 ;
  assign y169 = ~n549 ;
  assign y170 = ~n552 ;
  assign y171 = n556 ;
  assign y172 = ~1'b0 ;
  assign y173 = ~n559 ;
  assign y174 = ~n560 ;
  assign y175 = n567 ;
  assign y176 = n571 ;
  assign y177 = ~n572 ;
  assign y178 = ~n574 ;
  assign y179 = ~n577 ;
  assign y180 = n578 ;
  assign y181 = n582 ;
  assign y182 = ~1'b0 ;
  assign y183 = n588 ;
  assign y184 = n591 ;
  assign y185 = n595 ;
  assign y186 = ~n597 ;
  assign y187 = ~1'b0 ;
  assign y188 = n600 ;
  assign y189 = n603 ;
  assign y190 = ~n604 ;
  assign y191 = n341 ;
  assign y192 = ~n606 ;
  assign y193 = n610 ;
  assign y194 = ~1'b0 ;
  assign y195 = ~n335 ;
  assign y196 = ~n612 ;
  assign y197 = n617 ;
  assign y198 = ~n620 ;
  assign y199 = ~n629 ;
  assign y200 = ~n630 ;
  assign y201 = n635 ;
  assign y202 = ~n638 ;
  assign y203 = ~n639 ;
  assign y204 = ~n640 ;
  assign y205 = ~n649 ;
  assign y206 = ~n651 ;
  assign y207 = n652 ;
  assign y208 = n656 ;
  assign y209 = n660 ;
  assign y210 = ~n672 ;
  assign y211 = n673 ;
  assign y212 = ~1'b0 ;
  assign y213 = ~n697 ;
  assign y214 = ~1'b0 ;
  assign y215 = ~n699 ;
  assign y216 = n702 ;
  assign y217 = ~1'b0 ;
  assign y218 = ~n703 ;
  assign y219 = ~n706 ;
  assign y220 = n718 ;
  assign y221 = n723 ;
  assign y222 = ~1'b0 ;
  assign y223 = ~1'b0 ;
  assign y224 = ~1'b0 ;
  assign y225 = n727 ;
  assign y226 = n729 ;
  assign y227 = ~n736 ;
  assign y228 = n738 ;
  assign y229 = ~n740 ;
  assign y230 = n745 ;
  assign y231 = n748 ;
  assign y232 = n754 ;
  assign y233 = n764 ;
  assign y234 = n769 ;
  assign y235 = ~1'b0 ;
  assign y236 = n774 ;
  assign y237 = ~1'b0 ;
  assign y238 = ~n783 ;
  assign y239 = n790 ;
  assign y240 = n794 ;
  assign y241 = ~n797 ;
  assign y242 = ~n800 ;
  assign y243 = n803 ;
  assign y244 = ~n804 ;
  assign y245 = ~1'b0 ;
  assign y246 = n806 ;
  assign y247 = n808 ;
  assign y248 = ~n809 ;
  assign y249 = ~n811 ;
  assign y250 = ~n814 ;
  assign y251 = ~1'b0 ;
  assign y252 = ~n817 ;
  assign y253 = n823 ;
  assign y254 = ~n831 ;
  assign y255 = ~1'b0 ;
  assign y256 = ~n832 ;
  assign y257 = ~n840 ;
  assign y258 = n841 ;
  assign y259 = n845 ;
  assign y260 = ~n848 ;
  assign y261 = ~n856 ;
  assign y262 = ~1'b0 ;
  assign y263 = ~n857 ;
  assign y264 = ~1'b0 ;
  assign y265 = ~n860 ;
  assign y266 = ~n861 ;
  assign y267 = ~n863 ;
  assign y268 = ~1'b0 ;
  assign y269 = n864 ;
  assign y270 = ~1'b0 ;
  assign y271 = n873 ;
  assign y272 = n879 ;
  assign y273 = ~n884 ;
  assign y274 = ~n885 ;
  assign y275 = ~n887 ;
  assign y276 = ~1'b0 ;
  assign y277 = n890 ;
  assign y278 = n891 ;
  assign y279 = ~n894 ;
  assign y280 = ~n901 ;
  assign y281 = ~1'b0 ;
  assign y282 = ~1'b0 ;
  assign y283 = ~n902 ;
  assign y284 = ~n905 ;
  assign y285 = n909 ;
  assign y286 = ~n913 ;
  assign y287 = n914 ;
  assign y288 = ~n917 ;
  assign y289 = ~n923 ;
  assign y290 = ~1'b0 ;
  assign y291 = n927 ;
  assign y292 = ~n929 ;
  assign y293 = ~1'b0 ;
  assign y294 = n931 ;
  assign y295 = ~n944 ;
  assign y296 = ~1'b0 ;
  assign y297 = ~1'b0 ;
  assign y298 = n945 ;
  assign y299 = ~n956 ;
  assign y300 = ~n957 ;
  assign y301 = ~1'b0 ;
  assign y302 = ~n958 ;
  assign y303 = ~n962 ;
  assign y304 = ~n970 ;
  assign y305 = ~n976 ;
  assign y306 = n979 ;
  assign y307 = ~n980 ;
  assign y308 = ~1'b0 ;
  assign y309 = n982 ;
  assign y310 = ~1'b0 ;
  assign y311 = n983 ;
  assign y312 = n990 ;
  assign y313 = n991 ;
  assign y314 = n993 ;
  assign y315 = n1006 ;
  assign y316 = ~n1010 ;
  assign y317 = n1015 ;
  assign y318 = n1018 ;
  assign y319 = ~n1019 ;
  assign y320 = ~n1026 ;
  assign y321 = ~n1028 ;
  assign y322 = n1031 ;
  assign y323 = ~n1035 ;
  assign y324 = ~1'b0 ;
  assign y325 = ~n1037 ;
  assign y326 = ~n1038 ;
  assign y327 = ~n1039 ;
  assign y328 = ~1'b0 ;
  assign y329 = ~n1047 ;
  assign y330 = n1050 ;
  assign y331 = ~n1051 ;
  assign y332 = n1054 ;
  assign y333 = n1055 ;
  assign y334 = ~1'b0 ;
  assign y335 = n1057 ;
  assign y336 = n1061 ;
  assign y337 = ~n1071 ;
  assign y338 = n1073 ;
  assign y339 = n1074 ;
  assign y340 = x73 ;
  assign y341 = ~1'b0 ;
  assign y342 = ~n1076 ;
  assign y343 = n1077 ;
  assign y344 = ~n1084 ;
  assign y345 = ~n1096 ;
  assign y346 = n1098 ;
  assign y347 = ~n1100 ;
  assign y348 = n1104 ;
  assign y349 = ~1'b0 ;
  assign y350 = n1110 ;
  assign y351 = n1111 ;
  assign y352 = n1116 ;
  assign y353 = ~n1118 ;
  assign y354 = ~n1123 ;
  assign y355 = ~n1144 ;
  assign y356 = ~n1145 ;
  assign y357 = ~1'b0 ;
  assign y358 = ~n1150 ;
  assign y359 = n1152 ;
  assign y360 = ~1'b0 ;
  assign y361 = n1154 ;
  assign y362 = n1162 ;
  assign y363 = ~n1170 ;
  assign y364 = ~n1176 ;
  assign y365 = ~1'b0 ;
  assign y366 = n1185 ;
  assign y367 = ~1'b0 ;
  assign y368 = n1190 ;
  assign y369 = n1194 ;
  assign y370 = ~1'b0 ;
  assign y371 = n1196 ;
  assign y372 = n402 ;
  assign y373 = n1200 ;
  assign y374 = n1201 ;
  assign y375 = ~n1205 ;
  assign y376 = ~n1211 ;
  assign y377 = n1217 ;
  assign y378 = ~1'b0 ;
  assign y379 = ~n1219 ;
  assign y380 = n1224 ;
  assign y381 = n1225 ;
  assign y382 = n1232 ;
  assign y383 = ~n1236 ;
  assign y384 = n1239 ;
  assign y385 = ~n1240 ;
  assign y386 = ~n1244 ;
  assign y387 = n1246 ;
  assign y388 = ~n1248 ;
  assign y389 = ~n1250 ;
  assign y390 = n1260 ;
  assign y391 = n1265 ;
  assign y392 = ~n1267 ;
  assign y393 = n1270 ;
  assign y394 = ~n1286 ;
  assign y395 = n1291 ;
  assign y396 = ~1'b0 ;
  assign y397 = n1292 ;
  assign y398 = ~n1298 ;
  assign y399 = n1300 ;
  assign y400 = n1301 ;
  assign y401 = ~n1307 ;
  assign y402 = n1308 ;
  assign y403 = ~1'b0 ;
  assign y404 = n1318 ;
  assign y405 = ~n1321 ;
  assign y406 = n1326 ;
  assign y407 = n1327 ;
  assign y408 = ~1'b0 ;
  assign y409 = n1329 ;
  assign y410 = ~n1332 ;
  assign y411 = ~n1335 ;
  assign y412 = ~n1337 ;
  assign y413 = n1343 ;
  assign y414 = ~1'b0 ;
  assign y415 = ~n1345 ;
  assign y416 = ~1'b0 ;
  assign y417 = ~n1347 ;
  assign y418 = ~1'b0 ;
  assign y419 = ~1'b0 ;
  assign y420 = ~1'b0 ;
  assign y421 = n1349 ;
  assign y422 = ~n1350 ;
  assign y423 = ~1'b0 ;
  assign y424 = ~n1357 ;
  assign y425 = ~n1360 ;
  assign y426 = n1363 ;
  assign y427 = ~1'b0 ;
  assign y428 = ~n1364 ;
  assign y429 = ~n1372 ;
  assign y430 = ~n1377 ;
  assign y431 = ~n1378 ;
  assign y432 = ~n1385 ;
  assign y433 = ~n1386 ;
  assign y434 = ~1'b0 ;
  assign y435 = n1387 ;
  assign y436 = n1394 ;
  assign y437 = ~1'b0 ;
  assign y438 = ~n1401 ;
  assign y439 = n1402 ;
  assign y440 = n1403 ;
  assign y441 = n1409 ;
  assign y442 = ~n1415 ;
  assign y443 = ~1'b0 ;
  assign y444 = n1416 ;
  assign y445 = ~n1420 ;
  assign y446 = ~1'b0 ;
  assign y447 = ~1'b0 ;
  assign y448 = n1424 ;
  assign y449 = ~1'b0 ;
  assign y450 = ~n1429 ;
  assign y451 = ~n1430 ;
  assign y452 = ~n1434 ;
  assign y453 = ~n1442 ;
  assign y454 = n1444 ;
  assign y455 = ~n1447 ;
  assign y456 = 1'b0 ;
  assign y457 = ~1'b0 ;
  assign y458 = n1453 ;
  assign y459 = n1454 ;
  assign y460 = ~1'b0 ;
  assign y461 = ~n1463 ;
  assign y462 = ~n1470 ;
  assign y463 = n1476 ;
  assign y464 = ~n1327 ;
  assign y465 = n1478 ;
  assign y466 = ~n1481 ;
  assign y467 = 1'b0 ;
  assign y468 = ~1'b0 ;
  assign y469 = ~n1482 ;
  assign y470 = n1486 ;
  assign y471 = ~n1489 ;
  assign y472 = ~1'b0 ;
  assign y473 = n1493 ;
  assign y474 = ~n1494 ;
  assign y475 = ~n1503 ;
  assign y476 = ~n1505 ;
  assign y477 = n1508 ;
  assign y478 = n1510 ;
  assign y479 = n1516 ;
  assign y480 = ~n1519 ;
  assign y481 = n1522 ;
  assign y482 = ~n1524 ;
  assign y483 = ~n1525 ;
  assign y484 = n1529 ;
  assign y485 = ~n1532 ;
  assign y486 = n1538 ;
  assign y487 = n1540 ;
  assign y488 = x182 ;
  assign y489 = ~1'b0 ;
  assign y490 = n1542 ;
  assign y491 = n1543 ;
  assign y492 = ~x150 ;
  assign y493 = n1552 ;
  assign y494 = ~n1554 ;
  assign y495 = ~n1555 ;
  assign y496 = ~n1557 ;
  assign y497 = n1559 ;
  assign y498 = 1'b0 ;
  assign y499 = n1563 ;
  assign y500 = n1564 ;
  assign y501 = n1569 ;
  assign y502 = ~n1570 ;
  assign y503 = ~n1574 ;
  assign y504 = ~1'b0 ;
  assign y505 = ~n1578 ;
  assign y506 = ~1'b0 ;
  assign y507 = ~n1582 ;
  assign y508 = ~1'b0 ;
  assign y509 = ~n1583 ;
  assign y510 = ~n1585 ;
  assign y511 = ~n1592 ;
  assign y512 = ~n1595 ;
  assign y513 = ~n1597 ;
  assign y514 = n1598 ;
  assign y515 = ~n1600 ;
  assign y516 = n1606 ;
  assign y517 = ~n1609 ;
  assign y518 = ~n1618 ;
  assign y519 = ~1'b0 ;
  assign y520 = ~1'b0 ;
  assign y521 = ~1'b0 ;
  assign y522 = n1620 ;
  assign y523 = ~n1624 ;
  assign y524 = n1628 ;
  assign y525 = n1630 ;
  assign y526 = ~n1637 ;
  assign y527 = n1655 ;
  assign y528 = ~1'b0 ;
  assign y529 = ~n1658 ;
  assign y530 = ~n1661 ;
  assign y531 = n1664 ;
  assign y532 = n1667 ;
  assign y533 = n1671 ;
  assign y534 = ~n1672 ;
  assign y535 = n1675 ;
  assign y536 = ~1'b0 ;
  assign y537 = ~1'b0 ;
  assign y538 = ~n1682 ;
  assign y539 = n1684 ;
  assign y540 = ~n1688 ;
  assign y541 = ~n1694 ;
  assign y542 = x159 ;
  assign y543 = ~n1695 ;
  assign y544 = n1696 ;
  assign y545 = n1702 ;
  assign y546 = n1705 ;
  assign y547 = ~n1719 ;
  assign y548 = ~n1722 ;
  assign y549 = n1723 ;
  assign y550 = n1727 ;
  assign y551 = n1728 ;
  assign y552 = ~n1742 ;
  assign y553 = ~n1744 ;
  assign y554 = ~1'b0 ;
  assign y555 = ~n1746 ;
  assign y556 = ~1'b0 ;
  assign y557 = ~n1748 ;
  assign y558 = n1749 ;
  assign y559 = n1752 ;
  assign y560 = ~1'b0 ;
  assign y561 = ~n1755 ;
  assign y562 = ~n1758 ;
  assign y563 = n1761 ;
  assign y564 = ~n1765 ;
  assign y565 = ~n256 ;
  assign y566 = n1773 ;
  assign y567 = ~n1775 ;
  assign y568 = n1788 ;
  assign y569 = ~1'b0 ;
  assign y570 = ~1'b0 ;
  assign y571 = ~n1806 ;
  assign y572 = ~1'b0 ;
  assign y573 = n1812 ;
  assign y574 = n1830 ;
  assign y575 = n1838 ;
  assign y576 = ~1'b0 ;
  assign y577 = 1'b0 ;
  assign y578 = n1845 ;
  assign y579 = n1847 ;
  assign y580 = n1848 ;
  assign y581 = n1849 ;
  assign y582 = ~1'b0 ;
  assign y583 = ~n1852 ;
  assign y584 = ~n1859 ;
  assign y585 = ~1'b0 ;
  assign y586 = ~1'b0 ;
  assign y587 = n1862 ;
  assign y588 = ~n1870 ;
  assign y589 = x184 ;
  assign y590 = ~n1879 ;
  assign y591 = ~1'b0 ;
  assign y592 = ~1'b0 ;
  assign y593 = ~n1882 ;
  assign y594 = ~n1885 ;
  assign y595 = ~n1886 ;
  assign y596 = ~n1896 ;
  assign y597 = n1902 ;
  assign y598 = n1907 ;
  assign y599 = ~n1912 ;
  assign y600 = n1913 ;
  assign y601 = ~n1922 ;
  assign y602 = n1249 ;
  assign y603 = n1927 ;
  assign y604 = ~1'b0 ;
  assign y605 = ~1'b0 ;
  assign y606 = ~n1930 ;
  assign y607 = ~n1933 ;
  assign y608 = ~1'b0 ;
  assign y609 = ~1'b0 ;
  assign y610 = ~n1937 ;
  assign y611 = n1940 ;
  assign y612 = ~1'b0 ;
  assign y613 = n1946 ;
  assign y614 = ~n1948 ;
  assign y615 = ~n1950 ;
  assign y616 = ~n1951 ;
  assign y617 = n1953 ;
  assign y618 = ~1'b0 ;
  assign y619 = ~n1961 ;
  assign y620 = n1963 ;
  assign y621 = ~n1964 ;
  assign y622 = n1969 ;
  assign y623 = ~n1972 ;
  assign y624 = ~1'b0 ;
  assign y625 = ~n1980 ;
  assign y626 = ~n1983 ;
  assign y627 = ~n1991 ;
  assign y628 = n1994 ;
  assign y629 = ~n1998 ;
  assign y630 = ~1'b0 ;
  assign y631 = n1999 ;
  assign y632 = ~n2003 ;
  assign y633 = ~n2007 ;
  assign y634 = ~n2016 ;
  assign y635 = ~n2023 ;
  assign y636 = ~1'b0 ;
  assign y637 = ~1'b0 ;
  assign y638 = ~n2024 ;
  assign y639 = n2025 ;
  assign y640 = n2026 ;
  assign y641 = ~1'b0 ;
  assign y642 = ~n2033 ;
  assign y643 = ~1'b0 ;
  assign y644 = n2035 ;
  assign y645 = n2043 ;
  assign y646 = ~n2048 ;
  assign y647 = ~n2050 ;
  assign y648 = n2059 ;
  assign y649 = ~n2062 ;
  assign y650 = ~n2077 ;
  assign y651 = ~n2082 ;
  assign y652 = ~n2085 ;
  assign y653 = ~n2086 ;
  assign y654 = n2094 ;
  assign y655 = n2095 ;
  assign y656 = n2098 ;
  assign y657 = ~n2100 ;
  assign y658 = ~n2103 ;
  assign y659 = n2111 ;
  assign y660 = n2113 ;
  assign y661 = n2114 ;
  assign y662 = ~n2116 ;
  assign y663 = ~n2123 ;
  assign y664 = ~n2131 ;
  assign y665 = ~n2135 ;
  assign y666 = ~n2138 ;
  assign y667 = ~1'b0 ;
  assign y668 = ~n2140 ;
  assign y669 = ~1'b0 ;
  assign y670 = n2142 ;
  assign y671 = ~n2144 ;
  assign y672 = n2145 ;
  assign y673 = n2146 ;
  assign y674 = n2150 ;
  assign y675 = ~n2154 ;
  assign y676 = n2155 ;
  assign y677 = ~1'b0 ;
  assign y678 = ~n2159 ;
  assign y679 = ~n2171 ;
  assign y680 = ~n2172 ;
  assign y681 = ~1'b0 ;
  assign y682 = n2173 ;
  assign y683 = ~n2176 ;
  assign y684 = n2178 ;
  assign y685 = ~n2179 ;
  assign y686 = ~n2183 ;
  assign y687 = n2186 ;
  assign y688 = n2189 ;
  assign y689 = ~n2196 ;
  assign y690 = ~n574 ;
  assign y691 = n2197 ;
  assign y692 = ~1'b0 ;
  assign y693 = n1980 ;
  assign y694 = ~n2209 ;
  assign y695 = n2217 ;
  assign y696 = n2219 ;
  assign y697 = ~1'b0 ;
  assign y698 = ~n2225 ;
  assign y699 = ~n1955 ;
  assign y700 = ~n2226 ;
  assign y701 = n2229 ;
  assign y702 = n2231 ;
  assign y703 = n2233 ;
  assign y704 = n2243 ;
  assign y705 = ~n2248 ;
  assign y706 = ~1'b0 ;
  assign y707 = ~n2250 ;
  assign y708 = ~n2253 ;
  assign y709 = ~n2255 ;
  assign y710 = ~n2262 ;
  assign y711 = ~n2263 ;
  assign y712 = n2268 ;
  assign y713 = ~n1110 ;
  assign y714 = n2270 ;
  assign y715 = ~n2274 ;
  assign y716 = ~n2275 ;
  assign y717 = n2282 ;
  assign y718 = ~n2284 ;
  assign y719 = ~n2287 ;
  assign y720 = ~n2295 ;
  assign y721 = 1'b0 ;
  assign y722 = ~n2302 ;
  assign y723 = ~1'b0 ;
  assign y724 = n2304 ;
  assign y725 = n2305 ;
  assign y726 = n2307 ;
  assign y727 = n2308 ;
  assign y728 = n2314 ;
  assign y729 = ~n2315 ;
  assign y730 = ~n2317 ;
  assign y731 = ~1'b0 ;
  assign y732 = n2319 ;
  assign y733 = n2328 ;
  assign y734 = ~n2329 ;
  assign y735 = n2331 ;
  assign y736 = ~1'b0 ;
  assign y737 = n2332 ;
  assign y738 = ~n2333 ;
  assign y739 = ~n2336 ;
  assign y740 = n2340 ;
  assign y741 = ~n2341 ;
  assign y742 = ~1'b0 ;
  assign y743 = ~1'b0 ;
  assign y744 = ~1'b0 ;
  assign y745 = ~n2342 ;
  assign y746 = ~n2344 ;
  assign y747 = ~n2346 ;
  assign y748 = ~n2347 ;
  assign y749 = ~n2350 ;
  assign y750 = n1778 ;
  assign y751 = ~n2352 ;
  assign y752 = ~1'b0 ;
  assign y753 = ~1'b0 ;
  assign y754 = ~n2354 ;
  assign y755 = ~n2356 ;
  assign y756 = ~n2357 ;
  assign y757 = n2358 ;
  assign y758 = ~n2359 ;
  assign y759 = n2362 ;
  assign y760 = ~n2363 ;
  assign y761 = ~x226 ;
  assign y762 = n2369 ;
  assign y763 = n2373 ;
  assign y764 = ~n2374 ;
  assign y765 = n2375 ;
  assign y766 = ~n2385 ;
  assign y767 = ~1'b0 ;
  assign y768 = ~n2386 ;
  assign y769 = n2389 ;
  assign y770 = n2390 ;
  assign y771 = ~n2391 ;
  assign y772 = n2396 ;
  assign y773 = n2397 ;
  assign y774 = ~1'b0 ;
  assign y775 = ~n2406 ;
  assign y776 = n2407 ;
  assign y777 = ~n2409 ;
  assign y778 = ~1'b0 ;
  assign y779 = ~1'b0 ;
  assign y780 = ~1'b0 ;
  assign y781 = ~n2411 ;
  assign y782 = ~n2421 ;
  assign y783 = ~n1576 ;
  assign y784 = ~n2423 ;
  assign y785 = n2427 ;
  assign y786 = ~1'b0 ;
  assign y787 = n2431 ;
  assign y788 = n2440 ;
  assign y789 = ~n2445 ;
  assign y790 = ~n2450 ;
  assign y791 = ~n2451 ;
  assign y792 = ~1'b0 ;
  assign y793 = n1203 ;
  assign y794 = ~n2463 ;
  assign y795 = ~n2465 ;
  assign y796 = ~n2469 ;
  assign y797 = ~n2472 ;
  assign y798 = ~1'b0 ;
  assign y799 = ~n2473 ;
  assign y800 = ~n2478 ;
  assign y801 = n2479 ;
  assign y802 = ~1'b0 ;
  assign y803 = ~n2484 ;
  assign y804 = ~n519 ;
  assign y805 = ~n2486 ;
  assign y806 = n2493 ;
  assign y807 = ~n2494 ;
  assign y808 = n2498 ;
  assign y809 = n2499 ;
  assign y810 = n2500 ;
  assign y811 = ~n2506 ;
  assign y812 = ~1'b0 ;
  assign y813 = ~1'b0 ;
  assign y814 = n2515 ;
  assign y815 = ~1'b0 ;
  assign y816 = n2516 ;
  assign y817 = ~n2526 ;
  assign y818 = ~1'b0 ;
  assign y819 = n2527 ;
  assign y820 = ~n2534 ;
  assign y821 = x103 ;
  assign y822 = ~n2538 ;
  assign y823 = ~1'b0 ;
  assign y824 = ~n2541 ;
  assign y825 = n2542 ;
  assign y826 = n2548 ;
  assign y827 = ~n2549 ;
  assign y828 = ~1'b0 ;
  assign y829 = ~n2555 ;
  assign y830 = ~1'b0 ;
  assign y831 = ~1'b0 ;
  assign y832 = ~n2565 ;
  assign y833 = ~1'b0 ;
  assign y834 = ~1'b0 ;
  assign y835 = n2568 ;
  assign y836 = 1'b0 ;
  assign y837 = n2573 ;
  assign y838 = ~1'b0 ;
  assign y839 = ~n2577 ;
  assign y840 = ~1'b0 ;
  assign y841 = n2578 ;
  assign y842 = ~n2580 ;
  assign y843 = n932 ;
  assign y844 = n2585 ;
  assign y845 = ~1'b0 ;
  assign y846 = ~n2586 ;
  assign y847 = ~n2590 ;
  assign y848 = n2595 ;
  assign y849 = ~n2598 ;
  assign y850 = ~1'b0 ;
  assign y851 = n2607 ;
  assign y852 = n2613 ;
  assign y853 = n2614 ;
  assign y854 = ~n2628 ;
  assign y855 = ~n2280 ;
  assign y856 = ~n2636 ;
  assign y857 = ~1'b0 ;
  assign y858 = n2640 ;
  assign y859 = n2643 ;
  assign y860 = ~n2647 ;
  assign y861 = ~1'b0 ;
  assign y862 = ~n2650 ;
  assign y863 = ~n1350 ;
  assign y864 = n2653 ;
  assign y865 = n2654 ;
  assign y866 = ~1'b0 ;
  assign y867 = ~1'b0 ;
  assign y868 = ~n2658 ;
  assign y869 = ~1'b0 ;
  assign y870 = n2661 ;
  assign y871 = n2663 ;
  assign y872 = n2667 ;
  assign y873 = n2670 ;
  assign y874 = n2671 ;
  assign y875 = ~1'b0 ;
  assign y876 = n2672 ;
  assign y877 = ~1'b0 ;
  assign y878 = n2683 ;
  assign y879 = n2688 ;
  assign y880 = ~1'b0 ;
  assign y881 = n2691 ;
  assign y882 = ~n2693 ;
  assign y883 = ~n2695 ;
  assign y884 = ~n2697 ;
  assign y885 = n2702 ;
  assign y886 = ~n2703 ;
  assign y887 = ~n2708 ;
  assign y888 = ~n2711 ;
  assign y889 = n2712 ;
  assign y890 = ~n2713 ;
  assign y891 = n2714 ;
  assign y892 = ~n2715 ;
  assign y893 = n2720 ;
  assign y894 = ~n2721 ;
  assign y895 = ~n2722 ;
  assign y896 = ~n2723 ;
  assign y897 = ~n2727 ;
  assign y898 = ~1'b0 ;
  assign y899 = ~n2729 ;
  assign y900 = ~n2737 ;
  assign y901 = ~n2748 ;
  assign y902 = ~1'b0 ;
  assign y903 = ~1'b0 ;
  assign y904 = ~n2750 ;
  assign y905 = ~1'b0 ;
  assign y906 = ~1'b0 ;
  assign y907 = ~1'b0 ;
  assign y908 = n2755 ;
  assign y909 = ~n2759 ;
  assign y910 = ~n2762 ;
  assign y911 = ~n2766 ;
  assign y912 = n2774 ;
  assign y913 = ~n2777 ;
  assign y914 = ~n2778 ;
  assign y915 = n2779 ;
  assign y916 = ~n2781 ;
  assign y917 = ~n2788 ;
  assign y918 = ~n2791 ;
  assign y919 = ~n2794 ;
  assign y920 = ~1'b0 ;
  assign y921 = n2800 ;
  assign y922 = ~1'b0 ;
  assign y923 = ~n2804 ;
  assign y924 = n2807 ;
  assign y925 = n2812 ;
  assign y926 = ~n2817 ;
  assign y927 = n2818 ;
  assign y928 = n2827 ;
  assign y929 = n2828 ;
  assign y930 = n2830 ;
  assign y931 = n2831 ;
  assign y932 = n2832 ;
  assign y933 = ~n2836 ;
  assign y934 = ~1'b0 ;
  assign y935 = ~1'b0 ;
  assign y936 = n2837 ;
  assign y937 = ~n2841 ;
  assign y938 = ~n2845 ;
  assign y939 = ~n2846 ;
  assign y940 = ~1'b0 ;
  assign y941 = ~n2849 ;
  assign y942 = ~n2850 ;
  assign y943 = ~n2853 ;
  assign y944 = x159 ;
  assign y945 = n2854 ;
  assign y946 = n2857 ;
  assign y947 = ~n2861 ;
  assign y948 = n2863 ;
  assign y949 = ~n2865 ;
  assign y950 = ~n2874 ;
  assign y951 = ~n2879 ;
  assign y952 = ~1'b0 ;
  assign y953 = ~n2883 ;
  assign y954 = n2886 ;
  assign y955 = ~1'b0 ;
  assign y956 = ~1'b0 ;
  assign y957 = ~n2887 ;
  assign y958 = ~n2893 ;
  assign y959 = ~n2906 ;
  assign y960 = n2909 ;
  assign y961 = ~n2910 ;
  assign y962 = ~n2911 ;
  assign y963 = n2917 ;
  assign y964 = n2922 ;
  assign y965 = n2927 ;
  assign y966 = ~n2934 ;
  assign y967 = ~1'b0 ;
  assign y968 = ~n2937 ;
  assign y969 = n2938 ;
  assign y970 = ~n2943 ;
  assign y971 = n2946 ;
  assign y972 = ~n2948 ;
  assign y973 = n2951 ;
  assign y974 = n2954 ;
  assign y975 = n2959 ;
  assign y976 = n2962 ;
  assign y977 = ~n2967 ;
  assign y978 = ~n1655 ;
  assign y979 = ~n2968 ;
  assign y980 = ~n2972 ;
  assign y981 = n2978 ;
  assign y982 = ~n2980 ;
  assign y983 = ~n2985 ;
  assign y984 = ~1'b0 ;
  assign y985 = ~n2990 ;
  assign y986 = ~n2993 ;
  assign y987 = ~1'b0 ;
  assign y988 = ~n2997 ;
  assign y989 = ~n2998 ;
  assign y990 = ~1'b0 ;
  assign y991 = n3000 ;
  assign y992 = ~n3010 ;
  assign y993 = ~n3011 ;
  assign y994 = ~1'b0 ;
  assign y995 = ~n3014 ;
  assign y996 = n3017 ;
  assign y997 = ~n3023 ;
  assign y998 = ~n3033 ;
  assign y999 = n3036 ;
  assign y1000 = n3042 ;
  assign y1001 = n3044 ;
  assign y1002 = ~n3051 ;
  assign y1003 = ~n3063 ;
  assign y1004 = ~n3064 ;
  assign y1005 = n3065 ;
  assign y1006 = ~1'b0 ;
  assign y1007 = ~n3071 ;
  assign y1008 = ~1'b0 ;
  assign y1009 = ~n3075 ;
  assign y1010 = 1'b0 ;
  assign y1011 = ~n3079 ;
  assign y1012 = n3090 ;
  assign y1013 = ~n3095 ;
  assign y1014 = ~1'b0 ;
  assign y1015 = n3096 ;
  assign y1016 = n3097 ;
  assign y1017 = ~n3106 ;
  assign y1018 = n3107 ;
  assign y1019 = ~1'b0 ;
  assign y1020 = ~n3108 ;
  assign y1021 = ~n3112 ;
  assign y1022 = n3115 ;
  assign y1023 = ~1'b0 ;
  assign y1024 = n3121 ;
  assign y1025 = ~n3125 ;
  assign y1026 = n3133 ;
  assign y1027 = ~n3136 ;
  assign y1028 = ~n3139 ;
  assign y1029 = n3144 ;
  assign y1030 = ~n3147 ;
  assign y1031 = n3148 ;
  assign y1032 = ~1'b0 ;
  assign y1033 = n3150 ;
  assign y1034 = ~1'b0 ;
  assign y1035 = ~1'b0 ;
  assign y1036 = n3155 ;
  assign y1037 = ~n3163 ;
  assign y1038 = n3166 ;
  assign y1039 = ~n3168 ;
  assign y1040 = ~1'b0 ;
  assign y1041 = n3170 ;
  assign y1042 = ~n3173 ;
  assign y1043 = ~n3176 ;
  assign y1044 = ~1'b0 ;
  assign y1045 = n3194 ;
  assign y1046 = ~n2701 ;
  assign y1047 = ~1'b0 ;
  assign y1048 = n3200 ;
  assign y1049 = ~n3211 ;
  assign y1050 = ~n3213 ;
  assign y1051 = ~n3215 ;
  assign y1052 = n3216 ;
  assign y1053 = ~n3217 ;
  assign y1054 = ~1'b0 ;
  assign y1055 = n3219 ;
  assign y1056 = ~n3220 ;
  assign y1057 = n3222 ;
  assign y1058 = n3225 ;
  assign y1059 = ~n3227 ;
  assign y1060 = n3229 ;
  assign y1061 = n3236 ;
  assign y1062 = ~n3239 ;
  assign y1063 = n3245 ;
  assign y1064 = ~1'b0 ;
  assign y1065 = ~1'b0 ;
  assign y1066 = n3250 ;
  assign y1067 = n3256 ;
  assign y1068 = ~1'b0 ;
  assign y1069 = n3259 ;
  assign y1070 = n3260 ;
  assign y1071 = ~n3262 ;
  assign y1072 = ~1'b0 ;
  assign y1073 = ~n3281 ;
  assign y1074 = ~n3282 ;
  assign y1075 = ~n3288 ;
  assign y1076 = ~n3294 ;
  assign y1077 = n3297 ;
  assign y1078 = n3302 ;
  assign y1079 = ~n3304 ;
  assign y1080 = ~1'b0 ;
  assign y1081 = n3312 ;
  assign y1082 = ~1'b0 ;
  assign y1083 = ~n3314 ;
  assign y1084 = n3320 ;
  assign y1085 = ~n3321 ;
  assign y1086 = n3322 ;
  assign y1087 = ~n3324 ;
  assign y1088 = n3331 ;
  assign y1089 = ~n3335 ;
  assign y1090 = ~1'b0 ;
  assign y1091 = n3336 ;
  assign y1092 = ~n3341 ;
  assign y1093 = ~n3342 ;
  assign y1094 = n3344 ;
  assign y1095 = n3348 ;
  assign y1096 = ~1'b0 ;
  assign y1097 = n3360 ;
  assign y1098 = ~n3371 ;
  assign y1099 = n3383 ;
  assign y1100 = ~1'b0 ;
  assign y1101 = ~1'b0 ;
  assign y1102 = ~1'b0 ;
  assign y1103 = n3386 ;
  assign y1104 = n3389 ;
  assign y1105 = ~n3396 ;
  assign y1106 = ~1'b0 ;
  assign y1107 = ~n3401 ;
  assign y1108 = ~1'b0 ;
  assign y1109 = ~1'b0 ;
  assign y1110 = n3403 ;
  assign y1111 = n3404 ;
  assign y1112 = ~1'b0 ;
  assign y1113 = n3412 ;
  assign y1114 = n3414 ;
  assign y1115 = ~1'b0 ;
  assign y1116 = n3417 ;
  assign y1117 = ~1'b0 ;
  assign y1118 = n3418 ;
  assign y1119 = ~n3421 ;
  assign y1120 = ~n2541 ;
  assign y1121 = n3422 ;
  assign y1122 = ~1'b0 ;
  assign y1123 = ~n3425 ;
  assign y1124 = n3428 ;
  assign y1125 = n3433 ;
  assign y1126 = ~n3437 ;
  assign y1127 = ~1'b0 ;
  assign y1128 = n3440 ;
  assign y1129 = ~n3442 ;
  assign y1130 = n3086 ;
  assign y1131 = ~n3453 ;
  assign y1132 = n3457 ;
  assign y1133 = ~1'b0 ;
  assign y1134 = n3458 ;
  assign y1135 = ~1'b0 ;
  assign y1136 = n3463 ;
  assign y1137 = ~n3464 ;
  assign y1138 = ~1'b0 ;
  assign y1139 = ~1'b0 ;
  assign y1140 = ~n3466 ;
  assign y1141 = ~n1684 ;
  assign y1142 = ~1'b0 ;
  assign y1143 = n3469 ;
  assign y1144 = n3474 ;
  assign y1145 = ~1'b0 ;
  assign y1146 = ~n3487 ;
  assign y1147 = ~n3497 ;
  assign y1148 = n3508 ;
  assign y1149 = ~1'b0 ;
  assign y1150 = ~1'b0 ;
  assign y1151 = ~1'b0 ;
  assign y1152 = ~n3518 ;
  assign y1153 = ~1'b0 ;
  assign y1154 = ~n3525 ;
  assign y1155 = n3527 ;
  assign y1156 = ~n3531 ;
  assign y1157 = ~n3539 ;
  assign y1158 = n3540 ;
  assign y1159 = ~n3544 ;
  assign y1160 = ~1'b0 ;
  assign y1161 = n3547 ;
  assign y1162 = ~n3550 ;
  assign y1163 = ~n3556 ;
  assign y1164 = n3559 ;
  assign y1165 = n3564 ;
  assign y1166 = ~1'b0 ;
  assign y1167 = ~1'b0 ;
  assign y1168 = ~n3573 ;
  assign y1169 = n3578 ;
  assign y1170 = ~n3583 ;
  assign y1171 = ~n3587 ;
  assign y1172 = ~n3591 ;
  assign y1173 = n3593 ;
  assign y1174 = n2259 ;
  assign y1175 = ~1'b0 ;
  assign y1176 = ~n3595 ;
  assign y1177 = n3599 ;
  assign y1178 = ~n3600 ;
  assign y1179 = 1'b0 ;
  assign y1180 = ~n3602 ;
  assign y1181 = ~n3604 ;
  assign y1182 = n3608 ;
  assign y1183 = ~1'b0 ;
  assign y1184 = ~n3617 ;
  assign y1185 = ~n403 ;
  assign y1186 = ~n3619 ;
  assign y1187 = ~1'b0 ;
  assign y1188 = ~n3620 ;
  assign y1189 = ~1'b0 ;
  assign y1190 = ~n3622 ;
  assign y1191 = n3624 ;
  assign y1192 = n3629 ;
  assign y1193 = n3630 ;
  assign y1194 = ~n3638 ;
  assign y1195 = ~n3641 ;
  assign y1196 = ~n3646 ;
  assign y1197 = ~n3648 ;
  assign y1198 = n3652 ;
  assign y1199 = ~n3653 ;
  assign y1200 = ~1'b0 ;
  assign y1201 = ~1'b0 ;
  assign y1202 = n3658 ;
  assign y1203 = n292 ;
  assign y1204 = n3659 ;
  assign y1205 = ~n3661 ;
  assign y1206 = n3662 ;
  assign y1207 = ~n3666 ;
  assign y1208 = ~n3667 ;
  assign y1209 = n3669 ;
  assign y1210 = n1593 ;
  assign y1211 = ~n3675 ;
  assign y1212 = ~n3676 ;
  assign y1213 = ~1'b0 ;
  assign y1214 = ~n3685 ;
  assign y1215 = ~1'b0 ;
  assign y1216 = n3691 ;
  assign y1217 = ~n3694 ;
  assign y1218 = n3698 ;
  assign y1219 = ~1'b0 ;
  assign y1220 = ~n3702 ;
  assign y1221 = ~1'b0 ;
  assign y1222 = n3704 ;
  assign y1223 = n3707 ;
  assign y1224 = ~n3715 ;
  assign y1225 = n3721 ;
  assign y1226 = n3722 ;
  assign y1227 = n3724 ;
  assign y1228 = ~n3725 ;
  assign y1229 = ~1'b0 ;
  assign y1230 = ~n3726 ;
  assign y1231 = ~n3730 ;
  assign y1232 = 1'b0 ;
  assign y1233 = n3731 ;
  assign y1234 = ~n3740 ;
  assign y1235 = ~1'b0 ;
  assign y1236 = ~n3747 ;
  assign y1237 = ~n3751 ;
  assign y1238 = ~n3756 ;
  assign y1239 = ~n3764 ;
  assign y1240 = n3768 ;
  assign y1241 = n3771 ;
  assign y1242 = ~1'b0 ;
  assign y1243 = n3773 ;
  assign y1244 = ~n3779 ;
  assign y1245 = n3781 ;
  assign y1246 = ~n3782 ;
  assign y1247 = ~n3790 ;
  assign y1248 = ~n3791 ;
  assign y1249 = ~n3792 ;
  assign y1250 = n3795 ;
  assign y1251 = ~1'b0 ;
  assign y1252 = ~n3796 ;
  assign y1253 = ~1'b0 ;
  assign y1254 = ~n3806 ;
  assign y1255 = ~1'b0 ;
  assign y1256 = ~n3821 ;
  assign y1257 = ~n3823 ;
  assign y1258 = ~n898 ;
  assign y1259 = n3830 ;
  assign y1260 = ~n3836 ;
  assign y1261 = ~1'b0 ;
  assign y1262 = ~1'b0 ;
  assign y1263 = n3837 ;
  assign y1264 = ~n3024 ;
  assign y1265 = ~1'b0 ;
  assign y1266 = n3840 ;
  assign y1267 = ~1'b0 ;
  assign y1268 = ~n3842 ;
  assign y1269 = n3848 ;
  assign y1270 = ~1'b0 ;
  assign y1271 = n3853 ;
  assign y1272 = n3855 ;
  assign y1273 = n3859 ;
  assign y1274 = ~1'b0 ;
  assign y1275 = ~n3865 ;
  assign y1276 = ~n3869 ;
  assign y1277 = n3874 ;
  assign y1278 = ~1'b0 ;
  assign y1279 = ~n3880 ;
  assign y1280 = ~1'b0 ;
  assign y1281 = ~n3887 ;
  assign y1282 = ~n3889 ;
  assign y1283 = ~n3891 ;
  assign y1284 = ~n3899 ;
  assign y1285 = n3900 ;
  assign y1286 = ~n3907 ;
  assign y1287 = ~n3912 ;
  assign y1288 = ~n3919 ;
  assign y1289 = ~n3923 ;
  assign y1290 = ~n3926 ;
  assign y1291 = ~n3939 ;
  assign y1292 = n3941 ;
  assign y1293 = ~1'b0 ;
  assign y1294 = n3944 ;
  assign y1295 = ~n3949 ;
  assign y1296 = ~1'b0 ;
  assign y1297 = n3953 ;
  assign y1298 = n3959 ;
  assign y1299 = ~1'b0 ;
  assign y1300 = n3960 ;
  assign y1301 = ~n3963 ;
  assign y1302 = n3965 ;
  assign y1303 = ~n3966 ;
  assign y1304 = ~1'b0 ;
  assign y1305 = ~n3978 ;
  assign y1306 = ~1'b0 ;
  assign y1307 = ~n3980 ;
  assign y1308 = ~n3986 ;
  assign y1309 = ~1'b0 ;
  assign y1310 = ~1'b0 ;
  assign y1311 = ~n3987 ;
  assign y1312 = ~n3989 ;
  assign y1313 = ~n3990 ;
  assign y1314 = ~n3991 ;
  assign y1315 = n3995 ;
  assign y1316 = ~1'b0 ;
  assign y1317 = n3998 ;
  assign y1318 = ~n3999 ;
  assign y1319 = ~1'b0 ;
  assign y1320 = n4004 ;
  assign y1321 = n4005 ;
  assign y1322 = ~n4006 ;
  assign y1323 = n4008 ;
  assign y1324 = ~1'b0 ;
  assign y1325 = ~1'b0 ;
  assign y1326 = ~n4019 ;
  assign y1327 = ~n4031 ;
  assign y1328 = ~n4032 ;
  assign y1329 = n4036 ;
  assign y1330 = ~n4039 ;
  assign y1331 = ~1'b0 ;
  assign y1332 = n4043 ;
  assign y1333 = ~1'b0 ;
  assign y1334 = ~n4047 ;
  assign y1335 = n4048 ;
  assign y1336 = ~1'b0 ;
  assign y1337 = n4049 ;
  assign y1338 = ~1'b0 ;
  assign y1339 = n4050 ;
  assign y1340 = n4055 ;
  assign y1341 = ~n4056 ;
  assign y1342 = ~n4060 ;
  assign y1343 = n4065 ;
  assign y1344 = n4070 ;
  assign y1345 = n4074 ;
  assign y1346 = ~n4081 ;
  assign y1347 = n4083 ;
  assign y1348 = n4086 ;
  assign y1349 = ~1'b0 ;
  assign y1350 = n4088 ;
  assign y1351 = ~n4089 ;
  assign y1352 = ~n4090 ;
  assign y1353 = ~n4091 ;
  assign y1354 = n1463 ;
  assign y1355 = ~n4093 ;
  assign y1356 = n3381 ;
  assign y1357 = ~n4103 ;
  assign y1358 = ~n4104 ;
  assign y1359 = ~n4112 ;
  assign y1360 = ~1'b0 ;
  assign y1361 = n4113 ;
  assign y1362 = ~n4117 ;
  assign y1363 = n4121 ;
  assign y1364 = n4123 ;
  assign y1365 = n4127 ;
  assign y1366 = ~n4128 ;
  assign y1367 = n4129 ;
  assign y1368 = n4130 ;
  assign y1369 = 1'b0 ;
  assign y1370 = n4133 ;
  assign y1371 = n4138 ;
  assign y1372 = n4141 ;
  assign y1373 = n4144 ;
  assign y1374 = ~n4147 ;
  assign y1375 = n4153 ;
  assign y1376 = ~n4158 ;
  assign y1377 = ~n4168 ;
  assign y1378 = ~n4172 ;
  assign y1379 = n4174 ;
  assign y1380 = n4177 ;
  assign y1381 = ~n4182 ;
  assign y1382 = ~n4185 ;
  assign y1383 = ~n4189 ;
  assign y1384 = ~1'b0 ;
  assign y1385 = ~n4195 ;
  assign y1386 = n4198 ;
  assign y1387 = ~n4199 ;
  assign y1388 = n4209 ;
  assign y1389 = n4150 ;
  assign y1390 = n4212 ;
  assign y1391 = ~1'b0 ;
  assign y1392 = n4217 ;
  assign y1393 = n4220 ;
  assign y1394 = n4223 ;
  assign y1395 = ~n4227 ;
  assign y1396 = ~1'b0 ;
  assign y1397 = ~n4229 ;
  assign y1398 = n4230 ;
  assign y1399 = ~1'b0 ;
  assign y1400 = ~n4233 ;
  assign y1401 = ~1'b0 ;
  assign y1402 = ~n4236 ;
  assign y1403 = ~1'b0 ;
  assign y1404 = ~n4241 ;
  assign y1405 = n4243 ;
  assign y1406 = n4245 ;
  assign y1407 = n4251 ;
  assign y1408 = n4255 ;
  assign y1409 = n4256 ;
  assign y1410 = n4258 ;
  assign y1411 = n4261 ;
  assign y1412 = n4271 ;
  assign y1413 = ~n4273 ;
  assign y1414 = n4288 ;
  assign y1415 = n4294 ;
  assign y1416 = n4299 ;
  assign y1417 = n4301 ;
  assign y1418 = ~n4303 ;
  assign y1419 = ~n4307 ;
  assign y1420 = ~1'b0 ;
  assign y1421 = n4308 ;
  assign y1422 = n4310 ;
  assign y1423 = ~n4313 ;
  assign y1424 = ~n4321 ;
  assign y1425 = n4322 ;
  assign y1426 = ~n4324 ;
  assign y1427 = ~n449 ;
  assign y1428 = ~n4330 ;
  assign y1429 = n4333 ;
  assign y1430 = ~1'b0 ;
  assign y1431 = n4334 ;
  assign y1432 = n4336 ;
  assign y1433 = ~n4346 ;
  assign y1434 = ~1'b0 ;
  assign y1435 = n4347 ;
  assign y1436 = n4352 ;
  assign y1437 = ~n4359 ;
  assign y1438 = ~n4361 ;
  assign y1439 = n4363 ;
  assign y1440 = ~1'b0 ;
  assign y1441 = ~n4364 ;
  assign y1442 = ~n4370 ;
  assign y1443 = ~n4372 ;
  assign y1444 = ~n4374 ;
  assign y1445 = n4379 ;
  assign y1446 = n4386 ;
  assign y1447 = ~n4388 ;
  assign y1448 = n4389 ;
  assign y1449 = ~n4394 ;
  assign y1450 = n4396 ;
  assign y1451 = ~1'b0 ;
  assign y1452 = ~n4397 ;
  assign y1453 = ~n4400 ;
  assign y1454 = ~n4404 ;
  assign y1455 = n4411 ;
  assign y1456 = n4414 ;
  assign y1457 = ~1'b0 ;
  assign y1458 = ~n4419 ;
  assign y1459 = ~1'b0 ;
  assign y1460 = n4422 ;
  assign y1461 = ~n4424 ;
  assign y1462 = n4426 ;
  assign y1463 = ~1'b0 ;
  assign y1464 = ~1'b0 ;
  assign y1465 = ~n4427 ;
  assign y1466 = n4433 ;
  assign y1467 = ~1'b0 ;
  assign y1468 = n4434 ;
  assign y1469 = ~n4437 ;
  assign y1470 = ~n4438 ;
  assign y1471 = n4439 ;
  assign y1472 = n4444 ;
  assign y1473 = n4446 ;
  assign y1474 = ~n4447 ;
  assign y1475 = ~n4448 ;
  assign y1476 = ~1'b0 ;
  assign y1477 = ~n4450 ;
  assign y1478 = ~1'b0 ;
  assign y1479 = ~n4451 ;
  assign y1480 = n4457 ;
  assign y1481 = ~n4461 ;
  assign y1482 = ~1'b0 ;
  assign y1483 = ~n4462 ;
  assign y1484 = ~1'b0 ;
  assign y1485 = ~n4465 ;
  assign y1486 = 1'b0 ;
  assign y1487 = ~n4468 ;
  assign y1488 = ~1'b0 ;
  assign y1489 = ~n4472 ;
  assign y1490 = ~1'b0 ;
  assign y1491 = n4473 ;
  assign y1492 = n4481 ;
  assign y1493 = n4484 ;
  assign y1494 = ~n4485 ;
  assign y1495 = n4487 ;
  assign y1496 = ~n4489 ;
  assign y1497 = ~n4490 ;
  assign y1498 = ~n4499 ;
  assign y1499 = ~n4505 ;
  assign y1500 = ~1'b0 ;
  assign y1501 = ~1'b0 ;
  assign y1502 = ~1'b0 ;
  assign y1503 = n4506 ;
  assign y1504 = n1542 ;
  assign y1505 = n4508 ;
  assign y1506 = ~n4515 ;
  assign y1507 = ~1'b0 ;
  assign y1508 = ~n4517 ;
  assign y1509 = ~n4523 ;
  assign y1510 = ~n4525 ;
  assign y1511 = n4527 ;
  assign y1512 = ~n4532 ;
  assign y1513 = ~n4533 ;
  assign y1514 = ~n4536 ;
  assign y1515 = n4537 ;
  assign y1516 = n4542 ;
  assign y1517 = n4544 ;
  assign y1518 = ~1'b0 ;
  assign y1519 = ~n4547 ;
  assign y1520 = ~n4548 ;
  assign y1521 = ~n4550 ;
  assign y1522 = n4552 ;
  assign y1523 = ~1'b0 ;
  assign y1524 = ~n4553 ;
  assign y1525 = ~n4555 ;
  assign y1526 = ~n4561 ;
  assign y1527 = ~n4567 ;
  assign y1528 = ~n4578 ;
  assign y1529 = n4580 ;
  assign y1530 = ~n4587 ;
  assign y1531 = ~1'b0 ;
  assign y1532 = ~n4589 ;
  assign y1533 = ~1'b0 ;
  assign y1534 = ~n4597 ;
  assign y1535 = ~n4600 ;
  assign y1536 = ~n4601 ;
  assign y1537 = n4606 ;
  assign y1538 = ~1'b0 ;
  assign y1539 = n4616 ;
  assign y1540 = ~n4628 ;
  assign y1541 = ~n4630 ;
  assign y1542 = ~n4633 ;
  assign y1543 = ~n4637 ;
  assign y1544 = ~n4638 ;
  assign y1545 = ~n4642 ;
  assign y1546 = ~1'b0 ;
  assign y1547 = ~1'b0 ;
  assign y1548 = ~n4646 ;
  assign y1549 = ~n4652 ;
  assign y1550 = ~1'b0 ;
  assign y1551 = ~n4659 ;
  assign y1552 = ~n4666 ;
  assign y1553 = ~n4672 ;
  assign y1554 = n4676 ;
  assign y1555 = n4677 ;
  assign y1556 = ~1'b0 ;
  assign y1557 = ~1'b0 ;
  assign y1558 = n4678 ;
  assign y1559 = ~n4686 ;
  assign y1560 = ~n4696 ;
  assign y1561 = ~1'b0 ;
  assign y1562 = ~n4697 ;
  assign y1563 = ~1'b0 ;
  assign y1564 = ~n4698 ;
  assign y1565 = n4700 ;
  assign y1566 = n4701 ;
  assign y1567 = n4703 ;
  assign y1568 = n4707 ;
  assign y1569 = ~n4711 ;
  assign y1570 = ~1'b0 ;
  assign y1571 = ~1'b0 ;
  assign y1572 = ~n4712 ;
  assign y1573 = n4714 ;
  assign y1574 = n4715 ;
  assign y1575 = n4717 ;
  assign y1576 = n4722 ;
  assign y1577 = n4724 ;
  assign y1578 = n4731 ;
  assign y1579 = n4733 ;
  assign y1580 = ~n4735 ;
  assign y1581 = ~1'b0 ;
  assign y1582 = ~1'b0 ;
  assign y1583 = n4738 ;
  assign y1584 = n4744 ;
  assign y1585 = n4745 ;
  assign y1586 = n4756 ;
  assign y1587 = ~n4758 ;
  assign y1588 = ~n4766 ;
  assign y1589 = n4773 ;
  assign y1590 = ~n4783 ;
  assign y1591 = ~1'b0 ;
  assign y1592 = n3516 ;
  assign y1593 = ~n4784 ;
  assign y1594 = ~1'b0 ;
  assign y1595 = n4790 ;
  assign y1596 = n4792 ;
  assign y1597 = n4797 ;
  assign y1598 = ~n4803 ;
  assign y1599 = n4804 ;
  assign y1600 = ~n4807 ;
  assign y1601 = ~n4809 ;
  assign y1602 = n4812 ;
  assign y1603 = n4816 ;
  assign y1604 = ~n4826 ;
  assign y1605 = ~n4827 ;
  assign y1606 = ~n4832 ;
  assign y1607 = ~1'b0 ;
  assign y1608 = n4833 ;
  assign y1609 = ~n4835 ;
  assign y1610 = ~n4836 ;
  assign y1611 = ~n4840 ;
  assign y1612 = n4844 ;
  assign y1613 = ~n4847 ;
  assign y1614 = ~n4848 ;
  assign y1615 = ~n4852 ;
  assign y1616 = ~n4854 ;
  assign y1617 = ~1'b0 ;
  assign y1618 = ~n4855 ;
  assign y1619 = ~n2223 ;
  assign y1620 = n4870 ;
  assign y1621 = n4872 ;
  assign y1622 = ~1'b0 ;
  assign y1623 = n4881 ;
  assign y1624 = n4883 ;
  assign y1625 = ~1'b0 ;
  assign y1626 = ~n4886 ;
  assign y1627 = ~n4889 ;
  assign y1628 = ~n4890 ;
  assign y1629 = n4898 ;
  assign y1630 = ~n4906 ;
  assign y1631 = ~n4912 ;
  assign y1632 = ~n4916 ;
  assign y1633 = ~n4917 ;
  assign y1634 = ~1'b0 ;
  assign y1635 = ~n4919 ;
  assign y1636 = ~1'b0 ;
  assign y1637 = ~1'b0 ;
  assign y1638 = n4920 ;
  assign y1639 = ~n4927 ;
  assign y1640 = ~1'b0 ;
  assign y1641 = n4929 ;
  assign y1642 = ~n4941 ;
  assign y1643 = ~1'b0 ;
  assign y1644 = ~n4943 ;
  assign y1645 = ~n4947 ;
  assign y1646 = ~n4953 ;
  assign y1647 = n4954 ;
  assign y1648 = ~n4955 ;
  assign y1649 = n4961 ;
  assign y1650 = n4978 ;
  assign y1651 = ~n4981 ;
  assign y1652 = n4984 ;
  assign y1653 = ~n4986 ;
  assign y1654 = n4987 ;
  assign y1655 = ~1'b0 ;
  assign y1656 = n3766 ;
  assign y1657 = n4989 ;
  assign y1658 = ~1'b0 ;
  assign y1659 = ~n4992 ;
  assign y1660 = ~n5001 ;
  assign y1661 = n5007 ;
  assign y1662 = ~n5009 ;
  assign y1663 = n5015 ;
  assign y1664 = ~n5018 ;
  assign y1665 = ~n5020 ;
  assign y1666 = n5022 ;
  assign y1667 = ~1'b0 ;
  assign y1668 = n5025 ;
  assign y1669 = ~n5032 ;
  assign y1670 = n5039 ;
  assign y1671 = n5044 ;
  assign y1672 = ~n5047 ;
  assign y1673 = ~n5049 ;
  assign y1674 = n5055 ;
  assign y1675 = n5062 ;
  assign y1676 = n5073 ;
  assign y1677 = ~n5076 ;
  assign y1678 = ~n5077 ;
  assign y1679 = ~n5079 ;
  assign y1680 = ~1'b0 ;
  assign y1681 = ~n5081 ;
  assign y1682 = ~n5090 ;
  assign y1683 = ~1'b0 ;
  assign y1684 = ~1'b0 ;
  assign y1685 = ~n3097 ;
  assign y1686 = n5093 ;
  assign y1687 = ~1'b0 ;
  assign y1688 = ~n5095 ;
  assign y1689 = ~1'b0 ;
  assign y1690 = ~1'b0 ;
  assign y1691 = n5101 ;
  assign y1692 = n5102 ;
  assign y1693 = ~n5104 ;
  assign y1694 = ~n5108 ;
  assign y1695 = ~n5117 ;
  assign y1696 = n5119 ;
  assign y1697 = ~n5121 ;
  assign y1698 = ~1'b0 ;
  assign y1699 = ~n5124 ;
  assign y1700 = ~n5126 ;
  assign y1701 = ~n5129 ;
  assign y1702 = n5131 ;
  assign y1703 = ~1'b0 ;
  assign y1704 = n5135 ;
  assign y1705 = n5137 ;
  assign y1706 = n5149 ;
  assign y1707 = ~1'b0 ;
  assign y1708 = ~n5158 ;
  assign y1709 = ~n5165 ;
  assign y1710 = ~1'b0 ;
  assign y1711 = n5173 ;
  assign y1712 = n5175 ;
  assign y1713 = ~n5187 ;
  assign y1714 = ~1'b0 ;
  assign y1715 = ~n5191 ;
  assign y1716 = ~n5197 ;
  assign y1717 = ~n5198 ;
  assign y1718 = n1107 ;
  assign y1719 = ~n5201 ;
  assign y1720 = ~n5204 ;
  assign y1721 = ~1'b0 ;
  assign y1722 = ~1'b0 ;
  assign y1723 = n5209 ;
  assign y1724 = n5215 ;
  assign y1725 = ~n5219 ;
  assign y1726 = n5223 ;
  assign y1727 = ~n5228 ;
  assign y1728 = ~n5232 ;
  assign y1729 = ~n5236 ;
  assign y1730 = n5239 ;
  assign y1731 = n5242 ;
  assign y1732 = n5244 ;
  assign y1733 = ~1'b0 ;
  assign y1734 = n5258 ;
  assign y1735 = n5262 ;
  assign y1736 = ~n5272 ;
  assign y1737 = n5279 ;
  assign y1738 = n5281 ;
  assign y1739 = ~1'b0 ;
  assign y1740 = n5290 ;
  assign y1741 = ~1'b0 ;
  assign y1742 = n5291 ;
  assign y1743 = n5292 ;
  assign y1744 = ~1'b0 ;
  assign y1745 = ~n5300 ;
  assign y1746 = ~n5305 ;
  assign y1747 = ~n5306 ;
  assign y1748 = n5308 ;
  assign y1749 = n5313 ;
  assign y1750 = n5316 ;
  assign y1751 = n5322 ;
  assign y1752 = ~n5325 ;
  assign y1753 = ~n5330 ;
  assign y1754 = n5333 ;
  assign y1755 = ~n5335 ;
  assign y1756 = ~n5342 ;
  assign y1757 = ~1'b0 ;
  assign y1758 = 1'b0 ;
  assign y1759 = ~n5345 ;
  assign y1760 = ~n5347 ;
  assign y1761 = ~n5349 ;
  assign y1762 = ~n5357 ;
  assign y1763 = n5361 ;
  assign y1764 = ~n5367 ;
  assign y1765 = ~n5371 ;
  assign y1766 = ~1'b0 ;
  assign y1767 = n5374 ;
  assign y1768 = n3390 ;
  assign y1769 = ~n5384 ;
  assign y1770 = ~n5385 ;
  assign y1771 = ~n5386 ;
  assign y1772 = ~n5387 ;
  assign y1773 = ~n5388 ;
  assign y1774 = ~1'b0 ;
  assign y1775 = ~n5395 ;
  assign y1776 = n5396 ;
  assign y1777 = ~n5398 ;
  assign y1778 = n5404 ;
  assign y1779 = ~1'b0 ;
  assign y1780 = ~n5406 ;
  assign y1781 = n5408 ;
  assign y1782 = ~n5415 ;
  assign y1783 = ~1'b0 ;
  assign y1784 = ~n5416 ;
  assign y1785 = ~n5419 ;
  assign y1786 = ~1'b0 ;
  assign y1787 = n3578 ;
  assign y1788 = ~1'b0 ;
  assign y1789 = ~1'b0 ;
  assign y1790 = n5420 ;
  assign y1791 = n5422 ;
  assign y1792 = ~n5430 ;
  assign y1793 = n5436 ;
  assign y1794 = ~n1145 ;
  assign y1795 = ~n1051 ;
  assign y1796 = ~n5437 ;
  assign y1797 = n5445 ;
  assign y1798 = ~1'b0 ;
  assign y1799 = ~n5447 ;
  assign y1800 = n5449 ;
  assign y1801 = ~n5453 ;
  assign y1802 = ~1'b0 ;
  assign y1803 = ~n5454 ;
  assign y1804 = n5459 ;
  assign y1805 = ~n5460 ;
  assign y1806 = ~1'b0 ;
  assign y1807 = n5463 ;
  assign y1808 = ~1'b0 ;
  assign y1809 = ~1'b0 ;
  assign y1810 = ~n5468 ;
  assign y1811 = ~n5471 ;
  assign y1812 = n5472 ;
  assign y1813 = n5473 ;
  assign y1814 = n5479 ;
  assign y1815 = ~n5484 ;
  assign y1816 = n5486 ;
  assign y1817 = n5495 ;
  assign y1818 = ~n5501 ;
  assign y1819 = ~n5504 ;
  assign y1820 = ~n5505 ;
  assign y1821 = ~n5509 ;
  assign y1822 = ~n5516 ;
  assign y1823 = n5518 ;
  assign y1824 = ~n5524 ;
  assign y1825 = ~n5532 ;
  assign y1826 = ~1'b0 ;
  assign y1827 = ~n5534 ;
  assign y1828 = n5535 ;
  assign y1829 = ~1'b0 ;
  assign y1830 = ~1'b0 ;
  assign y1831 = ~n5539 ;
  assign y1832 = ~n5544 ;
  assign y1833 = ~n5546 ;
  assign y1834 = n5552 ;
  assign y1835 = ~n5553 ;
  assign y1836 = ~n5556 ;
  assign y1837 = ~n5564 ;
  assign y1838 = ~1'b0 ;
  assign y1839 = ~n5569 ;
  assign y1840 = ~n5578 ;
  assign y1841 = ~1'b0 ;
  assign y1842 = ~n5591 ;
  assign y1843 = n5592 ;
  assign y1844 = n5599 ;
  assign y1845 = n5602 ;
  assign y1846 = ~n5603 ;
  assign y1847 = ~n5215 ;
  assign y1848 = n5606 ;
  assign y1849 = n5608 ;
  assign y1850 = ~n5611 ;
  assign y1851 = n5613 ;
  assign y1852 = n5077 ;
  assign y1853 = n5615 ;
  assign y1854 = ~n5616 ;
  assign y1855 = ~n5619 ;
  assign y1856 = ~1'b0 ;
  assign y1857 = ~1'b0 ;
  assign y1858 = n5622 ;
  assign y1859 = n5623 ;
  assign y1860 = n5625 ;
  assign y1861 = n5626 ;
  assign y1862 = n5632 ;
  assign y1863 = ~n5638 ;
  assign y1864 = n5641 ;
  assign y1865 = ~1'b0 ;
  assign y1866 = ~n5642 ;
  assign y1867 = ~n5643 ;
  assign y1868 = n5646 ;
  assign y1869 = ~1'b0 ;
  assign y1870 = n5649 ;
  assign y1871 = ~n5650 ;
  assign y1872 = ~n5659 ;
  assign y1873 = ~1'b0 ;
  assign y1874 = n5662 ;
  assign y1875 = ~n5666 ;
  assign y1876 = ~1'b0 ;
  assign y1877 = ~1'b0 ;
  assign y1878 = ~n5670 ;
  assign y1879 = n5674 ;
  assign y1880 = n5675 ;
  assign y1881 = ~n5676 ;
  assign y1882 = ~n5686 ;
  assign y1883 = n5689 ;
  assign y1884 = ~n5690 ;
  assign y1885 = ~n5697 ;
  assign y1886 = n5699 ;
  assign y1887 = 1'b0 ;
  assign y1888 = n5702 ;
  assign y1889 = ~1'b0 ;
  assign y1890 = ~n5704 ;
  assign y1891 = n5709 ;
  assign y1892 = ~n5721 ;
  assign y1893 = ~1'b0 ;
  assign y1894 = n5726 ;
  assign y1895 = ~n2386 ;
  assign y1896 = n5739 ;
  assign y1897 = ~n5742 ;
  assign y1898 = ~n5746 ;
  assign y1899 = ~n5748 ;
  assign y1900 = n3599 ;
  assign y1901 = n5749 ;
  assign y1902 = n5751 ;
  assign y1903 = n5752 ;
  assign y1904 = ~1'b0 ;
  assign y1905 = ~1'b0 ;
  assign y1906 = ~n5755 ;
  assign y1907 = n2892 ;
  assign y1908 = ~n5756 ;
  assign y1909 = n5770 ;
  assign y1910 = ~n5775 ;
  assign y1911 = ~1'b0 ;
  assign y1912 = ~n5784 ;
  assign y1913 = n5792 ;
  assign y1914 = n5793 ;
  assign y1915 = ~n5795 ;
  assign y1916 = ~n5796 ;
  assign y1917 = ~n5798 ;
  assign y1918 = ~n5806 ;
  assign y1919 = ~1'b0 ;
  assign y1920 = ~n5814 ;
  assign y1921 = ~1'b0 ;
  assign y1922 = n5817 ;
  assign y1923 = n5821 ;
  assign y1924 = ~n5823 ;
  assign y1925 = n5824 ;
  assign y1926 = n5825 ;
  assign y1927 = ~n5828 ;
  assign y1928 = ~1'b0 ;
  assign y1929 = ~1'b0 ;
  assign y1930 = ~1'b0 ;
  assign y1931 = ~n5832 ;
  assign y1932 = n5834 ;
  assign y1933 = ~1'b0 ;
  assign y1934 = n5836 ;
  assign y1935 = ~1'b0 ;
  assign y1936 = n5838 ;
  assign y1937 = ~n5841 ;
  assign y1938 = n5844 ;
  assign y1939 = ~n5848 ;
  assign y1940 = n5850 ;
  assign y1941 = n5856 ;
  assign y1942 = n5858 ;
  assign y1943 = ~n5859 ;
  assign y1944 = n5860 ;
  assign y1945 = ~n5865 ;
  assign y1946 = n5867 ;
  assign y1947 = n5869 ;
  assign y1948 = ~1'b0 ;
  assign y1949 = n5870 ;
  assign y1950 = n5873 ;
  assign y1951 = n5874 ;
  assign y1952 = n5877 ;
  assign y1953 = ~n5712 ;
  assign y1954 = ~n604 ;
  assign y1955 = ~n5878 ;
  assign y1956 = n5882 ;
  assign y1957 = ~n5886 ;
  assign y1958 = n5893 ;
  assign y1959 = ~n5894 ;
  assign y1960 = ~1'b0 ;
  assign y1961 = n5895 ;
  assign y1962 = ~n5898 ;
  assign y1963 = ~n5899 ;
  assign y1964 = n5901 ;
  assign y1965 = n5911 ;
  assign y1966 = n5912 ;
  assign y1967 = ~1'b0 ;
  assign y1968 = n5918 ;
  assign y1969 = n5922 ;
  assign y1970 = n5933 ;
  assign y1971 = ~n4528 ;
  assign y1972 = n5944 ;
  assign y1973 = n5945 ;
  assign y1974 = n5950 ;
  assign y1975 = ~n5952 ;
  assign y1976 = ~n5954 ;
  assign y1977 = n5958 ;
  assign y1978 = ~1'b0 ;
  assign y1979 = n5959 ;
  assign y1980 = ~n5963 ;
  assign y1981 = ~1'b0 ;
  assign y1982 = 1'b0 ;
  assign y1983 = n5969 ;
  assign y1984 = ~1'b0 ;
  assign y1985 = ~n5973 ;
  assign y1986 = x155 ;
  assign y1987 = n5976 ;
  assign y1988 = ~1'b0 ;
  assign y1989 = ~1'b0 ;
  assign y1990 = ~n5978 ;
  assign y1991 = 1'b0 ;
  assign y1992 = n5982 ;
  assign y1993 = n5989 ;
  assign y1994 = n5990 ;
  assign y1995 = ~1'b0 ;
  assign y1996 = ~n5993 ;
  assign y1997 = ~n5998 ;
  assign y1998 = n5999 ;
  assign y1999 = n6003 ;
  assign y2000 = ~n6008 ;
  assign y2001 = ~1'b0 ;
  assign y2002 = n6010 ;
  assign y2003 = n2573 ;
  assign y2004 = n6011 ;
  assign y2005 = n6012 ;
  assign y2006 = n6014 ;
  assign y2007 = ~1'b0 ;
  assign y2008 = ~n6019 ;
  assign y2009 = ~n6020 ;
  assign y2010 = n6021 ;
  assign y2011 = ~n6028 ;
  assign y2012 = ~1'b0 ;
  assign y2013 = ~1'b0 ;
  assign y2014 = ~n6029 ;
  assign y2015 = ~n6038 ;
  assign y2016 = ~n6039 ;
  assign y2017 = ~n6041 ;
  assign y2018 = ~n6045 ;
  assign y2019 = ~n6048 ;
  assign y2020 = ~n6052 ;
  assign y2021 = ~1'b0 ;
  assign y2022 = n6056 ;
  assign y2023 = ~1'b0 ;
  assign y2024 = ~n6058 ;
  assign y2025 = n6060 ;
  assign y2026 = ~n6066 ;
  assign y2027 = ~n6070 ;
  assign y2028 = ~n6074 ;
  assign y2029 = ~1'b0 ;
  assign y2030 = n6078 ;
  assign y2031 = n6080 ;
  assign y2032 = n6085 ;
  assign y2033 = n6091 ;
  assign y2034 = n6093 ;
  assign y2035 = ~1'b0 ;
  assign y2036 = n6094 ;
  assign y2037 = ~1'b0 ;
  assign y2038 = ~1'b0 ;
  assign y2039 = n6098 ;
  assign y2040 = ~n6099 ;
  assign y2041 = ~n6100 ;
  assign y2042 = ~1'b0 ;
  assign y2043 = n6107 ;
  assign y2044 = n6109 ;
  assign y2045 = ~n6110 ;
  assign y2046 = ~n6111 ;
  assign y2047 = ~n6118 ;
  assign y2048 = n6119 ;
  assign y2049 = ~n6124 ;
  assign y2050 = ~1'b0 ;
  assign y2051 = n6132 ;
  assign y2052 = ~n6135 ;
  assign y2053 = n6140 ;
  assign y2054 = n6153 ;
  assign y2055 = 1'b0 ;
  assign y2056 = n6154 ;
  assign y2057 = ~n6159 ;
  assign y2058 = ~n6164 ;
  assign y2059 = ~1'b0 ;
  assign y2060 = ~1'b0 ;
  assign y2061 = n6171 ;
  assign y2062 = n6172 ;
  assign y2063 = ~n6175 ;
  assign y2064 = n6185 ;
  assign y2065 = n6190 ;
  assign y2066 = ~1'b0 ;
  assign y2067 = ~n6195 ;
  assign y2068 = n6202 ;
  assign y2069 = ~n6204 ;
  assign y2070 = ~n6205 ;
  assign y2071 = n6213 ;
  assign y2072 = ~n6218 ;
  assign y2073 = ~n6221 ;
  assign y2074 = n6222 ;
  assign y2075 = ~1'b0 ;
  assign y2076 = ~n6223 ;
  assign y2077 = ~n6225 ;
  assign y2078 = ~n6227 ;
  assign y2079 = ~n6230 ;
  assign y2080 = ~1'b0 ;
  assign y2081 = ~n6231 ;
  assign y2082 = ~1'b0 ;
  assign y2083 = ~n6234 ;
  assign y2084 = ~n6239 ;
  assign y2085 = n6242 ;
  assign y2086 = ~n6244 ;
  assign y2087 = ~n6254 ;
  assign y2088 = n6255 ;
  assign y2089 = n6257 ;
  assign y2090 = n6261 ;
  assign y2091 = ~1'b0 ;
  assign y2092 = n6262 ;
  assign y2093 = n6267 ;
  assign y2094 = ~n6272 ;
  assign y2095 = n6276 ;
  assign y2096 = ~1'b0 ;
  assign y2097 = ~1'b0 ;
  assign y2098 = n6282 ;
  assign y2099 = n6284 ;
  assign y2100 = n6290 ;
  assign y2101 = ~1'b0 ;
  assign y2102 = n6291 ;
  assign y2103 = n6292 ;
  assign y2104 = n5475 ;
  assign y2105 = ~n6296 ;
  assign y2106 = ~n6297 ;
  assign y2107 = ~n6300 ;
  assign y2108 = ~n6307 ;
  assign y2109 = n6308 ;
  assign y2110 = ~1'b0 ;
  assign y2111 = ~n6313 ;
  assign y2112 = n6314 ;
  assign y2113 = n6315 ;
  assign y2114 = n6318 ;
  assign y2115 = ~n6324 ;
  assign y2116 = ~n6334 ;
  assign y2117 = n6335 ;
  assign y2118 = ~n6338 ;
  assign y2119 = ~n6347 ;
  assign y2120 = ~n6350 ;
  assign y2121 = ~n6353 ;
  assign y2122 = n6355 ;
  assign y2123 = ~1'b0 ;
  assign y2124 = n6356 ;
  assign y2125 = ~1'b0 ;
  assign y2126 = 1'b0 ;
  assign y2127 = ~n6357 ;
  assign y2128 = ~1'b0 ;
  assign y2129 = ~n6358 ;
  assign y2130 = n6362 ;
  assign y2131 = n6367 ;
  assign y2132 = ~n6374 ;
  assign y2133 = n6379 ;
  assign y2134 = ~n6384 ;
  assign y2135 = ~1'b0 ;
  assign y2136 = ~n6385 ;
  assign y2137 = ~n6386 ;
  assign y2138 = ~1'b0 ;
  assign y2139 = n6390 ;
  assign y2140 = ~n6392 ;
  assign y2141 = n6394 ;
  assign y2142 = ~n6395 ;
  assign y2143 = n6402 ;
  assign y2144 = ~n6406 ;
  assign y2145 = ~n6410 ;
  assign y2146 = n6414 ;
  assign y2147 = n6417 ;
  assign y2148 = ~1'b0 ;
  assign y2149 = ~n6424 ;
  assign y2150 = ~n6437 ;
  assign y2151 = ~n6438 ;
  assign y2152 = ~1'b0 ;
  assign y2153 = ~1'b0 ;
  assign y2154 = n6445 ;
  assign y2155 = n6446 ;
  assign y2156 = n6447 ;
  assign y2157 = ~n6458 ;
  assign y2158 = n3657 ;
  assign y2159 = ~1'b0 ;
  assign y2160 = n6459 ;
  assign y2161 = ~n6468 ;
  assign y2162 = ~n6474 ;
  assign y2163 = n6476 ;
  assign y2164 = ~1'b0 ;
  assign y2165 = ~n6477 ;
  assign y2166 = ~n6480 ;
  assign y2167 = n6485 ;
  assign y2168 = n6486 ;
  assign y2169 = n6489 ;
  assign y2170 = ~1'b0 ;
  assign y2171 = ~n6491 ;
  assign y2172 = ~n6497 ;
  assign y2173 = n6502 ;
  assign y2174 = ~n6504 ;
  assign y2175 = ~1'b0 ;
  assign y2176 = n6507 ;
  assign y2177 = ~1'b0 ;
  assign y2178 = n6509 ;
  assign y2179 = n6512 ;
  assign y2180 = ~1'b0 ;
  assign y2181 = ~1'b0 ;
  assign y2182 = ~1'b0 ;
  assign y2183 = n6516 ;
  assign y2184 = ~1'b0 ;
  assign y2185 = n6520 ;
  assign y2186 = ~n6526 ;
  assign y2187 = ~n6527 ;
  assign y2188 = ~n6531 ;
  assign y2189 = n6533 ;
  assign y2190 = n6536 ;
  assign y2191 = ~n6538 ;
  assign y2192 = n6547 ;
  assign y2193 = n6549 ;
  assign y2194 = n6551 ;
  assign y2195 = ~n6565 ;
  assign y2196 = ~n6567 ;
  assign y2197 = ~1'b0 ;
  assign y2198 = n6568 ;
  assign y2199 = ~n6569 ;
  assign y2200 = n6581 ;
  assign y2201 = ~n6587 ;
  assign y2202 = ~n6588 ;
  assign y2203 = ~n6589 ;
  assign y2204 = n2005 ;
  assign y2205 = n6591 ;
  assign y2206 = n6592 ;
  assign y2207 = n6594 ;
  assign y2208 = n6599 ;
  assign y2209 = n1265 ;
  assign y2210 = ~n6602 ;
  assign y2211 = n6606 ;
  assign y2212 = ~1'b0 ;
  assign y2213 = ~n6607 ;
  assign y2214 = n6608 ;
  assign y2215 = ~n6609 ;
  assign y2216 = n6618 ;
  assign y2217 = n6621 ;
  assign y2218 = ~n6624 ;
  assign y2219 = ~n6628 ;
  assign y2220 = ~n1487 ;
  assign y2221 = ~1'b0 ;
  assign y2222 = ~n6629 ;
  assign y2223 = ~n6632 ;
  assign y2224 = ~n6643 ;
  assign y2225 = ~n3802 ;
  assign y2226 = n6645 ;
  assign y2227 = ~1'b0 ;
  assign y2228 = n6656 ;
  assign y2229 = n6661 ;
  assign y2230 = n6662 ;
  assign y2231 = n6669 ;
  assign y2232 = ~1'b0 ;
  assign y2233 = ~n6670 ;
  assign y2234 = ~1'b0 ;
  assign y2235 = ~n6673 ;
  assign y2236 = n2317 ;
  assign y2237 = ~n6675 ;
  assign y2238 = ~n6678 ;
  assign y2239 = n6681 ;
  assign y2240 = ~n6683 ;
  assign y2241 = n6684 ;
  assign y2242 = n6692 ;
  assign y2243 = ~n6697 ;
  assign y2244 = ~n6698 ;
  assign y2245 = n6701 ;
  assign y2246 = n6703 ;
  assign y2247 = n6708 ;
  assign y2248 = n6710 ;
  assign y2249 = n6715 ;
  assign y2250 = n6716 ;
  assign y2251 = ~1'b0 ;
  assign y2252 = ~1'b0 ;
  assign y2253 = ~1'b0 ;
  assign y2254 = n6718 ;
  assign y2255 = ~n6719 ;
  assign y2256 = ~n6721 ;
  assign y2257 = n6722 ;
  assign y2258 = n6730 ;
  assign y2259 = n6732 ;
  assign y2260 = ~n6737 ;
  assign y2261 = ~n6740 ;
  assign y2262 = n6742 ;
  assign y2263 = n6744 ;
  assign y2264 = ~1'b0 ;
  assign y2265 = ~n6748 ;
  assign y2266 = n6750 ;
  assign y2267 = ~1'b0 ;
  assign y2268 = ~n6753 ;
  assign y2269 = n1527 ;
  assign y2270 = ~n6759 ;
  assign y2271 = ~n6761 ;
  assign y2272 = n6763 ;
  assign y2273 = n6738 ;
  assign y2274 = n6772 ;
  assign y2275 = ~n6773 ;
  assign y2276 = ~1'b0 ;
  assign y2277 = n6774 ;
  assign y2278 = ~1'b0 ;
  assign y2279 = ~1'b0 ;
  assign y2280 = ~n6781 ;
  assign y2281 = ~n6782 ;
  assign y2282 = ~1'b0 ;
  assign y2283 = ~n6789 ;
  assign y2284 = ~n6794 ;
  assign y2285 = ~n6799 ;
  assign y2286 = ~n6802 ;
  assign y2287 = ~1'b0 ;
  assign y2288 = ~1'b0 ;
  assign y2289 = n6805 ;
  assign y2290 = n6807 ;
  assign y2291 = n6811 ;
  assign y2292 = ~n6815 ;
  assign y2293 = ~1'b0 ;
  assign y2294 = ~1'b0 ;
  assign y2295 = ~n6816 ;
  assign y2296 = ~n6821 ;
  assign y2297 = n6829 ;
  assign y2298 = n6832 ;
  assign y2299 = ~n6842 ;
  assign y2300 = ~n6843 ;
  assign y2301 = ~n6855 ;
  assign y2302 = n6856 ;
  assign y2303 = ~n6858 ;
  assign y2304 = ~n6860 ;
  assign y2305 = n6870 ;
  assign y2306 = ~1'b0 ;
  assign y2307 = n6874 ;
  assign y2308 = ~n6875 ;
  assign y2309 = n4703 ;
  assign y2310 = ~n6876 ;
  assign y2311 = n6879 ;
  assign y2312 = ~n6886 ;
  assign y2313 = n6891 ;
  assign y2314 = ~n6899 ;
  assign y2315 = n6903 ;
  assign y2316 = ~n6910 ;
  assign y2317 = n6917 ;
  assign y2318 = ~n6922 ;
  assign y2319 = ~1'b0 ;
  assign y2320 = ~1'b0 ;
  assign y2321 = n6930 ;
  assign y2322 = ~n6931 ;
  assign y2323 = ~n6934 ;
  assign y2324 = n6938 ;
  assign y2325 = ~n6940 ;
  assign y2326 = n6950 ;
  assign y2327 = ~1'b0 ;
  assign y2328 = n6954 ;
  assign y2329 = ~n6962 ;
  assign y2330 = ~1'b0 ;
  assign y2331 = ~x143 ;
  assign y2332 = ~n6968 ;
  assign y2333 = n6973 ;
  assign y2334 = ~1'b0 ;
  assign y2335 = n6979 ;
  assign y2336 = ~1'b0 ;
  assign y2337 = ~n6980 ;
  assign y2338 = ~1'b0 ;
  assign y2339 = ~n6986 ;
  assign y2340 = ~n6988 ;
  assign y2341 = ~n6990 ;
  assign y2342 = ~1'b0 ;
  assign y2343 = ~n6991 ;
  assign y2344 = ~n6993 ;
  assign y2345 = n6995 ;
  assign y2346 = n6997 ;
  assign y2347 = n6998 ;
  assign y2348 = ~n7008 ;
  assign y2349 = ~1'b0 ;
  assign y2350 = ~n7009 ;
  assign y2351 = ~n7016 ;
  assign y2352 = n7027 ;
  assign y2353 = n7029 ;
  assign y2354 = n7030 ;
  assign y2355 = ~n7032 ;
  assign y2356 = ~n7034 ;
  assign y2357 = ~1'b0 ;
  assign y2358 = ~n7045 ;
  assign y2359 = ~n7049 ;
  assign y2360 = n7051 ;
  assign y2361 = ~1'b0 ;
  assign y2362 = n7063 ;
  assign y2363 = ~1'b0 ;
  assign y2364 = ~n7064 ;
  assign y2365 = ~1'b0 ;
  assign y2366 = ~n7071 ;
  assign y2367 = 1'b0 ;
  assign y2368 = ~n7072 ;
  assign y2369 = ~n7073 ;
  assign y2370 = ~1'b0 ;
  assign y2371 = n7076 ;
  assign y2372 = ~1'b0 ;
  assign y2373 = n7085 ;
  assign y2374 = n7086 ;
  assign y2375 = n7087 ;
  assign y2376 = n7094 ;
  assign y2377 = ~n7101 ;
  assign y2378 = n7102 ;
  assign y2379 = n7104 ;
  assign y2380 = n7106 ;
  assign y2381 = n7108 ;
  assign y2382 = n7110 ;
  assign y2383 = ~1'b0 ;
  assign y2384 = ~n7117 ;
  assign y2385 = n3640 ;
  assign y2386 = ~n7122 ;
  assign y2387 = ~1'b0 ;
  assign y2388 = 1'b0 ;
  assign y2389 = n7125 ;
  assign y2390 = ~1'b0 ;
  assign y2391 = n7130 ;
  assign y2392 = ~n7134 ;
  assign y2393 = n7135 ;
  assign y2394 = ~n7136 ;
  assign y2395 = n7138 ;
  assign y2396 = n7145 ;
  assign y2397 = ~1'b0 ;
  assign y2398 = ~n7149 ;
  assign y2399 = n7152 ;
  assign y2400 = n7154 ;
  assign y2401 = n7159 ;
  assign y2402 = ~n7160 ;
  assign y2403 = n7165 ;
  assign y2404 = ~n7167 ;
  assign y2405 = ~1'b0 ;
  assign y2406 = ~1'b0 ;
  assign y2407 = ~n7171 ;
  assign y2408 = n7174 ;
  assign y2409 = n7176 ;
  assign y2410 = ~1'b0 ;
  assign y2411 = ~n7181 ;
  assign y2412 = n7187 ;
  assign y2413 = n7190 ;
  assign y2414 = ~n7202 ;
  assign y2415 = ~1'b0 ;
  assign y2416 = ~n7209 ;
  assign y2417 = n7210 ;
  assign y2418 = ~1'b0 ;
  assign y2419 = n7212 ;
  assign y2420 = ~1'b0 ;
  assign y2421 = ~n7214 ;
  assign y2422 = n7223 ;
  assign y2423 = n7230 ;
  assign y2424 = ~n7234 ;
  assign y2425 = n7236 ;
  assign y2426 = ~n7237 ;
  assign y2427 = n7250 ;
  assign y2428 = n7259 ;
  assign y2429 = ~n7269 ;
  assign y2430 = n7276 ;
  assign y2431 = n7277 ;
  assign y2432 = ~n7280 ;
  assign y2433 = n7291 ;
  assign y2434 = ~1'b0 ;
  assign y2435 = ~1'b0 ;
  assign y2436 = n7295 ;
  assign y2437 = ~n7298 ;
  assign y2438 = ~n7299 ;
  assign y2439 = n7300 ;
  assign y2440 = n7303 ;
  assign y2441 = ~1'b0 ;
  assign y2442 = ~1'b0 ;
  assign y2443 = ~n7304 ;
  assign y2444 = ~n7307 ;
  assign y2445 = n7308 ;
  assign y2446 = ~n7309 ;
  assign y2447 = ~1'b0 ;
  assign y2448 = ~n7311 ;
  assign y2449 = ~n7316 ;
  assign y2450 = ~1'b0 ;
  assign y2451 = ~n7319 ;
  assign y2452 = ~n7324 ;
  assign y2453 = ~n7331 ;
  assign y2454 = ~n7334 ;
  assign y2455 = ~n7336 ;
  assign y2456 = n3512 ;
  assign y2457 = ~n7340 ;
  assign y2458 = ~n7344 ;
  assign y2459 = n7346 ;
  assign y2460 = ~n7348 ;
  assign y2461 = n7351 ;
  assign y2462 = n7356 ;
  assign y2463 = n7361 ;
  assign y2464 = n6296 ;
  assign y2465 = ~n7364 ;
  assign y2466 = ~n7368 ;
  assign y2467 = ~n7373 ;
  assign y2468 = ~1'b0 ;
  assign y2469 = ~n7375 ;
  assign y2470 = ~1'b0 ;
  assign y2471 = ~1'b0 ;
  assign y2472 = ~n7378 ;
  assign y2473 = n7380 ;
  assign y2474 = n7381 ;
  assign y2475 = n7384 ;
  assign y2476 = ~n7385 ;
  assign y2477 = ~1'b0 ;
  assign y2478 = n7393 ;
  assign y2479 = ~n7394 ;
  assign y2480 = ~n7402 ;
  assign y2481 = ~n7408 ;
  assign y2482 = ~n7410 ;
  assign y2483 = ~n7415 ;
  assign y2484 = n7416 ;
  assign y2485 = ~n7420 ;
  assign y2486 = ~n7422 ;
  assign y2487 = n7427 ;
  assign y2488 = ~n7431 ;
  assign y2489 = ~n7436 ;
  assign y2490 = n7439 ;
  assign y2491 = n7440 ;
  assign y2492 = ~n7444 ;
  assign y2493 = ~n7446 ;
  assign y2494 = n7450 ;
  assign y2495 = n7452 ;
  assign y2496 = n7454 ;
  assign y2497 = ~n7456 ;
  assign y2498 = n7460 ;
  assign y2499 = ~n7462 ;
  assign y2500 = n7464 ;
  assign y2501 = ~1'b0 ;
  assign y2502 = ~n7465 ;
  assign y2503 = n7466 ;
  assign y2504 = n7470 ;
  assign y2505 = ~n7472 ;
  assign y2506 = 1'b0 ;
  assign y2507 = n7473 ;
  assign y2508 = ~n3007 ;
  assign y2509 = n7475 ;
  assign y2510 = ~n7476 ;
  assign y2511 = n7481 ;
  assign y2512 = n7485 ;
  assign y2513 = n7492 ;
  assign y2514 = ~n7493 ;
  assign y2515 = ~n7494 ;
  assign y2516 = ~n7502 ;
  assign y2517 = ~1'b0 ;
  assign y2518 = n7504 ;
  assign y2519 = ~n7508 ;
  assign y2520 = ~1'b0 ;
  assign y2521 = n7509 ;
  assign y2522 = ~n1840 ;
  assign y2523 = n7515 ;
  assign y2524 = ~n7519 ;
  assign y2525 = ~n7522 ;
  assign y2526 = ~1'b0 ;
  assign y2527 = ~n7523 ;
  assign y2528 = ~n7526 ;
  assign y2529 = n7529 ;
  assign y2530 = n7534 ;
  assign y2531 = ~n7536 ;
  assign y2532 = ~n7538 ;
  assign y2533 = n7542 ;
  assign y2534 = ~n7545 ;
  assign y2535 = ~n7546 ;
  assign y2536 = n7552 ;
  assign y2537 = n7559 ;
  assign y2538 = ~n7571 ;
  assign y2539 = ~n7575 ;
  assign y2540 = ~n7576 ;
  assign y2541 = ~n7577 ;
  assign y2542 = n7578 ;
  assign y2543 = ~n7581 ;
  assign y2544 = n7585 ;
  assign y2545 = ~1'b0 ;
  assign y2546 = n7590 ;
  assign y2547 = ~n7594 ;
  assign y2548 = ~n7595 ;
  assign y2549 = ~1'b0 ;
  assign y2550 = ~1'b0 ;
  assign y2551 = n7599 ;
  assign y2552 = n7601 ;
  assign y2553 = ~n7602 ;
  assign y2554 = ~1'b0 ;
  assign y2555 = n7608 ;
  assign y2556 = ~n7618 ;
  assign y2557 = ~n7622 ;
  assign y2558 = ~1'b0 ;
  assign y2559 = ~n7628 ;
  assign y2560 = ~1'b0 ;
  assign y2561 = n7634 ;
  assign y2562 = n7635 ;
  assign y2563 = ~n7647 ;
  assign y2564 = n7660 ;
  assign y2565 = n6865 ;
  assign y2566 = n7664 ;
  assign y2567 = ~1'b0 ;
  assign y2568 = ~n7667 ;
  assign y2569 = n7668 ;
  assign y2570 = n7670 ;
  assign y2571 = ~n7687 ;
  assign y2572 = ~1'b0 ;
  assign y2573 = ~n7692 ;
  assign y2574 = n7693 ;
  assign y2575 = ~n7694 ;
  assign y2576 = ~n7695 ;
  assign y2577 = n7696 ;
  assign y2578 = ~n7699 ;
  assign y2579 = ~n7701 ;
  assign y2580 = ~n7702 ;
  assign y2581 = ~1'b0 ;
  assign y2582 = ~1'b0 ;
  assign y2583 = ~n7703 ;
  assign y2584 = ~n7705 ;
  assign y2585 = ~n7708 ;
  assign y2586 = ~1'b0 ;
  assign y2587 = ~n7711 ;
  assign y2588 = ~n7720 ;
  assign y2589 = ~n7723 ;
  assign y2590 = n7731 ;
  assign y2591 = n7737 ;
  assign y2592 = ~n7744 ;
  assign y2593 = n7746 ;
  assign y2594 = n7754 ;
  assign y2595 = n7757 ;
  assign y2596 = ~n7758 ;
  assign y2597 = ~n7761 ;
  assign y2598 = ~1'b0 ;
  assign y2599 = ~n7765 ;
  assign y2600 = ~n7766 ;
  assign y2601 = n7770 ;
  assign y2602 = n7773 ;
  assign y2603 = ~n7775 ;
  assign y2604 = n7776 ;
  assign y2605 = ~n7782 ;
  assign y2606 = ~n7785 ;
  assign y2607 = n7790 ;
  assign y2608 = ~n7792 ;
  assign y2609 = ~1'b0 ;
  assign y2610 = ~n7794 ;
  assign y2611 = ~n5752 ;
  assign y2612 = n7800 ;
  assign y2613 = n7802 ;
  assign y2614 = n7808 ;
  assign y2615 = ~n7811 ;
  assign y2616 = n7815 ;
  assign y2617 = ~n7819 ;
  assign y2618 = ~n7829 ;
  assign y2619 = n7830 ;
  assign y2620 = ~n7833 ;
  assign y2621 = ~1'b0 ;
  assign y2622 = n7838 ;
  assign y2623 = ~1'b0 ;
  assign y2624 = ~n7842 ;
  assign y2625 = ~n7843 ;
  assign y2626 = ~n7845 ;
  assign y2627 = n7846 ;
  assign y2628 = ~n7852 ;
  assign y2629 = ~n7855 ;
  assign y2630 = n7857 ;
  assign y2631 = n7858 ;
  assign y2632 = ~1'b0 ;
  assign y2633 = ~1'b0 ;
  assign y2634 = n7862 ;
  assign y2635 = ~n7867 ;
  assign y2636 = ~n7869 ;
  assign y2637 = ~n7875 ;
  assign y2638 = n7877 ;
  assign y2639 = ~n7878 ;
  assign y2640 = ~n7881 ;
  assign y2641 = n7886 ;
  assign y2642 = ~n7888 ;
  assign y2643 = n7893 ;
  assign y2644 = 1'b0 ;
  assign y2645 = ~n7905 ;
  assign y2646 = ~n7906 ;
  assign y2647 = ~n7912 ;
  assign y2648 = ~n7923 ;
  assign y2649 = ~n7925 ;
  assign y2650 = ~n7927 ;
  assign y2651 = ~n7930 ;
  assign y2652 = ~1'b0 ;
  assign y2653 = n7938 ;
  assign y2654 = ~1'b0 ;
  assign y2655 = n7944 ;
  assign y2656 = n7957 ;
  assign y2657 = n7958 ;
  assign y2658 = ~n7959 ;
  assign y2659 = n7973 ;
  assign y2660 = ~n7974 ;
  assign y2661 = n7979 ;
  assign y2662 = ~n7982 ;
  assign y2663 = ~n7986 ;
  assign y2664 = ~n7988 ;
  assign y2665 = n7990 ;
  assign y2666 = ~n7992 ;
  assign y2667 = n8001 ;
  assign y2668 = n8003 ;
  assign y2669 = n8008 ;
  assign y2670 = n8009 ;
  assign y2671 = ~n8018 ;
  assign y2672 = n8023 ;
  assign y2673 = n8027 ;
  assign y2674 = n8032 ;
  assign y2675 = ~1'b0 ;
  assign y2676 = n8034 ;
  assign y2677 = ~n8042 ;
  assign y2678 = ~1'b0 ;
  assign y2679 = ~n8045 ;
  assign y2680 = ~n8048 ;
  assign y2681 = n8049 ;
  assign y2682 = n8054 ;
  assign y2683 = ~1'b0 ;
  assign y2684 = ~n8061 ;
  assign y2685 = ~1'b0 ;
  assign y2686 = n8063 ;
  assign y2687 = n8065 ;
  assign y2688 = ~1'b0 ;
  assign y2689 = ~1'b0 ;
  assign y2690 = ~n8066 ;
  assign y2691 = n8068 ;
  assign y2692 = ~1'b0 ;
  assign y2693 = ~n8071 ;
  assign y2694 = ~n8077 ;
  assign y2695 = n8078 ;
  assign y2696 = n8079 ;
  assign y2697 = ~n8085 ;
  assign y2698 = n8086 ;
  assign y2699 = n8089 ;
  assign y2700 = n8091 ;
  assign y2701 = n8092 ;
  assign y2702 = ~n8093 ;
  assign y2703 = n8094 ;
  assign y2704 = ~n8096 ;
  assign y2705 = n8099 ;
  assign y2706 = ~n8101 ;
  assign y2707 = ~n8108 ;
  assign y2708 = ~n8111 ;
  assign y2709 = n8117 ;
  assign y2710 = ~n8119 ;
  assign y2711 = ~n8120 ;
  assign y2712 = n8121 ;
  assign y2713 = ~n8134 ;
  assign y2714 = n8142 ;
  assign y2715 = n8144 ;
  assign y2716 = ~n8146 ;
  assign y2717 = ~1'b0 ;
  assign y2718 = ~n2645 ;
  assign y2719 = ~n8148 ;
  assign y2720 = n8159 ;
  assign y2721 = n8161 ;
  assign y2722 = n8169 ;
  assign y2723 = ~n8170 ;
  assign y2724 = n8173 ;
  assign y2725 = ~n8177 ;
  assign y2726 = ~1'b0 ;
  assign y2727 = n8186 ;
  assign y2728 = ~1'b0 ;
  assign y2729 = ~n8189 ;
  assign y2730 = n8196 ;
  assign y2731 = ~1'b0 ;
  assign y2732 = n8197 ;
  assign y2733 = n8200 ;
  assign y2734 = ~n8227 ;
  assign y2735 = ~1'b0 ;
  assign y2736 = n8234 ;
  assign y2737 = n8235 ;
  assign y2738 = ~1'b0 ;
  assign y2739 = ~1'b0 ;
  assign y2740 = ~n8237 ;
  assign y2741 = ~n8243 ;
  assign y2742 = n8246 ;
  assign y2743 = ~n8247 ;
  assign y2744 = ~n8249 ;
  assign y2745 = ~1'b0 ;
  assign y2746 = ~n8250 ;
  assign y2747 = n8252 ;
  assign y2748 = n5038 ;
  assign y2749 = ~1'b0 ;
  assign y2750 = n8255 ;
  assign y2751 = ~1'b0 ;
  assign y2752 = n8256 ;
  assign y2753 = n8257 ;
  assign y2754 = ~n8259 ;
  assign y2755 = ~1'b0 ;
  assign y2756 = n8272 ;
  assign y2757 = ~n8273 ;
  assign y2758 = ~1'b0 ;
  assign y2759 = ~n8275 ;
  assign y2760 = n8276 ;
  assign y2761 = n8280 ;
  assign y2762 = ~n8282 ;
  assign y2763 = n8284 ;
  assign y2764 = ~n8287 ;
  assign y2765 = ~1'b0 ;
  assign y2766 = n8288 ;
  assign y2767 = n8290 ;
  assign y2768 = n8294 ;
  assign y2769 = ~n8295 ;
  assign y2770 = ~n8301 ;
  assign y2771 = ~n8305 ;
  assign y2772 = ~1'b0 ;
  assign y2773 = n8306 ;
  assign y2774 = n4411 ;
  assign y2775 = n8310 ;
  assign y2776 = ~n8312 ;
  assign y2777 = ~1'b0 ;
  assign y2778 = n8318 ;
  assign y2779 = ~1'b0 ;
  assign y2780 = ~n8321 ;
  assign y2781 = n8323 ;
  assign y2782 = ~n8325 ;
  assign y2783 = ~1'b0 ;
  assign y2784 = n8331 ;
  assign y2785 = n8339 ;
  assign y2786 = n8341 ;
  assign y2787 = n8343 ;
  assign y2788 = n8348 ;
  assign y2789 = ~n8350 ;
  assign y2790 = ~n8351 ;
  assign y2791 = n8358 ;
  assign y2792 = n8360 ;
  assign y2793 = ~n8361 ;
  assign y2794 = ~n8362 ;
  assign y2795 = n8364 ;
  assign y2796 = n8367 ;
  assign y2797 = ~n8370 ;
  assign y2798 = ~n8380 ;
  assign y2799 = ~n8389 ;
  assign y2800 = ~n8390 ;
  assign y2801 = ~1'b0 ;
  assign y2802 = ~n8393 ;
  assign y2803 = ~1'b0 ;
  assign y2804 = ~n8394 ;
  assign y2805 = ~n8396 ;
  assign y2806 = n3688 ;
  assign y2807 = ~n8401 ;
  assign y2808 = ~n8412 ;
  assign y2809 = n6403 ;
  assign y2810 = ~n3097 ;
  assign y2811 = ~n8430 ;
  assign y2812 = ~1'b0 ;
  assign y2813 = ~1'b0 ;
  assign y2814 = n8435 ;
  assign y2815 = n8439 ;
  assign y2816 = ~n8448 ;
  assign y2817 = ~n8449 ;
  assign y2818 = ~1'b0 ;
  assign y2819 = n8451 ;
  assign y2820 = ~n8456 ;
  assign y2821 = ~n8460 ;
  assign y2822 = ~1'b0 ;
  assign y2823 = ~1'b0 ;
  assign y2824 = n8461 ;
  assign y2825 = ~n8467 ;
  assign y2826 = ~1'b0 ;
  assign y2827 = n8468 ;
  assign y2828 = ~n8469 ;
  assign y2829 = n8474 ;
  assign y2830 = ~n8475 ;
  assign y2831 = n8477 ;
  assign y2832 = ~n8480 ;
  assign y2833 = n8481 ;
  assign y2834 = ~n8484 ;
  assign y2835 = ~1'b0 ;
  assign y2836 = ~1'b0 ;
  assign y2837 = ~n8486 ;
  assign y2838 = ~1'b0 ;
  assign y2839 = ~n8491 ;
  assign y2840 = n8498 ;
  assign y2841 = ~n8504 ;
  assign y2842 = n8507 ;
  assign y2843 = ~1'b0 ;
  assign y2844 = ~n8511 ;
  assign y2845 = ~1'b0 ;
  assign y2846 = ~n4007 ;
  assign y2847 = ~n8520 ;
  assign y2848 = n8521 ;
  assign y2849 = n8524 ;
  assign y2850 = ~n8525 ;
  assign y2851 = n8527 ;
  assign y2852 = n8532 ;
  assign y2853 = n8534 ;
  assign y2854 = n8540 ;
  assign y2855 = ~1'b0 ;
  assign y2856 = n8543 ;
  assign y2857 = ~1'b0 ;
  assign y2858 = n8544 ;
  assign y2859 = ~1'b0 ;
  assign y2860 = ~1'b0 ;
  assign y2861 = ~n8545 ;
  assign y2862 = n1206 ;
  assign y2863 = n7772 ;
  assign y2864 = ~1'b0 ;
  assign y2865 = ~n8552 ;
  assign y2866 = n8559 ;
  assign y2867 = ~n8563 ;
  assign y2868 = ~1'b0 ;
  assign y2869 = ~1'b0 ;
  assign y2870 = n8567 ;
  assign y2871 = n8571 ;
  assign y2872 = ~n8573 ;
  assign y2873 = n8578 ;
  assign y2874 = ~n8584 ;
  assign y2875 = n8585 ;
  assign y2876 = ~n8591 ;
  assign y2877 = n8601 ;
  assign y2878 = ~1'b0 ;
  assign y2879 = ~1'b0 ;
  assign y2880 = ~1'b0 ;
  assign y2881 = n8613 ;
  assign y2882 = ~1'b0 ;
  assign y2883 = n1975 ;
  assign y2884 = ~n8620 ;
  assign y2885 = n8624 ;
  assign y2886 = ~1'b0 ;
  assign y2887 = n8629 ;
  assign y2888 = ~n8631 ;
  assign y2889 = ~n8634 ;
  assign y2890 = n8639 ;
  assign y2891 = ~n8640 ;
  assign y2892 = ~n8642 ;
  assign y2893 = ~n2282 ;
  assign y2894 = ~n8646 ;
  assign y2895 = n8651 ;
  assign y2896 = ~n8652 ;
  assign y2897 = ~n8653 ;
  assign y2898 = n8658 ;
  assign y2899 = ~n8659 ;
  assign y2900 = ~n8664 ;
  assign y2901 = ~1'b0 ;
  assign y2902 = n8669 ;
  assign y2903 = n8674 ;
  assign y2904 = n8678 ;
  assign y2905 = n8681 ;
  assign y2906 = n8683 ;
  assign y2907 = n8684 ;
  assign y2908 = ~n8685 ;
  assign y2909 = ~1'b0 ;
  assign y2910 = ~n8687 ;
  assign y2911 = ~n8688 ;
  assign y2912 = ~n8697 ;
  assign y2913 = ~1'b0 ;
  assign y2914 = ~1'b0 ;
  assign y2915 = n8705 ;
  assign y2916 = ~n8721 ;
  assign y2917 = n8724 ;
  assign y2918 = ~n8726 ;
  assign y2919 = ~n8727 ;
  assign y2920 = n2764 ;
  assign y2921 = ~1'b0 ;
  assign y2922 = ~n8731 ;
  assign y2923 = ~n8732 ;
  assign y2924 = n8733 ;
  assign y2925 = n8734 ;
  assign y2926 = ~n8736 ;
  assign y2927 = ~1'b0 ;
  assign y2928 = ~1'b0 ;
  assign y2929 = ~n8743 ;
  assign y2930 = ~n8748 ;
  assign y2931 = ~n8749 ;
  assign y2932 = ~1'b0 ;
  assign y2933 = ~n8750 ;
  assign y2934 = n8751 ;
  assign y2935 = n8753 ;
  assign y2936 = ~n8754 ;
  assign y2937 = n8756 ;
  assign y2938 = n8757 ;
  assign y2939 = ~n8758 ;
  assign y2940 = ~1'b0 ;
  assign y2941 = n8764 ;
  assign y2942 = ~n8771 ;
  assign y2943 = ~1'b0 ;
  assign y2944 = n8774 ;
  assign y2945 = ~n8776 ;
  assign y2946 = n8782 ;
  assign y2947 = ~n8783 ;
  assign y2948 = ~1'b0 ;
  assign y2949 = n8786 ;
  assign y2950 = n8788 ;
  assign y2951 = n8791 ;
  assign y2952 = n8792 ;
  assign y2953 = n8807 ;
  assign y2954 = ~1'b0 ;
  assign y2955 = ~n8812 ;
  assign y2956 = ~n2169 ;
  assign y2957 = n8816 ;
  assign y2958 = n8826 ;
  assign y2959 = n8827 ;
  assign y2960 = ~n8829 ;
  assign y2961 = ~n8830 ;
  assign y2962 = n8831 ;
  assign y2963 = ~n8833 ;
  assign y2964 = ~1'b0 ;
  assign y2965 = ~1'b0 ;
  assign y2966 = ~1'b0 ;
  assign y2967 = ~n8841 ;
  assign y2968 = ~n8843 ;
  assign y2969 = ~n8848 ;
  assign y2970 = ~n8853 ;
  assign y2971 = n8859 ;
  assign y2972 = ~n8863 ;
  assign y2973 = ~1'b0 ;
  assign y2974 = n8865 ;
  assign y2975 = ~n8867 ;
  assign y2976 = 1'b0 ;
  assign y2977 = ~n8869 ;
  assign y2978 = n8870 ;
  assign y2979 = ~1'b0 ;
  assign y2980 = ~1'b0 ;
  assign y2981 = ~1'b0 ;
  assign y2982 = n8873 ;
  assign y2983 = n8876 ;
  assign y2984 = ~n8878 ;
  assign y2985 = ~1'b0 ;
  assign y2986 = ~n8882 ;
  assign y2987 = n8887 ;
  assign y2988 = ~n8888 ;
  assign y2989 = 1'b0 ;
  assign y2990 = ~n8890 ;
  assign y2991 = n8893 ;
  assign y2992 = n8895 ;
  assign y2993 = ~n8897 ;
  assign y2994 = ~1'b0 ;
  assign y2995 = n8899 ;
  assign y2996 = ~n8904 ;
  assign y2997 = ~1'b0 ;
  assign y2998 = n8914 ;
  assign y2999 = ~n8918 ;
  assign y3000 = n8920 ;
  assign y3001 = ~n8923 ;
  assign y3002 = ~1'b0 ;
  assign y3003 = n8927 ;
  assign y3004 = ~n8930 ;
  assign y3005 = ~1'b0 ;
  assign y3006 = ~1'b0 ;
  assign y3007 = ~n8939 ;
  assign y3008 = n8941 ;
  assign y3009 = ~1'b0 ;
  assign y3010 = n8944 ;
  assign y3011 = ~n8945 ;
  assign y3012 = ~1'b0 ;
  assign y3013 = ~1'b0 ;
  assign y3014 = ~n4893 ;
  assign y3015 = ~n8946 ;
  assign y3016 = ~n8948 ;
  assign y3017 = n8967 ;
  assign y3018 = n8970 ;
  assign y3019 = ~1'b0 ;
  assign y3020 = n8973 ;
  assign y3021 = ~n8976 ;
  assign y3022 = ~n8979 ;
  assign y3023 = n8983 ;
  assign y3024 = n8989 ;
  assign y3025 = ~n8993 ;
  assign y3026 = n8995 ;
  assign y3027 = n9004 ;
  assign y3028 = ~n9012 ;
  assign y3029 = n9018 ;
  assign y3030 = n4332 ;
  assign y3031 = ~n9020 ;
  assign y3032 = n9024 ;
  assign y3033 = ~n9028 ;
  assign y3034 = ~n9035 ;
  assign y3035 = ~n9040 ;
  assign y3036 = n9041 ;
  assign y3037 = n9044 ;
  assign y3038 = ~n5153 ;
  assign y3039 = ~n9045 ;
  assign y3040 = ~n9047 ;
  assign y3041 = n9052 ;
  assign y3042 = ~n9056 ;
  assign y3043 = n9058 ;
  assign y3044 = ~1'b0 ;
  assign y3045 = n9059 ;
  assign y3046 = ~n9062 ;
  assign y3047 = n9063 ;
  assign y3048 = ~1'b0 ;
  assign y3049 = ~n9067 ;
  assign y3050 = ~1'b0 ;
  assign y3051 = ~n9070 ;
  assign y3052 = ~n9071 ;
  assign y3053 = ~n9074 ;
  assign y3054 = n3322 ;
  assign y3055 = ~n9075 ;
  assign y3056 = n9077 ;
  assign y3057 = n9078 ;
  assign y3058 = ~n9080 ;
  assign y3059 = ~n9081 ;
  assign y3060 = ~n9084 ;
  assign y3061 = ~n9092 ;
  assign y3062 = n9096 ;
  assign y3063 = n9100 ;
  assign y3064 = ~n9106 ;
  assign y3065 = n9108 ;
  assign y3066 = ~n9109 ;
  assign y3067 = n9110 ;
  assign y3068 = n9113 ;
  assign y3069 = ~1'b0 ;
  assign y3070 = ~n9117 ;
  assign y3071 = ~n9118 ;
  assign y3072 = ~n9120 ;
  assign y3073 = ~n6272 ;
  assign y3074 = ~1'b0 ;
  assign y3075 = n9121 ;
  assign y3076 = n9122 ;
  assign y3077 = ~n9123 ;
  assign y3078 = ~1'b0 ;
  assign y3079 = n9131 ;
  assign y3080 = ~n9132 ;
  assign y3081 = n9136 ;
  assign y3082 = ~1'b0 ;
  assign y3083 = ~n9143 ;
  assign y3084 = ~n9146 ;
  assign y3085 = n9148 ;
  assign y3086 = 1'b0 ;
  assign y3087 = n9155 ;
  assign y3088 = ~1'b0 ;
  assign y3089 = ~n9158 ;
  assign y3090 = ~1'b0 ;
  assign y3091 = n9159 ;
  assign y3092 = ~1'b0 ;
  assign y3093 = n3919 ;
  assign y3094 = ~n9160 ;
  assign y3095 = ~1'b0 ;
  assign y3096 = ~1'b0 ;
  assign y3097 = ~n9167 ;
  assign y3098 = n9170 ;
  assign y3099 = n9176 ;
  assign y3100 = ~n9180 ;
  assign y3101 = n9181 ;
  assign y3102 = ~n9185 ;
  assign y3103 = n9192 ;
  assign y3104 = ~n9196 ;
  assign y3105 = n9197 ;
  assign y3106 = ~n9210 ;
  assign y3107 = n9213 ;
  assign y3108 = ~n9215 ;
  assign y3109 = ~n9221 ;
  assign y3110 = n9224 ;
  assign y3111 = ~n9233 ;
  assign y3112 = ~n9236 ;
  assign y3113 = ~n9241 ;
  assign y3114 = ~1'b0 ;
  assign y3115 = ~n9245 ;
  assign y3116 = ~1'b0 ;
  assign y3117 = ~n9246 ;
  assign y3118 = ~1'b0 ;
  assign y3119 = n9248 ;
  assign y3120 = ~n9249 ;
  assign y3121 = n9258 ;
  assign y3122 = n9260 ;
  assign y3123 = ~n9261 ;
  assign y3124 = 1'b0 ;
  assign y3125 = ~n9264 ;
  assign y3126 = ~n9265 ;
  assign y3127 = n9268 ;
  assign y3128 = n9269 ;
  assign y3129 = n9271 ;
  assign y3130 = ~1'b0 ;
  assign y3131 = n9272 ;
  assign y3132 = n9274 ;
  assign y3133 = ~n9277 ;
  assign y3134 = n9278 ;
  assign y3135 = ~n9279 ;
  assign y3136 = n9280 ;
  assign y3137 = ~n9281 ;
  assign y3138 = ~n9286 ;
  assign y3139 = ~n9287 ;
  assign y3140 = ~1'b0 ;
  assign y3141 = ~1'b0 ;
  assign y3142 = ~n9290 ;
  assign y3143 = ~n6310 ;
  assign y3144 = ~1'b0 ;
  assign y3145 = n5859 ;
  assign y3146 = ~n9294 ;
  assign y3147 = ~n9300 ;
  assign y3148 = n9306 ;
  assign y3149 = ~n9308 ;
  assign y3150 = ~1'b0 ;
  assign y3151 = ~n9309 ;
  assign y3152 = n9316 ;
  assign y3153 = n9320 ;
  assign y3154 = ~n9325 ;
  assign y3155 = ~1'b0 ;
  assign y3156 = ~1'b0 ;
  assign y3157 = ~n9327 ;
  assign y3158 = n9330 ;
  assign y3159 = ~n9335 ;
  assign y3160 = ~n9338 ;
  assign y3161 = n9343 ;
  assign y3162 = ~1'b0 ;
  assign y3163 = n9344 ;
  assign y3164 = ~1'b0 ;
  assign y3165 = n9345 ;
  assign y3166 = n9349 ;
  assign y3167 = ~n9351 ;
  assign y3168 = n9354 ;
  assign y3169 = n9357 ;
  assign y3170 = ~1'b0 ;
  assign y3171 = ~n9359 ;
  assign y3172 = n9361 ;
  assign y3173 = ~1'b0 ;
  assign y3174 = ~n9371 ;
  assign y3175 = ~n9373 ;
  assign y3176 = ~n9375 ;
  assign y3177 = ~1'b0 ;
  assign y3178 = ~1'b0 ;
  assign y3179 = ~1'b0 ;
  assign y3180 = n9376 ;
  assign y3181 = ~n9377 ;
  assign y3182 = ~n9382 ;
  assign y3183 = ~n9386 ;
  assign y3184 = ~1'b0 ;
  assign y3185 = ~1'b0 ;
  assign y3186 = ~n9351 ;
  assign y3187 = n9392 ;
  assign y3188 = n9394 ;
  assign y3189 = ~n9396 ;
  assign y3190 = n9405 ;
  assign y3191 = n3237 ;
  assign y3192 = ~n9412 ;
  assign y3193 = ~n9413 ;
  assign y3194 = ~n9414 ;
  assign y3195 = n9419 ;
  assign y3196 = n9420 ;
  assign y3197 = n9423 ;
  assign y3198 = n9436 ;
  assign y3199 = ~n2427 ;
  assign y3200 = n9443 ;
  assign y3201 = ~n9444 ;
  assign y3202 = ~n9445 ;
  assign y3203 = ~n9451 ;
  assign y3204 = x123 ;
  assign y3205 = ~n9453 ;
  assign y3206 = n9459 ;
  assign y3207 = ~1'b0 ;
  assign y3208 = ~1'b0 ;
  assign y3209 = ~1'b0 ;
  assign y3210 = ~n9460 ;
  assign y3211 = n9463 ;
  assign y3212 = n9464 ;
  assign y3213 = ~n9472 ;
  assign y3214 = n9473 ;
  assign y3215 = ~n9474 ;
  assign y3216 = n9477 ;
  assign y3217 = ~n9488 ;
  assign y3218 = ~1'b0 ;
  assign y3219 = ~n9491 ;
  assign y3220 = ~n9492 ;
  assign y3221 = n1476 ;
  assign y3222 = n797 ;
  assign y3223 = ~n9496 ;
  assign y3224 = ~n9500 ;
  assign y3225 = ~n9501 ;
  assign y3226 = n9504 ;
  assign y3227 = ~n9506 ;
  assign y3228 = ~n9507 ;
  assign y3229 = ~1'b0 ;
  assign y3230 = ~n9510 ;
  assign y3231 = ~1'b0 ;
  assign y3232 = ~n9511 ;
  assign y3233 = ~n9512 ;
  assign y3234 = ~n9513 ;
  assign y3235 = ~1'b0 ;
  assign y3236 = ~1'b0 ;
  assign y3237 = ~n9517 ;
  assign y3238 = n9520 ;
  assign y3239 = n9522 ;
  assign y3240 = n9525 ;
  assign y3241 = ~n9527 ;
  assign y3242 = n9530 ;
  assign y3243 = ~1'b0 ;
  assign y3244 = ~n9534 ;
  assign y3245 = ~n9547 ;
  assign y3246 = ~1'b0 ;
  assign y3247 = ~n9554 ;
  assign y3248 = n9555 ;
  assign y3249 = ~n9558 ;
  assign y3250 = ~1'b0 ;
  assign y3251 = ~1'b0 ;
  assign y3252 = ~n9562 ;
  assign y3253 = ~1'b0 ;
  assign y3254 = ~n9563 ;
  assign y3255 = ~n9566 ;
  assign y3256 = ~n9567 ;
  assign y3257 = ~n9568 ;
  assign y3258 = n9571 ;
  assign y3259 = ~n9576 ;
  assign y3260 = ~1'b0 ;
  assign y3261 = ~1'b0 ;
  assign y3262 = ~n9577 ;
  assign y3263 = ~n9578 ;
  assign y3264 = ~n9590 ;
  assign y3265 = n9592 ;
  assign y3266 = ~n9593 ;
  assign y3267 = ~1'b0 ;
  assign y3268 = ~1'b0 ;
  assign y3269 = ~n9594 ;
  assign y3270 = n9599 ;
  assign y3271 = ~1'b0 ;
  assign y3272 = ~n9606 ;
  assign y3273 = n9607 ;
  assign y3274 = ~1'b0 ;
  assign y3275 = ~n9608 ;
  assign y3276 = n9612 ;
  assign y3277 = n9615 ;
  assign y3278 = n9617 ;
  assign y3279 = ~n9626 ;
  assign y3280 = ~1'b0 ;
  assign y3281 = ~1'b0 ;
  assign y3282 = ~n9630 ;
  assign y3283 = n9631 ;
  assign y3284 = ~1'b0 ;
  assign y3285 = n9640 ;
  assign y3286 = ~n9649 ;
  assign y3287 = n9650 ;
  assign y3288 = ~1'b0 ;
  assign y3289 = ~n9653 ;
  assign y3290 = n9654 ;
  assign y3291 = ~n9658 ;
  assign y3292 = ~1'b0 ;
  assign y3293 = n9660 ;
  assign y3294 = ~n9672 ;
  assign y3295 = ~n8983 ;
  assign y3296 = ~n9673 ;
  assign y3297 = ~n9675 ;
  assign y3298 = n9677 ;
  assign y3299 = ~n9692 ;
  assign y3300 = ~1'b0 ;
  assign y3301 = ~n9695 ;
  assign y3302 = ~n9698 ;
  assign y3303 = n9705 ;
  assign y3304 = ~n9712 ;
  assign y3305 = ~n9716 ;
  assign y3306 = n9717 ;
  assign y3307 = ~n9724 ;
  assign y3308 = n9731 ;
  assign y3309 = n9734 ;
  assign y3310 = ~n9735 ;
  assign y3311 = n9738 ;
  assign y3312 = ~1'b0 ;
  assign y3313 = ~n9741 ;
  assign y3314 = ~n9742 ;
  assign y3315 = ~1'b0 ;
  assign y3316 = ~1'b0 ;
  assign y3317 = n9746 ;
  assign y3318 = n9747 ;
  assign y3319 = n9749 ;
  assign y3320 = n9751 ;
  assign y3321 = ~n9756 ;
  assign y3322 = ~n9762 ;
  assign y3323 = ~n816 ;
  assign y3324 = n9767 ;
  assign y3325 = n9768 ;
  assign y3326 = n9779 ;
  assign y3327 = n9782 ;
  assign y3328 = ~1'b0 ;
  assign y3329 = ~n9783 ;
  assign y3330 = ~n9785 ;
  assign y3331 = n9787 ;
  assign y3332 = ~n9788 ;
  assign y3333 = n9792 ;
  assign y3334 = ~n9797 ;
  assign y3335 = ~n9809 ;
  assign y3336 = ~n9826 ;
  assign y3337 = ~n9827 ;
  assign y3338 = ~n9828 ;
  assign y3339 = n9444 ;
  assign y3340 = 1'b0 ;
  assign y3341 = ~n9829 ;
  assign y3342 = ~n9830 ;
  assign y3343 = ~1'b0 ;
  assign y3344 = ~n9834 ;
  assign y3345 = ~1'b0 ;
  assign y3346 = ~n9839 ;
  assign y3347 = n9842 ;
  assign y3348 = n9843 ;
  assign y3349 = ~1'b0 ;
  assign y3350 = n7580 ;
  assign y3351 = n9844 ;
  assign y3352 = n9845 ;
  assign y3353 = ~n9846 ;
  assign y3354 = n9849 ;
  assign y3355 = ~n9850 ;
  assign y3356 = ~n9852 ;
  assign y3357 = ~1'b0 ;
  assign y3358 = ~n9855 ;
  assign y3359 = ~1'b0 ;
  assign y3360 = ~1'b0 ;
  assign y3361 = ~n9858 ;
  assign y3362 = ~n9860 ;
  assign y3363 = n9864 ;
  assign y3364 = n9871 ;
  assign y3365 = n9872 ;
  assign y3366 = ~1'b0 ;
  assign y3367 = n9880 ;
  assign y3368 = n9886 ;
  assign y3369 = n9887 ;
  assign y3370 = n9889 ;
  assign y3371 = ~n9890 ;
  assign y3372 = ~1'b0 ;
  assign y3373 = ~n9891 ;
  assign y3374 = ~n9894 ;
  assign y3375 = ~1'b0 ;
  assign y3376 = ~n9896 ;
  assign y3377 = ~n9899 ;
  assign y3378 = n9902 ;
  assign y3379 = ~1'b0 ;
  assign y3380 = ~n5196 ;
  assign y3381 = n9904 ;
  assign y3382 = ~1'b0 ;
  assign y3383 = ~n9910 ;
  assign y3384 = ~1'b0 ;
  assign y3385 = n9914 ;
  assign y3386 = n9918 ;
  assign y3387 = ~n9921 ;
  assign y3388 = n9928 ;
  assign y3389 = ~1'b0 ;
  assign y3390 = ~1'b0 ;
  assign y3391 = 1'b0 ;
  assign y3392 = ~1'b0 ;
  assign y3393 = ~n9932 ;
  assign y3394 = n9936 ;
  assign y3395 = n9939 ;
  assign y3396 = n9947 ;
  assign y3397 = n9955 ;
  assign y3398 = n9960 ;
  assign y3399 = ~n9961 ;
  assign y3400 = n9964 ;
  assign y3401 = ~n9978 ;
  assign y3402 = ~n9980 ;
  assign y3403 = ~n9981 ;
  assign y3404 = n9982 ;
  assign y3405 = n9983 ;
  assign y3406 = ~n9987 ;
  assign y3407 = n9990 ;
  assign y3408 = n9991 ;
  assign y3409 = ~n9992 ;
  assign y3410 = ~n9993 ;
  assign y3411 = ~1'b0 ;
  assign y3412 = n9995 ;
  assign y3413 = ~n9996 ;
  assign y3414 = ~1'b0 ;
  assign y3415 = n10000 ;
  assign y3416 = n10001 ;
  assign y3417 = ~n10020 ;
  assign y3418 = n10023 ;
  assign y3419 = ~n10026 ;
  assign y3420 = ~n10039 ;
  assign y3421 = ~1'b0 ;
  assign y3422 = ~n10042 ;
  assign y3423 = ~n10046 ;
  assign y3424 = ~n10058 ;
  assign y3425 = ~1'b0 ;
  assign y3426 = ~1'b0 ;
  assign y3427 = ~n10059 ;
  assign y3428 = n10061 ;
  assign y3429 = n10064 ;
  assign y3430 = n10065 ;
  assign y3431 = ~n10068 ;
  assign y3432 = ~1'b0 ;
  assign y3433 = n10070 ;
  assign y3434 = n10071 ;
  assign y3435 = ~1'b0 ;
  assign y3436 = ~n10072 ;
  assign y3437 = ~n10078 ;
  assign y3438 = ~1'b0 ;
  assign y3439 = ~1'b0 ;
  assign y3440 = n10082 ;
  assign y3441 = ~n10088 ;
  assign y3442 = ~n10090 ;
  assign y3443 = ~n10091 ;
  assign y3444 = n10093 ;
  assign y3445 = ~n10101 ;
  assign y3446 = 1'b0 ;
  assign y3447 = ~1'b0 ;
  assign y3448 = ~n5500 ;
  assign y3449 = ~n10104 ;
  assign y3450 = n10113 ;
  assign y3451 = ~n10121 ;
  assign y3452 = n10124 ;
  assign y3453 = n10125 ;
  assign y3454 = ~1'b0 ;
  assign y3455 = ~1'b0 ;
  assign y3456 = ~1'b0 ;
  assign y3457 = n10130 ;
  assign y3458 = ~n10135 ;
  assign y3459 = ~n10137 ;
  assign y3460 = ~n10139 ;
  assign y3461 = n10147 ;
  assign y3462 = ~1'b0 ;
  assign y3463 = n10150 ;
  assign y3464 = ~n10152 ;
  assign y3465 = ~n10153 ;
  assign y3466 = n10154 ;
  assign y3467 = ~1'b0 ;
  assign y3468 = ~1'b0 ;
  assign y3469 = n10155 ;
  assign y3470 = ~n10157 ;
  assign y3471 = n10164 ;
  assign y3472 = ~n10167 ;
  assign y3473 = ~n10168 ;
  assign y3474 = ~1'b0 ;
  assign y3475 = n10170 ;
  assign y3476 = ~n10174 ;
  assign y3477 = n10178 ;
  assign y3478 = ~n10183 ;
  assign y3479 = n10190 ;
  assign y3480 = n10193 ;
  assign y3481 = ~n10196 ;
  assign y3482 = ~n10199 ;
  assign y3483 = ~1'b0 ;
  assign y3484 = ~n10200 ;
  assign y3485 = ~1'b0 ;
  assign y3486 = ~1'b0 ;
  assign y3487 = ~n10218 ;
  assign y3488 = ~n10221 ;
  assign y3489 = n10224 ;
  assign y3490 = ~1'b0 ;
  assign y3491 = ~n10232 ;
  assign y3492 = ~n10234 ;
  assign y3493 = ~1'b0 ;
  assign y3494 = ~n10239 ;
  assign y3495 = ~n10242 ;
  assign y3496 = n10245 ;
  assign y3497 = n571 ;
  assign y3498 = n6915 ;
  assign y3499 = ~n10247 ;
  assign y3500 = ~1'b0 ;
  assign y3501 = ~n10248 ;
  assign y3502 = n10250 ;
  assign y3503 = ~n10255 ;
  assign y3504 = ~n10257 ;
  assign y3505 = ~1'b0 ;
  assign y3506 = n10258 ;
  assign y3507 = ~n10260 ;
  assign y3508 = ~n10261 ;
  assign y3509 = ~1'b0 ;
  assign y3510 = n10266 ;
  assign y3511 = n10275 ;
  assign y3512 = n10286 ;
  assign y3513 = n10294 ;
  assign y3514 = n10299 ;
  assign y3515 = ~n10301 ;
  assign y3516 = ~n1227 ;
  assign y3517 = n10304 ;
  assign y3518 = n10309 ;
  assign y3519 = n10310 ;
  assign y3520 = ~n10313 ;
  assign y3521 = n5975 ;
  assign y3522 = n8858 ;
  assign y3523 = ~1'b0 ;
  assign y3524 = ~n10315 ;
  assign y3525 = n10318 ;
  assign y3526 = ~n10320 ;
  assign y3527 = n10322 ;
  assign y3528 = n10330 ;
  assign y3529 = ~1'b0 ;
  assign y3530 = n10332 ;
  assign y3531 = ~1'b0 ;
  assign y3532 = ~n10337 ;
  assign y3533 = ~n10342 ;
  assign y3534 = ~n10345 ;
  assign y3535 = ~1'b0 ;
  assign y3536 = ~n10353 ;
  assign y3537 = ~n10355 ;
  assign y3538 = n10357 ;
  assign y3539 = n10360 ;
  assign y3540 = n10363 ;
  assign y3541 = ~1'b0 ;
  assign y3542 = ~1'b0 ;
  assign y3543 = ~n10366 ;
  assign y3544 = n10371 ;
  assign y3545 = 1'b0 ;
  assign y3546 = n10377 ;
  assign y3547 = n10378 ;
  assign y3548 = ~1'b0 ;
  assign y3549 = n10381 ;
  assign y3550 = ~n10385 ;
  assign y3551 = n10391 ;
  assign y3552 = n2083 ;
  assign y3553 = n10408 ;
  assign y3554 = ~n10411 ;
  assign y3555 = n10414 ;
  assign y3556 = ~n10417 ;
  assign y3557 = ~n10425 ;
  assign y3558 = 1'b0 ;
  assign y3559 = n10426 ;
  assign y3560 = n10437 ;
  assign y3561 = n10442 ;
  assign y3562 = ~n10457 ;
  assign y3563 = n10463 ;
  assign y3564 = n10472 ;
  assign y3565 = ~n10473 ;
  assign y3566 = ~1'b0 ;
  assign y3567 = n10476 ;
  assign y3568 = n10477 ;
  assign y3569 = ~n10478 ;
  assign y3570 = n10480 ;
  assign y3571 = ~n10484 ;
  assign y3572 = n10492 ;
  assign y3573 = n10497 ;
  assign y3574 = ~n10498 ;
  assign y3575 = ~1'b0 ;
  assign y3576 = ~n10504 ;
  assign y3577 = ~n10505 ;
  assign y3578 = n10506 ;
  assign y3579 = n10507 ;
  assign y3580 = n10510 ;
  assign y3581 = n10512 ;
  assign y3582 = n10515 ;
  assign y3583 = ~n4395 ;
  assign y3584 = n10516 ;
  assign y3585 = ~1'b0 ;
  assign y3586 = n10518 ;
  assign y3587 = ~n10519 ;
  assign y3588 = ~n10525 ;
  assign y3589 = ~n10528 ;
  assign y3590 = n10532 ;
  assign y3591 = ~n10535 ;
  assign y3592 = n10544 ;
  assign y3593 = n10545 ;
  assign y3594 = ~1'b0 ;
  assign y3595 = ~1'b0 ;
  assign y3596 = ~n10553 ;
  assign y3597 = n10558 ;
  assign y3598 = ~n10561 ;
  assign y3599 = ~1'b0 ;
  assign y3600 = n10562 ;
  assign y3601 = n10564 ;
  assign y3602 = n10565 ;
  assign y3603 = n10568 ;
  assign y3604 = n10570 ;
  assign y3605 = ~n10571 ;
  assign y3606 = ~1'b0 ;
  assign y3607 = n10575 ;
  assign y3608 = n10583 ;
  assign y3609 = ~1'b0 ;
  assign y3610 = ~1'b0 ;
  assign y3611 = n10584 ;
  assign y3612 = ~n10595 ;
  assign y3613 = n10600 ;
  assign y3614 = ~n10601 ;
  assign y3615 = ~n10604 ;
  assign y3616 = ~1'b0 ;
  assign y3617 = ~n10611 ;
  assign y3618 = ~n10616 ;
  assign y3619 = n10619 ;
  assign y3620 = ~1'b0 ;
  assign y3621 = ~n10622 ;
  assign y3622 = ~n10624 ;
  assign y3623 = ~n10636 ;
  assign y3624 = ~n10637 ;
  assign y3625 = ~1'b0 ;
  assign y3626 = n10644 ;
  assign y3627 = 1'b0 ;
  assign y3628 = ~n10645 ;
  assign y3629 = ~1'b0 ;
  assign y3630 = n10650 ;
  assign y3631 = ~1'b0 ;
  assign y3632 = n10655 ;
  assign y3633 = ~1'b0 ;
  assign y3634 = ~1'b0 ;
  assign y3635 = n10658 ;
  assign y3636 = ~n10659 ;
  assign y3637 = ~n10661 ;
  assign y3638 = n10670 ;
  assign y3639 = ~n10671 ;
  assign y3640 = ~n10672 ;
  assign y3641 = n10675 ;
  assign y3642 = ~n10682 ;
  assign y3643 = ~1'b0 ;
  assign y3644 = n10683 ;
  assign y3645 = n10685 ;
  assign y3646 = n10686 ;
  assign y3647 = n10692 ;
  assign y3648 = n10694 ;
  assign y3649 = ~n10703 ;
  assign y3650 = ~n10704 ;
  assign y3651 = ~n4045 ;
  assign y3652 = ~n10706 ;
  assign y3653 = n10707 ;
  assign y3654 = ~n10710 ;
  assign y3655 = ~n10712 ;
  assign y3656 = n10714 ;
  assign y3657 = ~n10716 ;
  assign y3658 = ~n10718 ;
  assign y3659 = n10722 ;
  assign y3660 = n10723 ;
  assign y3661 = n10726 ;
  assign y3662 = ~n10727 ;
  assign y3663 = ~n10729 ;
  assign y3664 = 1'b0 ;
  assign y3665 = ~n10731 ;
  assign y3666 = ~1'b0 ;
  assign y3667 = ~n10735 ;
  assign y3668 = n10736 ;
  assign y3669 = ~n9276 ;
  assign y3670 = ~n10737 ;
  assign y3671 = n10738 ;
  assign y3672 = n10740 ;
  assign y3673 = n1999 ;
  assign y3674 = n1885 ;
  assign y3675 = ~n10741 ;
  assign y3676 = ~n10742 ;
  assign y3677 = ~n10743 ;
  assign y3678 = n10747 ;
  assign y3679 = n10752 ;
  assign y3680 = ~1'b0 ;
  assign y3681 = n10759 ;
  assign y3682 = n8572 ;
  assign y3683 = ~n10765 ;
  assign y3684 = n4546 ;
  assign y3685 = n10768 ;
  assign y3686 = ~1'b0 ;
  assign y3687 = n10774 ;
  assign y3688 = ~n10776 ;
  assign y3689 = ~1'b0 ;
  assign y3690 = ~n10787 ;
  assign y3691 = n10799 ;
  assign y3692 = n10812 ;
  assign y3693 = ~n10818 ;
  assign y3694 = ~n10821 ;
  assign y3695 = ~n10822 ;
  assign y3696 = n7457 ;
  assign y3697 = ~1'b0 ;
  assign y3698 = n10825 ;
  assign y3699 = ~1'b0 ;
  assign y3700 = ~1'b0 ;
  assign y3701 = ~n10826 ;
  assign y3702 = ~n10832 ;
  assign y3703 = ~1'b0 ;
  assign y3704 = ~1'b0 ;
  assign y3705 = n10833 ;
  assign y3706 = ~n10834 ;
  assign y3707 = ~n10835 ;
  assign y3708 = n10838 ;
  assign y3709 = ~1'b0 ;
  assign y3710 = ~1'b0 ;
  assign y3711 = ~1'b0 ;
  assign y3712 = ~n10840 ;
  assign y3713 = ~n10841 ;
  assign y3714 = ~n10844 ;
  assign y3715 = ~1'b0 ;
  assign y3716 = n10845 ;
  assign y3717 = ~1'b0 ;
  assign y3718 = ~n10852 ;
  assign y3719 = n10853 ;
  assign y3720 = n10857 ;
  assign y3721 = ~n10859 ;
  assign y3722 = n10861 ;
  assign y3723 = ~n10866 ;
  assign y3724 = ~1'b0 ;
  assign y3725 = n10871 ;
  assign y3726 = ~n10881 ;
  assign y3727 = n10882 ;
  assign y3728 = ~1'b0 ;
  assign y3729 = n10885 ;
  assign y3730 = n10886 ;
  assign y3731 = ~1'b0 ;
  assign y3732 = ~1'b0 ;
  assign y3733 = ~n10894 ;
  assign y3734 = ~n10895 ;
  assign y3735 = n10899 ;
  assign y3736 = ~n10910 ;
  assign y3737 = ~1'b0 ;
  assign y3738 = n10913 ;
  assign y3739 = n10915 ;
  assign y3740 = n10918 ;
  assign y3741 = ~n10919 ;
  assign y3742 = ~n10921 ;
  assign y3743 = n10924 ;
  assign y3744 = n10926 ;
  assign y3745 = n10930 ;
  assign y3746 = ~n10931 ;
  assign y3747 = n10936 ;
  assign y3748 = ~n10938 ;
  assign y3749 = n10939 ;
  assign y3750 = ~1'b0 ;
  assign y3751 = ~n10943 ;
  assign y3752 = ~n10945 ;
  assign y3753 = ~n10948 ;
  assign y3754 = ~1'b0 ;
  assign y3755 = ~n10952 ;
  assign y3756 = ~n10957 ;
  assign y3757 = 1'b0 ;
  assign y3758 = n10966 ;
  assign y3759 = ~n10971 ;
  assign y3760 = ~n1613 ;
  assign y3761 = ~n10973 ;
  assign y3762 = ~n10974 ;
  assign y3763 = ~n10980 ;
  assign y3764 = ~n10986 ;
  assign y3765 = n10988 ;
  assign y3766 = n10994 ;
  assign y3767 = ~n10996 ;
  assign y3768 = ~n11000 ;
  assign y3769 = ~n11008 ;
  assign y3770 = n11012 ;
  assign y3771 = n11017 ;
  assign y3772 = ~1'b0 ;
  assign y3773 = ~n11019 ;
  assign y3774 = n11023 ;
  assign y3775 = ~1'b0 ;
  assign y3776 = n11025 ;
  assign y3777 = ~n11028 ;
  assign y3778 = n11029 ;
  assign y3779 = ~n11033 ;
  assign y3780 = n11037 ;
  assign y3781 = ~n11041 ;
  assign y3782 = ~1'b0 ;
  assign y3783 = n11050 ;
  assign y3784 = ~n11052 ;
  assign y3785 = n1688 ;
  assign y3786 = ~n1733 ;
  assign y3787 = n11055 ;
  assign y3788 = n11062 ;
  assign y3789 = n11064 ;
  assign y3790 = ~n11073 ;
  assign y3791 = ~1'b0 ;
  assign y3792 = 1'b0 ;
  assign y3793 = ~1'b0 ;
  assign y3794 = ~1'b0 ;
  assign y3795 = ~n11074 ;
  assign y3796 = ~n11082 ;
  assign y3797 = ~n11084 ;
  assign y3798 = n11087 ;
  assign y3799 = n11089 ;
  assign y3800 = n11091 ;
  assign y3801 = n11097 ;
  assign y3802 = n11103 ;
  assign y3803 = ~1'b0 ;
  assign y3804 = ~n11109 ;
  assign y3805 = n2367 ;
  assign y3806 = ~n11111 ;
  assign y3807 = n11114 ;
  assign y3808 = ~n11115 ;
  assign y3809 = ~n11121 ;
  assign y3810 = ~n11122 ;
  assign y3811 = ~1'b0 ;
  assign y3812 = ~1'b0 ;
  assign y3813 = n11131 ;
  assign y3814 = ~n11133 ;
  assign y3815 = ~1'b0 ;
  assign y3816 = ~1'b0 ;
  assign y3817 = ~n11137 ;
  assign y3818 = ~1'b0 ;
  assign y3819 = n11139 ;
  assign y3820 = ~1'b0 ;
  assign y3821 = ~1'b0 ;
  assign y3822 = n11142 ;
  assign y3823 = n11143 ;
  assign y3824 = ~n11146 ;
  assign y3825 = ~n11157 ;
  assign y3826 = ~1'b0 ;
  assign y3827 = ~1'b0 ;
  assign y3828 = ~1'b0 ;
  assign y3829 = n11159 ;
  assign y3830 = n11161 ;
  assign y3831 = n11162 ;
  assign y3832 = ~n11167 ;
  assign y3833 = n11169 ;
  assign y3834 = n11171 ;
  assign y3835 = ~n11174 ;
  assign y3836 = n11176 ;
  assign y3837 = ~n11180 ;
  assign y3838 = n11182 ;
  assign y3839 = ~n11189 ;
  assign y3840 = ~1'b0 ;
  assign y3841 = ~1'b0 ;
  assign y3842 = ~1'b0 ;
  assign y3843 = ~n11190 ;
  assign y3844 = ~n11191 ;
  assign y3845 = ~n11200 ;
  assign y3846 = n11206 ;
  assign y3847 = n11215 ;
  assign y3848 = ~n11223 ;
  assign y3849 = n11227 ;
  assign y3850 = ~n11230 ;
  assign y3851 = n11231 ;
  assign y3852 = ~1'b0 ;
  assign y3853 = ~1'b0 ;
  assign y3854 = n11236 ;
  assign y3855 = n11243 ;
  assign y3856 = ~n11245 ;
  assign y3857 = n8193 ;
  assign y3858 = ~n11248 ;
  assign y3859 = n11249 ;
  assign y3860 = n11254 ;
  assign y3861 = ~n11256 ;
  assign y3862 = n11258 ;
  assign y3863 = ~1'b0 ;
  assign y3864 = ~1'b0 ;
  assign y3865 = ~1'b0 ;
  assign y3866 = ~1'b0 ;
  assign y3867 = n11262 ;
  assign y3868 = ~1'b0 ;
  assign y3869 = ~1'b0 ;
  assign y3870 = ~1'b0 ;
  assign y3871 = ~n11264 ;
  assign y3872 = ~n11281 ;
  assign y3873 = ~n11284 ;
  assign y3874 = ~n11286 ;
  assign y3875 = n11290 ;
  assign y3876 = ~n11291 ;
  assign y3877 = ~1'b0 ;
  assign y3878 = ~n11296 ;
  assign y3879 = n11298 ;
  assign y3880 = ~n11303 ;
  assign y3881 = n11304 ;
  assign y3882 = n11308 ;
  assign y3883 = ~n11310 ;
  assign y3884 = ~n11311 ;
  assign y3885 = ~1'b0 ;
  assign y3886 = ~n11312 ;
  assign y3887 = n11317 ;
  assign y3888 = ~n11324 ;
  assign y3889 = n11325 ;
  assign y3890 = ~n11327 ;
  assign y3891 = ~n11328 ;
  assign y3892 = n8991 ;
  assign y3893 = ~n11329 ;
  assign y3894 = ~1'b0 ;
  assign y3895 = ~n11336 ;
  assign y3896 = n11338 ;
  assign y3897 = n11344 ;
  assign y3898 = ~n11348 ;
  assign y3899 = n11355 ;
  assign y3900 = ~n11357 ;
  assign y3901 = ~n11359 ;
  assign y3902 = ~n11361 ;
  assign y3903 = ~n11362 ;
  assign y3904 = ~n11367 ;
  assign y3905 = ~1'b0 ;
  assign y3906 = n11371 ;
  assign y3907 = ~1'b0 ;
  assign y3908 = ~n11373 ;
  assign y3909 = ~n11375 ;
  assign y3910 = ~n11379 ;
  assign y3911 = ~n11387 ;
  assign y3912 = n11390 ;
  assign y3913 = ~n11391 ;
  assign y3914 = ~1'b0 ;
  assign y3915 = ~n11392 ;
  assign y3916 = n11397 ;
  assign y3917 = n11401 ;
  assign y3918 = ~n11406 ;
  assign y3919 = ~1'b0 ;
  assign y3920 = ~n11409 ;
  assign y3921 = ~1'b0 ;
  assign y3922 = ~n11420 ;
  assign y3923 = ~1'b0 ;
  assign y3924 = 1'b0 ;
  assign y3925 = ~n11425 ;
  assign y3926 = n11429 ;
  assign y3927 = ~n11431 ;
  assign y3928 = ~n11440 ;
  assign y3929 = ~n11442 ;
  assign y3930 = n11444 ;
  assign y3931 = n11448 ;
  assign y3932 = n11452 ;
  assign y3933 = ~1'b0 ;
  assign y3934 = ~n11454 ;
  assign y3935 = ~n11456 ;
  assign y3936 = n11457 ;
  assign y3937 = ~n11465 ;
  assign y3938 = ~1'b0 ;
  assign y3939 = n11466 ;
  assign y3940 = ~n11477 ;
  assign y3941 = ~1'b0 ;
  assign y3942 = ~n11479 ;
  assign y3943 = ~n11480 ;
  assign y3944 = ~n11483 ;
  assign y3945 = ~n11486 ;
  assign y3946 = ~1'b0 ;
  assign y3947 = n11490 ;
  assign y3948 = n11491 ;
  assign y3949 = n11493 ;
  assign y3950 = n11499 ;
  assign y3951 = ~n11501 ;
  assign y3952 = ~1'b0 ;
  assign y3953 = ~n11504 ;
  assign y3954 = 1'b0 ;
  assign y3955 = ~n11505 ;
  assign y3956 = ~n11506 ;
  assign y3957 = n11510 ;
  assign y3958 = n2992 ;
  assign y3959 = ~n11519 ;
  assign y3960 = n11523 ;
  assign y3961 = n11529 ;
  assign y3962 = ~n11534 ;
  assign y3963 = n11536 ;
  assign y3964 = n11540 ;
  assign y3965 = ~n11549 ;
  assign y3966 = ~n11552 ;
  assign y3967 = n11555 ;
  assign y3968 = n4558 ;
  assign y3969 = n11562 ;
  assign y3970 = ~n11566 ;
  assign y3971 = n11570 ;
  assign y3972 = n11572 ;
  assign y3973 = ~n11575 ;
  assign y3974 = ~n11577 ;
  assign y3975 = ~1'b0 ;
  assign y3976 = n11578 ;
  assign y3977 = n11585 ;
  assign y3978 = ~n11586 ;
  assign y3979 = ~1'b0 ;
  assign y3980 = 1'b0 ;
  assign y3981 = ~n11588 ;
  assign y3982 = ~1'b0 ;
  assign y3983 = ~1'b0 ;
  assign y3984 = n11592 ;
  assign y3985 = ~1'b0 ;
  assign y3986 = ~n11601 ;
  assign y3987 = ~n11603 ;
  assign y3988 = n11604 ;
  assign y3989 = n11608 ;
  assign y3990 = ~1'b0 ;
  assign y3991 = ~1'b0 ;
  assign y3992 = ~n11610 ;
  assign y3993 = n11611 ;
  assign y3994 = ~n11612 ;
  assign y3995 = n11617 ;
  assign y3996 = ~n11618 ;
  assign y3997 = n11619 ;
  assign y3998 = ~n11624 ;
  assign y3999 = n11627 ;
  assign y4000 = ~n11631 ;
  assign y4001 = ~1'b0 ;
  assign y4002 = ~1'b0 ;
  assign y4003 = n11636 ;
  assign y4004 = 1'b0 ;
  assign y4005 = n11648 ;
  assign y4006 = ~n11649 ;
  assign y4007 = n11652 ;
  assign y4008 = ~n11655 ;
  assign y4009 = ~1'b0 ;
  assign y4010 = ~1'b0 ;
  assign y4011 = ~n11658 ;
  assign y4012 = ~n11666 ;
  assign y4013 = n11668 ;
  assign y4014 = n11669 ;
  assign y4015 = n11679 ;
  assign y4016 = ~n11682 ;
  assign y4017 = ~n11689 ;
  assign y4018 = ~1'b0 ;
  assign y4019 = n11692 ;
  assign y4020 = n11694 ;
  assign y4021 = ~n11697 ;
  assign y4022 = ~1'b0 ;
  assign y4023 = ~1'b0 ;
  assign y4024 = ~n11706 ;
  assign y4025 = ~n11710 ;
  assign y4026 = ~n11712 ;
  assign y4027 = n11716 ;
  assign y4028 = n11721 ;
  assign y4029 = n11722 ;
  assign y4030 = n11729 ;
  assign y4031 = ~n11731 ;
  assign y4032 = n11733 ;
  assign y4033 = n11736 ;
  assign y4034 = ~n11743 ;
  assign y4035 = ~1'b0 ;
  assign y4036 = n11744 ;
  assign y4037 = ~1'b0 ;
  assign y4038 = ~1'b0 ;
  assign y4039 = ~n11749 ;
  assign y4040 = ~1'b0 ;
  assign y4041 = ~n11756 ;
  assign y4042 = ~n11760 ;
  assign y4043 = ~1'b0 ;
  assign y4044 = ~n11766 ;
  assign y4045 = n11769 ;
  assign y4046 = ~n11775 ;
  assign y4047 = ~n11786 ;
  assign y4048 = ~n11788 ;
  assign y4049 = ~n11792 ;
  assign y4050 = ~n11793 ;
  assign y4051 = ~n11795 ;
  assign y4052 = ~1'b0 ;
  assign y4053 = ~1'b0 ;
  assign y4054 = ~n11801 ;
  assign y4055 = n11804 ;
  assign y4056 = n11808 ;
  assign y4057 = ~1'b0 ;
  assign y4058 = ~n11814 ;
  assign y4059 = ~1'b0 ;
  assign y4060 = n11819 ;
  assign y4061 = ~n11823 ;
  assign y4062 = n11835 ;
  assign y4063 = ~n11840 ;
  assign y4064 = n11841 ;
  assign y4065 = n11842 ;
  assign y4066 = n11846 ;
  assign y4067 = n11849 ;
  assign y4068 = ~n11854 ;
  assign y4069 = ~n11855 ;
  assign y4070 = ~n11856 ;
  assign y4071 = ~n11857 ;
  assign y4072 = ~n11858 ;
  assign y4073 = ~n11865 ;
  assign y4074 = ~1'b0 ;
  assign y4075 = ~n11866 ;
  assign y4076 = ~1'b0 ;
  assign y4077 = n11867 ;
  assign y4078 = ~1'b0 ;
  assign y4079 = ~1'b0 ;
  assign y4080 = n11877 ;
  assign y4081 = n11878 ;
  assign y4082 = ~1'b0 ;
  assign y4083 = ~n11884 ;
  assign y4084 = n11886 ;
  assign y4085 = x120 ;
  assign y4086 = n11890 ;
  assign y4087 = ~1'b0 ;
  assign y4088 = n11892 ;
  assign y4089 = n11898 ;
  assign y4090 = n11900 ;
  assign y4091 = ~1'b0 ;
  assign y4092 = ~n11907 ;
  assign y4093 = ~n11913 ;
  assign y4094 = n11915 ;
  assign y4095 = ~n11918 ;
  assign y4096 = n11921 ;
  assign y4097 = ~n11923 ;
  assign y4098 = n11926 ;
  assign y4099 = ~1'b0 ;
  assign y4100 = ~1'b0 ;
  assign y4101 = ~1'b0 ;
  assign y4102 = n11934 ;
  assign y4103 = ~n3866 ;
  assign y4104 = n11938 ;
  assign y4105 = ~1'b0 ;
  assign y4106 = n11941 ;
  assign y4107 = ~1'b0 ;
  assign y4108 = n11944 ;
  assign y4109 = ~1'b0 ;
  assign y4110 = ~1'b0 ;
  assign y4111 = ~n11949 ;
  assign y4112 = n11951 ;
  assign y4113 = n11954 ;
  assign y4114 = ~1'b0 ;
  assign y4115 = n11955 ;
  assign y4116 = ~1'b0 ;
  assign y4117 = ~n9308 ;
  assign y4118 = n11957 ;
  assign y4119 = n11959 ;
  assign y4120 = ~n11963 ;
  assign y4121 = ~n11968 ;
  assign y4122 = ~n11973 ;
  assign y4123 = n11974 ;
  assign y4124 = ~n11976 ;
  assign y4125 = n11984 ;
  assign y4126 = n11987 ;
  assign y4127 = n11990 ;
  assign y4128 = n12003 ;
  assign y4129 = ~1'b0 ;
  assign y4130 = ~n12008 ;
  assign y4131 = n12010 ;
  assign y4132 = n8533 ;
  assign y4133 = ~n12012 ;
  assign y4134 = ~n12022 ;
  assign y4135 = ~n12023 ;
  assign y4136 = n12024 ;
  assign y4137 = n12032 ;
  assign y4138 = ~1'b0 ;
  assign y4139 = ~n12040 ;
  assign y4140 = n12041 ;
  assign y4141 = ~n12042 ;
  assign y4142 = ~n12045 ;
  assign y4143 = ~n12049 ;
  assign y4144 = ~1'b0 ;
  assign y4145 = n12051 ;
  assign y4146 = ~n12053 ;
  assign y4147 = n12059 ;
  assign y4148 = ~n12064 ;
  assign y4149 = ~1'b0 ;
  assign y4150 = n12065 ;
  assign y4151 = ~n12076 ;
  assign y4152 = ~n12082 ;
  assign y4153 = ~n12087 ;
  assign y4154 = ~n12091 ;
  assign y4155 = ~n12097 ;
  assign y4156 = n12100 ;
  assign y4157 = ~n12104 ;
  assign y4158 = ~n12107 ;
  assign y4159 = ~n12111 ;
  assign y4160 = n12112 ;
  assign y4161 = n12113 ;
  assign y4162 = ~1'b0 ;
  assign y4163 = n12114 ;
  assign y4164 = n12121 ;
  assign y4165 = n12123 ;
  assign y4166 = ~1'b0 ;
  assign y4167 = n12127 ;
  assign y4168 = ~1'b0 ;
  assign y4169 = ~n12131 ;
  assign y4170 = ~n12137 ;
  assign y4171 = ~n12144 ;
  assign y4172 = ~n12149 ;
  assign y4173 = ~n12151 ;
  assign y4174 = n12152 ;
  assign y4175 = n12167 ;
  assign y4176 = n12168 ;
  assign y4177 = n12169 ;
  assign y4178 = ~1'b0 ;
  assign y4179 = ~n6846 ;
  assign y4180 = ~1'b0 ;
  assign y4181 = ~n12171 ;
  assign y4182 = ~n12172 ;
  assign y4183 = ~n12181 ;
  assign y4184 = ~n12186 ;
  assign y4185 = ~n12190 ;
  assign y4186 = n12191 ;
  assign y4187 = ~n11437 ;
  assign y4188 = n12200 ;
  assign y4189 = ~n12202 ;
  assign y4190 = ~n1108 ;
  assign y4191 = ~n12207 ;
  assign y4192 = ~n12209 ;
  assign y4193 = n12210 ;
  assign y4194 = ~n12215 ;
  assign y4195 = ~1'b0 ;
  assign y4196 = ~1'b0 ;
  assign y4197 = ~1'b0 ;
  assign y4198 = ~n12218 ;
  assign y4199 = ~n12227 ;
  assign y4200 = n12228 ;
  assign y4201 = n12230 ;
  assign y4202 = ~n12231 ;
  assign y4203 = n12233 ;
  assign y4204 = n12240 ;
  assign y4205 = ~n12242 ;
  assign y4206 = ~1'b0 ;
  assign y4207 = ~1'b0 ;
  assign y4208 = n12244 ;
  assign y4209 = ~n12246 ;
  assign y4210 = ~n12249 ;
  assign y4211 = ~1'b0 ;
  assign y4212 = ~n12250 ;
  assign y4213 = ~n12251 ;
  assign y4214 = ~n12255 ;
  assign y4215 = ~n12258 ;
  assign y4216 = ~1'b0 ;
  assign y4217 = ~n12261 ;
  assign y4218 = ~n12268 ;
  assign y4219 = n12269 ;
  assign y4220 = n12273 ;
  assign y4221 = n12274 ;
  assign y4222 = ~1'b0 ;
  assign y4223 = ~n12282 ;
  assign y4224 = n1154 ;
  assign y4225 = ~n12283 ;
  assign y4226 = ~n12284 ;
  assign y4227 = ~n12290 ;
  assign y4228 = n12292 ;
  assign y4229 = ~1'b0 ;
  assign y4230 = ~n5011 ;
  assign y4231 = n10258 ;
  assign y4232 = ~1'b0 ;
  assign y4233 = ~1'b0 ;
  assign y4234 = ~n12294 ;
  assign y4235 = ~n12297 ;
  assign y4236 = n12299 ;
  assign y4237 = ~n12300 ;
  assign y4238 = ~n12302 ;
  assign y4239 = ~1'b0 ;
  assign y4240 = ~1'b0 ;
  assign y4241 = ~n12306 ;
  assign y4242 = ~n12308 ;
  assign y4243 = n12311 ;
  assign y4244 = n12313 ;
  assign y4245 = ~n12318 ;
  assign y4246 = n12320 ;
  assign y4247 = ~1'b0 ;
  assign y4248 = ~n12324 ;
  assign y4249 = ~1'b0 ;
  assign y4250 = n12326 ;
  assign y4251 = n12327 ;
  assign y4252 = n12344 ;
  assign y4253 = n12346 ;
  assign y4254 = n12349 ;
  assign y4255 = n12351 ;
  assign y4256 = n12352 ;
  assign y4257 = ~1'b0 ;
  assign y4258 = n12357 ;
  assign y4259 = ~n12358 ;
  assign y4260 = ~n12360 ;
  assign y4261 = ~1'b0 ;
  assign y4262 = n12366 ;
  assign y4263 = n12367 ;
  assign y4264 = n12368 ;
  assign y4265 = ~1'b0 ;
  assign y4266 = n12369 ;
  assign y4267 = n12370 ;
  assign y4268 = n12372 ;
  assign y4269 = n12377 ;
  assign y4270 = n12380 ;
  assign y4271 = ~n12388 ;
  assign y4272 = n12389 ;
  assign y4273 = n12390 ;
  assign y4274 = ~n12391 ;
  assign y4275 = ~1'b0 ;
  assign y4276 = ~1'b0 ;
  assign y4277 = ~1'b0 ;
  assign y4278 = n12395 ;
  assign y4279 = ~1'b0 ;
  assign y4280 = ~n12396 ;
  assign y4281 = ~1'b0 ;
  assign y4282 = ~1'b0 ;
  assign y4283 = n12400 ;
  assign y4284 = ~n12402 ;
  assign y4285 = ~n857 ;
  assign y4286 = ~n12405 ;
  assign y4287 = n12411 ;
  assign y4288 = n12417 ;
  assign y4289 = ~n12419 ;
  assign y4290 = ~n12420 ;
  assign y4291 = n12430 ;
  assign y4292 = ~1'b0 ;
  assign y4293 = n12433 ;
  assign y4294 = 1'b0 ;
  assign y4295 = n12434 ;
  assign y4296 = n12438 ;
  assign y4297 = ~n12442 ;
  assign y4298 = n12460 ;
  assign y4299 = ~n12461 ;
  assign y4300 = n12470 ;
  assign y4301 = n12471 ;
  assign y4302 = n12472 ;
  assign y4303 = ~n12473 ;
  assign y4304 = ~n12478 ;
  assign y4305 = ~1'b0 ;
  assign y4306 = ~1'b0 ;
  assign y4307 = ~n12479 ;
  assign y4308 = ~n12480 ;
  assign y4309 = ~n12482 ;
  assign y4310 = n12483 ;
  assign y4311 = ~n12488 ;
  assign y4312 = ~n12491 ;
  assign y4313 = n12497 ;
  assign y4314 = ~n12505 ;
  assign y4315 = ~n12508 ;
  assign y4316 = n12512 ;
  assign y4317 = ~n12513 ;
  assign y4318 = n12515 ;
  assign y4319 = ~n12516 ;
  assign y4320 = ~1'b0 ;
  assign y4321 = n12527 ;
  assign y4322 = ~1'b0 ;
  assign y4323 = ~n12530 ;
  assign y4324 = ~n12532 ;
  assign y4325 = ~n12533 ;
  assign y4326 = n12534 ;
  assign y4327 = ~n12538 ;
  assign y4328 = ~n12539 ;
  assign y4329 = ~n12541 ;
  assign y4330 = ~1'b0 ;
  assign y4331 = n12546 ;
  assign y4332 = ~1'b0 ;
  assign y4333 = ~n1369 ;
  assign y4334 = n12549 ;
  assign y4335 = ~n12552 ;
  assign y4336 = ~1'b0 ;
  assign y4337 = n12558 ;
  assign y4338 = n12559 ;
  assign y4339 = ~n12561 ;
  assign y4340 = ~n12562 ;
  assign y4341 = n12564 ;
  assign y4342 = n12565 ;
  assign y4343 = n12576 ;
  assign y4344 = n12582 ;
  assign y4345 = ~1'b0 ;
  assign y4346 = n12584 ;
  assign y4347 = ~1'b0 ;
  assign y4348 = n2394 ;
  assign y4349 = ~n12595 ;
  assign y4350 = ~n9277 ;
  assign y4351 = ~n12600 ;
  assign y4352 = ~1'b0 ;
  assign y4353 = n12601 ;
  assign y4354 = ~n10145 ;
  assign y4355 = ~n12604 ;
  assign y4356 = n12606 ;
  assign y4357 = ~n12607 ;
  assign y4358 = n12609 ;
  assign y4359 = n12610 ;
  assign y4360 = n12617 ;
  assign y4361 = ~n12624 ;
  assign y4362 = n12629 ;
  assign y4363 = n12631 ;
  assign y4364 = ~n12633 ;
  assign y4365 = n12638 ;
  assign y4366 = ~n12640 ;
  assign y4367 = ~n12642 ;
  assign y4368 = n1463 ;
  assign y4369 = ~n12646 ;
  assign y4370 = ~n12651 ;
  assign y4371 = n12654 ;
  assign y4372 = ~n12659 ;
  assign y4373 = ~n12662 ;
  assign y4374 = ~1'b0 ;
  assign y4375 = n12664 ;
  assign y4376 = ~n12673 ;
  assign y4377 = ~1'b0 ;
  assign y4378 = ~1'b0 ;
  assign y4379 = ~n12675 ;
  assign y4380 = n12676 ;
  assign y4381 = n12679 ;
  assign y4382 = ~n12681 ;
  assign y4383 = ~n12682 ;
  assign y4384 = ~1'b0 ;
  assign y4385 = ~n12684 ;
  assign y4386 = n12689 ;
  assign y4387 = ~n12690 ;
  assign y4388 = n12693 ;
  assign y4389 = n12696 ;
  assign y4390 = ~n12703 ;
  assign y4391 = n12439 ;
  assign y4392 = ~n12704 ;
  assign y4393 = ~n12706 ;
  assign y4394 = n12707 ;
  assign y4395 = n12708 ;
  assign y4396 = n12713 ;
  assign y4397 = ~n12717 ;
  assign y4398 = ~n12721 ;
  assign y4399 = n12724 ;
  assign y4400 = n12728 ;
  assign y4401 = ~n12731 ;
  assign y4402 = ~n12734 ;
  assign y4403 = n12735 ;
  assign y4404 = n12736 ;
  assign y4405 = ~1'b0 ;
  assign y4406 = ~n12740 ;
  assign y4407 = ~1'b0 ;
  assign y4408 = ~1'b0 ;
  assign y4409 = n12742 ;
  assign y4410 = n12748 ;
  assign y4411 = ~1'b0 ;
  assign y4412 = n12756 ;
  assign y4413 = ~1'b0 ;
  assign y4414 = ~n12757 ;
  assign y4415 = ~n12758 ;
  assign y4416 = n12766 ;
  assign y4417 = ~1'b0 ;
  assign y4418 = ~n12769 ;
  assign y4419 = ~1'b0 ;
  assign y4420 = ~n12771 ;
  assign y4421 = n12775 ;
  assign y4422 = ~n12781 ;
  assign y4423 = ~n12782 ;
  assign y4424 = n12785 ;
  assign y4425 = ~n12788 ;
  assign y4426 = n12790 ;
  assign y4427 = ~n12796 ;
  assign y4428 = ~n2202 ;
  assign y4429 = ~n12797 ;
  assign y4430 = ~n5387 ;
  assign y4431 = ~1'b0 ;
  assign y4432 = ~n12799 ;
  assign y4433 = ~1'b0 ;
  assign y4434 = 1'b0 ;
  assign y4435 = ~1'b0 ;
  assign y4436 = n12800 ;
  assign y4437 = ~n12801 ;
  assign y4438 = ~n12809 ;
  assign y4439 = ~n12810 ;
  assign y4440 = n12811 ;
  assign y4441 = ~n12818 ;
  assign y4442 = ~n12823 ;
  assign y4443 = ~n12825 ;
  assign y4444 = n12827 ;
  assign y4445 = ~n12829 ;
  assign y4446 = n12831 ;
  assign y4447 = n12836 ;
  assign y4448 = n12837 ;
  assign y4449 = ~n12843 ;
  assign y4450 = n12845 ;
  assign y4451 = n12852 ;
  assign y4452 = n12854 ;
  assign y4453 = n12857 ;
  assign y4454 = ~1'b0 ;
  assign y4455 = ~n12860 ;
  assign y4456 = ~1'b0 ;
  assign y4457 = ~n12865 ;
  assign y4458 = 1'b0 ;
  assign y4459 = ~n12867 ;
  assign y4460 = n12870 ;
  assign y4461 = n12873 ;
  assign y4462 = ~1'b0 ;
  assign y4463 = ~n12879 ;
  assign y4464 = n12882 ;
  assign y4465 = ~n12883 ;
  assign y4466 = n12887 ;
  assign y4467 = ~1'b0 ;
  assign y4468 = n12891 ;
  assign y4469 = n12901 ;
  assign y4470 = ~1'b0 ;
  assign y4471 = n12903 ;
  assign y4472 = ~n12907 ;
  assign y4473 = ~n12909 ;
  assign y4474 = ~n12913 ;
  assign y4475 = n12914 ;
  assign y4476 = n12916 ;
  assign y4477 = n12918 ;
  assign y4478 = ~1'b0 ;
  assign y4479 = n12920 ;
  assign y4480 = n12921 ;
  assign y4481 = ~n12925 ;
  assign y4482 = n12931 ;
  assign y4483 = ~n12938 ;
  assign y4484 = n12948 ;
  assign y4485 = ~1'b0 ;
  assign y4486 = ~n12950 ;
  assign y4487 = n12955 ;
  assign y4488 = ~n12958 ;
  assign y4489 = ~1'b0 ;
  assign y4490 = n12959 ;
  assign y4491 = n12960 ;
  assign y4492 = ~n12963 ;
  assign y4493 = ~n12966 ;
  assign y4494 = ~n12967 ;
  assign y4495 = ~n12969 ;
  assign y4496 = ~n12970 ;
  assign y4497 = n12972 ;
  assign y4498 = ~n12980 ;
  assign y4499 = n12991 ;
  assign y4500 = ~n12998 ;
  assign y4501 = n12999 ;
  assign y4502 = ~n13002 ;
  assign y4503 = ~n10957 ;
  assign y4504 = n13004 ;
  assign y4505 = n13005 ;
  assign y4506 = n6512 ;
  assign y4507 = ~n13007 ;
  assign y4508 = n13014 ;
  assign y4509 = n13016 ;
  assign y4510 = ~n13021 ;
  assign y4511 = n13023 ;
  assign y4512 = ~n13024 ;
  assign y4513 = ~n13025 ;
  assign y4514 = n13028 ;
  assign y4515 = ~n13033 ;
  assign y4516 = ~n13036 ;
  assign y4517 = ~n13042 ;
  assign y4518 = n13047 ;
  assign y4519 = ~n13052 ;
  assign y4520 = n8106 ;
  assign y4521 = ~1'b0 ;
  assign y4522 = n13054 ;
  assign y4523 = n13060 ;
  assign y4524 = n13063 ;
  assign y4525 = ~n13069 ;
  assign y4526 = ~n13073 ;
  assign y4527 = n13076 ;
  assign y4528 = ~1'b0 ;
  assign y4529 = n13077 ;
  assign y4530 = ~n13085 ;
  assign y4531 = ~n13086 ;
  assign y4532 = ~n13087 ;
  assign y4533 = ~1'b0 ;
  assign y4534 = ~1'b0 ;
  assign y4535 = n13095 ;
  assign y4536 = ~n13108 ;
  assign y4537 = n13109 ;
  assign y4538 = ~n13115 ;
  assign y4539 = ~1'b0 ;
  assign y4540 = ~n13119 ;
  assign y4541 = n13126 ;
  assign y4542 = ~1'b0 ;
  assign y4543 = n13130 ;
  assign y4544 = ~n13133 ;
  assign y4545 = n13137 ;
  assign y4546 = ~1'b0 ;
  assign y4547 = ~n10525 ;
  assign y4548 = ~n13138 ;
  assign y4549 = ~n13142 ;
  assign y4550 = ~n13144 ;
  assign y4551 = n13147 ;
  assign y4552 = ~n13152 ;
  assign y4553 = ~n13160 ;
  assign y4554 = ~n13166 ;
  assign y4555 = n13167 ;
  assign y4556 = n13173 ;
  assign y4557 = n13174 ;
  assign y4558 = n13175 ;
  assign y4559 = ~1'b0 ;
  assign y4560 = ~n13176 ;
  assign y4561 = ~n13179 ;
  assign y4562 = ~1'b0 ;
  assign y4563 = n13180 ;
  assign y4564 = n13186 ;
  assign y4565 = ~n13187 ;
  assign y4566 = n13188 ;
  assign y4567 = 1'b0 ;
  assign y4568 = n13191 ;
  assign y4569 = ~n13200 ;
  assign y4570 = n13201 ;
  assign y4571 = n13204 ;
  assign y4572 = ~n13207 ;
  assign y4573 = n13208 ;
  assign y4574 = ~1'b0 ;
  assign y4575 = ~1'b0 ;
  assign y4576 = n13209 ;
  assign y4577 = ~n13210 ;
  assign y4578 = n13212 ;
  assign y4579 = n13214 ;
  assign y4580 = n13218 ;
  assign y4581 = ~1'b0 ;
  assign y4582 = n9276 ;
  assign y4583 = ~1'b0 ;
  assign y4584 = ~n13223 ;
  assign y4585 = ~n13233 ;
  assign y4586 = n13237 ;
  assign y4587 = ~n13239 ;
  assign y4588 = ~n13241 ;
  assign y4589 = ~n13243 ;
  assign y4590 = ~n13249 ;
  assign y4591 = n13250 ;
  assign y4592 = n13251 ;
  assign y4593 = ~n13254 ;
  assign y4594 = ~n13257 ;
  assign y4595 = n13259 ;
  assign y4596 = n13260 ;
  assign y4597 = ~n13265 ;
  assign y4598 = n12407 ;
  assign y4599 = ~n13268 ;
  assign y4600 = ~n13275 ;
  assign y4601 = ~n6001 ;
  assign y4602 = n13277 ;
  assign y4603 = ~n13280 ;
  assign y4604 = n13281 ;
  assign y4605 = n13283 ;
  assign y4606 = ~1'b0 ;
  assign y4607 = ~n13284 ;
  assign y4608 = ~n13285 ;
  assign y4609 = n13291 ;
  assign y4610 = n13293 ;
  assign y4611 = ~1'b0 ;
  assign y4612 = n13295 ;
  assign y4613 = ~1'b0 ;
  assign y4614 = n13299 ;
  assign y4615 = ~n13300 ;
  assign y4616 = ~n13303 ;
  assign y4617 = ~n12906 ;
  assign y4618 = ~1'b0 ;
  assign y4619 = ~n13304 ;
  assign y4620 = n13312 ;
  assign y4621 = n13316 ;
  assign y4622 = ~1'b0 ;
  assign y4623 = ~n13317 ;
  assign y4624 = n13319 ;
  assign y4625 = ~n13321 ;
  assign y4626 = ~n13324 ;
  assign y4627 = ~n13329 ;
  assign y4628 = ~1'b0 ;
  assign y4629 = ~n13331 ;
  assign y4630 = n13333 ;
  assign y4631 = ~n13340 ;
  assign y4632 = ~1'b0 ;
  assign y4633 = n13342 ;
  assign y4634 = n13344 ;
  assign y4635 = n13345 ;
  assign y4636 = ~n13350 ;
  assign y4637 = n13353 ;
  assign y4638 = n13354 ;
  assign y4639 = n13358 ;
  assign y4640 = n13359 ;
  assign y4641 = n13361 ;
  assign y4642 = ~n13362 ;
  assign y4643 = ~n13367 ;
  assign y4644 = n13376 ;
  assign y4645 = n13385 ;
  assign y4646 = ~n13388 ;
  assign y4647 = n13389 ;
  assign y4648 = ~n13391 ;
  assign y4649 = ~n13393 ;
  assign y4650 = n13397 ;
  assign y4651 = ~n13400 ;
  assign y4652 = n13404 ;
  assign y4653 = n13405 ;
  assign y4654 = ~n13411 ;
  assign y4655 = n13415 ;
  assign y4656 = ~n13416 ;
  assign y4657 = n13417 ;
  assign y4658 = ~1'b0 ;
  assign y4659 = n13418 ;
  assign y4660 = ~1'b0 ;
  assign y4661 = ~1'b0 ;
  assign y4662 = ~1'b0 ;
  assign y4663 = n13420 ;
  assign y4664 = ~n13422 ;
  assign y4665 = ~n13429 ;
  assign y4666 = ~n13432 ;
  assign y4667 = ~n13435 ;
  assign y4668 = n13436 ;
  assign y4669 = ~1'b0 ;
  assign y4670 = ~n13440 ;
  assign y4671 = ~n13443 ;
  assign y4672 = n13449 ;
  assign y4673 = ~n13450 ;
  assign y4674 = ~1'b0 ;
  assign y4675 = n13451 ;
  assign y4676 = n13459 ;
  assign y4677 = n13464 ;
  assign y4678 = n13465 ;
  assign y4679 = ~1'b0 ;
  assign y4680 = ~n13466 ;
  assign y4681 = ~n13468 ;
  assign y4682 = ~n9729 ;
  assign y4683 = ~n13477 ;
  assign y4684 = n13480 ;
  assign y4685 = n13485 ;
  assign y4686 = ~n13489 ;
  assign y4687 = ~1'b0 ;
  assign y4688 = ~1'b0 ;
  assign y4689 = n13493 ;
  assign y4690 = ~n13502 ;
  assign y4691 = n13505 ;
  assign y4692 = ~1'b0 ;
  assign y4693 = ~1'b0 ;
  assign y4694 = n13507 ;
  assign y4695 = n13516 ;
  assign y4696 = ~n13518 ;
  assign y4697 = ~n13524 ;
  assign y4698 = ~n13526 ;
  assign y4699 = n13527 ;
  assign y4700 = ~n13529 ;
  assign y4701 = ~n13531 ;
  assign y4702 = n13534 ;
  assign y4703 = ~n13537 ;
  assign y4704 = n13538 ;
  assign y4705 = n13543 ;
  assign y4706 = ~1'b0 ;
  assign y4707 = ~n13548 ;
  assign y4708 = n13550 ;
  assign y4709 = ~n13555 ;
  assign y4710 = ~n13556 ;
  assign y4711 = ~1'b0 ;
  assign y4712 = ~n13557 ;
  assign y4713 = n2001 ;
  assign y4714 = ~n13559 ;
  assign y4715 = n13560 ;
  assign y4716 = n13562 ;
  assign y4717 = ~n13563 ;
  assign y4718 = n12400 ;
  assign y4719 = n13571 ;
  assign y4720 = n13574 ;
  assign y4721 = ~1'b0 ;
  assign y4722 = ~n13579 ;
  assign y4723 = n13585 ;
  assign y4724 = ~1'b0 ;
  assign y4725 = ~n13592 ;
  assign y4726 = ~1'b0 ;
  assign y4727 = n13595 ;
  assign y4728 = ~n13600 ;
  assign y4729 = n13602 ;
  assign y4730 = n13603 ;
  assign y4731 = n13605 ;
  assign y4732 = ~n13607 ;
  assign y4733 = ~n13609 ;
  assign y4734 = ~n13610 ;
  assign y4735 = ~n13612 ;
  assign y4736 = n13616 ;
  assign y4737 = ~n13617 ;
  assign y4738 = n13621 ;
  assign y4739 = ~n12231 ;
  assign y4740 = n13622 ;
  assign y4741 = n13623 ;
  assign y4742 = n13626 ;
  assign y4743 = n4177 ;
  assign y4744 = n13627 ;
  assign y4745 = ~n1707 ;
  assign y4746 = ~n13633 ;
  assign y4747 = ~n13635 ;
  assign y4748 = ~1'b0 ;
  assign y4749 = ~n13643 ;
  assign y4750 = ~n13644 ;
  assign y4751 = ~n13649 ;
  assign y4752 = ~1'b0 ;
  assign y4753 = ~n13650 ;
  assign y4754 = n13654 ;
  assign y4755 = n13656 ;
  assign y4756 = ~1'b0 ;
  assign y4757 = ~n13658 ;
  assign y4758 = n13664 ;
  assign y4759 = n13667 ;
  assign y4760 = ~n13669 ;
  assign y4761 = ~1'b0 ;
  assign y4762 = ~n13672 ;
  assign y4763 = ~n13673 ;
  assign y4764 = ~n13677 ;
  assign y4765 = ~n13681 ;
  assign y4766 = n13684 ;
  assign y4767 = ~n13689 ;
  assign y4768 = n13691 ;
  assign y4769 = n13693 ;
  assign y4770 = ~n1250 ;
  assign y4771 = ~1'b0 ;
  assign y4772 = ~1'b0 ;
  assign y4773 = ~n13706 ;
  assign y4774 = ~n702 ;
  assign y4775 = n13715 ;
  assign y4776 = ~n13718 ;
  assign y4777 = ~1'b0 ;
  assign y4778 = n13734 ;
  assign y4779 = ~n13738 ;
  assign y4780 = n13745 ;
  assign y4781 = ~n13751 ;
  assign y4782 = n13753 ;
  assign y4783 = ~n13754 ;
  assign y4784 = ~1'b0 ;
  assign y4785 = ~n13758 ;
  assign y4786 = ~n13759 ;
  assign y4787 = n13762 ;
  assign y4788 = ~1'b0 ;
  assign y4789 = ~n13763 ;
  assign y4790 = n13770 ;
  assign y4791 = ~n13773 ;
  assign y4792 = ~n13776 ;
  assign y4793 = ~n13781 ;
  assign y4794 = n13788 ;
  assign y4795 = n13792 ;
  assign y4796 = ~1'b0 ;
  assign y4797 = ~n13793 ;
  assign y4798 = ~n13796 ;
  assign y4799 = ~n13800 ;
  assign y4800 = ~n13801 ;
  assign y4801 = n13803 ;
  assign y4802 = ~1'b0 ;
  assign y4803 = ~n13808 ;
  assign y4804 = ~n13810 ;
  assign y4805 = ~n13812 ;
  assign y4806 = ~n13813 ;
  assign y4807 = ~n13816 ;
  assign y4808 = ~n13820 ;
  assign y4809 = n13822 ;
  assign y4810 = ~n13823 ;
  assign y4811 = n3899 ;
  assign y4812 = ~n13826 ;
  assign y4813 = n13841 ;
  assign y4814 = ~n13842 ;
  assign y4815 = ~n13844 ;
  assign y4816 = ~n13854 ;
  assign y4817 = ~n13862 ;
  assign y4818 = n13867 ;
  assign y4819 = ~1'b0 ;
  assign y4820 = n13869 ;
  assign y4821 = ~1'b0 ;
  assign y4822 = ~n13875 ;
  assign y4823 = n13879 ;
  assign y4824 = n13883 ;
  assign y4825 = ~1'b0 ;
  assign y4826 = n13886 ;
  assign y4827 = ~1'b0 ;
  assign y4828 = ~1'b0 ;
  assign y4829 = ~n13887 ;
  assign y4830 = ~1'b0 ;
  assign y4831 = ~n13890 ;
  assign y4832 = n13891 ;
  assign y4833 = ~n13892 ;
  assign y4834 = n11501 ;
  assign y4835 = ~n13894 ;
  assign y4836 = n12091 ;
  assign y4837 = ~1'b0 ;
  assign y4838 = n13895 ;
  assign y4839 = ~n13897 ;
  assign y4840 = n13899 ;
  assign y4841 = n13902 ;
  assign y4842 = n13903 ;
  assign y4843 = ~n13905 ;
  assign y4844 = n13907 ;
  assign y4845 = n13910 ;
  assign y4846 = n13913 ;
  assign y4847 = ~1'b0 ;
  assign y4848 = ~n13915 ;
  assign y4849 = ~1'b0 ;
  assign y4850 = ~n13918 ;
  assign y4851 = ~n13921 ;
  assign y4852 = ~n13922 ;
  assign y4853 = n13923 ;
  assign y4854 = ~n13926 ;
  assign y4855 = ~n13937 ;
  assign y4856 = ~1'b0 ;
  assign y4857 = n13940 ;
  assign y4858 = ~n13943 ;
  assign y4859 = n13946 ;
  assign y4860 = ~n13949 ;
  assign y4861 = ~n13951 ;
  assign y4862 = n13956 ;
  assign y4863 = n13961 ;
  assign y4864 = n13964 ;
  assign y4865 = ~n13976 ;
  assign y4866 = ~n13987 ;
  assign y4867 = ~n13992 ;
  assign y4868 = ~n13993 ;
  assign y4869 = ~1'b0 ;
  assign y4870 = ~1'b0 ;
  assign y4871 = ~n13998 ;
  assign y4872 = ~n13999 ;
  assign y4873 = ~n14007 ;
  assign y4874 = ~n14010 ;
  assign y4875 = ~1'b0 ;
  assign y4876 = n14012 ;
  assign y4877 = ~n14017 ;
  assign y4878 = ~n14019 ;
  assign y4879 = n3667 ;
  assign y4880 = ~1'b0 ;
  assign y4881 = ~1'b0 ;
  assign y4882 = ~n14025 ;
  assign y4883 = n14027 ;
  assign y4884 = n14030 ;
  assign y4885 = ~n14034 ;
  assign y4886 = n14037 ;
  assign y4887 = n14041 ;
  assign y4888 = ~n14043 ;
  assign y4889 = ~n14044 ;
  assign y4890 = n14045 ;
  assign y4891 = ~1'b0 ;
  assign y4892 = ~n14046 ;
  assign y4893 = n14052 ;
  assign y4894 = n4356 ;
  assign y4895 = ~n14056 ;
  assign y4896 = ~1'b0 ;
  assign y4897 = ~1'b0 ;
  assign y4898 = ~1'b0 ;
  assign y4899 = ~n14058 ;
  assign y4900 = ~n14061 ;
  assign y4901 = ~n14064 ;
  assign y4902 = n14067 ;
  assign y4903 = ~n14075 ;
  assign y4904 = ~n14077 ;
  assign y4905 = ~n14078 ;
  assign y4906 = ~n14081 ;
  assign y4907 = ~1'b0 ;
  assign y4908 = ~n14083 ;
  assign y4909 = n14085 ;
  assign y4910 = ~1'b0 ;
  assign y4911 = n14086 ;
  assign y4912 = n11665 ;
  assign y4913 = n14088 ;
  assign y4914 = ~1'b0 ;
  assign y4915 = ~n14089 ;
  assign y4916 = ~n14096 ;
  assign y4917 = ~1'b0 ;
  assign y4918 = n14102 ;
  assign y4919 = ~1'b0 ;
  assign y4920 = n14107 ;
  assign y4921 = ~n14113 ;
  assign y4922 = n14117 ;
  assign y4923 = n14119 ;
  assign y4924 = ~n14122 ;
  assign y4925 = ~n14127 ;
  assign y4926 = n13166 ;
  assign y4927 = ~n14133 ;
  assign y4928 = ~1'b0 ;
  assign y4929 = ~1'b0 ;
  assign y4930 = n14137 ;
  assign y4931 = ~n11373 ;
  assign y4932 = ~n14140 ;
  assign y4933 = n14146 ;
  assign y4934 = ~1'b0 ;
  assign y4935 = n14155 ;
  assign y4936 = ~n14156 ;
  assign y4937 = n14161 ;
  assign y4938 = n14163 ;
  assign y4939 = n14166 ;
  assign y4940 = ~n14168 ;
  assign y4941 = ~n14169 ;
  assign y4942 = ~n14172 ;
  assign y4943 = ~n14173 ;
  assign y4944 = ~n14174 ;
  assign y4945 = ~1'b0 ;
  assign y4946 = ~1'b0 ;
  assign y4947 = n14176 ;
  assign y4948 = ~n14177 ;
  assign y4949 = ~n14179 ;
  assign y4950 = ~n14180 ;
  assign y4951 = ~1'b0 ;
  assign y4952 = ~n14182 ;
  assign y4953 = n14183 ;
  assign y4954 = n14188 ;
  assign y4955 = n6556 ;
  assign y4956 = ~n14198 ;
  assign y4957 = ~n14199 ;
  assign y4958 = n14201 ;
  assign y4959 = n14204 ;
  assign y4960 = ~n14205 ;
  assign y4961 = n1517 ;
  assign y4962 = ~n14212 ;
  assign y4963 = ~n14213 ;
  assign y4964 = n14219 ;
  assign y4965 = ~n14223 ;
  assign y4966 = ~n14225 ;
  assign y4967 = ~n14227 ;
  assign y4968 = ~1'b0 ;
  assign y4969 = ~n14232 ;
  assign y4970 = n14241 ;
  assign y4971 = ~1'b0 ;
  assign y4972 = n14242 ;
  assign y4973 = ~1'b0 ;
  assign y4974 = ~1'b0 ;
  assign y4975 = ~n14248 ;
  assign y4976 = n14251 ;
  assign y4977 = n14252 ;
  assign y4978 = ~n14253 ;
  assign y4979 = ~n14255 ;
  assign y4980 = ~n14259 ;
  assign y4981 = ~n14260 ;
  assign y4982 = n14264 ;
  assign y4983 = ~1'b0 ;
  assign y4984 = n14265 ;
  assign y4985 = ~n14266 ;
  assign y4986 = n14268 ;
  assign y4987 = ~n14279 ;
  assign y4988 = n891 ;
  assign y4989 = ~n14281 ;
  assign y4990 = ~n14282 ;
  assign y4991 = ~n14288 ;
  assign y4992 = n14291 ;
  assign y4993 = n14297 ;
  assign y4994 = ~n14302 ;
  assign y4995 = ~n14306 ;
  assign y4996 = ~n14307 ;
  assign y4997 = n14309 ;
  assign y4998 = n14315 ;
  assign y4999 = ~n14318 ;
  assign y5000 = n14325 ;
  assign y5001 = n11315 ;
  assign y5002 = ~n14327 ;
  assign y5003 = n14328 ;
  assign y5004 = n14329 ;
  assign y5005 = ~n14331 ;
  assign y5006 = ~n9139 ;
  assign y5007 = ~n14333 ;
  assign y5008 = ~n14337 ;
  assign y5009 = n14339 ;
  assign y5010 = n14342 ;
  assign y5011 = ~n14351 ;
  assign y5012 = n14352 ;
  assign y5013 = n14353 ;
  assign y5014 = ~n14355 ;
  assign y5015 = ~n14361 ;
  assign y5016 = n14364 ;
  assign y5017 = ~n14365 ;
  assign y5018 = n14376 ;
  assign y5019 = n14377 ;
  assign y5020 = ~n14380 ;
  assign y5021 = n14384 ;
  assign y5022 = n14397 ;
  assign y5023 = ~n14398 ;
  assign y5024 = ~1'b0 ;
  assign y5025 = n14400 ;
  assign y5026 = ~n14402 ;
  assign y5027 = ~n14403 ;
  assign y5028 = n14404 ;
  assign y5029 = ~n14405 ;
  assign y5030 = ~n14406 ;
  assign y5031 = n14408 ;
  assign y5032 = ~n14409 ;
  assign y5033 = ~1'b0 ;
  assign y5034 = ~n14415 ;
  assign y5035 = ~1'b0 ;
  assign y5036 = ~n14418 ;
  assign y5037 = n14421 ;
  assign y5038 = n14423 ;
  assign y5039 = n14429 ;
  assign y5040 = 1'b0 ;
  assign y5041 = n14433 ;
  assign y5042 = ~n14435 ;
  assign y5043 = ~n14437 ;
  assign y5044 = ~n14438 ;
  assign y5045 = n14443 ;
  assign y5046 = n14446 ;
  assign y5047 = ~n14453 ;
  assign y5048 = ~n14454 ;
  assign y5049 = ~n14456 ;
  assign y5050 = n14458 ;
  assign y5051 = ~n14460 ;
  assign y5052 = ~n14462 ;
  assign y5053 = 1'b0 ;
  assign y5054 = ~n14464 ;
  assign y5055 = ~1'b0 ;
  assign y5056 = ~n14470 ;
  assign y5057 = ~n14473 ;
  assign y5058 = n14475 ;
  assign y5059 = ~n14481 ;
  assign y5060 = ~1'b0 ;
  assign y5061 = ~1'b0 ;
  assign y5062 = ~n14482 ;
  assign y5063 = ~n14483 ;
  assign y5064 = n14484 ;
  assign y5065 = n14485 ;
  assign y5066 = n14486 ;
  assign y5067 = ~n14492 ;
  assign y5068 = n14496 ;
  assign y5069 = ~1'b0 ;
  assign y5070 = ~n14498 ;
  assign y5071 = n14500 ;
  assign y5072 = ~1'b0 ;
  assign y5073 = ~n14508 ;
  assign y5074 = 1'b0 ;
  assign y5075 = ~n6574 ;
  assign y5076 = n14509 ;
  assign y5077 = ~n14517 ;
  assign y5078 = ~n14519 ;
  assign y5079 = ~1'b0 ;
  assign y5080 = n14521 ;
  assign y5081 = ~n14524 ;
  assign y5082 = n14531 ;
  assign y5083 = ~n14533 ;
  assign y5084 = ~n14536 ;
  assign y5085 = ~1'b0 ;
  assign y5086 = ~1'b0 ;
  assign y5087 = ~n14537 ;
  assign y5088 = ~n14539 ;
  assign y5089 = ~n14540 ;
  assign y5090 = n14558 ;
  assign y5091 = n14562 ;
  assign y5092 = n14565 ;
  assign y5093 = n14566 ;
  assign y5094 = ~n14567 ;
  assign y5095 = ~n14568 ;
  assign y5096 = n14573 ;
  assign y5097 = n14577 ;
  assign y5098 = 1'b0 ;
  assign y5099 = ~n14580 ;
  assign y5100 = ~n14581 ;
  assign y5101 = ~1'b0 ;
  assign y5102 = n2469 ;
  assign y5103 = n14582 ;
  assign y5104 = ~1'b0 ;
  assign y5105 = ~1'b0 ;
  assign y5106 = 1'b0 ;
  assign y5107 = ~n14589 ;
  assign y5108 = n14596 ;
  assign y5109 = ~1'b0 ;
  assign y5110 = ~1'b0 ;
  assign y5111 = ~n14598 ;
  assign y5112 = n14599 ;
  assign y5113 = n14602 ;
  assign y5114 = ~n14604 ;
  assign y5115 = n14608 ;
  assign y5116 = ~n3960 ;
  assign y5117 = n14609 ;
  assign y5118 = n14615 ;
  assign y5119 = ~n14621 ;
  assign y5120 = n14625 ;
  assign y5121 = ~n14626 ;
  assign y5122 = ~1'b0 ;
  assign y5123 = ~1'b0 ;
  assign y5124 = ~n14627 ;
  assign y5125 = ~n14630 ;
  assign y5126 = ~1'b0 ;
  assign y5127 = ~n14635 ;
  assign y5128 = n14638 ;
  assign y5129 = n14641 ;
  assign y5130 = n14644 ;
  assign y5131 = ~n14646 ;
  assign y5132 = ~n14649 ;
  assign y5133 = n14657 ;
  assign y5134 = n14661 ;
  assign y5135 = ~n6054 ;
  assign y5136 = ~n14667 ;
  assign y5137 = n14673 ;
  assign y5138 = ~1'b0 ;
  assign y5139 = n14685 ;
  assign y5140 = ~n14688 ;
  assign y5141 = ~n14690 ;
  assign y5142 = ~1'b0 ;
  assign y5143 = ~1'b0 ;
  assign y5144 = ~n14705 ;
  assign y5145 = ~n14707 ;
  assign y5146 = ~n14708 ;
  assign y5147 = n14717 ;
  assign y5148 = n14719 ;
  assign y5149 = ~n14722 ;
  assign y5150 = ~n14724 ;
  assign y5151 = n14725 ;
  assign y5152 = n14728 ;
  assign y5153 = n14731 ;
  assign y5154 = ~n14732 ;
  assign y5155 = ~n14735 ;
  assign y5156 = ~n14743 ;
  assign y5157 = ~n14744 ;
  assign y5158 = ~n14746 ;
  assign y5159 = n14748 ;
  assign y5160 = ~n14751 ;
  assign y5161 = ~n14755 ;
  assign y5162 = ~n14756 ;
  assign y5163 = ~1'b0 ;
  assign y5164 = ~1'b0 ;
  assign y5165 = ~n14757 ;
  assign y5166 = ~n9707 ;
  assign y5167 = ~1'b0 ;
  assign y5168 = n14760 ;
  assign y5169 = ~n14762 ;
  assign y5170 = ~n14765 ;
  assign y5171 = ~n14768 ;
  assign y5172 = 1'b0 ;
  assign y5173 = ~1'b0 ;
  assign y5174 = ~n14770 ;
  assign y5175 = ~1'b0 ;
  assign y5176 = n14772 ;
  assign y5177 = ~n14776 ;
  assign y5178 = ~n14778 ;
  assign y5179 = ~n14779 ;
  assign y5180 = n14780 ;
  assign y5181 = ~1'b0 ;
  assign y5182 = n14782 ;
  assign y5183 = ~n14784 ;
  assign y5184 = ~1'b0 ;
  assign y5185 = ~n14786 ;
  assign y5186 = 1'b0 ;
  assign y5187 = n14790 ;
  assign y5188 = n14795 ;
  assign y5189 = ~n14801 ;
  assign y5190 = ~n14804 ;
  assign y5191 = n14810 ;
  assign y5192 = ~1'b0 ;
  assign y5193 = ~n14813 ;
  assign y5194 = ~n14816 ;
  assign y5195 = n14825 ;
  assign y5196 = n14833 ;
  assign y5197 = ~1'b0 ;
  assign y5198 = n14838 ;
  assign y5199 = n2520 ;
  assign y5200 = n13987 ;
  assign y5201 = n14840 ;
  assign y5202 = ~n14842 ;
  assign y5203 = n14845 ;
  assign y5204 = n14852 ;
  assign y5205 = ~1'b0 ;
  assign y5206 = ~n14858 ;
  assign y5207 = ~n14864 ;
  assign y5208 = n14874 ;
  assign y5209 = ~n14876 ;
  assign y5210 = ~n14877 ;
  assign y5211 = ~1'b0 ;
  assign y5212 = n14878 ;
  assign y5213 = ~n14880 ;
  assign y5214 = ~n14883 ;
  assign y5215 = ~1'b0 ;
  assign y5216 = n14891 ;
  assign y5217 = ~n14892 ;
  assign y5218 = ~n14895 ;
  assign y5219 = n14899 ;
  assign y5220 = n14900 ;
  assign y5221 = ~n14919 ;
  assign y5222 = ~1'b0 ;
  assign y5223 = n14927 ;
  assign y5224 = ~n14934 ;
  assign y5225 = n14941 ;
  assign y5226 = ~1'b0 ;
  assign y5227 = ~n14942 ;
  assign y5228 = ~n14944 ;
  assign y5229 = ~n14949 ;
  assign y5230 = n14955 ;
  assign y5231 = n14958 ;
  assign y5232 = n14961 ;
  assign y5233 = ~n14963 ;
  assign y5234 = ~1'b0 ;
  assign y5235 = ~n14971 ;
  assign y5236 = ~n14973 ;
  assign y5237 = ~1'b0 ;
  assign y5238 = ~1'b0 ;
  assign y5239 = n14977 ;
  assign y5240 = n14980 ;
  assign y5241 = ~n14982 ;
  assign y5242 = n14983 ;
  assign y5243 = ~n14986 ;
  assign y5244 = ~1'b0 ;
  assign y5245 = ~1'b0 ;
  assign y5246 = ~n14988 ;
  assign y5247 = n14989 ;
  assign y5248 = n14990 ;
  assign y5249 = ~n14995 ;
  assign y5250 = ~1'b0 ;
  assign y5251 = ~1'b0 ;
  assign y5252 = n14998 ;
  assign y5253 = n15000 ;
  assign y5254 = ~n15006 ;
  assign y5255 = ~n15007 ;
  assign y5256 = ~n2080 ;
  assign y5257 = ~1'b0 ;
  assign y5258 = n15015 ;
  assign y5259 = n15017 ;
  assign y5260 = ~n15018 ;
  assign y5261 = ~n15020 ;
  assign y5262 = ~1'b0 ;
  assign y5263 = n15022 ;
  assign y5264 = ~n15024 ;
  assign y5265 = ~n15037 ;
  assign y5266 = ~n15042 ;
  assign y5267 = ~n15045 ;
  assign y5268 = n15050 ;
  assign y5269 = ~1'b0 ;
  assign y5270 = ~n15051 ;
  assign y5271 = ~n15056 ;
  assign y5272 = ~n15065 ;
  assign y5273 = ~n15070 ;
  assign y5274 = n15074 ;
  assign y5275 = ~n15082 ;
  assign y5276 = ~1'b0 ;
  assign y5277 = ~n1831 ;
  assign y5278 = n15083 ;
  assign y5279 = n15084 ;
  assign y5280 = ~n15088 ;
  assign y5281 = ~n15089 ;
  assign y5282 = ~n15090 ;
  assign y5283 = ~n15092 ;
  assign y5284 = n15093 ;
  assign y5285 = ~1'b0 ;
  assign y5286 = n15094 ;
  assign y5287 = ~1'b0 ;
  assign y5288 = n15095 ;
  assign y5289 = ~n15097 ;
  assign y5290 = n15099 ;
  assign y5291 = ~n15102 ;
  assign y5292 = n15106 ;
  assign y5293 = ~n15113 ;
  assign y5294 = n15116 ;
  assign y5295 = n2459 ;
  assign y5296 = n15120 ;
  assign y5297 = n15123 ;
  assign y5298 = ~n15126 ;
  assign y5299 = ~n15134 ;
  assign y5300 = ~n15136 ;
  assign y5301 = ~n15137 ;
  assign y5302 = ~1'b0 ;
  assign y5303 = ~n15142 ;
  assign y5304 = ~1'b0 ;
  assign y5305 = ~n15143 ;
  assign y5306 = n15147 ;
  assign y5307 = n15155 ;
  assign y5308 = ~n15157 ;
  assign y5309 = ~n15161 ;
  assign y5310 = ~n15164 ;
  assign y5311 = n15166 ;
  assign y5312 = ~n15167 ;
  assign y5313 = ~1'b0 ;
  assign y5314 = ~n15168 ;
  assign y5315 = n15169 ;
  assign y5316 = ~n15170 ;
  assign y5317 = n3837 ;
  assign y5318 = ~n15173 ;
  assign y5319 = ~n15175 ;
  assign y5320 = ~1'b0 ;
  assign y5321 = ~n15184 ;
  assign y5322 = ~n15187 ;
  assign y5323 = ~n15189 ;
  assign y5324 = n15192 ;
  assign y5325 = ~n15198 ;
  assign y5326 = ~n15202 ;
  assign y5327 = n15204 ;
  assign y5328 = ~n15205 ;
  assign y5329 = ~1'b0 ;
  assign y5330 = ~1'b0 ;
  assign y5331 = ~n15206 ;
  assign y5332 = ~n15210 ;
  assign y5333 = ~1'b0 ;
  assign y5334 = n15217 ;
  assign y5335 = n15223 ;
  assign y5336 = ~1'b0 ;
  assign y5337 = n15224 ;
  assign y5338 = n15230 ;
  assign y5339 = ~n15244 ;
  assign y5340 = ~n15248 ;
  assign y5341 = n15254 ;
  assign y5342 = n15255 ;
  assign y5343 = ~1'b0 ;
  assign y5344 = n15258 ;
  assign y5345 = ~n15261 ;
  assign y5346 = ~n15270 ;
  assign y5347 = n15271 ;
  assign y5348 = ~n15272 ;
  assign y5349 = n15274 ;
  assign y5350 = ~n4332 ;
  assign y5351 = ~n15275 ;
  assign y5352 = ~n15276 ;
  assign y5353 = ~n15279 ;
  assign y5354 = ~1'b0 ;
  assign y5355 = n15285 ;
  assign y5356 = ~n15288 ;
  assign y5357 = n15289 ;
  assign y5358 = n15293 ;
  assign y5359 = ~n15294 ;
  assign y5360 = ~1'b0 ;
  assign y5361 = ~1'b0 ;
  assign y5362 = ~n6170 ;
  assign y5363 = ~1'b0 ;
  assign y5364 = n15295 ;
  assign y5365 = ~n15296 ;
  assign y5366 = ~n15299 ;
  assign y5367 = ~1'b0 ;
  assign y5368 = ~n15303 ;
  assign y5369 = ~1'b0 ;
  assign y5370 = ~n15306 ;
  assign y5371 = ~n15307 ;
  assign y5372 = n15309 ;
  assign y5373 = n15315 ;
  assign y5374 = n15321 ;
  assign y5375 = n15323 ;
  assign y5376 = n15326 ;
  assign y5377 = n15327 ;
  assign y5378 = n15330 ;
  assign y5379 = ~n15333 ;
  assign y5380 = ~1'b0 ;
  assign y5381 = ~n15338 ;
  assign y5382 = ~n15341 ;
  assign y5383 = ~n15342 ;
  assign y5384 = ~1'b0 ;
  assign y5385 = ~n15345 ;
  assign y5386 = ~n15350 ;
  assign y5387 = ~n15357 ;
  assign y5388 = n15364 ;
  assign y5389 = ~1'b0 ;
  assign y5390 = n15368 ;
  assign y5391 = ~n15369 ;
  assign y5392 = ~1'b0 ;
  assign y5393 = n15373 ;
  assign y5394 = n15375 ;
  assign y5395 = ~n15380 ;
  assign y5396 = ~n15382 ;
  assign y5397 = n15383 ;
  assign y5398 = ~n15384 ;
  assign y5399 = n15385 ;
  assign y5400 = ~1'b0 ;
  assign y5401 = ~1'b0 ;
  assign y5402 = n15387 ;
  assign y5403 = n15388 ;
  assign y5404 = n15390 ;
  assign y5405 = ~n15393 ;
  assign y5406 = n15395 ;
  assign y5407 = ~1'b0 ;
  assign y5408 = n15403 ;
  assign y5409 = ~n15405 ;
  assign y5410 = ~n15406 ;
  assign y5411 = ~1'b0 ;
  assign y5412 = n15409 ;
  assign y5413 = ~n15413 ;
  assign y5414 = ~n15417 ;
  assign y5415 = n15420 ;
  assign y5416 = 1'b0 ;
  assign y5417 = ~n15423 ;
  assign y5418 = ~n652 ;
  assign y5419 = n15424 ;
  assign y5420 = ~n15432 ;
  assign y5421 = ~n15435 ;
  assign y5422 = ~1'b0 ;
  assign y5423 = n15440 ;
  assign y5424 = n15442 ;
  assign y5425 = n15447 ;
  assign y5426 = n7775 ;
  assign y5427 = n15450 ;
  assign y5428 = ~n15451 ;
  assign y5429 = n15455 ;
  assign y5430 = ~1'b0 ;
  assign y5431 = ~1'b0 ;
  assign y5432 = ~n15456 ;
  assign y5433 = n15457 ;
  assign y5434 = ~n15459 ;
  assign y5435 = n15461 ;
  assign y5436 = ~1'b0 ;
  assign y5437 = ~n15464 ;
  assign y5438 = n15466 ;
  assign y5439 = ~1'b0 ;
  assign y5440 = ~1'b0 ;
  assign y5441 = n15472 ;
  assign y5442 = n15474 ;
  assign y5443 = n15475 ;
  assign y5444 = n15477 ;
  assign y5445 = n15480 ;
  assign y5446 = n15484 ;
  assign y5447 = ~n15487 ;
  assign y5448 = n15490 ;
  assign y5449 = n15491 ;
  assign y5450 = n15493 ;
  assign y5451 = ~n15494 ;
  assign y5452 = ~n5950 ;
  assign y5453 = ~n15496 ;
  assign y5454 = n15497 ;
  assign y5455 = ~n15501 ;
  assign y5456 = n15503 ;
  assign y5457 = ~n15504 ;
  assign y5458 = n15506 ;
  assign y5459 = n15508 ;
  assign y5460 = ~1'b0 ;
  assign y5461 = ~n15511 ;
  assign y5462 = n9234 ;
  assign y5463 = n15512 ;
  assign y5464 = ~n15514 ;
  assign y5465 = ~n15516 ;
  assign y5466 = n15525 ;
  assign y5467 = ~n15528 ;
  assign y5468 = n15530 ;
  assign y5469 = n15532 ;
  assign y5470 = n15535 ;
  assign y5471 = ~n15537 ;
  assign y5472 = ~1'b0 ;
  assign y5473 = ~n15543 ;
  assign y5474 = ~n15545 ;
  assign y5475 = ~n15546 ;
  assign y5476 = ~n15549 ;
  assign y5477 = ~n15553 ;
  assign y5478 = ~n15555 ;
  assign y5479 = n15556 ;
  assign y5480 = n15557 ;
  assign y5481 = ~1'b0 ;
  assign y5482 = n15560 ;
  assign y5483 = ~n15563 ;
  assign y5484 = n15564 ;
  assign y5485 = ~n15569 ;
  assign y5486 = ~n15580 ;
  assign y5487 = ~n15582 ;
  assign y5488 = ~n15589 ;
  assign y5489 = ~n15591 ;
  assign y5490 = ~n15592 ;
  assign y5491 = ~n15597 ;
  assign y5492 = n1647 ;
  assign y5493 = ~n15599 ;
  assign y5494 = ~1'b0 ;
  assign y5495 = n15603 ;
  assign y5496 = ~n15609 ;
  assign y5497 = n15611 ;
  assign y5498 = ~n15614 ;
  assign y5499 = ~n15615 ;
  assign y5500 = ~n15618 ;
  assign y5501 = ~1'b0 ;
  assign y5502 = n15619 ;
  assign y5503 = ~n15620 ;
  assign y5504 = n15626 ;
  assign y5505 = n15628 ;
  assign y5506 = ~n15634 ;
  assign y5507 = ~1'b0 ;
  assign y5508 = ~1'b0 ;
  assign y5509 = ~n15636 ;
  assign y5510 = n15649 ;
  assign y5511 = n15650 ;
  assign y5512 = n15651 ;
  assign y5513 = n15652 ;
  assign y5514 = ~1'b0 ;
  assign y5515 = ~n15654 ;
  assign y5516 = ~n15658 ;
  assign y5517 = n15662 ;
  assign y5518 = ~n15665 ;
  assign y5519 = ~n15669 ;
  assign y5520 = n15674 ;
  assign y5521 = ~1'b0 ;
  assign y5522 = n15684 ;
  assign y5523 = ~n15690 ;
  assign y5524 = ~n15698 ;
  assign y5525 = ~n15701 ;
  assign y5526 = n8526 ;
  assign y5527 = ~n15706 ;
  assign y5528 = ~1'b0 ;
  assign y5529 = n15709 ;
  assign y5530 = ~1'b0 ;
  assign y5531 = ~n15715 ;
  assign y5532 = ~1'b0 ;
  assign y5533 = n15718 ;
  assign y5534 = n15725 ;
  assign y5535 = ~n15732 ;
  assign y5536 = n15735 ;
  assign y5537 = ~1'b0 ;
  assign y5538 = ~1'b0 ;
  assign y5539 = ~n3138 ;
  assign y5540 = ~n15736 ;
  assign y5541 = ~n15738 ;
  assign y5542 = ~n15743 ;
  assign y5543 = ~n15749 ;
  assign y5544 = ~n6231 ;
  assign y5545 = ~1'b0 ;
  assign y5546 = ~n15751 ;
  assign y5547 = ~n15752 ;
  assign y5548 = n15754 ;
  assign y5549 = ~n15756 ;
  assign y5550 = n15757 ;
  assign y5551 = ~n15763 ;
  assign y5552 = n15765 ;
  assign y5553 = n15768 ;
  assign y5554 = n15774 ;
  assign y5555 = n15776 ;
  assign y5556 = n15779 ;
  assign y5557 = ~n15780 ;
  assign y5558 = ~n15784 ;
  assign y5559 = ~n15790 ;
  assign y5560 = n15157 ;
  assign y5561 = n15792 ;
  assign y5562 = ~n15794 ;
  assign y5563 = ~1'b0 ;
  assign y5564 = ~1'b0 ;
  assign y5565 = n15795 ;
  assign y5566 = n1234 ;
  assign y5567 = n15796 ;
  assign y5568 = n15798 ;
  assign y5569 = n15806 ;
  assign y5570 = ~n15811 ;
  assign y5571 = n15815 ;
  assign y5572 = ~n15821 ;
  assign y5573 = n15823 ;
  assign y5574 = n15825 ;
  assign y5575 = ~n15827 ;
  assign y5576 = n15829 ;
  assign y5577 = ~n15835 ;
  assign y5578 = ~n15836 ;
  assign y5579 = ~n15843 ;
  assign y5580 = ~1'b0 ;
  assign y5581 = n15844 ;
  assign y5582 = n1862 ;
  assign y5583 = n15846 ;
  assign y5584 = n15848 ;
  assign y5585 = n15855 ;
  assign y5586 = ~1'b0 ;
  assign y5587 = n15858 ;
  assign y5588 = ~n15860 ;
  assign y5589 = ~n15863 ;
  assign y5590 = ~n15871 ;
  assign y5591 = ~n15872 ;
  assign y5592 = ~n15875 ;
  assign y5593 = ~n15880 ;
  assign y5594 = n15883 ;
  assign y5595 = ~n15884 ;
  assign y5596 = ~n15888 ;
  assign y5597 = ~n15891 ;
  assign y5598 = ~n15894 ;
  assign y5599 = ~n15902 ;
  assign y5600 = n15903 ;
  assign y5601 = ~1'b0 ;
  assign y5602 = ~n15906 ;
  assign y5603 = ~1'b0 ;
  assign y5604 = n15907 ;
  assign y5605 = n15912 ;
  assign y5606 = n15916 ;
  assign y5607 = n15920 ;
  assign y5608 = ~n15926 ;
  assign y5609 = 1'b0 ;
  assign y5610 = n15932 ;
  assign y5611 = ~n15939 ;
  assign y5612 = ~n15940 ;
  assign y5613 = ~n15943 ;
  assign y5614 = ~n15946 ;
  assign y5615 = ~1'b0 ;
  assign y5616 = ~n15947 ;
  assign y5617 = ~1'b0 ;
  assign y5618 = n15950 ;
  assign y5619 = n15951 ;
  assign y5620 = n15957 ;
  assign y5621 = ~n15974 ;
  assign y5622 = n15988 ;
  assign y5623 = ~1'b0 ;
  assign y5624 = ~1'b0 ;
  assign y5625 = ~n15994 ;
  assign y5626 = ~n15999 ;
  assign y5627 = ~n16003 ;
  assign y5628 = n16006 ;
  assign y5629 = n16019 ;
  assign y5630 = ~n7599 ;
  assign y5631 = n16021 ;
  assign y5632 = ~n16024 ;
  assign y5633 = n16029 ;
  assign y5634 = n16032 ;
  assign y5635 = ~n16033 ;
  assign y5636 = n4243 ;
  assign y5637 = ~1'b0 ;
  assign y5638 = ~n16034 ;
  assign y5639 = ~n16036 ;
  assign y5640 = n16038 ;
  assign y5641 = ~n16040 ;
  assign y5642 = ~n16042 ;
  assign y5643 = ~n16048 ;
  assign y5644 = ~n16049 ;
  assign y5645 = ~n16058 ;
  assign y5646 = n16064 ;
  assign y5647 = ~n16068 ;
  assign y5648 = ~n16069 ;
  assign y5649 = ~n16078 ;
  assign y5650 = ~1'b0 ;
  assign y5651 = ~n16089 ;
  assign y5652 = n16090 ;
  assign y5653 = ~n16092 ;
  assign y5654 = ~n16093 ;
  assign y5655 = ~n16099 ;
  assign y5656 = ~n16100 ;
  assign y5657 = ~1'b0 ;
  assign y5658 = n16105 ;
  assign y5659 = ~1'b0 ;
  assign y5660 = ~n16106 ;
  assign y5661 = n16109 ;
  assign y5662 = ~n16117 ;
  assign y5663 = ~n16120 ;
  assign y5664 = ~1'b0 ;
  assign y5665 = n16124 ;
  assign y5666 = ~n16125 ;
  assign y5667 = n16126 ;
  assign y5668 = ~1'b0 ;
  assign y5669 = ~1'b0 ;
  assign y5670 = ~n16133 ;
  assign y5671 = n16135 ;
  assign y5672 = ~n5062 ;
  assign y5673 = ~1'b0 ;
  assign y5674 = n16136 ;
  assign y5675 = ~n16140 ;
  assign y5676 = 1'b0 ;
  assign y5677 = n13481 ;
  assign y5678 = n16146 ;
  assign y5679 = ~1'b0 ;
  assign y5680 = ~n16147 ;
  assign y5681 = ~n16150 ;
  assign y5682 = ~n16152 ;
  assign y5683 = ~n13698 ;
  assign y5684 = n16155 ;
  assign y5685 = n16157 ;
  assign y5686 = n16159 ;
  assign y5687 = n7876 ;
  assign y5688 = n16163 ;
  assign y5689 = n16165 ;
  assign y5690 = ~n16168 ;
  assign y5691 = ~n16173 ;
  assign y5692 = ~1'b0 ;
  assign y5693 = n16177 ;
  assign y5694 = ~n16189 ;
  assign y5695 = ~1'b0 ;
  assign y5696 = n16194 ;
  assign y5697 = ~n16199 ;
  assign y5698 = ~1'b0 ;
  assign y5699 = ~n16204 ;
  assign y5700 = ~n16206 ;
  assign y5701 = n16207 ;
  assign y5702 = n16211 ;
  assign y5703 = ~n16216 ;
  assign y5704 = ~n16220 ;
  assign y5705 = n16229 ;
  assign y5706 = n16231 ;
  assign y5707 = ~n16232 ;
  assign y5708 = ~1'b0 ;
  assign y5709 = n16233 ;
  assign y5710 = ~1'b0 ;
  assign y5711 = ~1'b0 ;
  assign y5712 = n16234 ;
  assign y5713 = ~n16238 ;
  assign y5714 = ~n16239 ;
  assign y5715 = n16247 ;
  assign y5716 = ~n16250 ;
  assign y5717 = ~n16254 ;
  assign y5718 = ~1'b0 ;
  assign y5719 = n16256 ;
  assign y5720 = ~1'b0 ;
  assign y5721 = ~1'b0 ;
  assign y5722 = n16258 ;
  assign y5723 = ~n16263 ;
  assign y5724 = ~n16265 ;
  assign y5725 = n16266 ;
  assign y5726 = n16271 ;
  assign y5727 = n16277 ;
  assign y5728 = ~n16278 ;
  assign y5729 = ~1'b0 ;
  assign y5730 = n16281 ;
  assign y5731 = ~n16282 ;
  assign y5732 = ~1'b0 ;
  assign y5733 = ~n16284 ;
  assign y5734 = ~n16289 ;
  assign y5735 = n16290 ;
  assign y5736 = ~1'b0 ;
  assign y5737 = ~1'b0 ;
  assign y5738 = n16293 ;
  assign y5739 = ~n16294 ;
  assign y5740 = ~n16296 ;
  assign y5741 = n16298 ;
  assign y5742 = ~n16299 ;
  assign y5743 = n16300 ;
  assign y5744 = n7850 ;
  assign y5745 = ~1'b0 ;
  assign y5746 = n16303 ;
  assign y5747 = n16306 ;
  assign y5748 = n16309 ;
  assign y5749 = n16312 ;
  assign y5750 = n16313 ;
  assign y5751 = n16315 ;
  assign y5752 = ~n16317 ;
  assign y5753 = n16320 ;
  assign y5754 = n16321 ;
  assign y5755 = ~n16323 ;
  assign y5756 = ~n16327 ;
  assign y5757 = n16330 ;
  assign y5758 = ~1'b0 ;
  assign y5759 = n16336 ;
  assign y5760 = n16337 ;
  assign y5761 = n16340 ;
  assign y5762 = n16346 ;
  assign y5763 = ~1'b0 ;
  assign y5764 = n16352 ;
  assign y5765 = ~n16354 ;
  assign y5766 = ~n16358 ;
  assign y5767 = n16362 ;
  assign y5768 = ~n16363 ;
  assign y5769 = ~n16368 ;
  assign y5770 = ~n16378 ;
  assign y5771 = ~n16383 ;
  assign y5772 = n16385 ;
  assign y5773 = ~1'b0 ;
  assign y5774 = ~n16387 ;
  assign y5775 = n16388 ;
  assign y5776 = ~n16391 ;
  assign y5777 = ~n16392 ;
  assign y5778 = ~1'b0 ;
  assign y5779 = ~1'b0 ;
  assign y5780 = n16394 ;
  assign y5781 = n16397 ;
  assign y5782 = n16404 ;
  assign y5783 = ~n16405 ;
  assign y5784 = ~n16407 ;
  assign y5785 = n16408 ;
  assign y5786 = n16410 ;
  assign y5787 = ~n16412 ;
  assign y5788 = n16418 ;
  assign y5789 = ~n16420 ;
  assign y5790 = ~n16423 ;
  assign y5791 = ~n16430 ;
  assign y5792 = ~1'b0 ;
  assign y5793 = ~1'b0 ;
  assign y5794 = n16433 ;
  assign y5795 = ~n16434 ;
  assign y5796 = n16436 ;
  assign y5797 = ~n440 ;
  assign y5798 = ~n16437 ;
  assign y5799 = n16440 ;
  assign y5800 = n4449 ;
  assign y5801 = ~1'b0 ;
  assign y5802 = ~n16441 ;
  assign y5803 = ~n16447 ;
  assign y5804 = ~n16449 ;
  assign y5805 = ~1'b0 ;
  assign y5806 = n16450 ;
  assign y5807 = ~1'b0 ;
  assign y5808 = ~1'b0 ;
  assign y5809 = n16454 ;
  assign y5810 = ~n16455 ;
  assign y5811 = n16456 ;
  assign y5812 = n16470 ;
  assign y5813 = ~n16476 ;
  assign y5814 = n16477 ;
  assign y5815 = ~1'b0 ;
  assign y5816 = n16480 ;
  assign y5817 = ~1'b0 ;
  assign y5818 = ~n16482 ;
  assign y5819 = ~n16483 ;
  assign y5820 = ~n16485 ;
  assign y5821 = ~n16489 ;
  assign y5822 = n16490 ;
  assign y5823 = ~n16496 ;
  assign y5824 = n16499 ;
  assign y5825 = ~n16500 ;
  assign y5826 = ~n16431 ;
  assign y5827 = ~1'b0 ;
  assign y5828 = ~n16505 ;
  assign y5829 = ~n16508 ;
  assign y5830 = ~n16510 ;
  assign y5831 = ~n16514 ;
  assign y5832 = ~1'b0 ;
  assign y5833 = ~1'b0 ;
  assign y5834 = ~n9485 ;
  assign y5835 = ~n16518 ;
  assign y5836 = ~1'b0 ;
  assign y5837 = ~n16520 ;
  assign y5838 = ~n16524 ;
  assign y5839 = ~n16527 ;
  assign y5840 = ~n16528 ;
  assign y5841 = ~n16529 ;
  assign y5842 = n16530 ;
  assign y5843 = ~1'b0 ;
  assign y5844 = ~1'b0 ;
  assign y5845 = ~n16533 ;
  assign y5846 = ~n16535 ;
  assign y5847 = ~n16539 ;
  assign y5848 = ~n16542 ;
  assign y5849 = ~1'b0 ;
  assign y5850 = ~1'b0 ;
  assign y5851 = n16544 ;
  assign y5852 = n12607 ;
  assign y5853 = n16545 ;
  assign y5854 = ~1'b0 ;
  assign y5855 = ~n16546 ;
  assign y5856 = ~n16551 ;
  assign y5857 = ~n16553 ;
  assign y5858 = n16568 ;
  assign y5859 = n1465 ;
  assign y5860 = n16571 ;
  assign y5861 = ~1'b0 ;
  assign y5862 = n16575 ;
  assign y5863 = n16576 ;
  assign y5864 = ~1'b0 ;
  assign y5865 = ~n16577 ;
  assign y5866 = ~n16578 ;
  assign y5867 = ~n16589 ;
  assign y5868 = n16593 ;
  assign y5869 = n16594 ;
  assign y5870 = n16598 ;
  assign y5871 = ~1'b0 ;
  assign y5872 = n16601 ;
  assign y5873 = n16610 ;
  assign y5874 = n16611 ;
  assign y5875 = ~n16612 ;
  assign y5876 = ~1'b0 ;
  assign y5877 = ~n16622 ;
  assign y5878 = ~n16623 ;
  assign y5879 = n16628 ;
  assign y5880 = n16633 ;
  assign y5881 = n16638 ;
  assign y5882 = ~1'b0 ;
  assign y5883 = ~1'b0 ;
  assign y5884 = ~1'b0 ;
  assign y5885 = n16642 ;
  assign y5886 = n16647 ;
  assign y5887 = ~1'b0 ;
  assign y5888 = n16650 ;
  assign y5889 = n16653 ;
  assign y5890 = ~1'b0 ;
  assign y5891 = ~n16654 ;
  assign y5892 = n16660 ;
  assign y5893 = ~n16661 ;
  assign y5894 = n7102 ;
  assign y5895 = n16675 ;
  assign y5896 = n16678 ;
  assign y5897 = n16681 ;
  assign y5898 = n16684 ;
  assign y5899 = n16685 ;
  assign y5900 = n16688 ;
  assign y5901 = ~1'b0 ;
  assign y5902 = n16689 ;
  assign y5903 = n16691 ;
  assign y5904 = ~n5606 ;
  assign y5905 = ~n16693 ;
  assign y5906 = n16704 ;
  assign y5907 = n16711 ;
  assign y5908 = ~n16720 ;
  assign y5909 = ~n16722 ;
  assign y5910 = ~n16726 ;
  assign y5911 = n16730 ;
  assign y5912 = n16734 ;
  assign y5913 = ~1'b0 ;
  assign y5914 = n16742 ;
  assign y5915 = ~n16746 ;
  assign y5916 = ~1'b0 ;
  assign y5917 = n16748 ;
  assign y5918 = n16749 ;
  assign y5919 = ~n16751 ;
  assign y5920 = ~1'b0 ;
  assign y5921 = n16756 ;
  assign y5922 = n16758 ;
  assign y5923 = n16761 ;
  assign y5924 = ~n16763 ;
  assign y5925 = n16770 ;
  assign y5926 = ~n16771 ;
  assign y5927 = ~n16785 ;
  assign y5928 = ~n16789 ;
  assign y5929 = n16790 ;
  assign y5930 = n16794 ;
  assign y5931 = ~n16795 ;
  assign y5932 = ~1'b0 ;
  assign y5933 = n16796 ;
  assign y5934 = ~1'b0 ;
  assign y5935 = ~1'b0 ;
  assign y5936 = ~1'b0 ;
  assign y5937 = n16802 ;
  assign y5938 = ~n16804 ;
  assign y5939 = ~n16807 ;
  assign y5940 = ~1'b0 ;
  assign y5941 = ~n16816 ;
  assign y5942 = n16817 ;
  assign y5943 = ~n16819 ;
  assign y5944 = ~n16825 ;
  assign y5945 = ~n16829 ;
  assign y5946 = n16833 ;
  assign y5947 = ~n16836 ;
  assign y5948 = n16839 ;
  assign y5949 = n16849 ;
  assign y5950 = ~n16851 ;
  assign y5951 = ~n16854 ;
  assign y5952 = n16857 ;
  assign y5953 = ~1'b0 ;
  assign y5954 = ~1'b0 ;
  assign y5955 = ~1'b0 ;
  assign y5956 = n16859 ;
  assign y5957 = ~n16861 ;
  assign y5958 = ~n16865 ;
  assign y5959 = ~n16872 ;
  assign y5960 = ~n16880 ;
  assign y5961 = ~1'b0 ;
  assign y5962 = ~1'b0 ;
  assign y5963 = n16882 ;
  assign y5964 = n16885 ;
  assign y5965 = ~1'b0 ;
  assign y5966 = ~n16889 ;
  assign y5967 = ~1'b0 ;
  assign y5968 = n16891 ;
  assign y5969 = ~n16892 ;
  assign y5970 = n16893 ;
  assign y5971 = ~n16897 ;
  assign y5972 = n16901 ;
  assign y5973 = ~n16903 ;
  assign y5974 = ~n16905 ;
  assign y5975 = ~n16906 ;
  assign y5976 = n16907 ;
  assign y5977 = ~n15568 ;
  assign y5978 = ~1'b0 ;
  assign y5979 = n16909 ;
  assign y5980 = ~n16914 ;
  assign y5981 = ~n16915 ;
  assign y5982 = n16929 ;
  assign y5983 = ~n16931 ;
  assign y5984 = n16932 ;
  assign y5985 = n13626 ;
  assign y5986 = ~1'b0 ;
  assign y5987 = ~1'b0 ;
  assign y5988 = ~n16940 ;
  assign y5989 = n16943 ;
  assign y5990 = ~n16945 ;
  assign y5991 = ~n16953 ;
  assign y5992 = ~n16958 ;
  assign y5993 = ~n16962 ;
  assign y5994 = ~n16965 ;
  assign y5995 = n16966 ;
  assign y5996 = ~n16968 ;
  assign y5997 = n16970 ;
  assign y5998 = ~n16973 ;
  assign y5999 = n16976 ;
  assign y6000 = n16978 ;
  assign y6001 = ~n14138 ;
  assign y6002 = ~n16987 ;
  assign y6003 = n16994 ;
  assign y6004 = n17004 ;
  assign y6005 = ~n17006 ;
  assign y6006 = ~n17011 ;
  assign y6007 = ~n17014 ;
  assign y6008 = ~n17017 ;
  assign y6009 = ~1'b0 ;
  assign y6010 = ~n17020 ;
  assign y6011 = n17022 ;
  assign y6012 = 1'b0 ;
  assign y6013 = n17023 ;
  assign y6014 = ~n17025 ;
  assign y6015 = ~n17027 ;
  assign y6016 = ~n17029 ;
  assign y6017 = n17038 ;
  assign y6018 = n17043 ;
  assign y6019 = n17044 ;
  assign y6020 = ~1'b0 ;
  assign y6021 = n17045 ;
  assign y6022 = ~n17047 ;
  assign y6023 = ~1'b0 ;
  assign y6024 = ~1'b0 ;
  assign y6025 = ~1'b0 ;
  assign y6026 = n17053 ;
  assign y6027 = n17055 ;
  assign y6028 = ~1'b0 ;
  assign y6029 = n17059 ;
  assign y6030 = ~n17063 ;
  assign y6031 = n17066 ;
  assign y6032 = ~1'b0 ;
  assign y6033 = ~n17067 ;
  assign y6034 = ~1'b0 ;
  assign y6035 = ~1'b0 ;
  assign y6036 = ~n17068 ;
  assign y6037 = n17069 ;
  assign y6038 = ~n17072 ;
  assign y6039 = ~1'b0 ;
  assign y6040 = ~n17074 ;
  assign y6041 = n17075 ;
  assign y6042 = ~n17078 ;
  assign y6043 = ~n17080 ;
  assign y6044 = n17081 ;
  assign y6045 = ~n17084 ;
  assign y6046 = ~n17088 ;
  assign y6047 = n13920 ;
  assign y6048 = ~n17095 ;
  assign y6049 = ~n17099 ;
  assign y6050 = ~n17101 ;
  assign y6051 = n17107 ;
  assign y6052 = ~n17108 ;
  assign y6053 = n17117 ;
  assign y6054 = n17126 ;
  assign y6055 = ~1'b0 ;
  assign y6056 = n17128 ;
  assign y6057 = ~1'b0 ;
  assign y6058 = n17131 ;
  assign y6059 = ~n17133 ;
  assign y6060 = ~n6706 ;
  assign y6061 = n17137 ;
  assign y6062 = ~n17138 ;
  assign y6063 = n17142 ;
  assign y6064 = ~1'b0 ;
  assign y6065 = ~1'b0 ;
  assign y6066 = ~n17147 ;
  assign y6067 = ~n17148 ;
  assign y6068 = ~n17150 ;
  assign y6069 = n17152 ;
  assign y6070 = n5996 ;
  assign y6071 = ~n17153 ;
  assign y6072 = n17155 ;
  assign y6073 = n17156 ;
  assign y6074 = n17159 ;
  assign y6075 = n17165 ;
  assign y6076 = ~n17166 ;
  assign y6077 = ~n17171 ;
  assign y6078 = ~1'b0 ;
  assign y6079 = 1'b0 ;
  assign y6080 = ~n17172 ;
  assign y6081 = ~n17182 ;
  assign y6082 = ~n17187 ;
  assign y6083 = ~1'b0 ;
  assign y6084 = n17189 ;
  assign y6085 = ~n17192 ;
  assign y6086 = ~n8043 ;
  assign y6087 = ~1'b0 ;
  assign y6088 = n17193 ;
  assign y6089 = n17196 ;
  assign y6090 = n17197 ;
  assign y6091 = ~n17201 ;
  assign y6092 = ~n17204 ;
  assign y6093 = ~n17211 ;
  assign y6094 = ~n17214 ;
  assign y6095 = ~n17221 ;
  assign y6096 = ~1'b0 ;
  assign y6097 = ~1'b0 ;
  assign y6098 = n17224 ;
  assign y6099 = n17225 ;
  assign y6100 = ~1'b0 ;
  assign y6101 = ~n17227 ;
  assign y6102 = ~n17229 ;
  assign y6103 = ~n17231 ;
  assign y6104 = n17238 ;
  assign y6105 = n17239 ;
  assign y6106 = n17242 ;
  assign y6107 = ~1'b0 ;
  assign y6108 = ~n17243 ;
  assign y6109 = ~1'b0 ;
  assign y6110 = n17245 ;
  assign y6111 = ~n17248 ;
  assign y6112 = ~n17259 ;
  assign y6113 = ~n17261 ;
  assign y6114 = ~1'b0 ;
  assign y6115 = ~1'b0 ;
  assign y6116 = ~n17263 ;
  assign y6117 = n17266 ;
  assign y6118 = ~1'b0 ;
  assign y6119 = ~n17270 ;
  assign y6120 = n17271 ;
  assign y6121 = n17276 ;
  assign y6122 = ~n17281 ;
  assign y6123 = ~1'b0 ;
  assign y6124 = n3746 ;
  assign y6125 = ~n17287 ;
  assign y6126 = n17288 ;
  assign y6127 = ~n17289 ;
  assign y6128 = ~n17297 ;
  assign y6129 = n17306 ;
  assign y6130 = n17308 ;
  assign y6131 = ~n17311 ;
  assign y6132 = n17314 ;
  assign y6133 = ~1'b0 ;
  assign y6134 = n17317 ;
  assign y6135 = ~1'b0 ;
  assign y6136 = ~n17320 ;
  assign y6137 = ~n17322 ;
  assign y6138 = ~n17324 ;
  assign y6139 = ~n17325 ;
  assign y6140 = ~1'b0 ;
  assign y6141 = ~1'b0 ;
  assign y6142 = n17329 ;
  assign y6143 = n17331 ;
  assign y6144 = ~n17332 ;
  assign y6145 = ~n17334 ;
  assign y6146 = ~1'b0 ;
  assign y6147 = ~n17337 ;
  assign y6148 = ~n17344 ;
  assign y6149 = n17349 ;
  assign y6150 = ~1'b0 ;
  assign y6151 = ~n17350 ;
  assign y6152 = n17352 ;
  assign y6153 = n17356 ;
  assign y6154 = ~n17357 ;
  assign y6155 = n17358 ;
  assign y6156 = ~n17359 ;
  assign y6157 = ~n17362 ;
  assign y6158 = ~1'b0 ;
  assign y6159 = n17364 ;
  assign y6160 = 1'b0 ;
  assign y6161 = ~1'b0 ;
  assign y6162 = ~n17368 ;
  assign y6163 = n17369 ;
  assign y6164 = n17370 ;
  assign y6165 = n17372 ;
  assign y6166 = ~n17373 ;
  assign y6167 = ~1'b0 ;
  assign y6168 = n17376 ;
  assign y6169 = ~1'b0 ;
  assign y6170 = n17377 ;
  assign y6171 = ~1'b0 ;
  assign y6172 = n17386 ;
  assign y6173 = ~1'b0 ;
  assign y6174 = 1'b0 ;
  assign y6175 = n17389 ;
  assign y6176 = n17391 ;
  assign y6177 = n17392 ;
  assign y6178 = n17396 ;
  assign y6179 = ~1'b0 ;
  assign y6180 = n17399 ;
  assign y6181 = ~1'b0 ;
  assign y6182 = ~n17409 ;
  assign y6183 = ~n17413 ;
  assign y6184 = n17418 ;
  assign y6185 = ~n17420 ;
  assign y6186 = ~1'b0 ;
  assign y6187 = n17422 ;
  assign y6188 = ~n17424 ;
  assign y6189 = ~n17425 ;
  assign y6190 = n2818 ;
  assign y6191 = ~n17436 ;
  assign y6192 = ~n17438 ;
  assign y6193 = ~n17440 ;
  assign y6194 = n17448 ;
  assign y6195 = ~n17454 ;
  assign y6196 = n17457 ;
  assign y6197 = n17460 ;
  assign y6198 = n17462 ;
  assign y6199 = ~1'b0 ;
  assign y6200 = n17464 ;
  assign y6201 = ~n17469 ;
  assign y6202 = n17470 ;
  assign y6203 = ~n5931 ;
  assign y6204 = ~1'b0 ;
  assign y6205 = n17473 ;
  assign y6206 = ~1'b0 ;
  assign y6207 = n17475 ;
  assign y6208 = ~n17477 ;
  assign y6209 = ~1'b0 ;
  assign y6210 = n17479 ;
  assign y6211 = ~n17484 ;
  assign y6212 = n17488 ;
  assign y6213 = ~n17489 ;
  assign y6214 = ~n17498 ;
  assign y6215 = ~n17499 ;
  assign y6216 = ~n17503 ;
  assign y6217 = ~n17505 ;
  assign y6218 = ~n4326 ;
  assign y6219 = ~1'b0 ;
  assign y6220 = n17506 ;
  assign y6221 = ~1'b0 ;
  assign y6222 = ~n17508 ;
  assign y6223 = n17511 ;
  assign y6224 = n17515 ;
  assign y6225 = ~n17518 ;
  assign y6226 = ~1'b0 ;
  assign y6227 = ~1'b0 ;
  assign y6228 = ~1'b0 ;
  assign y6229 = n17521 ;
  assign y6230 = n17529 ;
  assign y6231 = ~n17533 ;
  assign y6232 = ~n17539 ;
  assign y6233 = ~n17541 ;
  assign y6234 = ~n17546 ;
  assign y6235 = ~1'b0 ;
  assign y6236 = n17547 ;
  assign y6237 = n17550 ;
  assign y6238 = ~1'b0 ;
  assign y6239 = n17555 ;
  assign y6240 = ~n17557 ;
  assign y6241 = ~n17558 ;
  assign y6242 = ~n17560 ;
  assign y6243 = ~n17561 ;
  assign y6244 = ~n17562 ;
  assign y6245 = n17568 ;
  assign y6246 = ~n17570 ;
  assign y6247 = ~n17576 ;
  assign y6248 = ~n17583 ;
  assign y6249 = n17585 ;
  assign y6250 = ~n17591 ;
  assign y6251 = ~n17593 ;
  assign y6252 = n17594 ;
  assign y6253 = n17597 ;
  assign y6254 = n17600 ;
  assign y6255 = ~n17604 ;
  assign y6256 = n17606 ;
  assign y6257 = ~n17608 ;
  assign y6258 = n17613 ;
  assign y6259 = 1'b0 ;
  assign y6260 = ~n17614 ;
  assign y6261 = n17616 ;
  assign y6262 = ~n17618 ;
  assign y6263 = ~n17623 ;
  assign y6264 = ~1'b0 ;
  assign y6265 = ~n17627 ;
  assign y6266 = ~n17628 ;
  assign y6267 = ~1'b0 ;
  assign y6268 = n17630 ;
  assign y6269 = n15661 ;
  assign y6270 = ~n17632 ;
  assign y6271 = n17633 ;
  assign y6272 = ~n17638 ;
  assign y6273 = ~n17642 ;
  assign y6274 = n10191 ;
  assign y6275 = ~n17643 ;
  assign y6276 = ~n17645 ;
  assign y6277 = ~n17646 ;
  assign y6278 = ~n17658 ;
  assign y6279 = n17665 ;
  assign y6280 = n17666 ;
  assign y6281 = ~n932 ;
  assign y6282 = n17670 ;
  assign y6283 = ~1'b0 ;
  assign y6284 = ~1'b0 ;
  assign y6285 = n17678 ;
  assign y6286 = ~n17681 ;
  assign y6287 = n17682 ;
  assign y6288 = ~n17689 ;
  assign y6289 = n17690 ;
  assign y6290 = ~n17695 ;
  assign y6291 = n17697 ;
  assign y6292 = n17700 ;
  assign y6293 = ~1'b0 ;
  assign y6294 = ~n17707 ;
  assign y6295 = n17708 ;
  assign y6296 = n17711 ;
  assign y6297 = ~n17723 ;
  assign y6298 = ~n17726 ;
  assign y6299 = ~n17729 ;
  assign y6300 = ~n17735 ;
  assign y6301 = n17739 ;
  assign y6302 = ~1'b0 ;
  assign y6303 = ~n17740 ;
  assign y6304 = ~n17744 ;
  assign y6305 = ~n17748 ;
  assign y6306 = ~1'b0 ;
  assign y6307 = ~n17750 ;
  assign y6308 = 1'b0 ;
  assign y6309 = n17754 ;
  assign y6310 = ~n17755 ;
  assign y6311 = ~n17756 ;
  assign y6312 = ~1'b0 ;
  assign y6313 = ~n17764 ;
  assign y6314 = n17778 ;
  assign y6315 = ~n17786 ;
  assign y6316 = ~1'b0 ;
  assign y6317 = ~1'b0 ;
  assign y6318 = n17792 ;
  assign y6319 = n17797 ;
  assign y6320 = ~n17798 ;
  assign y6321 = n17801 ;
  assign y6322 = ~n17803 ;
  assign y6323 = ~n17812 ;
  assign y6324 = ~1'b0 ;
  assign y6325 = n17819 ;
  assign y6326 = n17820 ;
  assign y6327 = ~n17824 ;
  assign y6328 = ~n17827 ;
  assign y6329 = n17828 ;
  assign y6330 = ~n17830 ;
  assign y6331 = n17831 ;
  assign y6332 = n17835 ;
  assign y6333 = ~1'b0 ;
  assign y6334 = ~n17836 ;
  assign y6335 = ~1'b0 ;
  assign y6336 = ~n17838 ;
  assign y6337 = ~n17839 ;
  assign y6338 = ~n17840 ;
  assign y6339 = n17842 ;
  assign y6340 = ~n17844 ;
  assign y6341 = n17845 ;
  assign y6342 = n17848 ;
  assign y6343 = ~1'b0 ;
  assign y6344 = n17849 ;
  assign y6345 = ~n17857 ;
  assign y6346 = n17865 ;
  assign y6347 = ~n17868 ;
  assign y6348 = n17872 ;
  assign y6349 = n17875 ;
  assign y6350 = ~n17878 ;
  assign y6351 = ~n17884 ;
  assign y6352 = n17885 ;
  assign y6353 = n17889 ;
  assign y6354 = ~n17890 ;
  assign y6355 = n17904 ;
  assign y6356 = ~1'b0 ;
  assign y6357 = 1'b0 ;
  assign y6358 = ~n17910 ;
  assign y6359 = ~n17917 ;
  assign y6360 = ~1'b0 ;
  assign y6361 = n17924 ;
  assign y6362 = ~n17925 ;
  assign y6363 = ~n17929 ;
  assign y6364 = ~1'b0 ;
  assign y6365 = ~n17936 ;
  assign y6366 = n17938 ;
  assign y6367 = ~n17941 ;
  assign y6368 = n17942 ;
  assign y6369 = n17949 ;
  assign y6370 = ~1'b0 ;
  assign y6371 = 1'b0 ;
  assign y6372 = ~1'b0 ;
  assign y6373 = ~n17951 ;
  assign y6374 = n17955 ;
  assign y6375 = n17963 ;
  assign y6376 = n17964 ;
  assign y6377 = ~n17968 ;
  assign y6378 = n17976 ;
  assign y6379 = n17978 ;
  assign y6380 = ~n17984 ;
  assign y6381 = ~n17985 ;
  assign y6382 = 1'b0 ;
  assign y6383 = ~1'b0 ;
  assign y6384 = n5072 ;
  assign y6385 = ~n17991 ;
  assign y6386 = ~1'b0 ;
  assign y6387 = ~n17997 ;
  assign y6388 = ~n18007 ;
  assign y6389 = ~n18010 ;
  assign y6390 = ~n18012 ;
  assign y6391 = ~1'b0 ;
  assign y6392 = n18013 ;
  assign y6393 = ~n18017 ;
  assign y6394 = n18021 ;
  assign y6395 = n18023 ;
  assign y6396 = n18025 ;
  assign y6397 = ~n18030 ;
  assign y6398 = n18034 ;
  assign y6399 = ~n18036 ;
  assign y6400 = ~1'b0 ;
  assign y6401 = n18037 ;
  assign y6402 = ~1'b0 ;
  assign y6403 = n18039 ;
  assign y6404 = n18040 ;
  assign y6405 = ~n18042 ;
  assign y6406 = ~n18051 ;
  assign y6407 = ~n18059 ;
  assign y6408 = ~1'b0 ;
  assign y6409 = n18062 ;
  assign y6410 = ~n18063 ;
  assign y6411 = ~n18065 ;
  assign y6412 = ~1'b0 ;
  assign y6413 = ~n18068 ;
  assign y6414 = ~n18070 ;
  assign y6415 = ~n1935 ;
  assign y6416 = n18073 ;
  assign y6417 = n2515 ;
  assign y6418 = ~n18075 ;
  assign y6419 = n18081 ;
  assign y6420 = ~1'b0 ;
  assign y6421 = ~n18084 ;
  assign y6422 = n18090 ;
  assign y6423 = n18095 ;
  assign y6424 = n17279 ;
  assign y6425 = ~1'b0 ;
  assign y6426 = ~n18096 ;
  assign y6427 = n18097 ;
  assign y6428 = ~n18104 ;
  assign y6429 = ~n18107 ;
  assign y6430 = ~n10121 ;
  assign y6431 = n18111 ;
  assign y6432 = n18115 ;
  assign y6433 = n18120 ;
  assign y6434 = ~1'b0 ;
  assign y6435 = ~n18124 ;
  assign y6436 = n18125 ;
  assign y6437 = n18126 ;
  assign y6438 = n8774 ;
  assign y6439 = ~1'b0 ;
  assign y6440 = ~n18129 ;
  assign y6441 = n18132 ;
  assign y6442 = ~n18136 ;
  assign y6443 = ~1'b0 ;
  assign y6444 = ~n18137 ;
  assign y6445 = n18143 ;
  assign y6446 = ~1'b0 ;
  assign y6447 = ~n18144 ;
  assign y6448 = ~n18149 ;
  assign y6449 = n18153 ;
  assign y6450 = n18158 ;
  assign y6451 = ~n18160 ;
  assign y6452 = n18161 ;
  assign y6453 = ~n18162 ;
  assign y6454 = ~1'b0 ;
  assign y6455 = n18164 ;
  assign y6456 = n12656 ;
  assign y6457 = ~n18166 ;
  assign y6458 = n7545 ;
  assign y6459 = ~n18167 ;
  assign y6460 = n18168 ;
  assign y6461 = ~n18170 ;
  assign y6462 = n18171 ;
  assign y6463 = n8719 ;
  assign y6464 = ~n18172 ;
  assign y6465 = n18174 ;
  assign y6466 = n18177 ;
  assign y6467 = n18178 ;
  assign y6468 = ~n18180 ;
  assign y6469 = ~n18181 ;
  assign y6470 = ~n18186 ;
  assign y6471 = ~n18187 ;
  assign y6472 = n18190 ;
  assign y6473 = ~n18191 ;
  assign y6474 = ~n18196 ;
  assign y6475 = ~n18198 ;
  assign y6476 = ~n18200 ;
  assign y6477 = ~n18202 ;
  assign y6478 = ~n18204 ;
  assign y6479 = ~n18206 ;
  assign y6480 = ~n18209 ;
  assign y6481 = ~n18211 ;
  assign y6482 = n15778 ;
  assign y6483 = n18214 ;
  assign y6484 = n18229 ;
  assign y6485 = n18233 ;
  assign y6486 = ~n18235 ;
  assign y6487 = n18236 ;
  assign y6488 = ~1'b0 ;
  assign y6489 = ~n18239 ;
  assign y6490 = ~n18242 ;
  assign y6491 = ~1'b0 ;
  assign y6492 = n18247 ;
  assign y6493 = ~n18248 ;
  assign y6494 = n18251 ;
  assign y6495 = n18253 ;
  assign y6496 = n18257 ;
  assign y6497 = ~n18259 ;
  assign y6498 = n18260 ;
  assign y6499 = ~1'b0 ;
  assign y6500 = ~n18268 ;
  assign y6501 = n18274 ;
  assign y6502 = ~n18277 ;
  assign y6503 = n18284 ;
  assign y6504 = n18287 ;
  assign y6505 = n18296 ;
  assign y6506 = ~1'b0 ;
  assign y6507 = ~n18297 ;
  assign y6508 = ~n18299 ;
  assign y6509 = n18300 ;
  assign y6510 = ~1'b0 ;
  assign y6511 = ~n18312 ;
  assign y6512 = n18313 ;
  assign y6513 = ~n18317 ;
  assign y6514 = ~n18318 ;
  assign y6515 = ~n18319 ;
  assign y6516 = n18323 ;
  assign y6517 = ~n18326 ;
  assign y6518 = ~n18329 ;
  assign y6519 = ~n18333 ;
  assign y6520 = ~n18337 ;
  assign y6521 = n18342 ;
  assign y6522 = n18343 ;
  assign y6523 = n18345 ;
  assign y6524 = ~n18349 ;
  assign y6525 = n18352 ;
  assign y6526 = ~n18353 ;
  assign y6527 = n18356 ;
  assign y6528 = ~n18359 ;
  assign y6529 = 1'b0 ;
  assign y6530 = n18363 ;
  assign y6531 = ~1'b0 ;
  assign y6532 = n18368 ;
  assign y6533 = n18371 ;
  assign y6534 = n18376 ;
  assign y6535 = n18382 ;
  assign y6536 = n18383 ;
  assign y6537 = n18388 ;
  assign y6538 = ~n18390 ;
  assign y6539 = n18396 ;
  assign y6540 = ~n18398 ;
  assign y6541 = ~n18399 ;
  assign y6542 = n18400 ;
  assign y6543 = ~n18402 ;
  assign y6544 = ~n11159 ;
  assign y6545 = n18403 ;
  assign y6546 = n18406 ;
  assign y6547 = n18407 ;
  assign y6548 = ~n18412 ;
  assign y6549 = 1'b0 ;
  assign y6550 = ~n18415 ;
  assign y6551 = n18420 ;
  assign y6552 = ~n18423 ;
  assign y6553 = n18425 ;
  assign y6554 = ~1'b0 ;
  assign y6555 = ~n18429 ;
  assign y6556 = ~n18433 ;
  assign y6557 = n18436 ;
  assign y6558 = n18438 ;
  assign y6559 = ~n18441 ;
  assign y6560 = n18444 ;
  assign y6561 = n18452 ;
  assign y6562 = n18459 ;
  assign y6563 = n18463 ;
  assign y6564 = ~n18464 ;
  assign y6565 = n18465 ;
  assign y6566 = ~n18468 ;
  assign y6567 = n18474 ;
  assign y6568 = ~n18475 ;
  assign y6569 = ~n18477 ;
  assign y6570 = n18480 ;
  assign y6571 = ~n18487 ;
  assign y6572 = n18489 ;
  assign y6573 = n18491 ;
  assign y6574 = n18494 ;
  assign y6575 = ~n18505 ;
  assign y6576 = n18506 ;
  assign y6577 = ~1'b0 ;
  assign y6578 = n18513 ;
  assign y6579 = ~1'b0 ;
  assign y6580 = ~n18515 ;
  assign y6581 = ~1'b0 ;
  assign y6582 = n18520 ;
  assign y6583 = ~n18523 ;
  assign y6584 = ~n18526 ;
  assign y6585 = ~1'b0 ;
  assign y6586 = ~1'b0 ;
  assign y6587 = ~1'b0 ;
  assign y6588 = ~n18533 ;
  assign y6589 = ~n18534 ;
  assign y6590 = ~n18535 ;
  assign y6591 = ~n18537 ;
  assign y6592 = n18541 ;
  assign y6593 = n18547 ;
  assign y6594 = n18549 ;
  assign y6595 = ~n18553 ;
  assign y6596 = n17343 ;
  assign y6597 = ~n18555 ;
  assign y6598 = n18558 ;
  assign y6599 = ~n18562 ;
  assign y6600 = ~n18566 ;
  assign y6601 = ~1'b0 ;
  assign y6602 = ~1'b0 ;
  assign y6603 = n9553 ;
  assign y6604 = ~1'b0 ;
  assign y6605 = ~1'b0 ;
  assign y6606 = n3050 ;
  assign y6607 = ~1'b0 ;
  assign y6608 = ~n18567 ;
  assign y6609 = n18571 ;
  assign y6610 = n3690 ;
  assign y6611 = ~n18582 ;
  assign y6612 = n10208 ;
  assign y6613 = ~1'b0 ;
  assign y6614 = n18583 ;
  assign y6615 = ~1'b0 ;
  assign y6616 = n18585 ;
  assign y6617 = n18589 ;
  assign y6618 = ~1'b0 ;
  assign y6619 = n18590 ;
  assign y6620 = ~n18596 ;
  assign y6621 = n18601 ;
  assign y6622 = ~n18606 ;
  assign y6623 = ~n18610 ;
  assign y6624 = n18620 ;
  assign y6625 = n18625 ;
  assign y6626 = ~n18627 ;
  assign y6627 = n18629 ;
  assign y6628 = n18633 ;
  assign y6629 = ~1'b0 ;
  assign y6630 = ~n18637 ;
  assign y6631 = ~1'b0 ;
  assign y6632 = n18644 ;
  assign y6633 = ~1'b0 ;
  assign y6634 = n12136 ;
  assign y6635 = ~n18645 ;
  assign y6636 = n18650 ;
  assign y6637 = ~n18658 ;
  assign y6638 = ~1'b0 ;
  assign y6639 = ~n18662 ;
  assign y6640 = n18664 ;
  assign y6641 = ~1'b0 ;
  assign y6642 = ~n18665 ;
  assign y6643 = ~1'b0 ;
  assign y6644 = ~1'b0 ;
  assign y6645 = ~n18670 ;
  assign y6646 = ~1'b0 ;
  assign y6647 = ~n18679 ;
  assign y6648 = n18681 ;
  assign y6649 = ~1'b0 ;
  assign y6650 = n18683 ;
  assign y6651 = ~n18686 ;
  assign y6652 = ~1'b0 ;
  assign y6653 = ~n18689 ;
  assign y6654 = ~n18692 ;
  assign y6655 = ~1'b0 ;
  assign y6656 = n18698 ;
  assign y6657 = ~1'b0 ;
  assign y6658 = n18707 ;
  assign y6659 = ~n18708 ;
  assign y6660 = ~n18715 ;
  assign y6661 = ~1'b0 ;
  assign y6662 = ~n18716 ;
  assign y6663 = n18720 ;
  assign y6664 = n18721 ;
  assign y6665 = ~n18725 ;
  assign y6666 = n18731 ;
  assign y6667 = ~1'b0 ;
  assign y6668 = ~n18733 ;
  assign y6669 = n18737 ;
  assign y6670 = ~1'b0 ;
  assign y6671 = n18739 ;
  assign y6672 = ~n18744 ;
  assign y6673 = ~n18750 ;
  assign y6674 = ~1'b0 ;
  assign y6675 = ~n18751 ;
  assign y6676 = ~n18757 ;
  assign y6677 = ~n18758 ;
  assign y6678 = ~1'b0 ;
  assign y6679 = ~1'b0 ;
  assign y6680 = ~n18759 ;
  assign y6681 = ~n3471 ;
  assign y6682 = ~1'b0 ;
  assign y6683 = ~n18762 ;
  assign y6684 = n18771 ;
  assign y6685 = n18772 ;
  assign y6686 = ~n18778 ;
  assign y6687 = ~1'b0 ;
  assign y6688 = n14157 ;
  assign y6689 = n18780 ;
  assign y6690 = ~1'b0 ;
  assign y6691 = ~n18782 ;
  assign y6692 = ~n18784 ;
  assign y6693 = ~n18788 ;
  assign y6694 = ~n18790 ;
  assign y6695 = n18800 ;
  assign y6696 = n18801 ;
  assign y6697 = ~n18806 ;
  assign y6698 = ~1'b0 ;
  assign y6699 = ~n18810 ;
  assign y6700 = ~n18813 ;
  assign y6701 = ~n18816 ;
  assign y6702 = n18822 ;
  assign y6703 = ~n18828 ;
  assign y6704 = ~1'b0 ;
  assign y6705 = ~1'b0 ;
  assign y6706 = n18832 ;
  assign y6707 = n18833 ;
  assign y6708 = n18839 ;
  assign y6709 = ~1'b0 ;
  assign y6710 = ~1'b0 ;
  assign y6711 = ~1'b0 ;
  assign y6712 = n18846 ;
  assign y6713 = n18849 ;
  assign y6714 = ~1'b0 ;
  assign y6715 = ~n18852 ;
  assign y6716 = ~n18853 ;
  assign y6717 = ~n18854 ;
  assign y6718 = ~n18858 ;
  assign y6719 = ~1'b0 ;
  assign y6720 = n18860 ;
  assign y6721 = n18870 ;
  assign y6722 = ~n18872 ;
  assign y6723 = ~1'b0 ;
  assign y6724 = ~1'b0 ;
  assign y6725 = n18875 ;
  assign y6726 = ~1'b0 ;
  assign y6727 = n18877 ;
  assign y6728 = ~n18879 ;
  assign y6729 = ~1'b0 ;
  assign y6730 = n18880 ;
  assign y6731 = ~n18881 ;
  assign y6732 = ~1'b0 ;
  assign y6733 = ~n18882 ;
  assign y6734 = n18887 ;
  assign y6735 = n18889 ;
  assign y6736 = ~n18894 ;
  assign y6737 = ~n18895 ;
  assign y6738 = ~n18899 ;
  assign y6739 = n18900 ;
  assign y6740 = ~n18905 ;
  assign y6741 = n18907 ;
  assign y6742 = ~n18911 ;
  assign y6743 = ~n18913 ;
  assign y6744 = ~n18914 ;
  assign y6745 = ~n18918 ;
  assign y6746 = n18919 ;
  assign y6747 = ~n18922 ;
  assign y6748 = ~1'b0 ;
  assign y6749 = n18923 ;
  assign y6750 = ~n18927 ;
  assign y6751 = ~1'b0 ;
  assign y6752 = ~n18929 ;
  assign y6753 = ~n18933 ;
  assign y6754 = ~n18935 ;
  assign y6755 = n18941 ;
  assign y6756 = ~n15085 ;
  assign y6757 = ~n18942 ;
  assign y6758 = ~n18946 ;
  assign y6759 = ~n1243 ;
  assign y6760 = ~n18948 ;
  assign y6761 = ~n18952 ;
  assign y6762 = n18955 ;
  assign y6763 = ~1'b0 ;
  assign y6764 = n18956 ;
  assign y6765 = ~n18958 ;
  assign y6766 = ~n18962 ;
  assign y6767 = ~1'b0 ;
  assign y6768 = ~1'b0 ;
  assign y6769 = n18965 ;
  assign y6770 = ~1'b0 ;
  assign y6771 = ~1'b0 ;
  assign y6772 = ~n18968 ;
  assign y6773 = n18969 ;
  assign y6774 = ~n18971 ;
  assign y6775 = n18974 ;
  assign y6776 = ~n18978 ;
  assign y6777 = ~1'b0 ;
  assign y6778 = ~1'b0 ;
  assign y6779 = ~n18979 ;
  assign y6780 = ~n18987 ;
  assign y6781 = ~n1882 ;
  assign y6782 = n18991 ;
  assign y6783 = ~1'b0 ;
  assign y6784 = ~n18995 ;
  assign y6785 = ~1'b0 ;
  assign y6786 = ~1'b0 ;
  assign y6787 = n18999 ;
  assign y6788 = ~n19001 ;
  assign y6789 = n19005 ;
  assign y6790 = ~1'b0 ;
  assign y6791 = n19009 ;
  assign y6792 = n19015 ;
  assign y6793 = ~n19016 ;
  assign y6794 = ~n19019 ;
  assign y6795 = n19021 ;
  assign y6796 = n19023 ;
  assign y6797 = n1206 ;
  assign y6798 = ~n19025 ;
  assign y6799 = ~n19026 ;
  assign y6800 = ~n19027 ;
  assign y6801 = n19033 ;
  assign y6802 = n19034 ;
  assign y6803 = ~n19050 ;
  assign y6804 = ~1'b0 ;
  assign y6805 = ~n19054 ;
  assign y6806 = ~n19055 ;
  assign y6807 = ~1'b0 ;
  assign y6808 = n19056 ;
  assign y6809 = n19058 ;
  assign y6810 = n19059 ;
  assign y6811 = n19061 ;
  assign y6812 = ~1'b0 ;
  assign y6813 = ~n19064 ;
  assign y6814 = n19065 ;
  assign y6815 = n19066 ;
  assign y6816 = n9010 ;
  assign y6817 = ~1'b0 ;
  assign y6818 = n19072 ;
  assign y6819 = n2766 ;
  assign y6820 = ~n19075 ;
  assign y6821 = n19079 ;
  assign y6822 = ~n19085 ;
  assign y6823 = n19089 ;
  assign y6824 = ~n19094 ;
  assign y6825 = n19095 ;
  assign y6826 = ~1'b0 ;
  assign y6827 = n19096 ;
  assign y6828 = n19097 ;
  assign y6829 = ~n6287 ;
  assign y6830 = ~n19098 ;
  assign y6831 = ~1'b0 ;
  assign y6832 = ~n19101 ;
  assign y6833 = ~n19105 ;
  assign y6834 = n19108 ;
  assign y6835 = ~n19109 ;
  assign y6836 = n19110 ;
  assign y6837 = n19117 ;
  assign y6838 = ~n19118 ;
  assign y6839 = n19129 ;
  assign y6840 = n19132 ;
  assign y6841 = ~n19135 ;
  assign y6842 = ~n19136 ;
  assign y6843 = ~n19137 ;
  assign y6844 = ~n19140 ;
  assign y6845 = ~1'b0 ;
  assign y6846 = n797 ;
  assign y6847 = n19141 ;
  assign y6848 = n19144 ;
  assign y6849 = ~n19148 ;
  assign y6850 = ~n19150 ;
  assign y6851 = ~n19151 ;
  assign y6852 = n19152 ;
  assign y6853 = n19155 ;
  assign y6854 = n19158 ;
  assign y6855 = ~n19161 ;
  assign y6856 = ~1'b0 ;
  assign y6857 = ~n19164 ;
  assign y6858 = ~n19165 ;
  assign y6859 = ~n19166 ;
  assign y6860 = ~n19169 ;
  assign y6861 = ~n19181 ;
  assign y6862 = ~n19184 ;
  assign y6863 = ~1'b0 ;
  assign y6864 = n19192 ;
  assign y6865 = n19194 ;
  assign y6866 = ~n19195 ;
  assign y6867 = ~n19200 ;
  assign y6868 = ~1'b0 ;
  assign y6869 = ~n19202 ;
  assign y6870 = n19203 ;
  assign y6871 = ~n19204 ;
  assign y6872 = ~1'b0 ;
  assign y6873 = ~n19209 ;
  assign y6874 = ~1'b0 ;
  assign y6875 = n19210 ;
  assign y6876 = ~n19213 ;
  assign y6877 = ~n19216 ;
  assign y6878 = n19217 ;
  assign y6879 = ~1'b0 ;
  assign y6880 = n19225 ;
  assign y6881 = n19230 ;
  assign y6882 = ~n19231 ;
  assign y6883 = ~n19232 ;
  assign y6884 = n19235 ;
  assign y6885 = ~n19244 ;
  assign y6886 = n19246 ;
  assign y6887 = ~n19254 ;
  assign y6888 = n2326 ;
  assign y6889 = ~1'b0 ;
  assign y6890 = ~1'b0 ;
  assign y6891 = ~n19261 ;
  assign y6892 = ~n19262 ;
  assign y6893 = ~n19264 ;
  assign y6894 = ~n19266 ;
  assign y6895 = ~n19268 ;
  assign y6896 = n19273 ;
  assign y6897 = ~1'b0 ;
  assign y6898 = ~1'b0 ;
  assign y6899 = n19280 ;
  assign y6900 = ~1'b0 ;
  assign y6901 = n19285 ;
  assign y6902 = ~n19286 ;
  assign y6903 = ~1'b0 ;
  assign y6904 = ~n19289 ;
  assign y6905 = ~n19299 ;
  assign y6906 = ~1'b0 ;
  assign y6907 = ~n19301 ;
  assign y6908 = ~1'b0 ;
  assign y6909 = n19302 ;
  assign y6910 = ~1'b0 ;
  assign y6911 = ~1'b0 ;
  assign y6912 = ~n19304 ;
  assign y6913 = ~n19305 ;
  assign y6914 = ~n19306 ;
  assign y6915 = ~1'b0 ;
  assign y6916 = ~1'b0 ;
  assign y6917 = n19307 ;
  assign y6918 = ~1'b0 ;
  assign y6919 = n19317 ;
  assign y6920 = ~n19327 ;
  assign y6921 = ~n19328 ;
  assign y6922 = ~1'b0 ;
  assign y6923 = n19331 ;
  assign y6924 = x85 ;
  assign y6925 = ~n19334 ;
  assign y6926 = ~n19336 ;
  assign y6927 = ~n19339 ;
  assign y6928 = n19340 ;
  assign y6929 = ~n19343 ;
  assign y6930 = n19348 ;
  assign y6931 = ~n19350 ;
  assign y6932 = ~1'b0 ;
  assign y6933 = ~1'b0 ;
  assign y6934 = ~n19354 ;
  assign y6935 = n19355 ;
  assign y6936 = ~1'b0 ;
  assign y6937 = n19361 ;
  assign y6938 = ~n19364 ;
  assign y6939 = n19368 ;
  assign y6940 = n19370 ;
  assign y6941 = ~n19373 ;
  assign y6942 = ~1'b0 ;
  assign y6943 = ~1'b0 ;
  assign y6944 = n19377 ;
  assign y6945 = ~n19378 ;
  assign y6946 = ~1'b0 ;
  assign y6947 = ~1'b0 ;
  assign y6948 = ~n15180 ;
  assign y6949 = ~1'b0 ;
  assign y6950 = ~n19379 ;
  assign y6951 = ~n19381 ;
  assign y6952 = ~1'b0 ;
  assign y6953 = ~1'b0 ;
  assign y6954 = ~1'b0 ;
  assign y6955 = ~1'b0 ;
  assign y6956 = n19391 ;
  assign y6957 = ~1'b0 ;
  assign y6958 = ~n19396 ;
  assign y6959 = n19401 ;
  assign y6960 = ~n19405 ;
  assign y6961 = n19407 ;
  assign y6962 = n19413 ;
  assign y6963 = ~n19414 ;
  assign y6964 = ~1'b0 ;
  assign y6965 = ~n19416 ;
  assign y6966 = n19420 ;
  assign y6967 = n19422 ;
  assign y6968 = ~n19425 ;
  assign y6969 = ~n19426 ;
  assign y6970 = ~n19436 ;
  assign y6971 = n19438 ;
  assign y6972 = ~1'b0 ;
  assign y6973 = ~n19441 ;
  assign y6974 = n19447 ;
  assign y6975 = n19454 ;
  assign y6976 = ~1'b0 ;
  assign y6977 = n19458 ;
  assign y6978 = ~n19459 ;
  assign y6979 = n19463 ;
  assign y6980 = n19466 ;
  assign y6981 = n19470 ;
  assign y6982 = ~n19471 ;
  assign y6983 = ~n19472 ;
  assign y6984 = ~1'b0 ;
  assign y6985 = ~1'b0 ;
  assign y6986 = n19475 ;
  assign y6987 = n19478 ;
  assign y6988 = n19480 ;
  assign y6989 = n19483 ;
  assign y6990 = n19488 ;
  assign y6991 = n19493 ;
  assign y6992 = ~n19496 ;
  assign y6993 = n19497 ;
  assign y6994 = ~1'b0 ;
  assign y6995 = n19499 ;
  assign y6996 = ~n19502 ;
  assign y6997 = n17694 ;
  assign y6998 = n19503 ;
  assign y6999 = ~n19507 ;
  assign y7000 = ~1'b0 ;
  assign y7001 = n19515 ;
  assign y7002 = n19516 ;
  assign y7003 = ~n19518 ;
  assign y7004 = ~1'b0 ;
  assign y7005 = ~1'b0 ;
  assign y7006 = n19523 ;
  assign y7007 = ~n19527 ;
  assign y7008 = ~n19528 ;
  assign y7009 = ~n19533 ;
  assign y7010 = ~n19535 ;
  assign y7011 = n19537 ;
  assign y7012 = n571 ;
  assign y7013 = n19539 ;
  assign y7014 = n19540 ;
  assign y7015 = x230 ;
  assign y7016 = n19542 ;
  assign y7017 = ~1'b0 ;
  assign y7018 = ~n19544 ;
  assign y7019 = ~n19549 ;
  assign y7020 = n19552 ;
  assign y7021 = ~1'b0 ;
  assign y7022 = ~n19560 ;
  assign y7023 = n19562 ;
  assign y7024 = n19563 ;
  assign y7025 = n19566 ;
  assign y7026 = n19569 ;
  assign y7027 = n19573 ;
  assign y7028 = ~1'b0 ;
  assign y7029 = ~n19584 ;
  assign y7030 = ~n19595 ;
  assign y7031 = n2760 ;
  assign y7032 = ~1'b0 ;
  assign y7033 = ~n19601 ;
  assign y7034 = ~n19607 ;
  assign y7035 = ~n19609 ;
  assign y7036 = ~n19617 ;
  assign y7037 = ~n19622 ;
  assign y7038 = ~1'b0 ;
  assign y7039 = ~n19630 ;
  assign y7040 = n19631 ;
  assign y7041 = ~n15044 ;
  assign y7042 = n19632 ;
  assign y7043 = ~n19633 ;
  assign y7044 = n19636 ;
  assign y7045 = 1'b0 ;
  assign y7046 = n19643 ;
  assign y7047 = n19651 ;
  assign y7048 = n19654 ;
  assign y7049 = ~1'b0 ;
  assign y7050 = ~1'b0 ;
  assign y7051 = ~n19661 ;
  assign y7052 = ~n19662 ;
  assign y7053 = ~n19665 ;
  assign y7054 = n19670 ;
  assign y7055 = ~1'b0 ;
  assign y7056 = ~1'b0 ;
  assign y7057 = ~n19671 ;
  assign y7058 = ~1'b0 ;
  assign y7059 = n19673 ;
  assign y7060 = ~n10031 ;
  assign y7061 = n19683 ;
  assign y7062 = ~n19685 ;
  assign y7063 = n19686 ;
  assign y7064 = n19689 ;
  assign y7065 = ~1'b0 ;
  assign y7066 = n11920 ;
  assign y7067 = ~n19690 ;
  assign y7068 = ~1'b0 ;
  assign y7069 = ~1'b0 ;
  assign y7070 = n19691 ;
  assign y7071 = ~n19695 ;
  assign y7072 = ~n19697 ;
  assign y7073 = ~n19698 ;
  assign y7074 = ~1'b0 ;
  assign y7075 = ~n19699 ;
  assign y7076 = ~n19715 ;
  assign y7077 = ~n19717 ;
  assign y7078 = n19718 ;
  assign y7079 = ~n19726 ;
  assign y7080 = ~n19727 ;
  assign y7081 = n19730 ;
  assign y7082 = ~n19734 ;
  assign y7083 = ~n19735 ;
  assign y7084 = ~1'b0 ;
  assign y7085 = ~1'b0 ;
  assign y7086 = ~n19738 ;
  assign y7087 = n19739 ;
  assign y7088 = n19743 ;
  assign y7089 = ~n19748 ;
  assign y7090 = ~n19750 ;
  assign y7091 = n19753 ;
  assign y7092 = ~n19755 ;
  assign y7093 = ~n19758 ;
  assign y7094 = ~1'b0 ;
  assign y7095 = ~1'b0 ;
  assign y7096 = n19759 ;
  assign y7097 = ~n19762 ;
  assign y7098 = ~n19763 ;
  assign y7099 = n19764 ;
  assign y7100 = n19767 ;
  assign y7101 = n19769 ;
  assign y7102 = ~1'b0 ;
  assign y7103 = ~1'b0 ;
  assign y7104 = ~n19770 ;
  assign y7105 = n19773 ;
  assign y7106 = ~n19777 ;
  assign y7107 = n19779 ;
  assign y7108 = n19782 ;
  assign y7109 = ~n19784 ;
  assign y7110 = ~n19785 ;
  assign y7111 = ~1'b0 ;
  assign y7112 = n19787 ;
  assign y7113 = ~1'b0 ;
  assign y7114 = n19791 ;
  assign y7115 = ~n19792 ;
  assign y7116 = ~1'b0 ;
  assign y7117 = ~1'b0 ;
  assign y7118 = ~1'b0 ;
  assign y7119 = n19793 ;
  assign y7120 = n19796 ;
  assign y7121 = n19798 ;
  assign y7122 = ~1'b0 ;
  assign y7123 = ~1'b0 ;
  assign y7124 = ~n19801 ;
  assign y7125 = ~n19805 ;
  assign y7126 = n19809 ;
  assign y7127 = ~n19811 ;
  assign y7128 = 1'b0 ;
  assign y7129 = n19816 ;
  assign y7130 = n7707 ;
  assign y7131 = n19818 ;
  assign y7132 = n19824 ;
  assign y7133 = ~n19827 ;
  assign y7134 = ~1'b0 ;
  assign y7135 = ~1'b0 ;
  assign y7136 = n19828 ;
  assign y7137 = ~n19830 ;
  assign y7138 = n19831 ;
  assign y7139 = n19835 ;
  assign y7140 = ~1'b0 ;
  assign y7141 = ~n19836 ;
  assign y7142 = ~n19837 ;
  assign y7143 = n19842 ;
  assign y7144 = ~n19844 ;
  assign y7145 = ~1'b0 ;
  assign y7146 = ~n19846 ;
  assign y7147 = ~1'b0 ;
  assign y7148 = n12305 ;
  assign y7149 = ~n19847 ;
  assign y7150 = ~n19848 ;
  assign y7151 = ~1'b0 ;
  assign y7152 = ~1'b0 ;
  assign y7153 = ~n19857 ;
  assign y7154 = ~1'b0 ;
  assign y7155 = ~n19859 ;
  assign y7156 = ~n19865 ;
  assign y7157 = ~n19868 ;
  assign y7158 = ~n19871 ;
  assign y7159 = n19872 ;
  assign y7160 = ~n19874 ;
  assign y7161 = n19878 ;
  assign y7162 = ~n19879 ;
  assign y7163 = ~1'b0 ;
  assign y7164 = ~n19880 ;
  assign y7165 = n19882 ;
  assign y7166 = ~1'b0 ;
  assign y7167 = ~n19884 ;
  assign y7168 = n19885 ;
  assign y7169 = ~n19888 ;
  assign y7170 = n19892 ;
  assign y7171 = n18668 ;
  assign y7172 = n19893 ;
  assign y7173 = ~n19895 ;
  assign y7174 = n19896 ;
  assign y7175 = n19898 ;
  assign y7176 = n19901 ;
  assign y7177 = ~1'b0 ;
  assign y7178 = n19906 ;
  assign y7179 = n19910 ;
  assign y7180 = n19912 ;
  assign y7181 = ~n19914 ;
  assign y7182 = n19869 ;
  assign y7183 = n19920 ;
  assign y7184 = ~n19921 ;
  assign y7185 = n19924 ;
  assign y7186 = ~1'b0 ;
  assign y7187 = n19928 ;
  assign y7188 = n19931 ;
  assign y7189 = n15094 ;
  assign y7190 = n19934 ;
  assign y7191 = ~1'b0 ;
  assign y7192 = ~n19945 ;
  assign y7193 = n19946 ;
  assign y7194 = n3062 ;
  assign y7195 = ~n19947 ;
  assign y7196 = ~n19950 ;
  assign y7197 = ~n19952 ;
  assign y7198 = n19955 ;
  assign y7199 = ~n19958 ;
  assign y7200 = n19961 ;
  assign y7201 = n19962 ;
  assign y7202 = ~1'b0 ;
  assign y7203 = ~n19964 ;
  assign y7204 = n11327 ;
  assign y7205 = ~1'b0 ;
  assign y7206 = n19965 ;
  assign y7207 = ~n19971 ;
  assign y7208 = n19972 ;
  assign y7209 = ~1'b0 ;
  assign y7210 = n19973 ;
  assign y7211 = ~n19974 ;
  assign y7212 = ~n19976 ;
  assign y7213 = ~n19977 ;
  assign y7214 = n19988 ;
  assign y7215 = ~n19989 ;
  assign y7216 = ~1'b0 ;
  assign y7217 = ~1'b0 ;
  assign y7218 = ~n19990 ;
  assign y7219 = n19992 ;
  assign y7220 = ~n19995 ;
  assign y7221 = ~1'b0 ;
  assign y7222 = n19997 ;
  assign y7223 = ~1'b0 ;
  assign y7224 = ~n19998 ;
  assign y7225 = ~1'b0 ;
  assign y7226 = n20000 ;
  assign y7227 = ~n7873 ;
  assign y7228 = ~n20003 ;
  assign y7229 = n20005 ;
  assign y7230 = ~n20011 ;
  assign y7231 = ~1'b0 ;
  assign y7232 = n20012 ;
  assign y7233 = ~n20015 ;
  assign y7234 = ~1'b0 ;
  assign y7235 = ~n20028 ;
  assign y7236 = n20029 ;
  assign y7237 = n20036 ;
  assign y7238 = ~n20038 ;
  assign y7239 = ~1'b0 ;
  assign y7240 = n20039 ;
  assign y7241 = ~1'b0 ;
  assign y7242 = ~n20042 ;
  assign y7243 = ~1'b0 ;
  assign y7244 = n20043 ;
  assign y7245 = ~n20052 ;
  assign y7246 = ~n20054 ;
  assign y7247 = 1'b0 ;
  assign y7248 = ~1'b0 ;
  assign y7249 = n20056 ;
  assign y7250 = ~n20057 ;
  assign y7251 = n20060 ;
  assign y7252 = ~n20063 ;
  assign y7253 = n20068 ;
  assign y7254 = ~n20069 ;
  assign y7255 = n20070 ;
  assign y7256 = ~n20078 ;
  assign y7257 = ~n20080 ;
  assign y7258 = n20081 ;
  assign y7259 = n20084 ;
  assign y7260 = ~1'b0 ;
  assign y7261 = n20085 ;
  assign y7262 = n20090 ;
  assign y7263 = ~n20093 ;
  assign y7264 = n20094 ;
  assign y7265 = n19065 ;
  assign y7266 = n20096 ;
  assign y7267 = n20101 ;
  assign y7268 = n20103 ;
  assign y7269 = n20105 ;
  assign y7270 = ~n20110 ;
  assign y7271 = ~n20112 ;
  assign y7272 = ~1'b0 ;
  assign y7273 = n20114 ;
  assign y7274 = n20116 ;
  assign y7275 = ~n20121 ;
  assign y7276 = ~x250 ;
  assign y7277 = n20124 ;
  assign y7278 = ~1'b0 ;
  assign y7279 = ~1'b0 ;
  assign y7280 = ~n20127 ;
  assign y7281 = n20130 ;
  assign y7282 = n20132 ;
  assign y7283 = ~n20136 ;
  assign y7284 = ~1'b0 ;
  assign y7285 = ~n10271 ;
  assign y7286 = n20138 ;
  assign y7287 = ~n20140 ;
  assign y7288 = ~n20151 ;
  assign y7289 = n20152 ;
  assign y7290 = ~n20153 ;
  assign y7291 = ~n20156 ;
  assign y7292 = n20160 ;
  assign y7293 = ~n20163 ;
  assign y7294 = ~1'b0 ;
  assign y7295 = n20171 ;
  assign y7296 = ~n20176 ;
  assign y7297 = n20178 ;
  assign y7298 = ~n20189 ;
  assign y7299 = ~n20190 ;
  assign y7300 = n20194 ;
  assign y7301 = ~n20197 ;
  assign y7302 = n20206 ;
  assign y7303 = ~1'b0 ;
  assign y7304 = n20207 ;
  assign y7305 = n20208 ;
  assign y7306 = n20210 ;
  assign y7307 = ~n20211 ;
  assign y7308 = ~1'b0 ;
  assign y7309 = ~n20222 ;
  assign y7310 = n20223 ;
  assign y7311 = ~n20227 ;
  assign y7312 = n3049 ;
  assign y7313 = ~n20230 ;
  assign y7314 = ~1'b0 ;
  assign y7315 = ~1'b0 ;
  assign y7316 = ~1'b0 ;
  assign y7317 = ~n20236 ;
  assign y7318 = ~1'b0 ;
  assign y7319 = ~1'b0 ;
  assign y7320 = ~1'b0 ;
  assign y7321 = ~n20242 ;
  assign y7322 = ~1'b0 ;
  assign y7323 = n20245 ;
  assign y7324 = n20246 ;
  assign y7325 = n20259 ;
  assign y7326 = n20261 ;
  assign y7327 = ~n20267 ;
  assign y7328 = ~n19026 ;
  assign y7329 = ~n20269 ;
  assign y7330 = ~n20280 ;
  assign y7331 = ~1'b0 ;
  assign y7332 = n20282 ;
  assign y7333 = n20285 ;
  assign y7334 = ~1'b0 ;
  assign y7335 = ~n20287 ;
  assign y7336 = ~1'b0 ;
  assign y7337 = ~1'b0 ;
  assign y7338 = n20288 ;
  assign y7339 = n20296 ;
  assign y7340 = n20299 ;
  assign y7341 = n2336 ;
  assign y7342 = ~n20303 ;
  assign y7343 = ~1'b0 ;
  assign y7344 = 1'b0 ;
  assign y7345 = ~n20307 ;
  assign y7346 = n6390 ;
  assign y7347 = ~1'b0 ;
  assign y7348 = ~n20308 ;
  assign y7349 = n20309 ;
  assign y7350 = n20312 ;
  assign y7351 = ~n20314 ;
  assign y7352 = ~n20318 ;
  assign y7353 = n20321 ;
  assign y7354 = ~n20324 ;
  assign y7355 = ~n20335 ;
  assign y7356 = ~n20337 ;
  assign y7357 = n20339 ;
  assign y7358 = n20340 ;
  assign y7359 = ~n20345 ;
  assign y7360 = ~1'b0 ;
  assign y7361 = ~n20348 ;
  assign y7362 = ~n20349 ;
  assign y7363 = n20363 ;
  assign y7364 = ~1'b0 ;
  assign y7365 = n1327 ;
  assign y7366 = n3843 ;
  assign y7367 = ~n20366 ;
  assign y7368 = n20367 ;
  assign y7369 = ~n20368 ;
  assign y7370 = ~n20371 ;
  assign y7371 = ~n20373 ;
  assign y7372 = ~n20375 ;
  assign y7373 = ~1'b0 ;
  assign y7374 = n20376 ;
  assign y7375 = n20380 ;
  assign y7376 = ~n10223 ;
  assign y7377 = ~n20381 ;
  assign y7378 = n20385 ;
  assign y7379 = ~n20387 ;
  assign y7380 = ~1'b0 ;
  assign y7381 = n20391 ;
  assign y7382 = ~n20393 ;
  assign y7383 = ~n20395 ;
  assign y7384 = n20397 ;
  assign y7385 = ~n20401 ;
  assign y7386 = n20406 ;
  assign y7387 = ~n20418 ;
  assign y7388 = ~n20420 ;
  assign y7389 = n17338 ;
  assign y7390 = ~n20422 ;
  assign y7391 = n20425 ;
  assign y7392 = ~n20429 ;
  assign y7393 = ~n20431 ;
  assign y7394 = ~n20437 ;
  assign y7395 = ~n20439 ;
  assign y7396 = ~n20440 ;
  assign y7397 = n20442 ;
  assign y7398 = ~1'b0 ;
  assign y7399 = ~1'b0 ;
  assign y7400 = n20445 ;
  assign y7401 = ~1'b0 ;
  assign y7402 = n20452 ;
  assign y7403 = n20458 ;
  assign y7404 = ~n20460 ;
  assign y7405 = ~n20467 ;
  assign y7406 = n20469 ;
  assign y7407 = n20474 ;
  assign y7408 = n20475 ;
  assign y7409 = ~n20476 ;
  assign y7410 = ~n20481 ;
  assign y7411 = ~1'b0 ;
  assign y7412 = ~1'b0 ;
  assign y7413 = ~n20483 ;
  assign y7414 = ~1'b0 ;
  assign y7415 = n20484 ;
  assign y7416 = ~n20487 ;
  assign y7417 = ~1'b0 ;
  assign y7418 = ~1'b0 ;
  assign y7419 = n20489 ;
  assign y7420 = n20491 ;
  assign y7421 = ~n20492 ;
  assign y7422 = ~n20498 ;
  assign y7423 = n20500 ;
  assign y7424 = ~1'b0 ;
  assign y7425 = n20506 ;
  assign y7426 = n20509 ;
  assign y7427 = ~n20520 ;
  assign y7428 = ~n20523 ;
  assign y7429 = ~n20528 ;
  assign y7430 = n20530 ;
  assign y7431 = n20532 ;
  assign y7432 = ~n20533 ;
  assign y7433 = ~n20539 ;
  assign y7434 = 1'b0 ;
  assign y7435 = n20541 ;
  assign y7436 = n20543 ;
  assign y7437 = ~1'b0 ;
  assign y7438 = ~n20545 ;
  assign y7439 = ~n20547 ;
  assign y7440 = n20550 ;
  assign y7441 = ~1'b0 ;
  assign y7442 = n20552 ;
  assign y7443 = ~1'b0 ;
  assign y7444 = ~n20565 ;
  assign y7445 = ~1'b0 ;
  assign y7446 = ~n20570 ;
  assign y7447 = n20571 ;
  assign y7448 = ~n20575 ;
  assign y7449 = n20576 ;
  assign y7450 = ~n20577 ;
  assign y7451 = ~n20578 ;
  assign y7452 = ~n20582 ;
  assign y7453 = n20587 ;
  assign y7454 = n20590 ;
  assign y7455 = n20593 ;
  assign y7456 = ~n20594 ;
  assign y7457 = ~n20595 ;
  assign y7458 = ~1'b0 ;
  assign y7459 = 1'b0 ;
  assign y7460 = n20598 ;
  assign y7461 = n20602 ;
  assign y7462 = ~n20607 ;
  assign y7463 = n20611 ;
  assign y7464 = n20615 ;
  assign y7465 = n20620 ;
  assign y7466 = n20621 ;
  assign y7467 = ~n20623 ;
  assign y7468 = ~n2804 ;
  assign y7469 = ~n20627 ;
  assign y7470 = ~n20632 ;
  assign y7471 = ~n20642 ;
  assign y7472 = ~n20643 ;
  assign y7473 = ~1'b0 ;
  assign y7474 = ~n20647 ;
  assign y7475 = n20649 ;
  assign y7476 = n20652 ;
  assign y7477 = n20656 ;
  assign y7478 = n20658 ;
  assign y7479 = n20666 ;
  assign y7480 = n20676 ;
  assign y7481 = n20681 ;
  assign y7482 = ~n20684 ;
  assign y7483 = ~1'b0 ;
  assign y7484 = n20687 ;
  assign y7485 = n20695 ;
  assign y7486 = n20707 ;
  assign y7487 = ~n20709 ;
  assign y7488 = n20711 ;
  assign y7489 = ~1'b0 ;
  assign y7490 = ~1'b0 ;
  assign y7491 = n20715 ;
  assign y7492 = n20718 ;
  assign y7493 = ~1'b0 ;
  assign y7494 = ~n6562 ;
  assign y7495 = ~1'b0 ;
  assign y7496 = ~n20721 ;
  assign y7497 = ~n20729 ;
  assign y7498 = ~n20733 ;
  assign y7499 = ~n20736 ;
  assign y7500 = ~1'b0 ;
  assign y7501 = ~n20740 ;
  assign y7502 = ~n20744 ;
  assign y7503 = n20746 ;
  assign y7504 = ~1'b0 ;
  assign y7505 = n20750 ;
  assign y7506 = ~1'b0 ;
  assign y7507 = n7325 ;
  assign y7508 = ~1'b0 ;
  assign y7509 = ~1'b0 ;
  assign y7510 = n20754 ;
  assign y7511 = ~1'b0 ;
  assign y7512 = ~n20757 ;
  assign y7513 = ~1'b0 ;
  assign y7514 = n20758 ;
  assign y7515 = ~n20760 ;
  assign y7516 = n20764 ;
  assign y7517 = n20767 ;
  assign y7518 = ~1'b0 ;
  assign y7519 = ~1'b0 ;
  assign y7520 = n20771 ;
  assign y7521 = n20776 ;
  assign y7522 = n20777 ;
  assign y7523 = ~n20783 ;
  assign y7524 = n20784 ;
  assign y7525 = ~n20792 ;
  assign y7526 = ~1'b0 ;
  assign y7527 = ~1'b0 ;
  assign y7528 = ~n20799 ;
  assign y7529 = ~n20800 ;
  assign y7530 = n20802 ;
  assign y7531 = 1'b0 ;
  assign y7532 = ~n20804 ;
  assign y7533 = n20810 ;
  assign y7534 = n19157 ;
  assign y7535 = ~n20811 ;
  assign y7536 = n20815 ;
  assign y7537 = ~n20816 ;
  assign y7538 = ~n20818 ;
  assign y7539 = n20823 ;
  assign y7540 = n20827 ;
  assign y7541 = n20832 ;
  assign y7542 = ~n20836 ;
  assign y7543 = n20845 ;
  assign y7544 = ~1'b0 ;
  assign y7545 = ~1'b0 ;
  assign y7546 = n20847 ;
  assign y7547 = n20856 ;
  assign y7548 = ~n20859 ;
  assign y7549 = ~1'b0 ;
  assign y7550 = n20862 ;
  assign y7551 = n20863 ;
  assign y7552 = ~1'b0 ;
  assign y7553 = ~1'b0 ;
  assign y7554 = n20881 ;
  assign y7555 = n20883 ;
  assign y7556 = ~n20884 ;
  assign y7557 = n20886 ;
  assign y7558 = n20891 ;
  assign y7559 = ~n20893 ;
  assign y7560 = n20894 ;
  assign y7561 = ~n20897 ;
  assign y7562 = n20904 ;
  assign y7563 = n20906 ;
  assign y7564 = ~n20907 ;
  assign y7565 = ~n20913 ;
  assign y7566 = ~1'b0 ;
  assign y7567 = ~1'b0 ;
  assign y7568 = ~1'b0 ;
  assign y7569 = n20915 ;
  assign y7570 = ~n20919 ;
  assign y7571 = ~n20922 ;
  assign y7572 = n20923 ;
  assign y7573 = ~n20925 ;
  assign y7574 = n20927 ;
  assign y7575 = n20929 ;
  assign y7576 = n20930 ;
  assign y7577 = ~n20932 ;
  assign y7578 = n20934 ;
  assign y7579 = n20935 ;
  assign y7580 = ~1'b0 ;
  assign y7581 = ~n20940 ;
  assign y7582 = n20942 ;
  assign y7583 = n20943 ;
  assign y7584 = ~n20946 ;
  assign y7585 = ~1'b0 ;
  assign y7586 = n20949 ;
  assign y7587 = n20953 ;
  assign y7588 = ~n13561 ;
  assign y7589 = ~1'b0 ;
  assign y7590 = ~1'b0 ;
  assign y7591 = ~n20960 ;
  assign y7592 = n20963 ;
  assign y7593 = ~1'b0 ;
  assign y7594 = ~1'b0 ;
  assign y7595 = ~1'b0 ;
  assign y7596 = ~1'b0 ;
  assign y7597 = ~n20968 ;
  assign y7598 = n20974 ;
  assign y7599 = ~1'b0 ;
  assign y7600 = n20975 ;
  assign y7601 = n20977 ;
  assign y7602 = n20981 ;
  assign y7603 = n20983 ;
  assign y7604 = ~n20985 ;
  assign y7605 = ~1'b0 ;
  assign y7606 = ~1'b0 ;
  assign y7607 = ~n20988 ;
  assign y7608 = ~n20990 ;
  assign y7609 = ~n20991 ;
  assign y7610 = 1'b0 ;
  assign y7611 = ~n20993 ;
  assign y7612 = ~n21006 ;
  assign y7613 = ~n21008 ;
  assign y7614 = ~n21012 ;
  assign y7615 = ~1'b0 ;
  assign y7616 = ~n21015 ;
  assign y7617 = ~n21017 ;
  assign y7618 = n21018 ;
  assign y7619 = n21019 ;
  assign y7620 = ~1'b0 ;
  assign y7621 = ~n21025 ;
  assign y7622 = n21030 ;
  assign y7623 = ~n21031 ;
  assign y7624 = n21037 ;
  assign y7625 = n21038 ;
  assign y7626 = ~n21040 ;
  assign y7627 = ~n21043 ;
  assign y7628 = ~n12041 ;
  assign y7629 = ~1'b0 ;
  assign y7630 = ~1'b0 ;
  assign y7631 = n21046 ;
  assign y7632 = ~n21049 ;
  assign y7633 = n21051 ;
  assign y7634 = ~n21053 ;
  assign y7635 = n21057 ;
  assign y7636 = ~1'b0 ;
  assign y7637 = n21064 ;
  assign y7638 = n21068 ;
  assign y7639 = ~n21073 ;
  assign y7640 = n21076 ;
  assign y7641 = ~n21077 ;
  assign y7642 = ~1'b0 ;
  assign y7643 = ~1'b0 ;
  assign y7644 = n8001 ;
  assign y7645 = ~n21080 ;
  assign y7646 = n21082 ;
  assign y7647 = ~1'b0 ;
  assign y7648 = ~n21089 ;
  assign y7649 = n21094 ;
  assign y7650 = ~n21095 ;
  assign y7651 = n21096 ;
  assign y7652 = ~n21098 ;
  assign y7653 = ~n21099 ;
  assign y7654 = ~1'b0 ;
  assign y7655 = ~1'b0 ;
  assign y7656 = n21102 ;
  assign y7657 = ~1'b0 ;
  assign y7658 = ~n21107 ;
  assign y7659 = n21109 ;
  assign y7660 = n21112 ;
  assign y7661 = ~1'b0 ;
  assign y7662 = n21113 ;
  assign y7663 = n21116 ;
  assign y7664 = ~n2068 ;
  assign y7665 = ~1'b0 ;
  assign y7666 = n21124 ;
  assign y7667 = n21128 ;
  assign y7668 = ~1'b0 ;
  assign y7669 = ~1'b0 ;
  assign y7670 = n21130 ;
  assign y7671 = ~n21131 ;
  assign y7672 = ~n21132 ;
  assign y7673 = ~1'b0 ;
  assign y7674 = ~1'b0 ;
  assign y7675 = n21133 ;
  assign y7676 = ~1'b0 ;
  assign y7677 = ~n21142 ;
  assign y7678 = n21144 ;
  assign y7679 = ~n21147 ;
  assign y7680 = ~n21155 ;
  assign y7681 = ~n21159 ;
  assign y7682 = ~1'b0 ;
  assign y7683 = n21161 ;
  assign y7684 = ~n21162 ;
  assign y7685 = n21168 ;
  assign y7686 = n21169 ;
  assign y7687 = n21171 ;
  assign y7688 = ~n21173 ;
  assign y7689 = ~n21174 ;
  assign y7690 = ~n21178 ;
  assign y7691 = n21182 ;
  assign y7692 = n21185 ;
  assign y7693 = n21192 ;
  assign y7694 = ~n21195 ;
  assign y7695 = ~n21207 ;
  assign y7696 = ~n21209 ;
  assign y7697 = ~1'b0 ;
  assign y7698 = n8012 ;
  assign y7699 = ~n21211 ;
  assign y7700 = ~n21212 ;
  assign y7701 = n8043 ;
  assign y7702 = ~n21215 ;
  assign y7703 = ~n21219 ;
  assign y7704 = ~1'b0 ;
  assign y7705 = n21222 ;
  assign y7706 = ~n21224 ;
  assign y7707 = n21227 ;
  assign y7708 = n21233 ;
  assign y7709 = n21243 ;
  assign y7710 = n21244 ;
  assign y7711 = n21245 ;
  assign y7712 = n21247 ;
  assign y7713 = n21249 ;
  assign y7714 = n21250 ;
  assign y7715 = ~n21253 ;
  assign y7716 = ~1'b0 ;
  assign y7717 = n21258 ;
  assign y7718 = ~1'b0 ;
  assign y7719 = ~n21268 ;
  assign y7720 = ~1'b0 ;
  assign y7721 = n21275 ;
  assign y7722 = ~n21281 ;
  assign y7723 = ~n1399 ;
  assign y7724 = n21283 ;
  assign y7725 = x177 ;
  assign y7726 = ~n21285 ;
  assign y7727 = ~n13324 ;
  assign y7728 = ~1'b0 ;
  assign y7729 = ~1'b0 ;
  assign y7730 = ~n15126 ;
  assign y7731 = ~1'b0 ;
  assign y7732 = ~n21287 ;
  assign y7733 = n21288 ;
  assign y7734 = ~1'b0 ;
  assign y7735 = ~n21291 ;
  assign y7736 = ~n21294 ;
  assign y7737 = n21296 ;
  assign y7738 = n21297 ;
  assign y7739 = ~n21301 ;
  assign y7740 = ~n21303 ;
  assign y7741 = n21308 ;
  assign y7742 = n21309 ;
  assign y7743 = ~1'b0 ;
  assign y7744 = n21310 ;
  assign y7745 = n21312 ;
  assign y7746 = ~n21323 ;
  assign y7747 = n21324 ;
  assign y7748 = n21327 ;
  assign y7749 = ~n21332 ;
  assign y7750 = n21334 ;
  assign y7751 = n21339 ;
  assign y7752 = n21340 ;
  assign y7753 = ~n21348 ;
  assign y7754 = ~1'b0 ;
  assign y7755 = ~n21352 ;
  assign y7756 = ~1'b0 ;
  assign y7757 = n21356 ;
  assign y7758 = n21358 ;
  assign y7759 = ~1'b0 ;
  assign y7760 = ~1'b0 ;
  assign y7761 = n21359 ;
  assign y7762 = ~n21364 ;
  assign y7763 = ~1'b0 ;
  assign y7764 = ~1'b0 ;
  assign y7765 = ~1'b0 ;
  assign y7766 = ~n21370 ;
  assign y7767 = ~n21373 ;
  assign y7768 = ~n3040 ;
  assign y7769 = ~n21377 ;
  assign y7770 = n21379 ;
  assign y7771 = ~n21388 ;
  assign y7772 = ~n21390 ;
  assign y7773 = n21392 ;
  assign y7774 = ~n21394 ;
  assign y7775 = n21402 ;
  assign y7776 = ~n21405 ;
  assign y7777 = n21406 ;
  assign y7778 = ~n21408 ;
  assign y7779 = ~n21410 ;
  assign y7780 = ~1'b0 ;
  assign y7781 = n21412 ;
  assign y7782 = ~n21413 ;
  assign y7783 = n21415 ;
  assign y7784 = n21417 ;
  assign y7785 = ~1'b0 ;
  assign y7786 = ~n21424 ;
  assign y7787 = ~n21425 ;
  assign y7788 = ~n21429 ;
  assign y7789 = n21434 ;
  assign y7790 = n21435 ;
  assign y7791 = ~n21442 ;
  assign y7792 = ~n21446 ;
  assign y7793 = ~n21448 ;
  assign y7794 = n21458 ;
  assign y7795 = ~n21461 ;
  assign y7796 = n21468 ;
  assign y7797 = n21470 ;
  assign y7798 = ~1'b0 ;
  assign y7799 = 1'b0 ;
  assign y7800 = ~n21472 ;
  assign y7801 = ~1'b0 ;
  assign y7802 = ~n21474 ;
  assign y7803 = ~n21476 ;
  assign y7804 = ~n21479 ;
  assign y7805 = ~n21482 ;
  assign y7806 = ~1'b0 ;
  assign y7807 = n21488 ;
  assign y7808 = ~1'b0 ;
  assign y7809 = ~1'b0 ;
  assign y7810 = n21490 ;
  assign y7811 = ~n21493 ;
  assign y7812 = ~n21498 ;
  assign y7813 = n21499 ;
  assign y7814 = n21501 ;
  assign y7815 = ~1'b0 ;
  assign y7816 = ~n21503 ;
  assign y7817 = ~n21517 ;
  assign y7818 = ~n21519 ;
  assign y7819 = n21520 ;
  assign y7820 = ~1'b0 ;
  assign y7821 = ~n21522 ;
  assign y7822 = ~1'b0 ;
  assign y7823 = n21523 ;
  assign y7824 = ~n21525 ;
  assign y7825 = n21526 ;
  assign y7826 = n21535 ;
  assign y7827 = n21537 ;
  assign y7828 = ~1'b0 ;
  assign y7829 = n21541 ;
  assign y7830 = n21542 ;
  assign y7831 = ~1'b0 ;
  assign y7832 = n21544 ;
  assign y7833 = n21547 ;
  assign y7834 = ~n21550 ;
  assign y7835 = n21552 ;
  assign y7836 = ~1'b0 ;
  assign y7837 = ~1'b0 ;
  assign y7838 = ~n21553 ;
  assign y7839 = ~n21558 ;
  assign y7840 = ~1'b0 ;
  assign y7841 = n21559 ;
  assign y7842 = ~1'b0 ;
  assign y7843 = n21568 ;
  assign y7844 = ~n21570 ;
  assign y7845 = ~1'b0 ;
  assign y7846 = ~n21575 ;
  assign y7847 = ~n21576 ;
  assign y7848 = n17078 ;
  assign y7849 = ~1'b0 ;
  assign y7850 = ~n21581 ;
  assign y7851 = ~n21584 ;
  assign y7852 = 1'b0 ;
  assign y7853 = ~n21586 ;
  assign y7854 = n21588 ;
  assign y7855 = ~1'b0 ;
  assign y7856 = ~n21589 ;
  assign y7857 = ~n21592 ;
  assign y7858 = n21597 ;
  assign y7859 = ~n21602 ;
  assign y7860 = ~n21607 ;
  assign y7861 = ~n21608 ;
  assign y7862 = n21609 ;
  assign y7863 = n21613 ;
  assign y7864 = n21616 ;
  assign y7865 = ~1'b0 ;
  assign y7866 = ~n21618 ;
  assign y7867 = ~n21620 ;
  assign y7868 = n21630 ;
  assign y7869 = ~n21632 ;
  assign y7870 = n21635 ;
  assign y7871 = ~n21641 ;
  assign y7872 = ~n21645 ;
  assign y7873 = n21649 ;
  assign y7874 = n21650 ;
  assign y7875 = ~n21654 ;
  assign y7876 = n21660 ;
  assign y7877 = n21662 ;
  assign y7878 = ~1'b0 ;
  assign y7879 = n21665 ;
  assign y7880 = ~n21667 ;
  assign y7881 = ~n21672 ;
  assign y7882 = ~n21673 ;
  assign y7883 = ~n21675 ;
  assign y7884 = ~n21676 ;
  assign y7885 = n21679 ;
  assign y7886 = n21680 ;
  assign y7887 = ~1'b0 ;
  assign y7888 = ~n21681 ;
  assign y7889 = n21686 ;
  assign y7890 = ~n21687 ;
  assign y7891 = n21689 ;
  assign y7892 = n21697 ;
  assign y7893 = n21704 ;
  assign y7894 = ~1'b0 ;
  assign y7895 = ~1'b0 ;
  assign y7896 = n21705 ;
  assign y7897 = n21711 ;
  assign y7898 = ~n21712 ;
  assign y7899 = n21713 ;
  assign y7900 = ~n21722 ;
  assign y7901 = n21726 ;
  assign y7902 = n21727 ;
  assign y7903 = ~n21731 ;
  assign y7904 = ~n21732 ;
  assign y7905 = ~n21733 ;
  assign y7906 = ~n21734 ;
  assign y7907 = n21736 ;
  assign y7908 = ~1'b0 ;
  assign y7909 = n21737 ;
  assign y7910 = ~n21739 ;
  assign y7911 = ~n21744 ;
  assign y7912 = n21745 ;
  assign y7913 = ~n21748 ;
  assign y7914 = ~n21751 ;
  assign y7915 = n21755 ;
  assign y7916 = n21758 ;
  assign y7917 = ~n21761 ;
  assign y7918 = n21766 ;
  assign y7919 = ~1'b0 ;
  assign y7920 = ~1'b0 ;
  assign y7921 = ~n21775 ;
  assign y7922 = n21778 ;
  assign y7923 = ~1'b0 ;
  assign y7924 = ~n21781 ;
  assign y7925 = n21785 ;
  assign y7926 = n21788 ;
  assign y7927 = ~1'b0 ;
  assign y7928 = ~n21791 ;
  assign y7929 = n21800 ;
  assign y7930 = ~n21802 ;
  assign y7931 = n21807 ;
  assign y7932 = ~n21818 ;
  assign y7933 = ~1'b0 ;
  assign y7934 = n21824 ;
  assign y7935 = n21825 ;
  assign y7936 = ~1'b0 ;
  assign y7937 = ~1'b0 ;
  assign y7938 = ~1'b0 ;
  assign y7939 = n21826 ;
  assign y7940 = ~n21831 ;
  assign y7941 = ~n21832 ;
  assign y7942 = n21839 ;
  assign y7943 = ~n21843 ;
  assign y7944 = ~n21846 ;
  assign y7945 = ~1'b0 ;
  assign y7946 = ~n21849 ;
  assign y7947 = n21853 ;
  assign y7948 = ~n21859 ;
  assign y7949 = ~n21860 ;
  assign y7950 = ~1'b0 ;
  assign y7951 = ~n21863 ;
  assign y7952 = n21864 ;
  assign y7953 = n21866 ;
  assign y7954 = n21867 ;
  assign y7955 = n21872 ;
  assign y7956 = ~1'b0 ;
  assign y7957 = n21877 ;
  assign y7958 = n21878 ;
  assign y7959 = ~1'b0 ;
  assign y7960 = ~n21879 ;
  assign y7961 = ~n21881 ;
  assign y7962 = ~n21883 ;
  assign y7963 = ~1'b0 ;
  assign y7964 = n21891 ;
  assign y7965 = n21902 ;
  assign y7966 = ~1'b0 ;
  assign y7967 = ~n21904 ;
  assign y7968 = ~n21906 ;
  assign y7969 = ~n21907 ;
  assign y7970 = ~n21909 ;
  assign y7971 = ~n21914 ;
  assign y7972 = ~n21915 ;
  assign y7973 = ~n21918 ;
  assign y7974 = n21923 ;
  assign y7975 = n21927 ;
  assign y7976 = ~1'b0 ;
  assign y7977 = ~n21930 ;
  assign y7978 = n21935 ;
  assign y7979 = n21936 ;
  assign y7980 = ~n21937 ;
  assign y7981 = n21938 ;
  assign y7982 = n21939 ;
  assign y7983 = ~n21942 ;
  assign y7984 = ~n7880 ;
  assign y7985 = n21946 ;
  assign y7986 = n21947 ;
  assign y7987 = ~n21952 ;
  assign y7988 = ~n21955 ;
  assign y7989 = ~1'b0 ;
  assign y7990 = n21959 ;
  assign y7991 = ~1'b0 ;
  assign y7992 = ~1'b0 ;
  assign y7993 = n21960 ;
  assign y7994 = ~1'b0 ;
  assign y7995 = 1'b0 ;
  assign y7996 = n21961 ;
  assign y7997 = ~n21964 ;
  assign y7998 = ~n21965 ;
  assign y7999 = ~1'b0 ;
  assign y8000 = n9353 ;
  assign y8001 = n21974 ;
  assign y8002 = n21975 ;
  assign y8003 = n21977 ;
  assign y8004 = n21981 ;
  assign y8005 = ~1'b0 ;
  assign y8006 = ~1'b0 ;
  assign y8007 = n21984 ;
  assign y8008 = n21985 ;
  assign y8009 = n21987 ;
  assign y8010 = ~n21992 ;
  assign y8011 = n21995 ;
  assign y8012 = ~1'b0 ;
  assign y8013 = ~n21999 ;
  assign y8014 = ~1'b0 ;
  assign y8015 = n22003 ;
  assign y8016 = ~n22007 ;
  assign y8017 = ~n22008 ;
  assign y8018 = n22009 ;
  assign y8019 = n22010 ;
  assign y8020 = n22014 ;
  assign y8021 = ~n22015 ;
  assign y8022 = ~1'b0 ;
  assign y8023 = n22020 ;
  assign y8024 = n22021 ;
  assign y8025 = n22022 ;
  assign y8026 = n22023 ;
  assign y8027 = ~1'b0 ;
  assign y8028 = n22024 ;
  assign y8029 = ~n22025 ;
  assign y8030 = n22027 ;
  assign y8031 = ~n22030 ;
  assign y8032 = ~1'b0 ;
  assign y8033 = ~1'b0 ;
  assign y8034 = n22031 ;
  assign y8035 = ~1'b0 ;
  assign y8036 = ~n22032 ;
  assign y8037 = 1'b0 ;
  assign y8038 = ~n22033 ;
  assign y8039 = n22045 ;
  assign y8040 = n22047 ;
  assign y8041 = n22052 ;
  assign y8042 = ~n22054 ;
  assign y8043 = ~n22058 ;
  assign y8044 = ~1'b0 ;
  assign y8045 = ~n22064 ;
  assign y8046 = n22066 ;
  assign y8047 = ~n22067 ;
  assign y8048 = ~1'b0 ;
  assign y8049 = n22069 ;
  assign y8050 = ~n22074 ;
  assign y8051 = ~n22077 ;
  assign y8052 = n22078 ;
  assign y8053 = ~n4827 ;
  assign y8054 = ~n22079 ;
  assign y8055 = n22080 ;
  assign y8056 = ~n22082 ;
  assign y8057 = ~1'b0 ;
  assign y8058 = n22085 ;
  assign y8059 = ~n22086 ;
  assign y8060 = n22087 ;
  assign y8061 = ~1'b0 ;
  assign y8062 = ~n22094 ;
  assign y8063 = ~n22096 ;
  assign y8064 = ~n22097 ;
  assign y8065 = ~n22101 ;
  assign y8066 = n22106 ;
  assign y8067 = ~1'b0 ;
  assign y8068 = ~n22110 ;
  assign y8069 = n22113 ;
  assign y8070 = ~1'b0 ;
  assign y8071 = n22114 ;
  assign y8072 = ~1'b0 ;
  assign y8073 = ~1'b0 ;
  assign y8074 = ~n22115 ;
  assign y8075 = ~1'b0 ;
  assign y8076 = n22128 ;
  assign y8077 = ~n22133 ;
  assign y8078 = ~n22135 ;
  assign y8079 = n22137 ;
  assign y8080 = ~n22139 ;
  assign y8081 = ~1'b0 ;
  assign y8082 = ~n22141 ;
  assign y8083 = ~n22142 ;
  assign y8084 = ~n14677 ;
  assign y8085 = ~n22145 ;
  assign y8086 = n22149 ;
  assign y8087 = ~1'b0 ;
  assign y8088 = n22157 ;
  assign y8089 = ~n12904 ;
  assign y8090 = ~1'b0 ;
  assign y8091 = ~1'b0 ;
  assign y8092 = ~n22162 ;
  assign y8093 = ~1'b0 ;
  assign y8094 = n22164 ;
  assign y8095 = n22166 ;
  assign y8096 = n22171 ;
  assign y8097 = n22177 ;
  assign y8098 = n22185 ;
  assign y8099 = n22186 ;
  assign y8100 = ~n22188 ;
  assign y8101 = ~n22189 ;
  assign y8102 = ~n22193 ;
  assign y8103 = ~1'b0 ;
  assign y8104 = n22195 ;
  assign y8105 = ~1'b0 ;
  assign y8106 = ~1'b0 ;
  assign y8107 = n22197 ;
  assign y8108 = n22198 ;
  assign y8109 = n22199 ;
  assign y8110 = n22204 ;
  assign y8111 = n22205 ;
  assign y8112 = ~n22207 ;
  assign y8113 = ~n22212 ;
  assign y8114 = ~1'b0 ;
  assign y8115 = ~1'b0 ;
  assign y8116 = ~1'b0 ;
  assign y8117 = ~n22213 ;
  assign y8118 = ~n22219 ;
  assign y8119 = ~n22225 ;
  assign y8120 = n22229 ;
  assign y8121 = n22231 ;
  assign y8122 = ~n22233 ;
  assign y8123 = ~1'b0 ;
  assign y8124 = ~1'b0 ;
  assign y8125 = ~n22234 ;
  assign y8126 = ~n22235 ;
  assign y8127 = n16067 ;
  assign y8128 = ~1'b0 ;
  assign y8129 = ~n22238 ;
  assign y8130 = n22240 ;
  assign y8131 = ~n22242 ;
  assign y8132 = ~n13077 ;
  assign y8133 = n22244 ;
  assign y8134 = n22246 ;
  assign y8135 = ~n22247 ;
  assign y8136 = ~n22251 ;
  assign y8137 = ~1'b0 ;
  assign y8138 = ~1'b0 ;
  assign y8139 = n22253 ;
  assign y8140 = n22263 ;
  assign y8141 = ~1'b0 ;
  assign y8142 = ~1'b0 ;
  assign y8143 = ~n22265 ;
  assign y8144 = ~1'b0 ;
  assign y8145 = ~n22266 ;
  assign y8146 = n22270 ;
  assign y8147 = n22271 ;
  assign y8148 = ~1'b0 ;
  assign y8149 = n22272 ;
  assign y8150 = n22273 ;
  assign y8151 = ~n22274 ;
  assign y8152 = ~n22276 ;
  assign y8153 = ~n22281 ;
  assign y8154 = ~n22285 ;
  assign y8155 = ~n22298 ;
  assign y8156 = n22300 ;
  assign y8157 = n22302 ;
  assign y8158 = 1'b0 ;
  assign y8159 = ~n22305 ;
  assign y8160 = ~n22308 ;
  assign y8161 = ~n22313 ;
  assign y8162 = ~n22317 ;
  assign y8163 = ~n2727 ;
  assign y8164 = ~1'b0 ;
  assign y8165 = ~1'b0 ;
  assign y8166 = ~n22318 ;
  assign y8167 = ~n22319 ;
  assign y8168 = ~n22324 ;
  assign y8169 = n22328 ;
  assign y8170 = ~n22332 ;
  assign y8171 = ~1'b0 ;
  assign y8172 = ~n22336 ;
  assign y8173 = ~n22342 ;
  assign y8174 = n22343 ;
  assign y8175 = n22344 ;
  assign y8176 = ~n22345 ;
  assign y8177 = n22348 ;
  assign y8178 = n22352 ;
  assign y8179 = ~1'b0 ;
  assign y8180 = ~n22357 ;
  assign y8181 = ~n22359 ;
  assign y8182 = ~1'b0 ;
  assign y8183 = ~n22362 ;
  assign y8184 = ~n22363 ;
  assign y8185 = ~n22364 ;
  assign y8186 = n22367 ;
  assign y8187 = n22369 ;
  assign y8188 = ~n22370 ;
  assign y8189 = n22374 ;
  assign y8190 = n22376 ;
  assign y8191 = ~n22379 ;
  assign y8192 = ~1'b0 ;
  assign y8193 = n22382 ;
  assign y8194 = ~n22385 ;
  assign y8195 = n22391 ;
  assign y8196 = n22395 ;
  assign y8197 = ~1'b0 ;
  assign y8198 = ~n22396 ;
  assign y8199 = n6865 ;
  assign y8200 = ~n22400 ;
  assign y8201 = ~1'b0 ;
  assign y8202 = ~n22402 ;
  assign y8203 = ~1'b0 ;
  assign y8204 = ~n22409 ;
  assign y8205 = ~n22419 ;
  assign y8206 = ~n22422 ;
  assign y8207 = ~n22427 ;
  assign y8208 = n22428 ;
  assign y8209 = ~1'b0 ;
  assign y8210 = ~1'b0 ;
  assign y8211 = n22436 ;
  assign y8212 = ~n22444 ;
  assign y8213 = n22445 ;
  assign y8214 = ~1'b0 ;
  assign y8215 = n22447 ;
  assign y8216 = ~n22449 ;
  assign y8217 = ~n22456 ;
  assign y8218 = ~1'b0 ;
  assign y8219 = n22458 ;
  assign y8220 = n22461 ;
  assign y8221 = n22463 ;
  assign y8222 = ~1'b0 ;
  assign y8223 = n22466 ;
  assign y8224 = ~1'b0 ;
  assign y8225 = ~1'b0 ;
  assign y8226 = ~n22468 ;
  assign y8227 = ~n22471 ;
  assign y8228 = ~n22474 ;
  assign y8229 = ~n22481 ;
  assign y8230 = ~n22483 ;
  assign y8231 = ~1'b0 ;
  assign y8232 = ~1'b0 ;
  assign y8233 = n22484 ;
  assign y8234 = ~n22489 ;
  assign y8235 = ~n22492 ;
  assign y8236 = n22494 ;
  assign y8237 = n22498 ;
  assign y8238 = n22502 ;
  assign y8239 = n22504 ;
  assign y8240 = n22506 ;
  assign y8241 = n22508 ;
  assign y8242 = n22511 ;
  assign y8243 = n22513 ;
  assign y8244 = n22525 ;
  assign y8245 = n22528 ;
  assign y8246 = n22531 ;
  assign y8247 = n22535 ;
  assign y8248 = ~n22537 ;
  assign y8249 = n22539 ;
  assign y8250 = n22543 ;
  assign y8251 = n22551 ;
  assign y8252 = n22560 ;
  assign y8253 = ~1'b0 ;
  assign y8254 = ~n22562 ;
  assign y8255 = ~1'b0 ;
  assign y8256 = n22563 ;
  assign y8257 = ~n22565 ;
  assign y8258 = n22566 ;
  assign y8259 = ~1'b0 ;
  assign y8260 = ~1'b0 ;
  assign y8261 = ~n22568 ;
  assign y8262 = ~n22573 ;
  assign y8263 = ~n22577 ;
  assign y8264 = n22579 ;
  assign y8265 = ~n22580 ;
  assign y8266 = n22582 ;
  assign y8267 = ~n22584 ;
  assign y8268 = ~n22585 ;
  assign y8269 = ~n22587 ;
  assign y8270 = ~n22589 ;
  assign y8271 = n22591 ;
  assign y8272 = ~n22596 ;
  assign y8273 = ~n22600 ;
  assign y8274 = n22601 ;
  assign y8275 = ~n22602 ;
  assign y8276 = n22608 ;
  assign y8277 = n22609 ;
  assign y8278 = ~1'b0 ;
  assign y8279 = ~n22626 ;
  assign y8280 = n22632 ;
  assign y8281 = ~n22634 ;
  assign y8282 = ~n22636 ;
  assign y8283 = n22637 ;
  assign y8284 = ~n22638 ;
  assign y8285 = ~n22640 ;
  assign y8286 = ~n22642 ;
  assign y8287 = ~n22646 ;
  assign y8288 = n22648 ;
  assign y8289 = ~n22650 ;
  assign y8290 = ~n22652 ;
  assign y8291 = ~1'b0 ;
  assign y8292 = n8734 ;
  assign y8293 = ~n22658 ;
  assign y8294 = ~n22659 ;
  assign y8295 = n22660 ;
  assign y8296 = n22661 ;
  assign y8297 = n22663 ;
  assign y8298 = ~n22665 ;
  assign y8299 = ~n22668 ;
  assign y8300 = ~1'b0 ;
  assign y8301 = n22669 ;
  assign y8302 = ~n2351 ;
  assign y8303 = ~n22671 ;
  assign y8304 = ~n22672 ;
  assign y8305 = ~n22674 ;
  assign y8306 = ~n22685 ;
  assign y8307 = ~n22698 ;
  assign y8308 = n22700 ;
  assign y8309 = ~n22702 ;
  assign y8310 = ~n22705 ;
  assign y8311 = ~n22708 ;
  assign y8312 = ~n22717 ;
  assign y8313 = n22719 ;
  assign y8314 = ~n22721 ;
  assign y8315 = ~n22727 ;
  assign y8316 = ~n22730 ;
  assign y8317 = n22732 ;
  assign y8318 = n22742 ;
  assign y8319 = n22744 ;
  assign y8320 = n22749 ;
  assign y8321 = ~n22751 ;
  assign y8322 = ~n22752 ;
  assign y8323 = ~1'b0 ;
  assign y8324 = ~1'b0 ;
  assign y8325 = n4581 ;
  assign y8326 = ~n22753 ;
  assign y8327 = ~1'b0 ;
  assign y8328 = n22760 ;
  assign y8329 = ~n22761 ;
  assign y8330 = ~n22762 ;
  assign y8331 = ~n22763 ;
  assign y8332 = n22771 ;
  assign y8333 = n22787 ;
  assign y8334 = ~1'b0 ;
  assign y8335 = ~n22791 ;
  assign y8336 = n22792 ;
  assign y8337 = ~n22793 ;
  assign y8338 = ~n22801 ;
  assign y8339 = ~n22804 ;
  assign y8340 = ~n22806 ;
  assign y8341 = n22807 ;
  assign y8342 = ~n22808 ;
  assign y8343 = n22813 ;
  assign y8344 = n22814 ;
  assign y8345 = ~n22819 ;
  assign y8346 = n22826 ;
  assign y8347 = n22834 ;
  assign y8348 = ~n22837 ;
  assign y8349 = ~n22838 ;
  assign y8350 = ~n22843 ;
  assign y8351 = ~n22848 ;
  assign y8352 = n22851 ;
  assign y8353 = n22859 ;
  assign y8354 = ~n22860 ;
  assign y8355 = ~n22863 ;
  assign y8356 = ~1'b0 ;
  assign y8357 = ~1'b0 ;
  assign y8358 = ~n22865 ;
  assign y8359 = ~n22866 ;
  assign y8360 = n22869 ;
  assign y8361 = n22877 ;
  assign y8362 = ~1'b0 ;
  assign y8363 = n22881 ;
  assign y8364 = ~n22884 ;
  assign y8365 = ~1'b0 ;
  assign y8366 = ~n22890 ;
  assign y8367 = ~n22893 ;
  assign y8368 = n22894 ;
  assign y8369 = ~1'b0 ;
  assign y8370 = ~n22900 ;
  assign y8371 = n15023 ;
  assign y8372 = n22902 ;
  assign y8373 = ~n22909 ;
  assign y8374 = ~1'b0 ;
  assign y8375 = ~n22911 ;
  assign y8376 = n22912 ;
  assign y8377 = ~n22914 ;
  assign y8378 = ~n22918 ;
  assign y8379 = ~1'b0 ;
  assign y8380 = n22921 ;
  assign y8381 = n22926 ;
  assign y8382 = n22931 ;
  assign y8383 = n22934 ;
  assign y8384 = ~1'b0 ;
  assign y8385 = ~1'b0 ;
  assign y8386 = ~n22937 ;
  assign y8387 = ~n22939 ;
  assign y8388 = n22941 ;
  assign y8389 = ~n22945 ;
  assign y8390 = n22947 ;
  assign y8391 = ~n22949 ;
  assign y8392 = ~1'b0 ;
  assign y8393 = ~n22951 ;
  assign y8394 = ~n22953 ;
  assign y8395 = n22960 ;
  assign y8396 = ~1'b0 ;
  assign y8397 = ~n22963 ;
  assign y8398 = ~1'b0 ;
  assign y8399 = ~1'b0 ;
  assign y8400 = n22964 ;
  assign y8401 = ~n22966 ;
  assign y8402 = ~n22968 ;
  assign y8403 = ~n22969 ;
  assign y8404 = ~1'b0 ;
  assign y8405 = ~n22970 ;
  assign y8406 = n22971 ;
  assign y8407 = n22972 ;
  assign y8408 = ~n22974 ;
  assign y8409 = n22977 ;
  assign y8410 = n22979 ;
  assign y8411 = n22983 ;
  assign y8412 = n22984 ;
  assign y8413 = ~n22986 ;
  assign y8414 = ~n22988 ;
  assign y8415 = ~n22989 ;
  assign y8416 = n22996 ;
  assign y8417 = ~1'b0 ;
  assign y8418 = n22998 ;
  assign y8419 = n23001 ;
  assign y8420 = ~n23007 ;
  assign y8421 = n23010 ;
  assign y8422 = ~1'b0 ;
  assign y8423 = n23015 ;
  assign y8424 = n23018 ;
  assign y8425 = ~n23020 ;
  assign y8426 = n23023 ;
  assign y8427 = n23025 ;
  assign y8428 = n23033 ;
  assign y8429 = ~1'b0 ;
  assign y8430 = n23041 ;
  assign y8431 = ~n23045 ;
  assign y8432 = n23047 ;
  assign y8433 = ~n23051 ;
  assign y8434 = 1'b0 ;
  assign y8435 = ~1'b0 ;
  assign y8436 = ~n23052 ;
  assign y8437 = ~n23060 ;
  assign y8438 = ~n23061 ;
  assign y8439 = 1'b0 ;
  assign y8440 = ~1'b0 ;
  assign y8441 = ~n23066 ;
  assign y8442 = n8764 ;
  assign y8443 = n23071 ;
  assign y8444 = ~1'b0 ;
  assign y8445 = ~n23076 ;
  assign y8446 = ~n23077 ;
  assign y8447 = ~n23078 ;
  assign y8448 = ~n23080 ;
  assign y8449 = n23088 ;
  assign y8450 = ~n23095 ;
  assign y8451 = n23096 ;
  assign y8452 = n23100 ;
  assign y8453 = n23104 ;
  assign y8454 = ~n23110 ;
  assign y8455 = n23112 ;
  assign y8456 = ~1'b0 ;
  assign y8457 = ~n23113 ;
  assign y8458 = ~n23114 ;
  assign y8459 = ~1'b0 ;
  assign y8460 = ~n23120 ;
  assign y8461 = ~n23124 ;
  assign y8462 = n23126 ;
  assign y8463 = ~n23129 ;
  assign y8464 = n23131 ;
  assign y8465 = n23133 ;
  assign y8466 = ~n23134 ;
  assign y8467 = ~n23136 ;
  assign y8468 = n23139 ;
  assign y8469 = ~1'b0 ;
  assign y8470 = ~n23142 ;
  assign y8471 = n23145 ;
  assign y8472 = ~n23146 ;
  assign y8473 = n23148 ;
  assign y8474 = ~n23150 ;
  assign y8475 = ~n23151 ;
  assign y8476 = n23153 ;
  assign y8477 = ~n10157 ;
  assign y8478 = ~1'b0 ;
  assign y8479 = ~n23155 ;
  assign y8480 = ~n23158 ;
  assign y8481 = ~n23161 ;
  assign y8482 = n365 ;
  assign y8483 = ~1'b0 ;
  assign y8484 = n23162 ;
  assign y8485 = ~1'b0 ;
  assign y8486 = ~1'b0 ;
  assign y8487 = n23171 ;
  assign y8488 = n23175 ;
  assign y8489 = ~n23178 ;
  assign y8490 = ~n23186 ;
  assign y8491 = ~n9156 ;
  assign y8492 = n23187 ;
  assign y8493 = ~n10900 ;
  assign y8494 = n23188 ;
  assign y8495 = ~1'b0 ;
  assign y8496 = n23190 ;
  assign y8497 = ~n23194 ;
  assign y8498 = ~n23200 ;
  assign y8499 = ~n23203 ;
  assign y8500 = ~1'b0 ;
  assign y8501 = ~n23205 ;
  assign y8502 = ~1'b0 ;
  assign y8503 = ~n23207 ;
  assign y8504 = n23208 ;
  assign y8505 = ~1'b0 ;
  assign y8506 = n23209 ;
  assign y8507 = n22108 ;
  assign y8508 = ~n23210 ;
  assign y8509 = ~n23213 ;
  assign y8510 = ~n23214 ;
  assign y8511 = ~n23218 ;
  assign y8512 = ~n23221 ;
  assign y8513 = n23225 ;
  assign y8514 = ~n23227 ;
  assign y8515 = ~n23235 ;
  assign y8516 = ~1'b0 ;
  assign y8517 = ~n23238 ;
  assign y8518 = ~n23241 ;
  assign y8519 = n23242 ;
  assign y8520 = ~n23248 ;
  assign y8521 = ~n12340 ;
  assign y8522 = ~n23251 ;
  assign y8523 = ~n23253 ;
  assign y8524 = ~n23255 ;
  assign y8525 = n23259 ;
  assign y8526 = ~n23260 ;
  assign y8527 = ~1'b0 ;
  assign y8528 = ~n23261 ;
  assign y8529 = ~n23267 ;
  assign y8530 = ~1'b0 ;
  assign y8531 = n23269 ;
  assign y8532 = n23272 ;
  assign y8533 = ~n23275 ;
  assign y8534 = ~n23278 ;
  assign y8535 = ~n23281 ;
  assign y8536 = ~n23285 ;
  assign y8537 = ~n23288 ;
  assign y8538 = ~1'b0 ;
  assign y8539 = ~n23290 ;
  assign y8540 = ~n23293 ;
  assign y8541 = ~n23295 ;
  assign y8542 = ~n4274 ;
  assign y8543 = n23302 ;
  assign y8544 = ~1'b0 ;
  assign y8545 = n23305 ;
  assign y8546 = ~n23307 ;
  assign y8547 = ~n23308 ;
  assign y8548 = n23309 ;
  assign y8549 = ~n23312 ;
  assign y8550 = ~n23313 ;
  assign y8551 = n23323 ;
  assign y8552 = ~1'b0 ;
  assign y8553 = ~1'b0 ;
  assign y8554 = n23325 ;
  assign y8555 = ~n23327 ;
  assign y8556 = n23329 ;
  assign y8557 = ~n23331 ;
  assign y8558 = n23332 ;
  assign y8559 = ~n23334 ;
  assign y8560 = ~1'b0 ;
  assign y8561 = n13656 ;
  assign y8562 = n23337 ;
  assign y8563 = n23341 ;
  assign y8564 = ~n23345 ;
  assign y8565 = ~n23352 ;
  assign y8566 = n23354 ;
  assign y8567 = ~1'b0 ;
  assign y8568 = n23357 ;
  assign y8569 = n23359 ;
  assign y8570 = n23360 ;
  assign y8571 = ~1'b0 ;
  assign y8572 = n23364 ;
  assign y8573 = ~n23365 ;
  assign y8574 = ~n23366 ;
  assign y8575 = 1'b0 ;
  assign y8576 = n23367 ;
  assign y8577 = ~n23368 ;
  assign y8578 = ~n23369 ;
  assign y8579 = ~1'b0 ;
  assign y8580 = n23372 ;
  assign y8581 = 1'b0 ;
  assign y8582 = ~n23378 ;
  assign y8583 = ~1'b0 ;
  assign y8584 = n23379 ;
  assign y8585 = ~1'b0 ;
  assign y8586 = ~1'b0 ;
  assign y8587 = n23381 ;
  assign y8588 = n23385 ;
  assign y8589 = ~n23390 ;
  assign y8590 = n23396 ;
  assign y8591 = n23398 ;
  assign y8592 = n23402 ;
  assign y8593 = ~n23407 ;
  assign y8594 = ~1'b0 ;
  assign y8595 = ~n23411 ;
  assign y8596 = ~n23413 ;
  assign y8597 = ~1'b0 ;
  assign y8598 = ~n23417 ;
  assign y8599 = n23420 ;
  assign y8600 = ~n23422 ;
  assign y8601 = n23423 ;
  assign y8602 = ~n23425 ;
  assign y8603 = n23426 ;
  assign y8604 = ~n23429 ;
  assign y8605 = n23432 ;
  assign y8606 = ~n23435 ;
  assign y8607 = ~1'b0 ;
  assign y8608 = ~1'b0 ;
  assign y8609 = n23437 ;
  assign y8610 = n23441 ;
  assign y8611 = ~n23442 ;
  assign y8612 = ~n23445 ;
  assign y8613 = ~n23450 ;
  assign y8614 = n23454 ;
  assign y8615 = n23459 ;
  assign y8616 = ~n23464 ;
  assign y8617 = ~1'b0 ;
  assign y8618 = n23465 ;
  assign y8619 = ~n23466 ;
  assign y8620 = ~n23472 ;
  assign y8621 = n23474 ;
  assign y8622 = ~1'b0 ;
  assign y8623 = n23475 ;
  assign y8624 = ~1'b0 ;
  assign y8625 = ~n23479 ;
  assign y8626 = ~n23484 ;
  assign y8627 = n2824 ;
  assign y8628 = n23489 ;
  assign y8629 = ~n23491 ;
  assign y8630 = ~n23493 ;
  assign y8631 = ~1'b0 ;
  assign y8632 = n23496 ;
  assign y8633 = ~n23500 ;
  assign y8634 = ~1'b0 ;
  assign y8635 = n23507 ;
  assign y8636 = ~n23520 ;
  assign y8637 = ~1'b0 ;
  assign y8638 = ~n10372 ;
  assign y8639 = ~n23521 ;
  assign y8640 = ~n23523 ;
  assign y8641 = n23528 ;
  assign y8642 = ~n23530 ;
  assign y8643 = ~1'b0 ;
  assign y8644 = ~n23533 ;
  assign y8645 = n23537 ;
  assign y8646 = n23543 ;
  assign y8647 = n23548 ;
  assign y8648 = ~1'b0 ;
  assign y8649 = ~n23553 ;
  assign y8650 = n23558 ;
  assign y8651 = n23561 ;
  assign y8652 = ~1'b0 ;
  assign y8653 = ~n23568 ;
  assign y8654 = n23570 ;
  assign y8655 = 1'b0 ;
  assign y8656 = n23573 ;
  assign y8657 = ~1'b0 ;
  assign y8658 = ~n23574 ;
  assign y8659 = ~1'b0 ;
  assign y8660 = n23575 ;
  assign y8661 = n23579 ;
  assign y8662 = ~n23581 ;
  assign y8663 = n23582 ;
  assign y8664 = n23585 ;
  assign y8665 = ~n23595 ;
  assign y8666 = n23596 ;
  assign y8667 = n23598 ;
  assign y8668 = n23600 ;
  assign y8669 = ~n485 ;
  assign y8670 = ~n23603 ;
  assign y8671 = ~n23607 ;
  assign y8672 = n23611 ;
  assign y8673 = ~n23613 ;
  assign y8674 = ~n23615 ;
  assign y8675 = ~n23621 ;
  assign y8676 = ~n1034 ;
  assign y8677 = ~1'b0 ;
  assign y8678 = ~n23627 ;
  assign y8679 = ~n23639 ;
  assign y8680 = ~n13696 ;
  assign y8681 = n23644 ;
  assign y8682 = ~1'b0 ;
  assign y8683 = ~1'b0 ;
  assign y8684 = n23645 ;
  assign y8685 = ~n23646 ;
  assign y8686 = 1'b0 ;
  assign y8687 = ~n23653 ;
  assign y8688 = ~n23655 ;
  assign y8689 = ~1'b0 ;
  assign y8690 = n23656 ;
  assign y8691 = ~n23658 ;
  assign y8692 = ~n23659 ;
  assign y8693 = n23661 ;
  assign y8694 = ~n23662 ;
  assign y8695 = ~n23664 ;
  assign y8696 = n23668 ;
  assign y8697 = ~1'b0 ;
  assign y8698 = n23672 ;
  assign y8699 = n23673 ;
  assign y8700 = n23678 ;
  assign y8701 = n23679 ;
  assign y8702 = 1'b0 ;
  assign y8703 = ~n23688 ;
  assign y8704 = n23689 ;
  assign y8705 = ~n23691 ;
  assign y8706 = n23693 ;
  assign y8707 = ~1'b0 ;
  assign y8708 = n23697 ;
  assign y8709 = n23698 ;
  assign y8710 = n23710 ;
  assign y8711 = ~n23713 ;
  assign y8712 = ~n23715 ;
  assign y8713 = n23717 ;
  assign y8714 = ~n23720 ;
  assign y8715 = ~n23723 ;
  assign y8716 = 1'b0 ;
  assign y8717 = ~1'b0 ;
  assign y8718 = ~1'b0 ;
  assign y8719 = n23724 ;
  assign y8720 = n23726 ;
  assign y8721 = ~n23728 ;
  assign y8722 = ~n23730 ;
  assign y8723 = ~n23731 ;
  assign y8724 = ~n23732 ;
  assign y8725 = ~n23733 ;
  assign y8726 = ~n23736 ;
  assign y8727 = ~n23746 ;
  assign y8728 = ~n23751 ;
  assign y8729 = ~n23754 ;
  assign y8730 = ~n23762 ;
  assign y8731 = ~1'b0 ;
  assign y8732 = n23765 ;
  assign y8733 = n11116 ;
  assign y8734 = n23766 ;
  assign y8735 = n23768 ;
  assign y8736 = n23775 ;
  assign y8737 = n23776 ;
  assign y8738 = n23778 ;
  assign y8739 = ~1'b0 ;
  assign y8740 = n23780 ;
  assign y8741 = n23782 ;
  assign y8742 = ~n23785 ;
  assign y8743 = ~n23787 ;
  assign y8744 = ~n23790 ;
  assign y8745 = ~n23793 ;
  assign y8746 = n23794 ;
  assign y8747 = n23801 ;
  assign y8748 = ~n23803 ;
  assign y8749 = n23804 ;
  assign y8750 = ~n2355 ;
  assign y8751 = ~n23805 ;
  assign y8752 = ~n23806 ;
  assign y8753 = n23811 ;
  assign y8754 = ~1'b0 ;
  assign y8755 = n23813 ;
  assign y8756 = n23815 ;
  assign y8757 = n23818 ;
  assign y8758 = n23823 ;
  assign y8759 = ~n23824 ;
  assign y8760 = ~n23826 ;
  assign y8761 = ~1'b0 ;
  assign y8762 = ~1'b0 ;
  assign y8763 = ~n23827 ;
  assign y8764 = ~1'b0 ;
  assign y8765 = n23828 ;
  assign y8766 = ~n23830 ;
  assign y8767 = n23833 ;
  assign y8768 = ~n23839 ;
  assign y8769 = 1'b0 ;
  assign y8770 = n23842 ;
  assign y8771 = ~n23848 ;
  assign y8772 = n23850 ;
  assign y8773 = ~n23851 ;
  assign y8774 = ~n2469 ;
  assign y8775 = ~n23859 ;
  assign y8776 = n5627 ;
  assign y8777 = n23861 ;
  assign y8778 = ~n23865 ;
  assign y8779 = ~n23869 ;
  assign y8780 = ~n23871 ;
  assign y8781 = n23877 ;
  assign y8782 = ~n2289 ;
  assign y8783 = 1'b0 ;
  assign y8784 = ~n23883 ;
  assign y8785 = n23886 ;
  assign y8786 = n23890 ;
  assign y8787 = n23891 ;
  assign y8788 = n23893 ;
  assign y8789 = ~n23895 ;
  assign y8790 = n23902 ;
  assign y8791 = ~1'b0 ;
  assign y8792 = ~n23905 ;
  assign y8793 = ~n23907 ;
  assign y8794 = n23910 ;
  assign y8795 = ~n23912 ;
  assign y8796 = ~1'b0 ;
  assign y8797 = n23918 ;
  assign y8798 = ~1'b0 ;
  assign y8799 = ~1'b0 ;
  assign y8800 = ~n23919 ;
  assign y8801 = n23921 ;
  assign y8802 = ~1'b0 ;
  assign y8803 = ~n23922 ;
  assign y8804 = ~n23928 ;
  assign y8805 = ~1'b0 ;
  assign y8806 = 1'b0 ;
  assign y8807 = n23929 ;
  assign y8808 = ~1'b0 ;
  assign y8809 = ~n23930 ;
  assign y8810 = ~1'b0 ;
  assign y8811 = ~n23935 ;
  assign y8812 = ~n23937 ;
  assign y8813 = ~1'b0 ;
  assign y8814 = ~1'b0 ;
  assign y8815 = ~1'b0 ;
  assign y8816 = ~n23938 ;
  assign y8817 = n23939 ;
  assign y8818 = ~n23942 ;
  assign y8819 = n23945 ;
  assign y8820 = n23947 ;
  assign y8821 = n23949 ;
  assign y8822 = ~n23951 ;
  assign y8823 = ~n23952 ;
  assign y8824 = ~1'b0 ;
  assign y8825 = n23956 ;
  assign y8826 = n17921 ;
  assign y8827 = ~n23957 ;
  assign y8828 = ~1'b0 ;
  assign y8829 = ~n23959 ;
  assign y8830 = ~n23975 ;
  assign y8831 = ~n23976 ;
  assign y8832 = n23977 ;
  assign y8833 = ~n23980 ;
  assign y8834 = ~n23982 ;
  assign y8835 = n23985 ;
  assign y8836 = ~n23987 ;
  assign y8837 = n23990 ;
  assign y8838 = n23993 ;
  assign y8839 = ~n23995 ;
  assign y8840 = ~1'b0 ;
  assign y8841 = ~n19479 ;
  assign y8842 = ~n23996 ;
  assign y8843 = ~n23998 ;
  assign y8844 = ~1'b0 ;
  assign y8845 = n24008 ;
  assign y8846 = 1'b0 ;
  assign y8847 = n24010 ;
  assign y8848 = ~1'b0 ;
  assign y8849 = ~n24016 ;
  assign y8850 = n24017 ;
  assign y8851 = ~n24020 ;
  assign y8852 = ~1'b0 ;
  assign y8853 = ~n24022 ;
  assign y8854 = ~1'b0 ;
  assign y8855 = ~1'b0 ;
  assign y8856 = n24027 ;
  assign y8857 = n24029 ;
  assign y8858 = n24030 ;
  assign y8859 = ~n24034 ;
  assign y8860 = ~n24038 ;
  assign y8861 = ~n24041 ;
  assign y8862 = n24043 ;
  assign y8863 = ~1'b0 ;
  assign y8864 = n24044 ;
  assign y8865 = ~n24045 ;
  assign y8866 = n24048 ;
  assign y8867 = ~n24050 ;
  assign y8868 = ~n24055 ;
  assign y8869 = n24063 ;
  assign y8870 = n24068 ;
  assign y8871 = ~n24074 ;
  assign y8872 = ~n24075 ;
  assign y8873 = ~n24081 ;
  assign y8874 = ~n24083 ;
  assign y8875 = ~1'b0 ;
  assign y8876 = ~n24090 ;
  assign y8877 = n24093 ;
  assign y8878 = n24098 ;
  assign y8879 = ~1'b0 ;
  assign y8880 = n24100 ;
  assign y8881 = ~1'b0 ;
  assign y8882 = n24101 ;
  assign y8883 = ~n24107 ;
  assign y8884 = ~1'b0 ;
  assign y8885 = ~n24109 ;
  assign y8886 = ~1'b0 ;
  assign y8887 = n24112 ;
  assign y8888 = ~1'b0 ;
  assign y8889 = n24119 ;
  assign y8890 = ~1'b0 ;
  assign y8891 = ~n24123 ;
  assign y8892 = ~n24124 ;
  assign y8893 = n24127 ;
  assign y8894 = ~n24128 ;
  assign y8895 = n24133 ;
  assign y8896 = n24135 ;
  assign y8897 = n9232 ;
  assign y8898 = n290 ;
  assign y8899 = 1'b0 ;
  assign y8900 = ~n24136 ;
  assign y8901 = ~1'b0 ;
  assign y8902 = n24137 ;
  assign y8903 = ~n24138 ;
  assign y8904 = ~n24139 ;
  assign y8905 = ~n24145 ;
  assign y8906 = n24152 ;
  assign y8907 = ~n24156 ;
  assign y8908 = n24160 ;
  assign y8909 = ~1'b0 ;
  assign y8910 = ~n24161 ;
  assign y8911 = n24162 ;
  assign y8912 = ~1'b0 ;
  assign y8913 = ~1'b0 ;
  assign y8914 = ~1'b0 ;
  assign y8915 = n24165 ;
  assign y8916 = ~1'b0 ;
  assign y8917 = ~1'b0 ;
  assign y8918 = ~n24170 ;
  assign y8919 = ~n24175 ;
  assign y8920 = ~n24178 ;
  assign y8921 = n24181 ;
  assign y8922 = 1'b0 ;
  assign y8923 = ~1'b0 ;
  assign y8924 = ~1'b0 ;
  assign y8925 = n24191 ;
  assign y8926 = n24199 ;
  assign y8927 = n292 ;
  assign y8928 = n24203 ;
  assign y8929 = ~x113 ;
  assign y8930 = ~n24205 ;
  assign y8931 = ~1'b0 ;
  assign y8932 = ~1'b0 ;
  assign y8933 = n20801 ;
  assign y8934 = n24208 ;
  assign y8935 = ~n24219 ;
  assign y8936 = n24220 ;
  assign y8937 = ~1'b0 ;
  assign y8938 = n24222 ;
  assign y8939 = n24224 ;
  assign y8940 = ~n24228 ;
  assign y8941 = ~n24234 ;
  assign y8942 = n24235 ;
  assign y8943 = ~n24240 ;
  assign y8944 = ~1'b0 ;
  assign y8945 = n24245 ;
  assign y8946 = n24246 ;
  assign y8947 = ~1'b0 ;
  assign y8948 = ~n24252 ;
  assign y8949 = n24253 ;
  assign y8950 = ~1'b0 ;
  assign y8951 = n24260 ;
  assign y8952 = n24262 ;
  assign y8953 = n24263 ;
  assign y8954 = ~n24266 ;
  assign y8955 = ~n24268 ;
  assign y8956 = ~1'b0 ;
  assign y8957 = n24269 ;
  assign y8958 = n24270 ;
  assign y8959 = n24277 ;
  assign y8960 = ~n24278 ;
  assign y8961 = ~1'b0 ;
  assign y8962 = ~n24281 ;
  assign y8963 = ~n24282 ;
  assign y8964 = ~1'b0 ;
  assign y8965 = ~1'b0 ;
  assign y8966 = 1'b0 ;
  assign y8967 = ~n24283 ;
  assign y8968 = ~n24286 ;
  assign y8969 = n24288 ;
  assign y8970 = ~1'b0 ;
  assign y8971 = ~n24290 ;
  assign y8972 = n24294 ;
  assign y8973 = n24295 ;
  assign y8974 = n24296 ;
  assign y8975 = ~n24298 ;
  assign y8976 = ~1'b0 ;
  assign y8977 = ~n24299 ;
  assign y8978 = ~n24302 ;
  assign y8979 = n24304 ;
  assign y8980 = n24308 ;
  assign y8981 = n24311 ;
  assign y8982 = ~n24313 ;
  assign y8983 = ~n24316 ;
  assign y8984 = ~n24318 ;
  assign y8985 = n24327 ;
  assign y8986 = n24329 ;
  assign y8987 = n24330 ;
  assign y8988 = ~n24331 ;
  assign y8989 = n24336 ;
  assign y8990 = n24340 ;
  assign y8991 = ~n24342 ;
  assign y8992 = n24348 ;
  assign y8993 = n24350 ;
  assign y8994 = ~1'b0 ;
  assign y8995 = ~n24353 ;
  assign y8996 = ~1'b0 ;
  assign y8997 = ~n24361 ;
  assign y8998 = ~1'b0 ;
  assign y8999 = ~n24365 ;
  assign y9000 = ~n24372 ;
  assign y9001 = n24376 ;
  assign y9002 = n24378 ;
  assign y9003 = ~1'b0 ;
  assign y9004 = ~n24381 ;
  assign y9005 = n24382 ;
  assign y9006 = ~1'b0 ;
  assign y9007 = ~n24385 ;
  assign y9008 = ~1'b0 ;
  assign y9009 = ~1'b0 ;
  assign y9010 = ~n24392 ;
  assign y9011 = n24393 ;
  assign y9012 = ~n24404 ;
  assign y9013 = n24405 ;
  assign y9014 = ~1'b0 ;
  assign y9015 = ~n24407 ;
  assign y9016 = ~1'b0 ;
  assign y9017 = n24409 ;
  assign y9018 = ~1'b0 ;
  assign y9019 = ~n24411 ;
  assign y9020 = ~n24417 ;
  assign y9021 = ~1'b0 ;
  assign y9022 = n24423 ;
  assign y9023 = ~n24425 ;
  assign y9024 = ~n24426 ;
  assign y9025 = n24427 ;
  assign y9026 = n24431 ;
  assign y9027 = ~n24433 ;
  assign y9028 = ~1'b0 ;
  assign y9029 = ~1'b0 ;
  assign y9030 = ~n24434 ;
  assign y9031 = n24439 ;
  assign y9032 = n24444 ;
  assign y9033 = ~1'b0 ;
  assign y9034 = ~1'b0 ;
  assign y9035 = n24452 ;
  assign y9036 = ~n24457 ;
  assign y9037 = n24458 ;
  assign y9038 = ~n24461 ;
  assign y9039 = ~n24465 ;
  assign y9040 = ~n24467 ;
  assign y9041 = n24469 ;
  assign y9042 = ~n24472 ;
  assign y9043 = ~1'b0 ;
  assign y9044 = ~1'b0 ;
  assign y9045 = n24479 ;
  assign y9046 = ~1'b0 ;
  assign y9047 = ~n24480 ;
  assign y9048 = n24482 ;
  assign y9049 = n24484 ;
  assign y9050 = n24486 ;
  assign y9051 = n24487 ;
  assign y9052 = n17072 ;
  assign y9053 = ~1'b0 ;
  assign y9054 = ~n24488 ;
  assign y9055 = ~n24492 ;
  assign y9056 = n24496 ;
  assign y9057 = n24499 ;
  assign y9058 = n24504 ;
  assign y9059 = ~n24507 ;
  assign y9060 = n24508 ;
  assign y9061 = ~n24510 ;
  assign y9062 = ~n24511 ;
  assign y9063 = n24512 ;
  assign y9064 = ~n5466 ;
  assign y9065 = ~1'b0 ;
  assign y9066 = n24513 ;
  assign y9067 = n24514 ;
  assign y9068 = n24515 ;
  assign y9069 = 1'b0 ;
  assign y9070 = ~1'b0 ;
  assign y9071 = n24516 ;
  assign y9072 = n24520 ;
  assign y9073 = n24524 ;
  assign y9074 = ~n24526 ;
  assign y9075 = n24529 ;
  assign y9076 = n24536 ;
  assign y9077 = n24538 ;
  assign y9078 = n24556 ;
  assign y9079 = ~n4240 ;
  assign y9080 = n24561 ;
  assign y9081 = n16106 ;
  assign y9082 = ~n24564 ;
  assign y9083 = ~n24565 ;
  assign y9084 = n12439 ;
  assign y9085 = ~n24567 ;
  assign y9086 = ~n24571 ;
  assign y9087 = ~1'b0 ;
  assign y9088 = ~n24580 ;
  assign y9089 = ~n24590 ;
  assign y9090 = ~n24592 ;
  assign y9091 = ~n24593 ;
  assign y9092 = ~n24594 ;
  assign y9093 = ~1'b0 ;
  assign y9094 = n24596 ;
  assign y9095 = ~n24601 ;
  assign y9096 = ~n24608 ;
  assign y9097 = ~n24609 ;
  assign y9098 = n24616 ;
  assign y9099 = ~n24617 ;
  assign y9100 = n20470 ;
  assign y9101 = n24620 ;
  assign y9102 = ~n24626 ;
  assign y9103 = n24627 ;
  assign y9104 = n24628 ;
  assign y9105 = ~1'b0 ;
  assign y9106 = ~1'b0 ;
  assign y9107 = ~n24631 ;
  assign y9108 = n24632 ;
  assign y9109 = ~n24633 ;
  assign y9110 = ~1'b0 ;
  assign y9111 = ~n24636 ;
  assign y9112 = n24644 ;
  assign y9113 = ~n24646 ;
  assign y9114 = ~1'b0 ;
  assign y9115 = ~1'b0 ;
  assign y9116 = n24648 ;
  assign y9117 = n24649 ;
  assign y9118 = n24650 ;
  assign y9119 = ~n24653 ;
  assign y9120 = ~n24655 ;
  assign y9121 = ~n24658 ;
  assign y9122 = ~1'b0 ;
  assign y9123 = ~n24660 ;
  assign y9124 = ~n24664 ;
  assign y9125 = ~1'b0 ;
  assign y9126 = ~n24667 ;
  assign y9127 = ~n24671 ;
  assign y9128 = n24673 ;
  assign y9129 = ~1'b0 ;
  assign y9130 = ~n24674 ;
  assign y9131 = n24676 ;
  assign y9132 = ~n6972 ;
  assign y9133 = ~n24680 ;
  assign y9134 = ~n24683 ;
  assign y9135 = ~n24687 ;
  assign y9136 = n24689 ;
  assign y9137 = ~1'b0 ;
  assign y9138 = ~1'b0 ;
  assign y9139 = ~1'b0 ;
  assign y9140 = n24693 ;
  assign y9141 = n24697 ;
  assign y9142 = ~n24703 ;
  assign y9143 = ~1'b0 ;
  assign y9144 = ~n24705 ;
  assign y9145 = ~1'b0 ;
  assign y9146 = ~1'b0 ;
  assign y9147 = ~n24712 ;
  assign y9148 = ~n24713 ;
  assign y9149 = ~n24714 ;
  assign y9150 = n5475 ;
  assign y9151 = n24716 ;
  assign y9152 = ~n24717 ;
  assign y9153 = ~1'b0 ;
  assign y9154 = ~n24720 ;
  assign y9155 = ~n24721 ;
  assign y9156 = ~n24724 ;
  assign y9157 = n24726 ;
  assign y9158 = n24727 ;
  assign y9159 = n24728 ;
  assign y9160 = ~n24729 ;
  assign y9161 = n24731 ;
  assign y9162 = n24733 ;
  assign y9163 = ~n24735 ;
  assign y9164 = ~n24740 ;
  assign y9165 = n24743 ;
  assign y9166 = ~n24744 ;
  assign y9167 = n24746 ;
  assign y9168 = ~n24752 ;
  assign y9169 = ~1'b0 ;
  assign y9170 = ~n24757 ;
  assign y9171 = ~n24760 ;
  assign y9172 = ~1'b0 ;
  assign y9173 = ~1'b0 ;
  assign y9174 = ~n24763 ;
  assign y9175 = ~n13040 ;
  assign y9176 = ~n24765 ;
  assign y9177 = ~n24766 ;
  assign y9178 = ~n24771 ;
  assign y9179 = ~n24773 ;
  assign y9180 = n24774 ;
  assign y9181 = ~n24776 ;
  assign y9182 = n24781 ;
  assign y9183 = ~n24786 ;
  assign y9184 = n24795 ;
  assign y9185 = ~n24799 ;
  assign y9186 = n24801 ;
  assign y9187 = n24803 ;
  assign y9188 = n24804 ;
  assign y9189 = n24809 ;
  assign y9190 = n24810 ;
  assign y9191 = ~n24811 ;
  assign y9192 = ~1'b0 ;
  assign y9193 = n24820 ;
  assign y9194 = ~1'b0 ;
  assign y9195 = n24821 ;
  assign y9196 = n24825 ;
  assign y9197 = n24827 ;
  assign y9198 = ~1'b0 ;
  assign y9199 = ~n24830 ;
  assign y9200 = n24832 ;
  assign y9201 = ~n4840 ;
  assign y9202 = ~n24836 ;
  assign y9203 = ~n24842 ;
  assign y9204 = ~n24844 ;
  assign y9205 = ~1'b0 ;
  assign y9206 = ~1'b0 ;
  assign y9207 = ~n1951 ;
  assign y9208 = n24847 ;
  assign y9209 = n24851 ;
  assign y9210 = ~n24852 ;
  assign y9211 = n24854 ;
  assign y9212 = ~1'b0 ;
  assign y9213 = ~1'b0 ;
  assign y9214 = n24856 ;
  assign y9215 = n24859 ;
  assign y9216 = n24865 ;
  assign y9217 = n24867 ;
  assign y9218 = ~1'b0 ;
  assign y9219 = n24869 ;
  assign y9220 = n24870 ;
  assign y9221 = n24871 ;
  assign y9222 = ~1'b0 ;
  assign y9223 = n24872 ;
  assign y9224 = n24873 ;
  assign y9225 = n24882 ;
  assign y9226 = ~n4685 ;
  assign y9227 = n24885 ;
  assign y9228 = ~1'b0 ;
  assign y9229 = ~n24889 ;
  assign y9230 = ~n24893 ;
  assign y9231 = n24894 ;
  assign y9232 = ~1'b0 ;
  assign y9233 = n24899 ;
  assign y9234 = ~n24901 ;
  assign y9235 = ~n24905 ;
  assign y9236 = n24906 ;
  assign y9237 = ~1'b0 ;
  assign y9238 = n24907 ;
  assign y9239 = ~n24909 ;
  assign y9240 = n24917 ;
  assign y9241 = ~n24918 ;
  assign y9242 = ~n4729 ;
  assign y9243 = n24921 ;
  assign y9244 = ~n24925 ;
  assign y9245 = n24926 ;
  assign y9246 = ~n24927 ;
  assign y9247 = n24930 ;
  assign y9248 = n24934 ;
  assign y9249 = ~n24936 ;
  assign y9250 = ~1'b0 ;
  assign y9251 = ~n24939 ;
  assign y9252 = n15417 ;
  assign y9253 = ~1'b0 ;
  assign y9254 = ~n24942 ;
  assign y9255 = ~1'b0 ;
  assign y9256 = n24943 ;
  assign y9257 = ~n24945 ;
  assign y9258 = n24948 ;
  assign y9259 = n24951 ;
  assign y9260 = n24957 ;
  assign y9261 = ~n24962 ;
  assign y9262 = n24964 ;
  assign y9263 = n24965 ;
  assign y9264 = n24966 ;
  assign y9265 = ~1'b0 ;
  assign y9266 = n24970 ;
  assign y9267 = ~1'b0 ;
  assign y9268 = ~n24972 ;
  assign y9269 = ~n24973 ;
  assign y9270 = n24979 ;
  assign y9271 = n24987 ;
  assign y9272 = ~n24988 ;
  assign y9273 = ~n24990 ;
  assign y9274 = ~1'b0 ;
  assign y9275 = ~n24992 ;
  assign y9276 = n24993 ;
  assign y9277 = n24994 ;
  assign y9278 = ~n25001 ;
  assign y9279 = n25008 ;
  assign y9280 = n25009 ;
  assign y9281 = n25013 ;
  assign y9282 = ~n25015 ;
  assign y9283 = n25018 ;
  assign y9284 = n25019 ;
  assign y9285 = ~1'b0 ;
  assign y9286 = ~1'b0 ;
  assign y9287 = ~1'b0 ;
  assign y9288 = ~n25023 ;
  assign y9289 = n25024 ;
  assign y9290 = ~n25026 ;
  assign y9291 = ~n25027 ;
  assign y9292 = n25028 ;
  assign y9293 = n25036 ;
  assign y9294 = ~1'b0 ;
  assign y9295 = ~n25038 ;
  assign y9296 = ~1'b0 ;
  assign y9297 = n25041 ;
  assign y9298 = n25043 ;
  assign y9299 = n25047 ;
  assign y9300 = n25048 ;
  assign y9301 = ~n25050 ;
  assign y9302 = n25051 ;
  assign y9303 = n5519 ;
  assign y9304 = ~n25053 ;
  assign y9305 = n25055 ;
  assign y9306 = ~n25056 ;
  assign y9307 = ~n25058 ;
  assign y9308 = n25060 ;
  assign y9309 = ~n25066 ;
  assign y9310 = ~1'b0 ;
  assign y9311 = n25071 ;
  assign y9312 = ~n25075 ;
  assign y9313 = ~n25076 ;
  assign y9314 = ~n25077 ;
  assign y9315 = n25085 ;
  assign y9316 = ~n25089 ;
  assign y9317 = n25090 ;
  assign y9318 = n25093 ;
  assign y9319 = ~n25099 ;
  assign y9320 = ~n25102 ;
  assign y9321 = ~n25105 ;
  assign y9322 = n25112 ;
  assign y9323 = ~n25116 ;
  assign y9324 = ~1'b0 ;
  assign y9325 = n25121 ;
  assign y9326 = ~n25125 ;
  assign y9327 = ~n25129 ;
  assign y9328 = ~1'b0 ;
  assign y9329 = ~n25133 ;
  assign y9330 = ~n25134 ;
  assign y9331 = n25135 ;
  assign y9332 = ~n25137 ;
  assign y9333 = ~n25140 ;
  assign y9334 = n25142 ;
  assign y9335 = ~n25143 ;
  assign y9336 = n25148 ;
  assign y9337 = n25150 ;
  assign y9338 = ~n25151 ;
  assign y9339 = n25152 ;
  assign y9340 = 1'b0 ;
  assign y9341 = n25154 ;
  assign y9342 = ~n25156 ;
  assign y9343 = ~n25157 ;
  assign y9344 = ~n25159 ;
  assign y9345 = ~n25167 ;
  assign y9346 = n25168 ;
  assign y9347 = ~n25173 ;
  assign y9348 = n25177 ;
  assign y9349 = n25178 ;
  assign y9350 = ~1'b0 ;
  assign y9351 = ~n25183 ;
  assign y9352 = ~n25186 ;
  assign y9353 = ~1'b0 ;
  assign y9354 = ~n25193 ;
  assign y9355 = ~1'b0 ;
  assign y9356 = ~1'b0 ;
  assign y9357 = n25195 ;
  assign y9358 = n25196 ;
  assign y9359 = ~n25198 ;
  assign y9360 = ~1'b0 ;
  assign y9361 = n25199 ;
  assign y9362 = ~1'b0 ;
  assign y9363 = n25205 ;
  assign y9364 = n25207 ;
  assign y9365 = ~n25208 ;
  assign y9366 = ~n25209 ;
  assign y9367 = ~1'b0 ;
  assign y9368 = ~n25212 ;
  assign y9369 = ~1'b0 ;
  assign y9370 = ~n25214 ;
  assign y9371 = ~n25226 ;
  assign y9372 = n25232 ;
  assign y9373 = ~n25234 ;
  assign y9374 = n25235 ;
  assign y9375 = n25236 ;
  assign y9376 = n25237 ;
  assign y9377 = ~n25241 ;
  assign y9378 = ~1'b0 ;
  assign y9379 = ~n25244 ;
  assign y9380 = n25245 ;
  assign y9381 = n25247 ;
  assign y9382 = n25248 ;
  assign y9383 = n25256 ;
  assign y9384 = n25262 ;
  assign y9385 = ~1'b0 ;
  assign y9386 = ~n25264 ;
  assign y9387 = n25265 ;
  assign y9388 = n25266 ;
  assign y9389 = ~1'b0 ;
  assign y9390 = n25268 ;
  assign y9391 = ~n25276 ;
  assign y9392 = n25278 ;
  assign y9393 = ~n25282 ;
  assign y9394 = ~n25284 ;
  assign y9395 = ~1'b0 ;
  assign y9396 = ~1'b0 ;
  assign y9397 = n25285 ;
  assign y9398 = n25287 ;
  assign y9399 = ~n5755 ;
  assign y9400 = ~n25289 ;
  assign y9401 = ~n25298 ;
  assign y9402 = ~1'b0 ;
  assign y9403 = ~n25300 ;
  assign y9404 = ~n25307 ;
  assign y9405 = n25311 ;
  assign y9406 = ~1'b0 ;
  assign y9407 = n8476 ;
  assign y9408 = ~1'b0 ;
  assign y9409 = ~n25317 ;
  assign y9410 = n25320 ;
  assign y9411 = n25321 ;
  assign y9412 = n25322 ;
  assign y9413 = ~n25331 ;
  assign y9414 = ~1'b0 ;
  assign y9415 = 1'b0 ;
  assign y9416 = n25332 ;
  assign y9417 = ~n25336 ;
  assign y9418 = ~n25343 ;
  assign y9419 = ~n25347 ;
  assign y9420 = n25358 ;
  assign y9421 = n5211 ;
  assign y9422 = n25360 ;
  assign y9423 = n25366 ;
  assign y9424 = n25371 ;
  assign y9425 = ~n25374 ;
  assign y9426 = ~n25378 ;
  assign y9427 = ~n4968 ;
  assign y9428 = ~n25382 ;
  assign y9429 = ~1'b0 ;
  assign y9430 = ~n25386 ;
  assign y9431 = ~n21508 ;
  assign y9432 = ~n5715 ;
  assign y9433 = n25388 ;
  assign y9434 = n25390 ;
  assign y9435 = n25391 ;
  assign y9436 = ~n658 ;
  assign y9437 = ~n25393 ;
  assign y9438 = n25398 ;
  assign y9439 = ~1'b0 ;
  assign y9440 = ~1'b0 ;
  assign y9441 = n14943 ;
  assign y9442 = n25399 ;
  assign y9443 = ~n25405 ;
  assign y9444 = n25411 ;
  assign y9445 = n21736 ;
  assign y9446 = n25412 ;
  assign y9447 = ~1'b0 ;
  assign y9448 = ~n25414 ;
  assign y9449 = n25416 ;
  assign y9450 = ~n25417 ;
  assign y9451 = n25424 ;
  assign y9452 = ~1'b0 ;
  assign y9453 = ~n25428 ;
  assign y9454 = n25432 ;
  assign y9455 = n21761 ;
  assign y9456 = ~1'b0 ;
  assign y9457 = n25440 ;
  assign y9458 = ~n25445 ;
  assign y9459 = ~1'b0 ;
  assign y9460 = ~1'b0 ;
  assign y9461 = ~1'b0 ;
  assign y9462 = n25448 ;
  assign y9463 = ~n25449 ;
  assign y9464 = n25453 ;
  assign y9465 = n25455 ;
  assign y9466 = ~n25458 ;
  assign y9467 = ~1'b0 ;
  assign y9468 = ~n25462 ;
  assign y9469 = n25463 ;
  assign y9470 = ~n25469 ;
  assign y9471 = n25471 ;
  assign y9472 = n25478 ;
  assign y9473 = ~1'b0 ;
  assign y9474 = n25479 ;
  assign y9475 = ~n25480 ;
  assign y9476 = ~n17372 ;
  assign y9477 = n25482 ;
  assign y9478 = ~1'b0 ;
  assign y9479 = n25488 ;
  assign y9480 = ~1'b0 ;
  assign y9481 = ~1'b0 ;
  assign y9482 = n25492 ;
  assign y9483 = ~n2192 ;
  assign y9484 = n25493 ;
  assign y9485 = ~n25494 ;
  assign y9486 = ~1'b0 ;
  assign y9487 = n25495 ;
  assign y9488 = ~n25499 ;
  assign y9489 = n25500 ;
  assign y9490 = n25501 ;
  assign y9491 = n25503 ;
  assign y9492 = ~n25504 ;
  assign y9493 = ~n25505 ;
  assign y9494 = ~n25507 ;
  assign y9495 = n25509 ;
  assign y9496 = ~1'b0 ;
  assign y9497 = n25514 ;
  assign y9498 = ~1'b0 ;
  assign y9499 = n25516 ;
  assign y9500 = ~n25522 ;
  assign y9501 = ~n25523 ;
  assign y9502 = ~n25525 ;
  assign y9503 = ~n25527 ;
  assign y9504 = ~n25536 ;
  assign y9505 = ~1'b0 ;
  assign y9506 = ~n25539 ;
  assign y9507 = n25540 ;
  assign y9508 = n25541 ;
  assign y9509 = ~n8658 ;
  assign y9510 = ~1'b0 ;
  assign y9511 = ~n25542 ;
  assign y9512 = ~1'b0 ;
  assign y9513 = ~1'b0 ;
  assign y9514 = ~n25544 ;
  assign y9515 = n25548 ;
  assign y9516 = n25550 ;
  assign y9517 = n25557 ;
  assign y9518 = ~1'b0 ;
  assign y9519 = ~n25560 ;
  assign y9520 = n25561 ;
  assign y9521 = ~1'b0 ;
  assign y9522 = ~n25566 ;
  assign y9523 = ~n25568 ;
  assign y9524 = ~n25571 ;
  assign y9525 = ~1'b0 ;
  assign y9526 = ~n25574 ;
  assign y9527 = ~1'b0 ;
  assign y9528 = ~1'b0 ;
  assign y9529 = ~n25575 ;
  assign y9530 = n25576 ;
  assign y9531 = ~1'b0 ;
  assign y9532 = ~n25578 ;
  assign y9533 = ~n25581 ;
  assign y9534 = ~n25589 ;
  assign y9535 = n25590 ;
  assign y9536 = ~1'b0 ;
  assign y9537 = ~1'b0 ;
  assign y9538 = ~n25591 ;
  assign y9539 = n25600 ;
  assign y9540 = ~n25601 ;
  assign y9541 = n25603 ;
  assign y9542 = ~n25606 ;
  assign y9543 = ~n25607 ;
  assign y9544 = ~n25611 ;
  assign y9545 = ~n25614 ;
  assign y9546 = n25616 ;
  assign y9547 = ~1'b0 ;
  assign y9548 = n25622 ;
  assign y9549 = ~n25623 ;
  assign y9550 = ~n15813 ;
  assign y9551 = ~n25629 ;
  assign y9552 = ~n25633 ;
  assign y9553 = n25638 ;
  assign y9554 = ~1'b0 ;
  assign y9555 = n25642 ;
  assign y9556 = n25643 ;
  assign y9557 = ~n25658 ;
  assign y9558 = n25661 ;
  assign y9559 = n25667 ;
  assign y9560 = n25669 ;
  assign y9561 = n25675 ;
  assign y9562 = n25679 ;
  assign y9563 = n25686 ;
  assign y9564 = ~n25692 ;
  assign y9565 = ~1'b0 ;
  assign y9566 = ~1'b0 ;
  assign y9567 = n25695 ;
  assign y9568 = n25706 ;
  assign y9569 = n25708 ;
  assign y9570 = n25709 ;
  assign y9571 = ~n25712 ;
  assign y9572 = ~n25713 ;
  assign y9573 = ~n25714 ;
  assign y9574 = ~n25716 ;
  assign y9575 = ~n25720 ;
  assign y9576 = ~n25722 ;
  assign y9577 = ~n25723 ;
  assign y9578 = ~1'b0 ;
  assign y9579 = ~1'b0 ;
  assign y9580 = ~n25724 ;
  assign y9581 = ~n25727 ;
  assign y9582 = ~n25733 ;
  assign y9583 = 1'b0 ;
  assign y9584 = n25734 ;
  assign y9585 = ~n25741 ;
  assign y9586 = 1'b0 ;
  assign y9587 = ~1'b0 ;
  assign y9588 = n25743 ;
  assign y9589 = n25744 ;
  assign y9590 = n25749 ;
  assign y9591 = ~1'b0 ;
  assign y9592 = ~1'b0 ;
  assign y9593 = n25750 ;
  assign y9594 = ~1'b0 ;
  assign y9595 = ~n25754 ;
  assign y9596 = ~n25757 ;
  assign y9597 = n25767 ;
  assign y9598 = n25770 ;
  assign y9599 = n25774 ;
  assign y9600 = n25775 ;
  assign y9601 = ~n25778 ;
  assign y9602 = ~1'b0 ;
  assign y9603 = ~1'b0 ;
  assign y9604 = ~n25780 ;
  assign y9605 = n25785 ;
  assign y9606 = ~n25792 ;
  assign y9607 = ~n25795 ;
  assign y9608 = ~n25797 ;
  assign y9609 = n25800 ;
  assign y9610 = n25801 ;
  assign y9611 = n25807 ;
  assign y9612 = ~n25811 ;
  assign y9613 = n25816 ;
  assign y9614 = ~n25820 ;
  assign y9615 = ~1'b0 ;
  assign y9616 = n25826 ;
  assign y9617 = n25827 ;
  assign y9618 = n25835 ;
  assign y9619 = n25836 ;
  assign y9620 = ~1'b0 ;
  assign y9621 = ~n25840 ;
  assign y9622 = ~n25843 ;
  assign y9623 = ~n25847 ;
  assign y9624 = n25858 ;
  assign y9625 = n25860 ;
  assign y9626 = ~n25861 ;
  assign y9627 = ~n25862 ;
  assign y9628 = ~n25865 ;
  assign y9629 = n25869 ;
  assign y9630 = ~1'b0 ;
  assign y9631 = ~1'b0 ;
  assign y9632 = n25876 ;
  assign y9633 = n25878 ;
  assign y9634 = ~n25882 ;
  assign y9635 = n25885 ;
  assign y9636 = n25887 ;
  assign y9637 = n25888 ;
  assign y9638 = ~n25896 ;
  assign y9639 = ~n25900 ;
  assign y9640 = n25902 ;
  assign y9641 = ~n25905 ;
  assign y9642 = n25919 ;
  assign y9643 = ~n25921 ;
  assign y9644 = ~n25922 ;
  assign y9645 = ~n25923 ;
  assign y9646 = ~n25926 ;
  assign y9647 = n25936 ;
  assign y9648 = ~n25939 ;
  assign y9649 = ~1'b0 ;
  assign y9650 = ~1'b0 ;
  assign y9651 = n6274 ;
  assign y9652 = n25944 ;
  assign y9653 = ~n18017 ;
  assign y9654 = ~n25946 ;
  assign y9655 = n2146 ;
  assign y9656 = ~n25948 ;
  assign y9657 = ~n25949 ;
  assign y9658 = ~1'b0 ;
  assign y9659 = ~n25951 ;
  assign y9660 = ~1'b0 ;
  assign y9661 = n25955 ;
  assign y9662 = ~n25956 ;
  assign y9663 = ~n25957 ;
  assign y9664 = ~1'b0 ;
  assign y9665 = ~1'b0 ;
  assign y9666 = ~n25962 ;
  assign y9667 = ~n25963 ;
  assign y9668 = n25965 ;
  assign y9669 = ~1'b0 ;
  assign y9670 = ~n25967 ;
  assign y9671 = ~n25975 ;
  assign y9672 = n25976 ;
  assign y9673 = n9594 ;
  assign y9674 = n25979 ;
  assign y9675 = 1'b0 ;
  assign y9676 = ~n25981 ;
  assign y9677 = ~n25983 ;
  assign y9678 = ~n25984 ;
  assign y9679 = n25989 ;
  assign y9680 = n25990 ;
  assign y9681 = ~n25994 ;
  assign y9682 = ~n26000 ;
  assign y9683 = n26005 ;
  assign y9684 = ~n26007 ;
  assign y9685 = ~n26010 ;
  assign y9686 = ~n26014 ;
  assign y9687 = ~1'b0 ;
  assign y9688 = ~1'b0 ;
  assign y9689 = ~1'b0 ;
  assign y9690 = n26015 ;
  assign y9691 = ~n26016 ;
  assign y9692 = ~n26019 ;
  assign y9693 = ~n26023 ;
  assign y9694 = ~n26026 ;
  assign y9695 = n3521 ;
  assign y9696 = ~n26027 ;
  assign y9697 = n26028 ;
  assign y9698 = n26029 ;
  assign y9699 = ~n26033 ;
  assign y9700 = n26036 ;
  assign y9701 = ~1'b0 ;
  assign y9702 = ~n26037 ;
  assign y9703 = ~n26038 ;
  assign y9704 = n26040 ;
  assign y9705 = n26041 ;
  assign y9706 = ~1'b0 ;
  assign y9707 = n26044 ;
  assign y9708 = n26046 ;
  assign y9709 = ~n26051 ;
  assign y9710 = n26052 ;
  assign y9711 = ~n26053 ;
  assign y9712 = ~1'b0 ;
  assign y9713 = ~n26057 ;
  assign y9714 = ~1'b0 ;
  assign y9715 = n26058 ;
  assign y9716 = n26059 ;
  assign y9717 = ~1'b0 ;
  assign y9718 = ~n26061 ;
  assign y9719 = n26062 ;
  assign y9720 = ~1'b0 ;
  assign y9721 = n26064 ;
  assign y9722 = ~1'b0 ;
  assign y9723 = n19728 ;
  assign y9724 = ~1'b0 ;
  assign y9725 = n26068 ;
  assign y9726 = n26069 ;
  assign y9727 = ~n26074 ;
  assign y9728 = ~n26076 ;
  assign y9729 = n26081 ;
  assign y9730 = n26088 ;
  assign y9731 = ~n26091 ;
  assign y9732 = ~n26098 ;
  assign y9733 = ~n26100 ;
  assign y9734 = ~n26106 ;
  assign y9735 = n26109 ;
  assign y9736 = ~n26110 ;
  assign y9737 = n26112 ;
  assign y9738 = ~n26113 ;
  assign y9739 = n26118 ;
  assign y9740 = n26121 ;
  assign y9741 = n26122 ;
  assign y9742 = ~n24143 ;
  assign y9743 = ~n26124 ;
  assign y9744 = n26126 ;
  assign y9745 = ~n26130 ;
  assign y9746 = ~1'b0 ;
  assign y9747 = n26139 ;
  assign y9748 = ~1'b0 ;
  assign y9749 = ~n26140 ;
  assign y9750 = ~1'b0 ;
  assign y9751 = ~1'b0 ;
  assign y9752 = ~n26145 ;
  assign y9753 = n26148 ;
  assign y9754 = ~1'b0 ;
  assign y9755 = ~1'b0 ;
  assign y9756 = n26155 ;
  assign y9757 = ~n26163 ;
  assign y9758 = ~1'b0 ;
  assign y9759 = n26166 ;
  assign y9760 = ~1'b0 ;
  assign y9761 = ~n26168 ;
  assign y9762 = n26169 ;
  assign y9763 = n26170 ;
  assign y9764 = n26174 ;
  assign y9765 = ~n26179 ;
  assign y9766 = n26180 ;
  assign y9767 = ~n26184 ;
  assign y9768 = ~n26187 ;
  assign y9769 = ~n26188 ;
  assign y9770 = ~n26195 ;
  assign y9771 = ~n26197 ;
  assign y9772 = ~n26199 ;
  assign y9773 = n26202 ;
  assign y9774 = ~n26203 ;
  assign y9775 = n26204 ;
  assign y9776 = ~1'b0 ;
  assign y9777 = n26212 ;
  assign y9778 = n26214 ;
  assign y9779 = n26217 ;
  assign y9780 = n26221 ;
  assign y9781 = ~n26223 ;
  assign y9782 = ~n26224 ;
  assign y9783 = ~n26226 ;
  assign y9784 = ~n26229 ;
  assign y9785 = n6287 ;
  assign y9786 = n26230 ;
  assign y9787 = ~1'b0 ;
  assign y9788 = n26237 ;
  assign y9789 = n26239 ;
  assign y9790 = n26242 ;
  assign y9791 = n26243 ;
  assign y9792 = n26246 ;
  assign y9793 = n26247 ;
  assign y9794 = n26257 ;
  assign y9795 = n26258 ;
  assign y9796 = n26260 ;
  assign y9797 = n26264 ;
  assign y9798 = ~n26265 ;
  assign y9799 = ~1'b0 ;
  assign y9800 = ~1'b0 ;
  assign y9801 = ~n4411 ;
  assign y9802 = ~n26267 ;
  assign y9803 = n26272 ;
  assign y9804 = n26275 ;
  assign y9805 = n26277 ;
  assign y9806 = n26279 ;
  assign y9807 = ~1'b0 ;
  assign y9808 = ~1'b0 ;
  assign y9809 = ~n26283 ;
  assign y9810 = ~1'b0 ;
  assign y9811 = n26286 ;
  assign y9812 = ~n26290 ;
  assign y9813 = n26291 ;
  assign y9814 = ~n26300 ;
  assign y9815 = n26302 ;
  assign y9816 = n26308 ;
  assign y9817 = ~n26314 ;
  assign y9818 = ~n26320 ;
  assign y9819 = n26323 ;
  assign y9820 = n26324 ;
  assign y9821 = ~n26327 ;
  assign y9822 = ~n26332 ;
  assign y9823 = n26335 ;
  assign y9824 = n26337 ;
  assign y9825 = ~1'b0 ;
  assign y9826 = n26338 ;
  assign y9827 = n26339 ;
  assign y9828 = n26341 ;
  assign y9829 = ~n26342 ;
  assign y9830 = ~1'b0 ;
  assign y9831 = ~1'b0 ;
  assign y9832 = ~n26345 ;
  assign y9833 = 1'b0 ;
  assign y9834 = n26350 ;
  assign y9835 = ~n26355 ;
  assign y9836 = ~1'b0 ;
  assign y9837 = ~n26360 ;
  assign y9838 = n26361 ;
  assign y9839 = n26363 ;
  assign y9840 = n26367 ;
  assign y9841 = n26375 ;
  assign y9842 = n26377 ;
  assign y9843 = ~n26378 ;
  assign y9844 = ~1'b0 ;
  assign y9845 = ~1'b0 ;
  assign y9846 = n26380 ;
  assign y9847 = ~1'b0 ;
  assign y9848 = ~1'b0 ;
  assign y9849 = ~n26385 ;
  assign y9850 = ~1'b0 ;
  assign y9851 = ~1'b0 ;
  assign y9852 = n26387 ;
  assign y9853 = n2614 ;
  assign y9854 = ~n26390 ;
  assign y9855 = ~n26392 ;
  assign y9856 = ~1'b0 ;
  assign y9857 = ~n26394 ;
  assign y9858 = n26396 ;
  assign y9859 = ~n26397 ;
  assign y9860 = ~n26401 ;
  assign y9861 = n26402 ;
  assign y9862 = ~n26405 ;
  assign y9863 = ~n26406 ;
  assign y9864 = ~1'b0 ;
  assign y9865 = n26409 ;
  assign y9866 = n26411 ;
  assign y9867 = ~n26417 ;
  assign y9868 = ~n26419 ;
  assign y9869 = ~n26421 ;
  assign y9870 = ~n26423 ;
  assign y9871 = ~n26425 ;
  assign y9872 = ~n26427 ;
  assign y9873 = n26428 ;
  assign y9874 = n26429 ;
  assign y9875 = n26430 ;
  assign y9876 = ~n26432 ;
  assign y9877 = ~n26433 ;
  assign y9878 = n26434 ;
  assign y9879 = ~n26440 ;
  assign y9880 = n26443 ;
  assign y9881 = n26448 ;
  assign y9882 = n26451 ;
  assign y9883 = n26453 ;
  assign y9884 = ~n26455 ;
  assign y9885 = ~n26460 ;
  assign y9886 = ~n20963 ;
  assign y9887 = n26462 ;
  assign y9888 = ~1'b0 ;
  assign y9889 = n3605 ;
  assign y9890 = ~1'b0 ;
  assign y9891 = ~n26465 ;
  assign y9892 = n26466 ;
  assign y9893 = ~n26468 ;
  assign y9894 = n26469 ;
  assign y9895 = ~n25522 ;
  assign y9896 = n26471 ;
  assign y9897 = ~1'b0 ;
  assign y9898 = n26475 ;
  assign y9899 = n26476 ;
  assign y9900 = n26478 ;
  assign y9901 = ~1'b0 ;
  assign y9902 = ~n26482 ;
  assign y9903 = ~n26485 ;
  assign y9904 = ~n26487 ;
  assign y9905 = ~n26489 ;
  assign y9906 = ~n26491 ;
  assign y9907 = ~n26493 ;
  assign y9908 = ~n26494 ;
  assign y9909 = n26501 ;
  assign y9910 = n26505 ;
  assign y9911 = n26507 ;
  assign y9912 = ~n26513 ;
  assign y9913 = ~n26514 ;
  assign y9914 = n26523 ;
  assign y9915 = n26524 ;
  assign y9916 = ~n26526 ;
  assign y9917 = 1'b0 ;
  assign y9918 = n26528 ;
  assign y9919 = ~1'b0 ;
  assign y9920 = n26529 ;
  assign y9921 = ~n26535 ;
  assign y9922 = n26537 ;
  assign y9923 = n26538 ;
  assign y9924 = ~1'b0 ;
  assign y9925 = n26542 ;
  assign y9926 = ~n26544 ;
  assign y9927 = n26552 ;
  assign y9928 = ~n26559 ;
  assign y9929 = ~n26562 ;
  assign y9930 = ~n26564 ;
  assign y9931 = ~1'b0 ;
  assign y9932 = n26565 ;
  assign y9933 = n26573 ;
  assign y9934 = n26575 ;
  assign y9935 = ~n26580 ;
  assign y9936 = ~n26585 ;
  assign y9937 = ~n26596 ;
  assign y9938 = ~n26598 ;
  assign y9939 = ~n26600 ;
  assign y9940 = n26601 ;
  assign y9941 = n26605 ;
  assign y9942 = ~n26615 ;
  assign y9943 = ~1'b0 ;
  assign y9944 = n26617 ;
  assign y9945 = ~n26620 ;
  assign y9946 = n26622 ;
  assign y9947 = ~1'b0 ;
  assign y9948 = ~n26623 ;
  assign y9949 = ~n26629 ;
  assign y9950 = ~1'b0 ;
  assign y9951 = ~n26632 ;
  assign y9952 = n26633 ;
  assign y9953 = n26634 ;
  assign y9954 = ~n26645 ;
  assign y9955 = ~1'b0 ;
  assign y9956 = n26647 ;
  assign y9957 = ~n26649 ;
  assign y9958 = ~n26650 ;
  assign y9959 = ~n26659 ;
  assign y9960 = ~n11711 ;
  assign y9961 = ~1'b0 ;
  assign y9962 = ~n26663 ;
  assign y9963 = n26667 ;
  assign y9964 = n26669 ;
  assign y9965 = n26670 ;
  assign y9966 = ~1'b0 ;
  assign y9967 = ~1'b0 ;
  assign y9968 = ~n26671 ;
  assign y9969 = ~n26673 ;
  assign y9970 = n26676 ;
  assign y9971 = ~n5377 ;
  assign y9972 = n26678 ;
  assign y9973 = n26679 ;
  assign y9974 = ~1'b0 ;
  assign y9975 = n26681 ;
  assign y9976 = ~n26682 ;
  assign y9977 = n26684 ;
  assign y9978 = n26685 ;
  assign y9979 = ~n26688 ;
  assign y9980 = ~n26690 ;
  assign y9981 = ~n26699 ;
  assign y9982 = n26701 ;
  assign y9983 = n26702 ;
  assign y9984 = ~1'b0 ;
  assign y9985 = ~1'b0 ;
  assign y9986 = n26704 ;
  assign y9987 = ~n26709 ;
  assign y9988 = ~n26715 ;
  assign y9989 = ~1'b0 ;
  assign y9990 = n26716 ;
  assign y9991 = ~n26728 ;
  assign y9992 = ~n26734 ;
  assign y9993 = ~n26737 ;
  assign y9994 = n26738 ;
  assign y9995 = ~n26739 ;
  assign y9996 = n26742 ;
  assign y9997 = ~n26744 ;
  assign y9998 = ~1'b0 ;
  assign y9999 = ~n26746 ;
  assign y10000 = n13251 ;
  assign y10001 = ~1'b0 ;
  assign y10002 = n26747 ;
  assign y10003 = n26748 ;
  assign y10004 = ~1'b0 ;
  assign y10005 = ~n26751 ;
  assign y10006 = n26753 ;
  assign y10007 = ~1'b0 ;
  assign y10008 = ~1'b0 ;
  assign y10009 = ~n26754 ;
  assign y10010 = ~n26757 ;
  assign y10011 = n26763 ;
  assign y10012 = ~n26767 ;
  assign y10013 = n26768 ;
  assign y10014 = ~n26774 ;
  assign y10015 = ~n26778 ;
  assign y10016 = ~n26781 ;
  assign y10017 = ~1'b0 ;
  assign y10018 = n26785 ;
  assign y10019 = ~1'b0 ;
  assign y10020 = n20159 ;
  assign y10021 = ~n26787 ;
  assign y10022 = ~n17471 ;
  assign y10023 = n26788 ;
  assign y10024 = ~n26789 ;
  assign y10025 = ~n26794 ;
  assign y10026 = ~n26796 ;
  assign y10027 = ~n26802 ;
  assign y10028 = n26803 ;
  assign y10029 = 1'b0 ;
  assign y10030 = ~n26804 ;
  assign y10031 = ~n26814 ;
  assign y10032 = ~n26816 ;
  assign y10033 = ~n26818 ;
  assign y10034 = n26820 ;
  assign y10035 = ~n26822 ;
  assign y10036 = n26835 ;
  assign y10037 = ~n26845 ;
  assign y10038 = n26850 ;
  assign y10039 = ~n26852 ;
  assign y10040 = ~1'b0 ;
  assign y10041 = ~n26854 ;
  assign y10042 = n26855 ;
  assign y10043 = n26860 ;
  assign y10044 = n26864 ;
  assign y10045 = n26868 ;
  assign y10046 = n26869 ;
  assign y10047 = ~n26870 ;
  assign y10048 = ~1'b0 ;
  assign y10049 = ~n26874 ;
  assign y10050 = ~1'b0 ;
  assign y10051 = ~1'b0 ;
  assign y10052 = n26879 ;
  assign y10053 = ~n26880 ;
  assign y10054 = ~n26883 ;
  assign y10055 = n26884 ;
  assign y10056 = ~n26891 ;
  assign y10057 = ~1'b0 ;
  assign y10058 = ~n26894 ;
  assign y10059 = n26896 ;
  assign y10060 = n26897 ;
  assign y10061 = n26898 ;
  assign y10062 = n26905 ;
  assign y10063 = ~n26908 ;
  assign y10064 = ~1'b0 ;
  assign y10065 = n23400 ;
  assign y10066 = n26914 ;
  assign y10067 = ~n26917 ;
  assign y10068 = ~n26919 ;
  assign y10069 = n26922 ;
  assign y10070 = n26923 ;
  assign y10071 = ~n26924 ;
  assign y10072 = n26926 ;
  assign y10073 = ~1'b0 ;
  assign y10074 = ~n26927 ;
  assign y10075 = n26928 ;
  assign y10076 = ~n26932 ;
  assign y10077 = ~1'b0 ;
  assign y10078 = ~n26935 ;
  assign y10079 = ~n26938 ;
  assign y10080 = ~n26940 ;
  assign y10081 = n26945 ;
  assign y10082 = ~n26950 ;
  assign y10083 = ~n26956 ;
  assign y10084 = ~1'b0 ;
  assign y10085 = n26959 ;
  assign y10086 = n26962 ;
  assign y10087 = ~n26964 ;
  assign y10088 = n26968 ;
  assign y10089 = n26970 ;
  assign y10090 = n26971 ;
  assign y10091 = ~n26975 ;
  assign y10092 = ~1'b0 ;
  assign y10093 = n26977 ;
  assign y10094 = ~1'b0 ;
  assign y10095 = ~n26978 ;
  assign y10096 = n26981 ;
  assign y10097 = ~n26985 ;
  assign y10098 = ~n26988 ;
  assign y10099 = n26989 ;
  assign y10100 = ~1'b0 ;
  assign y10101 = ~n26990 ;
  assign y10102 = ~n26998 ;
  assign y10103 = ~1'b0 ;
  assign y10104 = ~n27000 ;
  assign y10105 = ~1'b0 ;
  assign y10106 = ~n27002 ;
  assign y10107 = ~n27006 ;
  assign y10108 = ~n27009 ;
  assign y10109 = ~n27012 ;
  assign y10110 = n27019 ;
  assign y10111 = ~n27022 ;
  assign y10112 = n27023 ;
  assign y10113 = ~n9897 ;
  assign y10114 = ~1'b0 ;
  assign y10115 = ~1'b0 ;
  assign y10116 = ~n27028 ;
  assign y10117 = ~n27031 ;
  assign y10118 = n27036 ;
  assign y10119 = n27037 ;
  assign y10120 = ~1'b0 ;
  assign y10121 = n27039 ;
  assign y10122 = ~n27042 ;
  assign y10123 = n27045 ;
  assign y10124 = n27048 ;
  assign y10125 = n27051 ;
  assign y10126 = ~n27053 ;
  assign y10127 = ~n27055 ;
  assign y10128 = ~n27056 ;
  assign y10129 = ~n27061 ;
  assign y10130 = ~n27066 ;
  assign y10131 = ~n27069 ;
  assign y10132 = ~n27071 ;
  assign y10133 = ~n27075 ;
  assign y10134 = ~1'b0 ;
  assign y10135 = n27077 ;
  assign y10136 = n27080 ;
  assign y10137 = ~n27081 ;
  assign y10138 = n27086 ;
  assign y10139 = n27090 ;
  assign y10140 = ~n27091 ;
  assign y10141 = n27093 ;
  assign y10142 = ~n27104 ;
  assign y10143 = n27106 ;
  assign y10144 = n27109 ;
  assign y10145 = ~1'b0 ;
  assign y10146 = n27113 ;
  assign y10147 = ~n27118 ;
  assign y10148 = ~n27124 ;
  assign y10149 = ~n27126 ;
  assign y10150 = ~n27127 ;
  assign y10151 = ~n27132 ;
  assign y10152 = ~1'b0 ;
  assign y10153 = ~n27133 ;
  assign y10154 = n27134 ;
  assign y10155 = ~n27136 ;
  assign y10156 = ~1'b0 ;
  assign y10157 = ~n27137 ;
  assign y10158 = ~n27140 ;
  assign y10159 = ~n27142 ;
  assign y10160 = ~n27143 ;
  assign y10161 = ~1'b0 ;
  assign y10162 = n27145 ;
  assign y10163 = ~n27148 ;
  assign y10164 = ~n9986 ;
  assign y10165 = ~1'b0 ;
  assign y10166 = ~1'b0 ;
  assign y10167 = ~1'b0 ;
  assign y10168 = n27150 ;
  assign y10169 = n27154 ;
  assign y10170 = ~n27155 ;
  assign y10171 = ~n27159 ;
  assign y10172 = n27162 ;
  assign y10173 = ~1'b0 ;
  assign y10174 = n27163 ;
  assign y10175 = n27164 ;
  assign y10176 = n27167 ;
  assign y10177 = n27171 ;
  assign y10178 = ~n27172 ;
  assign y10179 = n27175 ;
  assign y10180 = ~n27181 ;
  assign y10181 = ~n27186 ;
  assign y10182 = ~n27195 ;
  assign y10183 = ~1'b0 ;
  assign y10184 = ~1'b0 ;
  assign y10185 = n27197 ;
  assign y10186 = ~n27202 ;
  assign y10187 = ~n27203 ;
  assign y10188 = ~1'b0 ;
  assign y10189 = ~n27204 ;
  assign y10190 = ~1'b0 ;
  assign y10191 = ~1'b0 ;
  assign y10192 = ~n27208 ;
  assign y10193 = ~1'b0 ;
  assign y10194 = ~n27212 ;
  assign y10195 = ~n4052 ;
  assign y10196 = ~1'b0 ;
  assign y10197 = ~1'b0 ;
  assign y10198 = ~1'b0 ;
  assign y10199 = ~n27213 ;
  assign y10200 = n27220 ;
  assign y10201 = ~n27228 ;
  assign y10202 = ~1'b0 ;
  assign y10203 = ~1'b0 ;
  assign y10204 = ~n27232 ;
  assign y10205 = ~n27235 ;
  assign y10206 = n27236 ;
  assign y10207 = n27237 ;
  assign y10208 = ~1'b0 ;
  assign y10209 = ~1'b0 ;
  assign y10210 = ~1'b0 ;
  assign y10211 = n27238 ;
  assign y10212 = n27241 ;
  assign y10213 = n27243 ;
  assign y10214 = n27245 ;
  assign y10215 = n3690 ;
  assign y10216 = ~n27250 ;
  assign y10217 = ~n27252 ;
  assign y10218 = n27253 ;
  assign y10219 = n27254 ;
  assign y10220 = ~n27257 ;
  assign y10221 = ~n27259 ;
  assign y10222 = n27262 ;
  assign y10223 = ~n27265 ;
  assign y10224 = ~1'b0 ;
  assign y10225 = ~n27267 ;
  assign y10226 = ~1'b0 ;
  assign y10227 = ~n27268 ;
  assign y10228 = ~n27271 ;
  assign y10229 = n27273 ;
  assign y10230 = n27275 ;
  assign y10231 = ~n27276 ;
  assign y10232 = ~n27285 ;
  assign y10233 = ~n27287 ;
  assign y10234 = ~n27288 ;
  assign y10235 = n27293 ;
  assign y10236 = n27301 ;
  assign y10237 = n27306 ;
  assign y10238 = ~1'b0 ;
  assign y10239 = n15528 ;
  assign y10240 = ~1'b0 ;
  assign y10241 = ~n27309 ;
  assign y10242 = ~1'b0 ;
  assign y10243 = n21864 ;
  assign y10244 = ~1'b0 ;
  assign y10245 = ~n27313 ;
  assign y10246 = ~n13250 ;
  assign y10247 = ~1'b0 ;
  assign y10248 = n27317 ;
  assign y10249 = ~1'b0 ;
  assign y10250 = ~n27323 ;
  assign y10251 = ~n27324 ;
  assign y10252 = ~1'b0 ;
  assign y10253 = n27329 ;
  assign y10254 = ~1'b0 ;
  assign y10255 = ~n27334 ;
  assign y10256 = n27337 ;
  assign y10257 = n27339 ;
  assign y10258 = ~n27343 ;
  assign y10259 = ~n27345 ;
  assign y10260 = ~1'b0 ;
  assign y10261 = ~n27348 ;
  assign y10262 = n27350 ;
  assign y10263 = n4679 ;
  assign y10264 = ~n27353 ;
  assign y10265 = ~1'b0 ;
  assign y10266 = n27354 ;
  assign y10267 = ~n27357 ;
  assign y10268 = n27358 ;
  assign y10269 = n27365 ;
  assign y10270 = n27366 ;
  assign y10271 = n27367 ;
  assign y10272 = ~n27369 ;
  assign y10273 = ~n27382 ;
  assign y10274 = n27389 ;
  assign y10275 = ~n27392 ;
  assign y10276 = ~n27395 ;
  assign y10277 = n27398 ;
  assign y10278 = ~n27401 ;
  assign y10279 = ~n27407 ;
  assign y10280 = n27409 ;
  assign y10281 = ~n27413 ;
  assign y10282 = n27421 ;
  assign y10283 = ~n27424 ;
  assign y10284 = n27430 ;
  assign y10285 = n27432 ;
  assign y10286 = ~n27436 ;
  assign y10287 = ~n27438 ;
  assign y10288 = ~n27440 ;
  assign y10289 = ~n27442 ;
  assign y10290 = ~n21980 ;
  assign y10291 = ~1'b0 ;
  assign y10292 = ~1'b0 ;
  assign y10293 = n27443 ;
  assign y10294 = ~1'b0 ;
  assign y10295 = n27444 ;
  assign y10296 = ~1'b0 ;
  assign y10297 = n27445 ;
  assign y10298 = ~n27451 ;
  assign y10299 = n27454 ;
  assign y10300 = n27456 ;
  assign y10301 = ~1'b0 ;
  assign y10302 = ~n27457 ;
  assign y10303 = ~n27460 ;
  assign y10304 = n27469 ;
  assign y10305 = ~n27472 ;
  assign y10306 = ~n27477 ;
  assign y10307 = ~n27478 ;
  assign y10308 = ~n27481 ;
  assign y10309 = ~n27482 ;
  assign y10310 = n27486 ;
  assign y10311 = ~1'b0 ;
  assign y10312 = n27487 ;
  assign y10313 = ~1'b0 ;
  assign y10314 = ~1'b0 ;
  assign y10315 = n27492 ;
  assign y10316 = n27494 ;
  assign y10317 = n27496 ;
  assign y10318 = n13828 ;
  assign y10319 = ~n27497 ;
  assign y10320 = n27498 ;
  assign y10321 = ~1'b0 ;
  assign y10322 = ~1'b0 ;
  assign y10323 = n27500 ;
  assign y10324 = n27503 ;
  assign y10325 = n27506 ;
  assign y10326 = n27510 ;
  assign y10327 = ~n27512 ;
  assign y10328 = n27516 ;
  assign y10329 = n27519 ;
  assign y10330 = n27521 ;
  assign y10331 = n27528 ;
  assign y10332 = n27534 ;
  assign y10333 = n27539 ;
  assign y10334 = ~n27542 ;
  assign y10335 = ~n4356 ;
  assign y10336 = n27546 ;
  assign y10337 = ~n27548 ;
  assign y10338 = ~n27550 ;
  assign y10339 = ~n27556 ;
  assign y10340 = n27559 ;
  assign y10341 = n27564 ;
  assign y10342 = ~n27569 ;
  assign y10343 = ~n27571 ;
  assign y10344 = ~n27575 ;
  assign y10345 = n27576 ;
  assign y10346 = ~1'b0 ;
  assign y10347 = n27578 ;
  assign y10348 = n27580 ;
  assign y10349 = n27583 ;
  assign y10350 = n27584 ;
  assign y10351 = n27589 ;
  assign y10352 = ~1'b0 ;
  assign y10353 = n27590 ;
  assign y10354 = ~n27591 ;
  assign y10355 = n27592 ;
  assign y10356 = ~1'b0 ;
  assign y10357 = ~1'b0 ;
  assign y10358 = ~1'b0 ;
  assign y10359 = ~n27599 ;
  assign y10360 = n789 ;
  assign y10361 = ~n27601 ;
  assign y10362 = n27606 ;
  assign y10363 = n27608 ;
  assign y10364 = ~1'b0 ;
  assign y10365 = ~n27616 ;
  assign y10366 = n27618 ;
  assign y10367 = n27621 ;
  assign y10368 = n27622 ;
  assign y10369 = ~n1769 ;
  assign y10370 = n27625 ;
  assign y10371 = ~1'b0 ;
  assign y10372 = n27630 ;
  assign y10373 = ~n27634 ;
  assign y10374 = n27638 ;
  assign y10375 = ~n27640 ;
  assign y10376 = n21026 ;
  assign y10377 = ~1'b0 ;
  assign y10378 = n27641 ;
  assign y10379 = n2874 ;
  assign y10380 = ~n27642 ;
  assign y10381 = ~1'b0 ;
  assign y10382 = n27643 ;
  assign y10383 = ~n27648 ;
  assign y10384 = ~n27650 ;
  assign y10385 = n27655 ;
  assign y10386 = n27658 ;
  assign y10387 = n19775 ;
  assign y10388 = ~1'b0 ;
  assign y10389 = n27661 ;
  assign y10390 = ~n27662 ;
  assign y10391 = ~n27673 ;
  assign y10392 = ~n27675 ;
  assign y10393 = ~n27676 ;
  assign y10394 = ~n27678 ;
  assign y10395 = ~1'b0 ;
  assign y10396 = n27680 ;
  assign y10397 = ~n27683 ;
  assign y10398 = n27688 ;
  assign y10399 = ~n27692 ;
  assign y10400 = n27696 ;
  assign y10401 = ~n27699 ;
  assign y10402 = ~n27701 ;
  assign y10403 = ~1'b0 ;
  assign y10404 = ~1'b0 ;
  assign y10405 = ~n27703 ;
  assign y10406 = n27704 ;
  assign y10407 = ~n27710 ;
  assign y10408 = ~1'b0 ;
  assign y10409 = n27711 ;
  assign y10410 = n27712 ;
  assign y10411 = ~1'b0 ;
  assign y10412 = ~n27714 ;
  assign y10413 = n27715 ;
  assign y10414 = ~n27717 ;
  assign y10415 = n27719 ;
  assign y10416 = ~n27721 ;
  assign y10417 = n8552 ;
  assign y10418 = ~n27728 ;
  assign y10419 = ~n27731 ;
  assign y10420 = n27738 ;
  assign y10421 = ~n27741 ;
  assign y10422 = n27742 ;
  assign y10423 = ~n27743 ;
  assign y10424 = ~n27748 ;
  assign y10425 = ~n3604 ;
  assign y10426 = ~n27752 ;
  assign y10427 = 1'b0 ;
  assign y10428 = n27754 ;
  assign y10429 = ~1'b0 ;
  assign y10430 = n27756 ;
  assign y10431 = ~n27759 ;
  assign y10432 = ~n27763 ;
  assign y10433 = ~n27765 ;
  assign y10434 = n27768 ;
  assign y10435 = ~n27773 ;
  assign y10436 = n27776 ;
  assign y10437 = ~n27777 ;
  assign y10438 = ~1'b0 ;
  assign y10439 = ~1'b0 ;
  assign y10440 = ~1'b0 ;
  assign y10441 = ~n27779 ;
  assign y10442 = ~n27781 ;
  assign y10443 = n27782 ;
  assign y10444 = n27785 ;
  assign y10445 = ~1'b0 ;
  assign y10446 = n27788 ;
  assign y10447 = n27791 ;
  assign y10448 = n27794 ;
  assign y10449 = ~n27803 ;
  assign y10450 = ~n27807 ;
  assign y10451 = n27811 ;
  assign y10452 = ~n27813 ;
  assign y10453 = n27819 ;
  assign y10454 = ~1'b0 ;
  assign y10455 = n27824 ;
  assign y10456 = ~n27826 ;
  assign y10457 = ~1'b0 ;
  assign y10458 = ~1'b0 ;
  assign y10459 = n27830 ;
  assign y10460 = n27833 ;
  assign y10461 = n27837 ;
  assign y10462 = n27840 ;
  assign y10463 = ~1'b0 ;
  assign y10464 = ~n27843 ;
  assign y10465 = ~1'b0 ;
  assign y10466 = n27844 ;
  assign y10467 = ~n27845 ;
  assign y10468 = ~n27849 ;
  assign y10469 = ~n27850 ;
  assign y10470 = ~n27854 ;
  assign y10471 = ~n27856 ;
  assign y10472 = ~n27858 ;
  assign y10473 = ~1'b0 ;
  assign y10474 = n27862 ;
  assign y10475 = n27863 ;
  assign y10476 = ~n27864 ;
  assign y10477 = ~1'b0 ;
  assign y10478 = n27869 ;
  assign y10479 = ~1'b0 ;
  assign y10480 = n27870 ;
  assign y10481 = n27873 ;
  assign y10482 = ~1'b0 ;
  assign y10483 = ~n27874 ;
  assign y10484 = ~1'b0 ;
  assign y10485 = ~n27876 ;
  assign y10486 = n27877 ;
  assign y10487 = n27881 ;
  assign y10488 = ~n27882 ;
  assign y10489 = ~1'b0 ;
  assign y10490 = n27884 ;
  assign y10491 = n27889 ;
  assign y10492 = n27896 ;
  assign y10493 = ~n27897 ;
  assign y10494 = ~1'b0 ;
  assign y10495 = n27899 ;
  assign y10496 = ~1'b0 ;
  assign y10497 = ~1'b0 ;
  assign y10498 = ~n27900 ;
  assign y10499 = ~n27901 ;
  assign y10500 = n27904 ;
  assign y10501 = n20429 ;
  assign y10502 = ~n27909 ;
  assign y10503 = ~n27914 ;
  assign y10504 = ~n27915 ;
  assign y10505 = n27918 ;
  assign y10506 = ~n27920 ;
  assign y10507 = ~1'b0 ;
  assign y10508 = ~1'b0 ;
  assign y10509 = n27924 ;
  assign y10510 = ~1'b0 ;
  assign y10511 = n27925 ;
  assign y10512 = ~1'b0 ;
  assign y10513 = ~n27929 ;
  assign y10514 = n8170 ;
  assign y10515 = ~1'b0 ;
  assign y10516 = n27931 ;
  assign y10517 = ~1'b0 ;
  assign y10518 = n27934 ;
  assign y10519 = ~n27944 ;
  assign y10520 = ~n27945 ;
  assign y10521 = n27947 ;
  assign y10522 = ~1'b0 ;
  assign y10523 = n27949 ;
  assign y10524 = ~1'b0 ;
  assign y10525 = n27952 ;
  assign y10526 = n27955 ;
  assign y10527 = n27956 ;
  assign y10528 = ~n27958 ;
  assign y10529 = ~n27959 ;
  assign y10530 = ~n25959 ;
  assign y10531 = n27966 ;
  assign y10532 = ~1'b0 ;
  assign y10533 = n27970 ;
  assign y10534 = n27979 ;
  assign y10535 = ~n27981 ;
  assign y10536 = n27982 ;
  assign y10537 = n27985 ;
  assign y10538 = ~n27988 ;
  assign y10539 = ~1'b0 ;
  assign y10540 = n27989 ;
  assign y10541 = ~n28001 ;
  assign y10542 = ~n28003 ;
  assign y10543 = ~1'b0 ;
  assign y10544 = ~n28004 ;
  assign y10545 = ~n28005 ;
  assign y10546 = ~1'b0 ;
  assign y10547 = ~n28008 ;
  assign y10548 = ~n28011 ;
  assign y10549 = n28013 ;
  assign y10550 = ~n28014 ;
  assign y10551 = ~n28015 ;
  assign y10552 = ~n28016 ;
  assign y10553 = ~1'b0 ;
  assign y10554 = ~n28030 ;
  assign y10555 = ~n28032 ;
  assign y10556 = ~n28034 ;
  assign y10557 = ~n28036 ;
  assign y10558 = n28040 ;
  assign y10559 = ~n28042 ;
  assign y10560 = n28047 ;
  assign y10561 = n28048 ;
  assign y10562 = n28052 ;
  assign y10563 = ~1'b0 ;
  assign y10564 = n28055 ;
  assign y10565 = ~n28057 ;
  assign y10566 = n28059 ;
  assign y10567 = ~n28060 ;
  assign y10568 = ~n28065 ;
  assign y10569 = n28067 ;
  assign y10570 = n28068 ;
  assign y10571 = n28072 ;
  assign y10572 = ~n28074 ;
  assign y10573 = ~n28080 ;
  assign y10574 = ~n28081 ;
  assign y10575 = n28087 ;
  assign y10576 = n28088 ;
  assign y10577 = ~n28091 ;
  assign y10578 = n28093 ;
  assign y10579 = n28094 ;
  assign y10580 = n28101 ;
  assign y10581 = ~1'b0 ;
  assign y10582 = n28103 ;
  assign y10583 = ~n28106 ;
  assign y10584 = n28108 ;
  assign y10585 = n28109 ;
  assign y10586 = n28111 ;
  assign y10587 = ~n28112 ;
  assign y10588 = n19943 ;
  assign y10589 = n28114 ;
  assign y10590 = ~n28115 ;
  assign y10591 = ~1'b0 ;
  assign y10592 = n28119 ;
  assign y10593 = ~n28123 ;
  assign y10594 = ~1'b0 ;
  assign y10595 = ~n28126 ;
  assign y10596 = ~n28134 ;
  assign y10597 = ~n28138 ;
  assign y10598 = ~1'b0 ;
  assign y10599 = n28141 ;
  assign y10600 = ~n28142 ;
  assign y10601 = 1'b0 ;
  assign y10602 = ~n28149 ;
  assign y10603 = n28150 ;
  assign y10604 = ~1'b0 ;
  assign y10605 = ~n28152 ;
  assign y10606 = n28158 ;
  assign y10607 = ~1'b0 ;
  assign y10608 = ~n28160 ;
  assign y10609 = n28161 ;
  assign y10610 = ~n28162 ;
  assign y10611 = ~n28163 ;
  assign y10612 = n28165 ;
  assign y10613 = ~n28169 ;
  assign y10614 = ~n28171 ;
  assign y10615 = ~n28173 ;
  assign y10616 = ~x71 ;
  assign y10617 = ~n28175 ;
  assign y10618 = ~n28176 ;
  assign y10619 = ~n28177 ;
  assign y10620 = ~1'b0 ;
  assign y10621 = 1'b0 ;
  assign y10622 = n28183 ;
  assign y10623 = ~n28193 ;
  assign y10624 = ~n28197 ;
  assign y10625 = n28199 ;
  assign y10626 = ~n28204 ;
  assign y10627 = ~n28205 ;
  assign y10628 = ~1'b0 ;
  assign y10629 = n28207 ;
  assign y10630 = ~1'b0 ;
  assign y10631 = n28212 ;
  assign y10632 = n28215 ;
  assign y10633 = n28221 ;
  assign y10634 = ~n28226 ;
  assign y10635 = n28228 ;
  assign y10636 = n28231 ;
  assign y10637 = n28232 ;
  assign y10638 = n28234 ;
  assign y10639 = ~1'b0 ;
  assign y10640 = ~n28238 ;
  assign y10641 = n28242 ;
  assign y10642 = ~n28251 ;
  assign y10643 = n28252 ;
  assign y10644 = ~n28257 ;
  assign y10645 = ~1'b0 ;
  assign y10646 = ~n28260 ;
  assign y10647 = ~n28266 ;
  assign y10648 = n28267 ;
  assign y10649 = ~1'b0 ;
  assign y10650 = ~n28268 ;
  assign y10651 = n28271 ;
  assign y10652 = ~1'b0 ;
  assign y10653 = ~n28272 ;
  assign y10654 = n28275 ;
  assign y10655 = ~n28284 ;
  assign y10656 = ~n28285 ;
  assign y10657 = ~n28289 ;
  assign y10658 = n28291 ;
  assign y10659 = ~n28297 ;
  assign y10660 = ~n28299 ;
  assign y10661 = ~n28301 ;
  assign y10662 = n25618 ;
  assign y10663 = ~n28302 ;
  assign y10664 = ~1'b0 ;
  assign y10665 = n28306 ;
  assign y10666 = n28310 ;
  assign y10667 = n28312 ;
  assign y10668 = n28315 ;
  assign y10669 = n28316 ;
  assign y10670 = n28318 ;
  assign y10671 = n28319 ;
  assign y10672 = ~n28323 ;
  assign y10673 = ~1'b0 ;
  assign y10674 = ~n28326 ;
  assign y10675 = ~1'b0 ;
  assign y10676 = ~n28327 ;
  assign y10677 = ~1'b0 ;
  assign y10678 = ~n28329 ;
  assign y10679 = ~n28334 ;
  assign y10680 = ~n28335 ;
  assign y10681 = n28336 ;
  assign y10682 = ~n28338 ;
  assign y10683 = ~n28339 ;
  assign y10684 = n28340 ;
  assign y10685 = n28341 ;
  assign y10686 = ~1'b0 ;
  assign y10687 = n28346 ;
  assign y10688 = ~n28347 ;
  assign y10689 = ~n28349 ;
  assign y10690 = n28350 ;
  assign y10691 = ~1'b0 ;
  assign y10692 = n28354 ;
  assign y10693 = ~1'b0 ;
  assign y10694 = ~1'b0 ;
  assign y10695 = n28360 ;
  assign y10696 = n6305 ;
  assign y10697 = 1'b0 ;
  assign y10698 = ~n28366 ;
  assign y10699 = ~n28369 ;
  assign y10700 = ~n28373 ;
  assign y10701 = ~n28376 ;
  assign y10702 = ~n28378 ;
  assign y10703 = n28380 ;
  assign y10704 = n28382 ;
  assign y10705 = ~1'b0 ;
  assign y10706 = ~1'b0 ;
  assign y10707 = ~n28387 ;
  assign y10708 = n28388 ;
  assign y10709 = x167 ;
  assign y10710 = n28391 ;
  assign y10711 = n28392 ;
  assign y10712 = ~n28398 ;
  assign y10713 = ~n28400 ;
  assign y10714 = ~n28405 ;
  assign y10715 = ~1'b0 ;
  assign y10716 = ~n28407 ;
  assign y10717 = n28408 ;
  assign y10718 = n28410 ;
  assign y10719 = ~1'b0 ;
  assign y10720 = ~1'b0 ;
  assign y10721 = n28411 ;
  assign y10722 = ~n28414 ;
  assign y10723 = n28415 ;
  assign y10724 = n28417 ;
  assign y10725 = ~n28418 ;
  assign y10726 = ~1'b0 ;
  assign y10727 = ~n28419 ;
  assign y10728 = n28421 ;
  assign y10729 = ~1'b0 ;
  assign y10730 = ~n28425 ;
  assign y10731 = ~n28428 ;
  assign y10732 = ~1'b0 ;
  assign y10733 = n28430 ;
  assign y10734 = ~n28431 ;
  assign y10735 = ~n28434 ;
  assign y10736 = n28435 ;
  assign y10737 = ~1'b0 ;
  assign y10738 = n28439 ;
  assign y10739 = n14398 ;
  assign y10740 = ~n28441 ;
  assign y10741 = ~n28442 ;
  assign y10742 = ~1'b0 ;
  assign y10743 = ~n28444 ;
  assign y10744 = n15733 ;
  assign y10745 = ~n2727 ;
  assign y10746 = ~n28445 ;
  assign y10747 = n28447 ;
  assign y10748 = n28449 ;
  assign y10749 = n28451 ;
  assign y10750 = ~n28454 ;
  assign y10751 = ~n28455 ;
  assign y10752 = n28460 ;
  assign y10753 = ~n28463 ;
  assign y10754 = ~1'b0 ;
  assign y10755 = ~n28465 ;
  assign y10756 = ~n28466 ;
  assign y10757 = ~n28467 ;
  assign y10758 = n28468 ;
  assign y10759 = ~n28472 ;
  assign y10760 = ~1'b0 ;
  assign y10761 = n28474 ;
  assign y10762 = ~n28475 ;
  assign y10763 = n28478 ;
  assign y10764 = ~n28479 ;
  assign y10765 = ~1'b0 ;
  assign y10766 = n28480 ;
  assign y10767 = ~1'b0 ;
  assign y10768 = n23952 ;
  assign y10769 = n28482 ;
  assign y10770 = n28485 ;
  assign y10771 = ~n28489 ;
  assign y10772 = n27367 ;
  assign y10773 = ~1'b0 ;
  assign y10774 = n28491 ;
  assign y10775 = ~n28492 ;
  assign y10776 = n28495 ;
  assign y10777 = ~n28503 ;
  assign y10778 = ~n28506 ;
  assign y10779 = ~n28509 ;
  assign y10780 = ~n28513 ;
  assign y10781 = ~n28516 ;
  assign y10782 = n28523 ;
  assign y10783 = n28524 ;
  assign y10784 = ~1'b0 ;
  assign y10785 = ~n24638 ;
  assign y10786 = n28529 ;
  assign y10787 = ~1'b0 ;
  assign y10788 = n28534 ;
  assign y10789 = n24219 ;
  assign y10790 = ~n28537 ;
  assign y10791 = n4397 ;
  assign y10792 = ~n28540 ;
  assign y10793 = n28545 ;
  assign y10794 = ~n28547 ;
  assign y10795 = ~n28548 ;
  assign y10796 = n28553 ;
  assign y10797 = ~n28554 ;
  assign y10798 = n28560 ;
  assign y10799 = ~n28566 ;
  assign y10800 = ~n20929 ;
  assign y10801 = n28568 ;
  assign y10802 = n28572 ;
  assign y10803 = ~1'b0 ;
  assign y10804 = ~n28578 ;
  assign y10805 = n28579 ;
  assign y10806 = ~n28585 ;
  assign y10807 = n5097 ;
  assign y10808 = n28587 ;
  assign y10809 = n6606 ;
  assign y10810 = ~n28588 ;
  assign y10811 = n28589 ;
  assign y10812 = ~n28590 ;
  assign y10813 = ~1'b0 ;
  assign y10814 = ~n28597 ;
  assign y10815 = ~n28598 ;
  assign y10816 = n28601 ;
  assign y10817 = ~n28605 ;
  assign y10818 = ~n28615 ;
  assign y10819 = ~1'b0 ;
  assign y10820 = n28618 ;
  assign y10821 = ~n28620 ;
  assign y10822 = ~n28621 ;
  assign y10823 = ~1'b0 ;
  assign y10824 = ~n28624 ;
  assign y10825 = ~1'b0 ;
  assign y10826 = n28626 ;
  assign y10827 = ~n28630 ;
  assign y10828 = ~1'b0 ;
  assign y10829 = ~1'b0 ;
  assign y10830 = ~n28634 ;
  assign y10831 = ~n28636 ;
  assign y10832 = n28640 ;
  assign y10833 = ~n28641 ;
  assign y10834 = n28645 ;
  assign y10835 = ~1'b0 ;
  assign y10836 = ~n28648 ;
  assign y10837 = ~1'b0 ;
  assign y10838 = ~n28652 ;
  assign y10839 = n28654 ;
  assign y10840 = ~n28656 ;
  assign y10841 = n28662 ;
  assign y10842 = 1'b0 ;
  assign y10843 = ~n28666 ;
  assign y10844 = n28669 ;
  assign y10845 = n28670 ;
  assign y10846 = n28672 ;
  assign y10847 = ~n15951 ;
  assign y10848 = ~n28679 ;
  assign y10849 = n28684 ;
  assign y10850 = ~n28694 ;
  assign y10851 = ~n28703 ;
  assign y10852 = ~1'b0 ;
  assign y10853 = ~n28706 ;
  assign y10854 = n28707 ;
  assign y10855 = ~n28715 ;
  assign y10856 = n28716 ;
  assign y10857 = ~n28721 ;
  assign y10858 = ~1'b0 ;
  assign y10859 = n20691 ;
  assign y10860 = ~1'b0 ;
  assign y10861 = ~1'b0 ;
  assign y10862 = ~1'b0 ;
  assign y10863 = ~n28723 ;
  assign y10864 = n28725 ;
  assign y10865 = n9560 ;
  assign y10866 = n28730 ;
  assign y10867 = n28732 ;
  assign y10868 = n28739 ;
  assign y10869 = ~n28741 ;
  assign y10870 = n28742 ;
  assign y10871 = n28743 ;
  assign y10872 = ~n28745 ;
  assign y10873 = n28748 ;
  assign y10874 = ~n28749 ;
  assign y10875 = ~n28751 ;
  assign y10876 = n28755 ;
  assign y10877 = n28757 ;
  assign y10878 = n28758 ;
  assign y10879 = n28759 ;
  assign y10880 = n28760 ;
  assign y10881 = ~n28770 ;
  assign y10882 = ~n28771 ;
  assign y10883 = ~1'b0 ;
  assign y10884 = ~n11509 ;
  assign y10885 = ~n28773 ;
  assign y10886 = ~1'b0 ;
  assign y10887 = ~n28774 ;
  assign y10888 = ~n28775 ;
  assign y10889 = ~1'b0 ;
  assign y10890 = n28778 ;
  assign y10891 = 1'b0 ;
  assign y10892 = ~n28782 ;
  assign y10893 = ~1'b0 ;
  assign y10894 = n28783 ;
  assign y10895 = ~n28785 ;
  assign y10896 = ~n28787 ;
  assign y10897 = n28790 ;
  assign y10898 = n28796 ;
  assign y10899 = ~1'b0 ;
  assign y10900 = ~n28798 ;
  assign y10901 = n28799 ;
  assign y10902 = n28805 ;
  assign y10903 = ~1'b0 ;
  assign y10904 = ~n28807 ;
  assign y10905 = ~1'b0 ;
  assign y10906 = n28808 ;
  assign y10907 = n28815 ;
  assign y10908 = ~1'b0 ;
  assign y10909 = ~1'b0 ;
  assign y10910 = ~1'b0 ;
  assign y10911 = ~1'b0 ;
  assign y10912 = ~n28817 ;
  assign y10913 = ~n28818 ;
  assign y10914 = ~n28822 ;
  assign y10915 = ~1'b0 ;
  assign y10916 = n28826 ;
  assign y10917 = ~n28829 ;
  assign y10918 = ~n28830 ;
  assign y10919 = ~n28832 ;
  assign y10920 = ~n28833 ;
  assign y10921 = n28835 ;
  assign y10922 = ~n28838 ;
  assign y10923 = n28839 ;
  assign y10924 = ~1'b0 ;
  assign y10925 = ~n28842 ;
  assign y10926 = n28844 ;
  assign y10927 = n28848 ;
  assign y10928 = ~1'b0 ;
  assign y10929 = n28849 ;
  assign y10930 = n28850 ;
  assign y10931 = ~n28852 ;
  assign y10932 = ~n28854 ;
  assign y10933 = ~1'b0 ;
  assign y10934 = ~n28859 ;
  assign y10935 = ~n13303 ;
  assign y10936 = n28860 ;
  assign y10937 = n28863 ;
  assign y10938 = ~n28867 ;
  assign y10939 = ~1'b0 ;
  assign y10940 = n28868 ;
  assign y10941 = ~n28869 ;
  assign y10942 = n28871 ;
  assign y10943 = n28877 ;
  assign y10944 = n28883 ;
  assign y10945 = ~1'b0 ;
  assign y10946 = ~1'b0 ;
  assign y10947 = ~n28885 ;
  assign y10948 = ~1'b0 ;
  assign y10949 = ~n28890 ;
  assign y10950 = ~n28891 ;
  assign y10951 = ~n28893 ;
  assign y10952 = ~n28895 ;
  assign y10953 = ~1'b0 ;
  assign y10954 = ~1'b0 ;
  assign y10955 = ~1'b0 ;
  assign y10956 = ~n28900 ;
  assign y10957 = n28909 ;
  assign y10958 = ~1'b0 ;
  assign y10959 = ~n28916 ;
  assign y10960 = n28920 ;
  assign y10961 = n28921 ;
  assign y10962 = n28924 ;
  assign y10963 = ~1'b0 ;
  assign y10964 = ~n28932 ;
  assign y10965 = n28933 ;
  assign y10966 = ~n28934 ;
  assign y10967 = ~n28936 ;
  assign y10968 = ~1'b0 ;
  assign y10969 = n28938 ;
  assign y10970 = ~n28943 ;
  assign y10971 = n28945 ;
  assign y10972 = ~n28946 ;
  assign y10973 = n28949 ;
  assign y10974 = ~n28950 ;
  assign y10975 = n28952 ;
  assign y10976 = n28953 ;
  assign y10977 = ~n28958 ;
  assign y10978 = ~n28960 ;
  assign y10979 = n28961 ;
  assign y10980 = n28962 ;
  assign y10981 = ~n28964 ;
  assign y10982 = n28971 ;
  assign y10983 = ~n28973 ;
  assign y10984 = ~n20015 ;
  assign y10985 = ~1'b0 ;
  assign y10986 = ~n28975 ;
  assign y10987 = n28976 ;
  assign y10988 = ~n28978 ;
  assign y10989 = n28980 ;
  assign y10990 = n28981 ;
  assign y10991 = n28984 ;
  assign y10992 = ~1'b0 ;
  assign y10993 = n28986 ;
  assign y10994 = n28990 ;
  assign y10995 = ~n28991 ;
  assign y10996 = ~n15888 ;
  assign y10997 = ~n28992 ;
  assign y10998 = ~1'b0 ;
  assign y10999 = ~n28994 ;
  assign y11000 = n29004 ;
  assign y11001 = n29005 ;
  assign y11002 = n29006 ;
  assign y11003 = ~n29009 ;
  assign y11004 = ~n29010 ;
  assign y11005 = n29013 ;
  assign y11006 = ~1'b0 ;
  assign y11007 = ~n29021 ;
  assign y11008 = ~n29024 ;
  assign y11009 = ~n29028 ;
  assign y11010 = ~n29030 ;
  assign y11011 = ~1'b0 ;
  assign y11012 = ~1'b0 ;
  assign y11013 = ~1'b0 ;
  assign y11014 = n29031 ;
  assign y11015 = ~n29032 ;
  assign y11016 = n29035 ;
  assign y11017 = ~n29039 ;
  assign y11018 = ~n29041 ;
  assign y11019 = ~n29044 ;
  assign y11020 = ~n29050 ;
  assign y11021 = n29054 ;
  assign y11022 = ~1'b0 ;
  assign y11023 = ~n29058 ;
  assign y11024 = ~n29064 ;
  assign y11025 = n29066 ;
  assign y11026 = ~1'b0 ;
  assign y11027 = ~n1084 ;
  assign y11028 = ~n29073 ;
  assign y11029 = n29074 ;
  assign y11030 = ~n29075 ;
  assign y11031 = n29081 ;
  assign y11032 = ~1'b0 ;
  assign y11033 = n29083 ;
  assign y11034 = n29085 ;
  assign y11035 = n29090 ;
  assign y11036 = ~n29094 ;
  assign y11037 = ~n29096 ;
  assign y11038 = n29104 ;
  assign y11039 = ~n29114 ;
  assign y11040 = n29116 ;
  assign y11041 = ~1'b0 ;
  assign y11042 = n29117 ;
  assign y11043 = ~n29122 ;
  assign y11044 = ~n29128 ;
  assign y11045 = ~n29131 ;
  assign y11046 = ~n29138 ;
  assign y11047 = ~1'b0 ;
  assign y11048 = ~n29139 ;
  assign y11049 = ~n29143 ;
  assign y11050 = ~n29147 ;
  assign y11051 = ~n29149 ;
  assign y11052 = ~n29152 ;
  assign y11053 = ~n29155 ;
  assign y11054 = ~n29162 ;
  assign y11055 = ~n29164 ;
  assign y11056 = n29165 ;
  assign y11057 = n29170 ;
  assign y11058 = n29173 ;
  assign y11059 = ~1'b0 ;
  assign y11060 = ~1'b0 ;
  assign y11061 = ~n29178 ;
  assign y11062 = n29179 ;
  assign y11063 = n29180 ;
  assign y11064 = n22941 ;
  assign y11065 = ~n29182 ;
  assign y11066 = ~n29185 ;
  assign y11067 = n6054 ;
  assign y11068 = n29187 ;
  assign y11069 = n29191 ;
  assign y11070 = ~1'b0 ;
  assign y11071 = n29198 ;
  assign y11072 = n29201 ;
  assign y11073 = n29202 ;
  assign y11074 = ~n13009 ;
  assign y11075 = ~n29203 ;
  assign y11076 = n29207 ;
  assign y11077 = n29214 ;
  assign y11078 = ~n29216 ;
  assign y11079 = n29218 ;
  assign y11080 = ~n29220 ;
  assign y11081 = ~1'b0 ;
  assign y11082 = ~1'b0 ;
  assign y11083 = ~n29222 ;
  assign y11084 = ~n29223 ;
  assign y11085 = ~n29226 ;
  assign y11086 = ~1'b0 ;
  assign y11087 = ~n29232 ;
  assign y11088 = ~n29234 ;
  assign y11089 = n29235 ;
  assign y11090 = n29236 ;
  assign y11091 = ~n29238 ;
  assign y11092 = ~1'b0 ;
  assign y11093 = n29242 ;
  assign y11094 = ~1'b0 ;
  assign y11095 = n29245 ;
  assign y11096 = n17422 ;
  assign y11097 = ~n29249 ;
  assign y11098 = ~n29250 ;
  assign y11099 = ~n29251 ;
  assign y11100 = ~n29252 ;
  assign y11101 = ~n29254 ;
  assign y11102 = ~1'b0 ;
  assign y11103 = ~n29258 ;
  assign y11104 = ~n29263 ;
  assign y11105 = n29276 ;
  assign y11106 = ~n29281 ;
  assign y11107 = n29282 ;
  assign y11108 = n29283 ;
  assign y11109 = ~1'b0 ;
  assign y11110 = ~n29284 ;
  assign y11111 = ~n29285 ;
  assign y11112 = ~1'b0 ;
  assign y11113 = 1'b0 ;
  assign y11114 = ~1'b0 ;
  assign y11115 = ~n29287 ;
  assign y11116 = ~n29289 ;
  assign y11117 = n29290 ;
  assign y11118 = ~n29296 ;
  assign y11119 = ~1'b0 ;
  assign y11120 = n29297 ;
  assign y11121 = ~n29304 ;
  assign y11122 = ~n29305 ;
  assign y11123 = ~n29306 ;
  assign y11124 = n29309 ;
  assign y11125 = ~1'b0 ;
  assign y11126 = ~n29311 ;
  assign y11127 = n29317 ;
  assign y11128 = ~n29324 ;
  assign y11129 = n29326 ;
  assign y11130 = n29330 ;
  assign y11131 = ~n29333 ;
  assign y11132 = ~1'b0 ;
  assign y11133 = n29336 ;
  assign y11134 = ~n29341 ;
  assign y11135 = ~n29342 ;
  assign y11136 = ~n29343 ;
  assign y11137 = ~n29345 ;
  assign y11138 = ~n29350 ;
  assign y11139 = n29355 ;
  assign y11140 = ~n29357 ;
  assign y11141 = ~n29358 ;
  assign y11142 = n29360 ;
  assign y11143 = ~n29361 ;
  assign y11144 = n29363 ;
  assign y11145 = ~n29364 ;
  assign y11146 = n29365 ;
  assign y11147 = n29366 ;
  assign y11148 = n29367 ;
  assign y11149 = n29369 ;
  assign y11150 = n29371 ;
  assign y11151 = n29375 ;
  assign y11152 = n29376 ;
  assign y11153 = n29378 ;
  assign y11154 = ~1'b0 ;
  assign y11155 = n29381 ;
  assign y11156 = ~n29384 ;
  assign y11157 = ~n29385 ;
  assign y11158 = n29387 ;
  assign y11159 = ~n29390 ;
  assign y11160 = ~n29393 ;
  assign y11161 = n29395 ;
  assign y11162 = ~1'b0 ;
  assign y11163 = ~1'b0 ;
  assign y11164 = n29396 ;
  assign y11165 = ~1'b0 ;
  assign y11166 = ~n29400 ;
  assign y11167 = n29405 ;
  assign y11168 = ~n29406 ;
  assign y11169 = n29411 ;
  assign y11170 = n29414 ;
  assign y11171 = n29415 ;
  assign y11172 = ~n29416 ;
  assign y11173 = ~n29417 ;
  assign y11174 = n29418 ;
  assign y11175 = ~n29014 ;
  assign y11176 = n14578 ;
  assign y11177 = n29419 ;
  assign y11178 = ~1'b0 ;
  assign y11179 = ~1'b0 ;
  assign y11180 = ~n29423 ;
  assign y11181 = n29429 ;
  assign y11182 = n29434 ;
  assign y11183 = ~n29436 ;
  assign y11184 = ~1'b0 ;
  assign y11185 = n29438 ;
  assign y11186 = 1'b0 ;
  assign y11187 = ~n29445 ;
  assign y11188 = n29446 ;
  assign y11189 = ~n16244 ;
  assign y11190 = ~1'b0 ;
  assign y11191 = ~1'b0 ;
  assign y11192 = n29447 ;
  assign y11193 = n29448 ;
  assign y11194 = ~n29450 ;
  assign y11195 = 1'b0 ;
  assign y11196 = ~1'b0 ;
  assign y11197 = ~n29451 ;
  assign y11198 = ~1'b0 ;
  assign y11199 = n29455 ;
  assign y11200 = n29458 ;
  assign y11201 = n29460 ;
  assign y11202 = n29467 ;
  assign y11203 = ~1'b0 ;
  assign y11204 = n29472 ;
  assign y11205 = ~1'b0 ;
  assign y11206 = n29475 ;
  assign y11207 = ~1'b0 ;
  assign y11208 = n29477 ;
  assign y11209 = ~1'b0 ;
  assign y11210 = ~n29482 ;
  assign y11211 = ~1'b0 ;
  assign y11212 = ~1'b0 ;
  assign y11213 = n29493 ;
  assign y11214 = ~n29494 ;
  assign y11215 = ~n29495 ;
  assign y11216 = ~n29496 ;
  assign y11217 = n29497 ;
  assign y11218 = ~1'b0 ;
  assign y11219 = n15996 ;
  assign y11220 = ~1'b0 ;
  assign y11221 = ~1'b0 ;
  assign y11222 = n29499 ;
  assign y11223 = n29500 ;
  assign y11224 = ~1'b0 ;
  assign y11225 = ~n12061 ;
  assign y11226 = n29503 ;
  assign y11227 = n29504 ;
  assign y11228 = ~n29505 ;
  assign y11229 = n29508 ;
  assign y11230 = ~1'b0 ;
  assign y11231 = ~n29509 ;
  assign y11232 = ~1'b0 ;
  assign y11233 = ~1'b0 ;
  assign y11234 = ~n29511 ;
  assign y11235 = ~1'b0 ;
  assign y11236 = n29514 ;
  assign y11237 = n29516 ;
  assign y11238 = n29523 ;
  assign y11239 = ~1'b0 ;
  assign y11240 = ~n29526 ;
  assign y11241 = n29527 ;
  assign y11242 = ~1'b0 ;
  assign y11243 = n29529 ;
  assign y11244 = n29530 ;
  assign y11245 = ~n29531 ;
  assign y11246 = ~n29533 ;
  assign y11247 = ~n29538 ;
  assign y11248 = ~n29545 ;
  assign y11249 = n29552 ;
  assign y11250 = n29554 ;
  assign y11251 = n29560 ;
  assign y11252 = ~n14831 ;
  assign y11253 = ~n5367 ;
  assign y11254 = n29561 ;
  assign y11255 = ~n29564 ;
  assign y11256 = n29569 ;
  assign y11257 = ~n29571 ;
  assign y11258 = ~1'b0 ;
  assign y11259 = ~n29577 ;
  assign y11260 = n29580 ;
  assign y11261 = ~1'b0 ;
  assign y11262 = n29581 ;
  assign y11263 = ~n29583 ;
  assign y11264 = ~n29592 ;
  assign y11265 = n29596 ;
  assign y11266 = n29599 ;
  assign y11267 = n29601 ;
  assign y11268 = n29604 ;
  assign y11269 = n29607 ;
  assign y11270 = ~1'b0 ;
  assign y11271 = n29608 ;
  assign y11272 = n5144 ;
  assign y11273 = ~n29609 ;
  assign y11274 = ~n29610 ;
  assign y11275 = ~n29616 ;
  assign y11276 = n29617 ;
  assign y11277 = ~n29618 ;
  assign y11278 = ~n29621 ;
  assign y11279 = ~n29623 ;
  assign y11280 = n14275 ;
  assign y11281 = ~1'b0 ;
  assign y11282 = ~n29632 ;
  assign y11283 = ~n29634 ;
  assign y11284 = n29637 ;
  assign y11285 = ~n29639 ;
  assign y11286 = ~n29643 ;
  assign y11287 = ~n29644 ;
  assign y11288 = n29658 ;
  assign y11289 = n29667 ;
  assign y11290 = n29669 ;
  assign y11291 = n29671 ;
  assign y11292 = n29672 ;
  assign y11293 = ~1'b0 ;
  assign y11294 = n29675 ;
  assign y11295 = n29677 ;
  assign y11296 = ~n29682 ;
  assign y11297 = n29688 ;
  assign y11298 = ~n29691 ;
  assign y11299 = ~n29693 ;
  assign y11300 = ~n29696 ;
  assign y11301 = n29701 ;
  assign y11302 = ~n29702 ;
  assign y11303 = ~n29703 ;
  assign y11304 = n29709 ;
  assign y11305 = ~n29711 ;
  assign y11306 = ~n29713 ;
  assign y11307 = ~n29717 ;
  assign y11308 = ~n29718 ;
  assign y11309 = ~1'b0 ;
  assign y11310 = ~n29720 ;
  assign y11311 = ~1'b0 ;
  assign y11312 = n29728 ;
  assign y11313 = n29731 ;
  assign y11314 = n29734 ;
  assign y11315 = ~1'b0 ;
  assign y11316 = ~1'b0 ;
  assign y11317 = ~n29735 ;
  assign y11318 = n14505 ;
  assign y11319 = ~n29737 ;
  assign y11320 = ~n29740 ;
  assign y11321 = n29744 ;
  assign y11322 = ~1'b0 ;
  assign y11323 = ~n29745 ;
  assign y11324 = ~n29749 ;
  assign y11325 = ~n29751 ;
  assign y11326 = ~n29754 ;
  assign y11327 = ~n29756 ;
  assign y11328 = n29757 ;
  assign y11329 = ~n29758 ;
  assign y11330 = ~n29760 ;
  assign y11331 = ~n29765 ;
  assign y11332 = ~n29766 ;
  assign y11333 = ~1'b0 ;
  assign y11334 = ~1'b0 ;
  assign y11335 = ~n29767 ;
  assign y11336 = ~1'b0 ;
  assign y11337 = n29771 ;
  assign y11338 = n29772 ;
  assign y11339 = ~1'b0 ;
  assign y11340 = ~1'b0 ;
  assign y11341 = ~n29778 ;
  assign y11342 = n29779 ;
  assign y11343 = n29780 ;
  assign y11344 = ~n29783 ;
  assign y11345 = ~1'b0 ;
  assign y11346 = ~n29785 ;
  assign y11347 = ~1'b0 ;
  assign y11348 = ~n29786 ;
  assign y11349 = n29789 ;
  assign y11350 = ~n29791 ;
  assign y11351 = n29793 ;
  assign y11352 = ~n29800 ;
  assign y11353 = n29801 ;
  assign y11354 = ~1'b0 ;
  assign y11355 = ~1'b0 ;
  assign y11356 = ~1'b0 ;
  assign y11357 = n29806 ;
  assign y11358 = n29814 ;
  assign y11359 = ~n29818 ;
  assign y11360 = n29820 ;
  assign y11361 = ~1'b0 ;
  assign y11362 = ~1'b0 ;
  assign y11363 = n5159 ;
  assign y11364 = ~n29828 ;
  assign y11365 = ~n29829 ;
  assign y11366 = n29830 ;
  assign y11367 = n29836 ;
  assign y11368 = ~1'b0 ;
  assign y11369 = n4034 ;
  assign y11370 = ~n29842 ;
  assign y11371 = n29843 ;
  assign y11372 = ~n29845 ;
  assign y11373 = ~n29847 ;
  assign y11374 = n29851 ;
  assign y11375 = ~n29855 ;
  assign y11376 = n29857 ;
  assign y11377 = ~n29858 ;
  assign y11378 = n29859 ;
  assign y11379 = ~n29861 ;
  assign y11380 = n29866 ;
  assign y11381 = n29695 ;
  assign y11382 = n29868 ;
  assign y11383 = ~n29870 ;
  assign y11384 = ~n29871 ;
  assign y11385 = 1'b0 ;
  assign y11386 = n29874 ;
  assign y11387 = ~n29881 ;
  assign y11388 = ~n29882 ;
  assign y11389 = ~1'b0 ;
  assign y11390 = ~1'b0 ;
  assign y11391 = ~n29885 ;
  assign y11392 = ~n29887 ;
  assign y11393 = n29889 ;
  assign y11394 = ~n29890 ;
  assign y11395 = n29899 ;
  assign y11396 = n29900 ;
  assign y11397 = n29902 ;
  assign y11398 = n29903 ;
  assign y11399 = ~1'b0 ;
  assign y11400 = n29907 ;
  assign y11401 = ~n29911 ;
  assign y11402 = n29915 ;
  assign y11403 = ~n29918 ;
  assign y11404 = n29920 ;
  assign y11405 = ~1'b0 ;
  assign y11406 = ~1'b0 ;
  assign y11407 = n3074 ;
  assign y11408 = n29924 ;
  assign y11409 = ~1'b0 ;
  assign y11410 = n29927 ;
  assign y11411 = ~n29930 ;
  assign y11412 = n29932 ;
  assign y11413 = n29933 ;
  assign y11414 = ~n29934 ;
  assign y11415 = ~n29936 ;
  assign y11416 = ~n29937 ;
  assign y11417 = ~n29940 ;
  assign y11418 = n29941 ;
  assign y11419 = n29943 ;
  assign y11420 = n29944 ;
  assign y11421 = n29948 ;
  assign y11422 = n29959 ;
  assign y11423 = n29962 ;
  assign y11424 = n29966 ;
  assign y11425 = ~1'b0 ;
  assign y11426 = n29973 ;
  assign y11427 = n29974 ;
  assign y11428 = ~n29975 ;
  assign y11429 = ~n29976 ;
  assign y11430 = ~n29978 ;
  assign y11431 = ~1'b0 ;
  assign y11432 = ~n29980 ;
  assign y11433 = n8850 ;
  assign y11434 = ~n29982 ;
  assign y11435 = ~n29984 ;
  assign y11436 = ~n29997 ;
  assign y11437 = n30006 ;
  assign y11438 = ~n30007 ;
  assign y11439 = ~n30008 ;
  assign y11440 = ~n30010 ;
  assign y11441 = n30011 ;
  assign y11442 = ~n30015 ;
  assign y11443 = ~1'b0 ;
  assign y11444 = ~n30018 ;
  assign y11445 = ~n30022 ;
  assign y11446 = ~n30024 ;
  assign y11447 = n30025 ;
  assign y11448 = ~n30028 ;
  assign y11449 = n30029 ;
  assign y11450 = ~1'b0 ;
  assign y11451 = n30035 ;
  assign y11452 = ~n30042 ;
  assign y11453 = ~n30046 ;
  assign y11454 = ~n30047 ;
  assign y11455 = ~n30048 ;
  assign y11456 = ~1'b0 ;
  assign y11457 = ~1'b0 ;
  assign y11458 = ~n30050 ;
  assign y11459 = 1'b0 ;
  assign y11460 = n30052 ;
  assign y11461 = ~n30054 ;
  assign y11462 = n30059 ;
  assign y11463 = ~1'b0 ;
  assign y11464 = ~n30060 ;
  assign y11465 = 1'b0 ;
  assign y11466 = n30063 ;
  assign y11467 = ~1'b0 ;
  assign y11468 = n30069 ;
  assign y11469 = n30070 ;
  assign y11470 = ~1'b0 ;
  assign y11471 = ~1'b0 ;
  assign y11472 = ~n30073 ;
  assign y11473 = n30074 ;
  assign y11474 = ~n30076 ;
  assign y11475 = ~n30082 ;
  assign y11476 = n30084 ;
  assign y11477 = ~n30085 ;
  assign y11478 = ~n30087 ;
  assign y11479 = n30089 ;
  assign y11480 = ~n30095 ;
  assign y11481 = ~n30096 ;
  assign y11482 = n30098 ;
  assign y11483 = ~1'b0 ;
  assign y11484 = 1'b0 ;
  assign y11485 = n30099 ;
  assign y11486 = n30100 ;
  assign y11487 = n30107 ;
  assign y11488 = ~1'b0 ;
  assign y11489 = ~n30110 ;
  assign y11490 = ~n30114 ;
  assign y11491 = ~1'b0 ;
  assign y11492 = ~n30126 ;
  assign y11493 = ~n30128 ;
  assign y11494 = ~1'b0 ;
  assign y11495 = ~1'b0 ;
  assign y11496 = n30136 ;
  assign y11497 = ~n30140 ;
  assign y11498 = n30141 ;
  assign y11499 = ~n30142 ;
  assign y11500 = n30147 ;
  assign y11501 = n30148 ;
  assign y11502 = ~1'b0 ;
  assign y11503 = n1328 ;
  assign y11504 = n21875 ;
  assign y11505 = n30149 ;
  assign y11506 = n30151 ;
  assign y11507 = n30153 ;
  assign y11508 = n30163 ;
  assign y11509 = ~n30164 ;
  assign y11510 = ~n30166 ;
  assign y11511 = ~n30167 ;
  assign y11512 = ~1'b0 ;
  assign y11513 = n30168 ;
  assign y11514 = n30171 ;
  assign y11515 = ~1'b0 ;
  assign y11516 = n30173 ;
  assign y11517 = ~n30174 ;
  assign y11518 = ~n30175 ;
  assign y11519 = n30176 ;
  assign y11520 = n30177 ;
  assign y11521 = ~1'b0 ;
  assign y11522 = n30179 ;
  assign y11523 = n30187 ;
  assign y11524 = ~n30189 ;
  assign y11525 = ~n30191 ;
  assign y11526 = ~n9925 ;
  assign y11527 = ~1'b0 ;
  assign y11528 = ~n30193 ;
  assign y11529 = ~n30198 ;
  assign y11530 = ~n30203 ;
  assign y11531 = n30207 ;
  assign y11532 = ~n30209 ;
  assign y11533 = ~n30210 ;
  assign y11534 = n30215 ;
  assign y11535 = ~n30224 ;
  assign y11536 = n30225 ;
  assign y11537 = n30227 ;
  assign y11538 = ~n30233 ;
  assign y11539 = ~n19930 ;
  assign y11540 = n30235 ;
  assign y11541 = ~n30237 ;
  assign y11542 = n28143 ;
  assign y11543 = ~n30239 ;
  assign y11544 = n30241 ;
  assign y11545 = ~1'b0 ;
  assign y11546 = ~1'b0 ;
  assign y11547 = n30242 ;
  assign y11548 = n30244 ;
  assign y11549 = ~n30249 ;
  assign y11550 = n30256 ;
  assign y11551 = n30257 ;
  assign y11552 = n30258 ;
  assign y11553 = ~1'b0 ;
  assign y11554 = ~1'b0 ;
  assign y11555 = ~1'b0 ;
  assign y11556 = ~1'b0 ;
  assign y11557 = n30262 ;
  assign y11558 = n30266 ;
  assign y11559 = ~n30267 ;
  assign y11560 = ~1'b0 ;
  assign y11561 = ~n30273 ;
  assign y11562 = n30278 ;
  assign y11563 = n30283 ;
  assign y11564 = ~n30290 ;
  assign y11565 = ~n30297 ;
  assign y11566 = ~n30301 ;
  assign y11567 = ~1'b0 ;
  assign y11568 = ~1'b0 ;
  assign y11569 = ~1'b0 ;
  assign y11570 = ~n30302 ;
  assign y11571 = ~n30303 ;
  assign y11572 = n30306 ;
  assign y11573 = n30307 ;
  assign y11574 = ~n30308 ;
  assign y11575 = ~n30309 ;
  assign y11576 = ~n30312 ;
  assign y11577 = n30313 ;
  assign y11578 = ~1'b0 ;
  assign y11579 = ~1'b0 ;
  assign y11580 = ~n30314 ;
  assign y11581 = ~n30316 ;
  assign y11582 = n30318 ;
  assign y11583 = ~n8813 ;
  assign y11584 = n30319 ;
  assign y11585 = n30321 ;
  assign y11586 = n30324 ;
  assign y11587 = n30331 ;
  assign y11588 = ~n30337 ;
  assign y11589 = ~1'b0 ;
  assign y11590 = ~1'b0 ;
  assign y11591 = ~1'b0 ;
  assign y11592 = ~1'b0 ;
  assign y11593 = ~1'b0 ;
  assign y11594 = ~1'b0 ;
  assign y11595 = n30342 ;
  assign y11596 = n30344 ;
  assign y11597 = n30345 ;
  assign y11598 = n30346 ;
  assign y11599 = n30352 ;
  assign y11600 = ~n30359 ;
  assign y11601 = n30360 ;
  assign y11602 = ~n30362 ;
  assign y11603 = n30363 ;
  assign y11604 = ~1'b0 ;
  assign y11605 = n30370 ;
  assign y11606 = ~n30372 ;
  assign y11607 = ~1'b0 ;
  assign y11608 = ~n30375 ;
  assign y11609 = ~n30377 ;
  assign y11610 = n30380 ;
  assign y11611 = ~1'b0 ;
  assign y11612 = ~1'b0 ;
  assign y11613 = n30383 ;
  assign y11614 = ~n30386 ;
  assign y11615 = ~n30388 ;
  assign y11616 = ~1'b0 ;
  assign y11617 = ~n30392 ;
  assign y11618 = n30394 ;
  assign y11619 = n30395 ;
  assign y11620 = n30402 ;
  assign y11621 = n30409 ;
  assign y11622 = ~n30410 ;
  assign y11623 = n30411 ;
  assign y11624 = n30416 ;
  assign y11625 = ~n30418 ;
  assign y11626 = ~1'b0 ;
  assign y11627 = n30424 ;
  assign y11628 = n30426 ;
  assign y11629 = n30428 ;
  assign y11630 = n30430 ;
  assign y11631 = ~1'b0 ;
  assign y11632 = ~1'b0 ;
  assign y11633 = n30432 ;
  assign y11634 = ~n30433 ;
  assign y11635 = ~n30435 ;
  assign y11636 = n30437 ;
  assign y11637 = n30438 ;
  assign y11638 = ~n30441 ;
  assign y11639 = n26531 ;
  assign y11640 = n21458 ;
  assign y11641 = n30444 ;
  assign y11642 = ~n30445 ;
  assign y11643 = ~n30453 ;
  assign y11644 = ~1'b0 ;
  assign y11645 = ~1'b0 ;
  assign y11646 = n30456 ;
  assign y11647 = ~n30460 ;
  assign y11648 = n30462 ;
  assign y11649 = ~n30463 ;
  assign y11650 = ~n30466 ;
  assign y11651 = ~n30470 ;
  assign y11652 = ~n30472 ;
  assign y11653 = ~1'b0 ;
  assign y11654 = ~n30477 ;
  assign y11655 = n30478 ;
  assign y11656 = ~1'b0 ;
  assign y11657 = ~n30481 ;
  assign y11658 = n30483 ;
  assign y11659 = ~n30484 ;
  assign y11660 = ~n30487 ;
  assign y11661 = n30490 ;
  assign y11662 = n30491 ;
  assign y11663 = n30496 ;
  assign y11664 = n30500 ;
  assign y11665 = n30503 ;
  assign y11666 = ~n30505 ;
  assign y11667 = ~n30507 ;
  assign y11668 = ~1'b0 ;
  assign y11669 = ~n30510 ;
  assign y11670 = ~n30512 ;
  assign y11671 = ~1'b0 ;
  assign y11672 = ~1'b0 ;
  assign y11673 = ~n30513 ;
  assign y11674 = ~n30514 ;
  assign y11675 = ~1'b0 ;
  assign y11676 = n9518 ;
  assign y11677 = n30517 ;
  assign y11678 = ~n30521 ;
  assign y11679 = n30524 ;
  assign y11680 = ~1'b0 ;
  assign y11681 = ~1'b0 ;
  assign y11682 = ~1'b0 ;
  assign y11683 = n30526 ;
  assign y11684 = ~1'b0 ;
  assign y11685 = ~n30529 ;
  assign y11686 = n30530 ;
  assign y11687 = ~n30532 ;
  assign y11688 = ~1'b0 ;
  assign y11689 = ~1'b0 ;
  assign y11690 = ~1'b0 ;
  assign y11691 = ~n30536 ;
  assign y11692 = n30539 ;
  assign y11693 = ~n15799 ;
  assign y11694 = ~1'b0 ;
  assign y11695 = ~1'b0 ;
  assign y11696 = ~n30542 ;
  assign y11697 = ~n30543 ;
  assign y11698 = n30544 ;
  assign y11699 = n30550 ;
  assign y11700 = ~1'b0 ;
  assign y11701 = ~n30555 ;
  assign y11702 = ~1'b0 ;
  assign y11703 = n30558 ;
  assign y11704 = ~n30563 ;
  assign y11705 = n30566 ;
  assign y11706 = ~n30567 ;
  assign y11707 = ~1'b0 ;
  assign y11708 = n30569 ;
  assign y11709 = n30577 ;
  assign y11710 = ~n30579 ;
  assign y11711 = ~n30583 ;
  assign y11712 = n30584 ;
  assign y11713 = ~n30585 ;
  assign y11714 = ~1'b0 ;
  assign y11715 = ~n30589 ;
  assign y11716 = n30590 ;
  assign y11717 = ~1'b0 ;
  assign y11718 = ~n24953 ;
  assign y11719 = ~n26531 ;
  assign y11720 = n30591 ;
  assign y11721 = ~n30593 ;
  assign y11722 = ~1'b0 ;
  assign y11723 = ~1'b0 ;
  assign y11724 = n30596 ;
  assign y11725 = ~n30597 ;
  assign y11726 = n8075 ;
  assign y11727 = ~n30602 ;
  assign y11728 = ~1'b0 ;
  assign y11729 = n30604 ;
  assign y11730 = ~1'b0 ;
  assign y11731 = n30606 ;
  assign y11732 = ~n30607 ;
  assign y11733 = ~1'b0 ;
  assign y11734 = n30613 ;
  assign y11735 = ~1'b0 ;
  assign y11736 = n30617 ;
  assign y11737 = n30619 ;
  assign y11738 = n30622 ;
  assign y11739 = ~n30625 ;
  assign y11740 = ~n30626 ;
  assign y11741 = ~n30627 ;
  assign y11742 = ~n30631 ;
  assign y11743 = ~n30635 ;
  assign y11744 = n30636 ;
  assign y11745 = ~n30637 ;
  assign y11746 = n30638 ;
  assign y11747 = ~n30640 ;
  assign y11748 = n30651 ;
  assign y11749 = n30653 ;
  assign y11750 = ~n30654 ;
  assign y11751 = n30656 ;
  assign y11752 = ~n30659 ;
  assign y11753 = n30661 ;
  assign y11754 = ~n30663 ;
  assign y11755 = n30670 ;
  assign y11756 = ~n30676 ;
  assign y11757 = ~n30678 ;
  assign y11758 = ~n30680 ;
  assign y11759 = ~1'b0 ;
  assign y11760 = n30681 ;
  assign y11761 = n30683 ;
  assign y11762 = n30687 ;
  assign y11763 = ~n30691 ;
  assign y11764 = n30696 ;
  assign y11765 = n30698 ;
  assign y11766 = ~1'b0 ;
  assign y11767 = ~n30702 ;
  assign y11768 = ~n30704 ;
  assign y11769 = ~1'b0 ;
  assign y11770 = ~n30705 ;
  assign y11771 = n30708 ;
  assign y11772 = ~n30711 ;
  assign y11773 = ~n30713 ;
  assign y11774 = ~n30715 ;
  assign y11775 = ~n30717 ;
  assign y11776 = ~n30720 ;
  assign y11777 = n30721 ;
  assign y11778 = ~n30726 ;
  assign y11779 = ~1'b0 ;
  assign y11780 = ~n30733 ;
  assign y11781 = ~n30738 ;
  assign y11782 = ~n30739 ;
  assign y11783 = ~n30752 ;
  assign y11784 = ~n30755 ;
  assign y11785 = n30758 ;
  assign y11786 = n30759 ;
  assign y11787 = ~1'b0 ;
  assign y11788 = ~1'b0 ;
  assign y11789 = n30760 ;
  assign y11790 = ~1'b0 ;
  assign y11791 = ~n30761 ;
  assign y11792 = ~n30767 ;
  assign y11793 = n30769 ;
  assign y11794 = ~n30770 ;
  assign y11795 = ~n30771 ;
  assign y11796 = n30773 ;
  assign y11797 = ~n30774 ;
  assign y11798 = ~1'b0 ;
  assign y11799 = n30776 ;
  assign y11800 = ~n30779 ;
  assign y11801 = n30783 ;
  assign y11802 = ~n30790 ;
  assign y11803 = ~n30794 ;
  assign y11804 = n30802 ;
  assign y11805 = n30805 ;
  assign y11806 = n30806 ;
  assign y11807 = ~n30809 ;
  assign y11808 = n30812 ;
  assign y11809 = n30816 ;
  assign y11810 = n30820 ;
  assign y11811 = ~n30823 ;
  assign y11812 = ~n30825 ;
  assign y11813 = ~n30828 ;
  assign y11814 = ~n22143 ;
  assign y11815 = n9596 ;
  assign y11816 = ~1'b0 ;
  assign y11817 = n30839 ;
  assign y11818 = ~n30841 ;
  assign y11819 = n30844 ;
  assign y11820 = ~1'b0 ;
  assign y11821 = n30847 ;
  assign y11822 = ~1'b0 ;
  assign y11823 = n30850 ;
  assign y11824 = n30854 ;
  assign y11825 = n30855 ;
  assign y11826 = n30857 ;
  assign y11827 = ~n30860 ;
  assign y11828 = ~n30861 ;
  assign y11829 = ~1'b0 ;
  assign y11830 = n30862 ;
  assign y11831 = ~n30864 ;
  assign y11832 = ~1'b0 ;
  assign y11833 = ~n30869 ;
  assign y11834 = n30870 ;
  assign y11835 = ~1'b0 ;
  assign y11836 = ~1'b0 ;
  assign y11837 = n30871 ;
  assign y11838 = n30873 ;
  assign y11839 = n30876 ;
  assign y11840 = n30878 ;
  assign y11841 = n30883 ;
  assign y11842 = ~n30887 ;
  assign y11843 = n30896 ;
  assign y11844 = ~1'b0 ;
  assign y11845 = ~n30904 ;
  assign y11846 = ~n30906 ;
  assign y11847 = ~n30907 ;
  assign y11848 = ~1'b0 ;
  assign y11849 = ~n30912 ;
  assign y11850 = ~1'b0 ;
  assign y11851 = ~1'b0 ;
  assign y11852 = n30914 ;
  assign y11853 = ~n22004 ;
  assign y11854 = ~n30916 ;
  assign y11855 = ~1'b0 ;
  assign y11856 = ~n30917 ;
  assign y11857 = ~n30919 ;
  assign y11858 = n30925 ;
  assign y11859 = ~n30931 ;
  assign y11860 = n30935 ;
  assign y11861 = n30939 ;
  assign y11862 = ~n30942 ;
  assign y11863 = n30945 ;
  assign y11864 = n30954 ;
  assign y11865 = ~1'b0 ;
  assign y11866 = n30959 ;
  assign y11867 = ~n30962 ;
  assign y11868 = n30966 ;
  assign y11869 = ~n30973 ;
  assign y11870 = ~n30977 ;
  assign y11871 = ~1'b0 ;
  assign y11872 = ~1'b0 ;
  assign y11873 = n30979 ;
  assign y11874 = ~n30981 ;
  assign y11875 = ~1'b0 ;
  assign y11876 = ~1'b0 ;
  assign y11877 = ~1'b0 ;
  assign y11878 = n30985 ;
  assign y11879 = n30989 ;
  assign y11880 = n6182 ;
  assign y11881 = n30998 ;
  assign y11882 = ~1'b0 ;
  assign y11883 = n30999 ;
  assign y11884 = ~n31007 ;
  assign y11885 = ~1'b0 ;
  assign y11886 = ~n31009 ;
  assign y11887 = ~n31011 ;
  assign y11888 = n31012 ;
  assign y11889 = ~n31015 ;
  assign y11890 = ~n31018 ;
  assign y11891 = n31021 ;
  assign y11892 = n31023 ;
  assign y11893 = ~n31026 ;
  assign y11894 = n31030 ;
  assign y11895 = n31031 ;
  assign y11896 = n31034 ;
  assign y11897 = ~1'b0 ;
  assign y11898 = n31038 ;
  assign y11899 = ~1'b0 ;
  assign y11900 = n31040 ;
  assign y11901 = n31046 ;
  assign y11902 = ~n31048 ;
  assign y11903 = ~n31049 ;
  assign y11904 = ~n31051 ;
  assign y11905 = ~n31052 ;
  assign y11906 = 1'b0 ;
  assign y11907 = ~1'b0 ;
  assign y11908 = ~1'b0 ;
  assign y11909 = n31063 ;
  assign y11910 = n31064 ;
  assign y11911 = ~1'b0 ;
  assign y11912 = n31068 ;
  assign y11913 = ~1'b0 ;
  assign y11914 = ~n31069 ;
  assign y11915 = ~n31070 ;
  assign y11916 = n31078 ;
  assign y11917 = n31079 ;
  assign y11918 = n31081 ;
  assign y11919 = n31082 ;
  assign y11920 = ~n31087 ;
  assign y11921 = ~1'b0 ;
  assign y11922 = ~1'b0 ;
  assign y11923 = n31095 ;
  assign y11924 = ~n31098 ;
  assign y11925 = n31105 ;
  assign y11926 = ~n31106 ;
  assign y11927 = ~1'b0 ;
  assign y11928 = ~1'b0 ;
  assign y11929 = ~n31110 ;
  assign y11930 = n31111 ;
  assign y11931 = ~n31115 ;
  assign y11932 = n31122 ;
  assign y11933 = n31123 ;
  assign y11934 = n31125 ;
  assign y11935 = ~1'b0 ;
  assign y11936 = ~1'b0 ;
  assign y11937 = ~n31127 ;
  assign y11938 = n31128 ;
  assign y11939 = ~n31130 ;
  assign y11940 = ~1'b0 ;
  assign y11941 = ~n31134 ;
  assign y11942 = ~1'b0 ;
  assign y11943 = ~n31142 ;
  assign y11944 = ~n31143 ;
  assign y11945 = n31144 ;
  assign y11946 = ~n31146 ;
  assign y11947 = ~n31148 ;
  assign y11948 = ~n31149 ;
  assign y11949 = ~n31153 ;
  assign y11950 = ~n31156 ;
  assign y11951 = n31158 ;
  assign y11952 = ~n5602 ;
  assign y11953 = ~1'b0 ;
  assign y11954 = n31159 ;
  assign y11955 = ~1'b0 ;
  assign y11956 = n31160 ;
  assign y11957 = n31162 ;
  assign y11958 = ~n19976 ;
  assign y11959 = ~1'b0 ;
  assign y11960 = ~n31166 ;
  assign y11961 = ~n31167 ;
  assign y11962 = ~n6370 ;
  assign y11963 = n31168 ;
  assign y11964 = n31170 ;
  assign y11965 = n31175 ;
  assign y11966 = ~n31177 ;
  assign y11967 = ~n31183 ;
  assign y11968 = n31184 ;
  assign y11969 = ~1'b0 ;
  assign y11970 = ~1'b0 ;
  assign y11971 = n31189 ;
  assign y11972 = n31190 ;
  assign y11973 = ~1'b0 ;
  assign y11974 = n31195 ;
  assign y11975 = n31197 ;
  assign y11976 = ~n31199 ;
  assign y11977 = n31202 ;
  assign y11978 = ~n31205 ;
  assign y11979 = ~n31212 ;
  assign y11980 = n31214 ;
  assign y11981 = ~1'b0 ;
  assign y11982 = ~1'b0 ;
  assign y11983 = ~1'b0 ;
  assign y11984 = ~n31215 ;
  assign y11985 = ~n31218 ;
  assign y11986 = ~n31222 ;
  assign y11987 = ~1'b0 ;
  assign y11988 = n31227 ;
  assign y11989 = ~1'b0 ;
  assign y11990 = ~n31229 ;
  assign y11991 = ~n31230 ;
  assign y11992 = n31231 ;
  assign y11993 = ~n31233 ;
  assign y11994 = n31235 ;
  assign y11995 = ~n31236 ;
  assign y11996 = n31237 ;
  assign y11997 = n31241 ;
  assign y11998 = ~n31242 ;
  assign y11999 = ~n31245 ;
  assign y12000 = ~n31247 ;
  assign y12001 = ~n31248 ;
  assign y12002 = ~n31251 ;
  assign y12003 = n31253 ;
  assign y12004 = ~n7592 ;
  assign y12005 = ~n31255 ;
  assign y12006 = ~n31256 ;
  assign y12007 = ~n31257 ;
  assign y12008 = ~n31259 ;
  assign y12009 = ~n31260 ;
  assign y12010 = ~1'b0 ;
  assign y12011 = ~n31269 ;
  assign y12012 = ~1'b0 ;
  assign y12013 = ~n31270 ;
  assign y12014 = n31272 ;
  assign y12015 = ~1'b0 ;
  assign y12016 = ~1'b0 ;
  assign y12017 = ~n31273 ;
  assign y12018 = ~n31276 ;
  assign y12019 = ~n31277 ;
  assign y12020 = n31281 ;
  assign y12021 = ~1'b0 ;
  assign y12022 = ~1'b0 ;
  assign y12023 = ~1'b0 ;
  assign y12024 = ~n7098 ;
  assign y12025 = n31285 ;
  assign y12026 = n31288 ;
  assign y12027 = ~n31289 ;
  assign y12028 = ~1'b0 ;
  assign y12029 = ~n31291 ;
  assign y12030 = ~1'b0 ;
  assign y12031 = ~1'b0 ;
  assign y12032 = n31296 ;
  assign y12033 = n31298 ;
  assign y12034 = n31305 ;
  assign y12035 = n31306 ;
  assign y12036 = ~n31307 ;
  assign y12037 = n31310 ;
  assign y12038 = ~1'b0 ;
  assign y12039 = n31317 ;
  assign y12040 = n31318 ;
  assign y12041 = ~n31325 ;
  assign y12042 = n31326 ;
  assign y12043 = n31327 ;
  assign y12044 = n27094 ;
  assign y12045 = ~n31329 ;
  assign y12046 = ~n31333 ;
  assign y12047 = ~n31337 ;
  assign y12048 = ~n31341 ;
  assign y12049 = ~n31344 ;
  assign y12050 = ~n31347 ;
  assign y12051 = ~n31351 ;
  assign y12052 = n31353 ;
  assign y12053 = n31360 ;
  assign y12054 = n31362 ;
  assign y12055 = ~n31363 ;
  assign y12056 = ~n31369 ;
  assign y12057 = ~n31372 ;
  assign y12058 = n31375 ;
  assign y12059 = ~n31376 ;
  assign y12060 = n31378 ;
  assign y12061 = ~1'b0 ;
  assign y12062 = ~n31380 ;
  assign y12063 = n31382 ;
  assign y12064 = ~n31384 ;
  assign y12065 = ~n31391 ;
  assign y12066 = ~n31396 ;
  assign y12067 = n31397 ;
  assign y12068 = ~n31399 ;
  assign y12069 = ~n31405 ;
  assign y12070 = ~1'b0 ;
  assign y12071 = 1'b0 ;
  assign y12072 = ~1'b0 ;
  assign y12073 = ~n31407 ;
  assign y12074 = ~n31408 ;
  assign y12075 = ~n31411 ;
  assign y12076 = n31412 ;
  assign y12077 = ~n31416 ;
  assign y12078 = ~1'b0 ;
  assign y12079 = ~1'b0 ;
  assign y12080 = ~n31423 ;
  assign y12081 = ~1'b0 ;
  assign y12082 = ~n31424 ;
  assign y12083 = n31428 ;
  assign y12084 = n31431 ;
  assign y12085 = ~1'b0 ;
  assign y12086 = n31435 ;
  assign y12087 = ~1'b0 ;
  assign y12088 = ~1'b0 ;
  assign y12089 = ~n31436 ;
  assign y12090 = n4405 ;
  assign y12091 = ~n31438 ;
  assign y12092 = ~1'b0 ;
  assign y12093 = ~n31442 ;
  assign y12094 = ~1'b0 ;
  assign y12095 = n17497 ;
  assign y12096 = ~n31446 ;
  assign y12097 = n31447 ;
  assign y12098 = ~n31452 ;
  assign y12099 = ~n31453 ;
  assign y12100 = n31454 ;
  assign y12101 = ~n31458 ;
  assign y12102 = n31460 ;
  assign y12103 = ~1'b0 ;
  assign y12104 = ~n31467 ;
  assign y12105 = ~1'b0 ;
  assign y12106 = ~n31469 ;
  assign y12107 = ~n31470 ;
  assign y12108 = n31473 ;
  assign y12109 = n31474 ;
  assign y12110 = ~n31478 ;
  assign y12111 = ~1'b0 ;
  assign y12112 = n31479 ;
  assign y12113 = ~n31480 ;
  assign y12114 = ~n31483 ;
  assign y12115 = n31484 ;
  assign y12116 = ~n31487 ;
  assign y12117 = n31489 ;
  assign y12118 = ~n31491 ;
  assign y12119 = n31494 ;
  assign y12120 = ~n31503 ;
  assign y12121 = n31505 ;
  assign y12122 = ~n31509 ;
  assign y12123 = ~n31511 ;
  assign y12124 = ~1'b0 ;
  assign y12125 = n31512 ;
  assign y12126 = ~n31514 ;
  assign y12127 = ~1'b0 ;
  assign y12128 = ~n31518 ;
  assign y12129 = ~n31519 ;
  assign y12130 = n31523 ;
  assign y12131 = n31526 ;
  assign y12132 = n31527 ;
  assign y12133 = n31529 ;
  assign y12134 = n31530 ;
  assign y12135 = ~n31531 ;
  assign y12136 = ~n31535 ;
  assign y12137 = n31542 ;
  assign y12138 = n31544 ;
  assign y12139 = n31546 ;
  assign y12140 = n31548 ;
  assign y12141 = ~n31551 ;
  assign y12142 = n31553 ;
  assign y12143 = ~n31563 ;
  assign y12144 = ~n31565 ;
  assign y12145 = n31566 ;
  assign y12146 = n31567 ;
  assign y12147 = ~1'b0 ;
  assign y12148 = ~n31569 ;
  assign y12149 = ~1'b0 ;
  assign y12150 = ~n31571 ;
  assign y12151 = n31572 ;
  assign y12152 = ~n31575 ;
  assign y12153 = n31579 ;
  assign y12154 = ~n31581 ;
  assign y12155 = ~1'b0 ;
  assign y12156 = ~n31586 ;
  assign y12157 = ~n31589 ;
  assign y12158 = n31593 ;
  assign y12159 = ~1'b0 ;
  assign y12160 = n31594 ;
  assign y12161 = n31596 ;
  assign y12162 = n31599 ;
  assign y12163 = n31600 ;
  assign y12164 = ~n31602 ;
  assign y12165 = ~1'b0 ;
  assign y12166 = ~n31606 ;
  assign y12167 = ~n31608 ;
  assign y12168 = n31610 ;
  assign y12169 = ~n31613 ;
  assign y12170 = ~n31614 ;
  assign y12171 = n31615 ;
  assign y12172 = ~n31617 ;
  assign y12173 = n31621 ;
  assign y12174 = ~n31622 ;
  assign y12175 = n31625 ;
  assign y12176 = ~n31626 ;
  assign y12177 = ~n31633 ;
  assign y12178 = n31636 ;
  assign y12179 = n31640 ;
  assign y12180 = ~n31641 ;
  assign y12181 = n31643 ;
  assign y12182 = n31651 ;
  assign y12183 = ~n31654 ;
  assign y12184 = n31656 ;
  assign y12185 = n31659 ;
  assign y12186 = ~1'b0 ;
  assign y12187 = n31661 ;
  assign y12188 = ~n31663 ;
  assign y12189 = ~n31668 ;
  assign y12190 = ~1'b0 ;
  assign y12191 = ~1'b0 ;
  assign y12192 = ~n31669 ;
  assign y12193 = n31672 ;
  assign y12194 = n31674 ;
  assign y12195 = ~n31676 ;
  assign y12196 = n31677 ;
  assign y12197 = ~1'b0 ;
  assign y12198 = ~n31679 ;
  assign y12199 = n31680 ;
  assign y12200 = n31689 ;
  assign y12201 = n31690 ;
  assign y12202 = ~n31691 ;
  assign y12203 = ~1'b0 ;
  assign y12204 = n31704 ;
  assign y12205 = ~n31705 ;
  assign y12206 = n31706 ;
  assign y12207 = n11363 ;
  assign y12208 = ~1'b0 ;
  assign y12209 = n31714 ;
  assign y12210 = ~n31716 ;
  assign y12211 = ~n31717 ;
  assign y12212 = ~n31721 ;
  assign y12213 = ~1'b0 ;
  assign y12214 = ~n31725 ;
  assign y12215 = n31726 ;
  assign y12216 = ~n31727 ;
  assign y12217 = ~n31731 ;
  assign y12218 = ~n31732 ;
  assign y12219 = ~n31736 ;
  assign y12220 = ~n31738 ;
  assign y12221 = ~n31739 ;
  assign y12222 = ~1'b0 ;
  assign y12223 = ~1'b0 ;
  assign y12224 = n31742 ;
  assign y12225 = ~n31745 ;
  assign y12226 = ~1'b0 ;
  assign y12227 = ~n31749 ;
  assign y12228 = n31753 ;
  assign y12229 = n31756 ;
  assign y12230 = ~1'b0 ;
  assign y12231 = n31757 ;
  assign y12232 = ~n31762 ;
  assign y12233 = n31768 ;
  assign y12234 = ~n31770 ;
  assign y12235 = n31774 ;
  assign y12236 = n19842 ;
  assign y12237 = ~n31775 ;
  assign y12238 = ~1'b0 ;
  assign y12239 = n31776 ;
  assign y12240 = ~n31777 ;
  assign y12241 = ~n31784 ;
  assign y12242 = n31785 ;
  assign y12243 = n31787 ;
  assign y12244 = ~n31792 ;
  assign y12245 = n31798 ;
  assign y12246 = ~n31804 ;
  assign y12247 = ~n31808 ;
  assign y12248 = ~1'b0 ;
  assign y12249 = ~1'b0 ;
  assign y12250 = ~1'b0 ;
  assign y12251 = ~n31809 ;
  assign y12252 = n31811 ;
  assign y12253 = ~1'b0 ;
  assign y12254 = ~n31814 ;
  assign y12255 = n31815 ;
  assign y12256 = ~n31816 ;
  assign y12257 = ~n31819 ;
  assign y12258 = ~n31822 ;
  assign y12259 = n31823 ;
  assign y12260 = ~1'b0 ;
  assign y12261 = n31827 ;
  assign y12262 = n31828 ;
  assign y12263 = n31834 ;
  assign y12264 = ~n31835 ;
  assign y12265 = n31840 ;
  assign y12266 = ~1'b0 ;
  assign y12267 = ~n31841 ;
  assign y12268 = ~1'b0 ;
  assign y12269 = ~n31842 ;
  assign y12270 = ~n31845 ;
  assign y12271 = ~n31846 ;
  assign y12272 = n31847 ;
  assign y12273 = ~n31851 ;
  assign y12274 = ~1'b0 ;
  assign y12275 = n31854 ;
  assign y12276 = n31856 ;
  assign y12277 = n31860 ;
  assign y12278 = ~1'b0 ;
  assign y12279 = ~n31866 ;
  assign y12280 = ~n31867 ;
  assign y12281 = n31869 ;
  assign y12282 = ~n31871 ;
  assign y12283 = ~n31873 ;
  assign y12284 = ~n31875 ;
  assign y12285 = ~n31876 ;
  assign y12286 = ~n31879 ;
  assign y12287 = n31881 ;
  assign y12288 = n31885 ;
  assign y12289 = ~1'b0 ;
  assign y12290 = n31887 ;
  assign y12291 = n31889 ;
  assign y12292 = n31890 ;
  assign y12293 = ~n31891 ;
  assign y12294 = ~1'b0 ;
  assign y12295 = n31893 ;
  assign y12296 = ~n31894 ;
  assign y12297 = ~n31895 ;
  assign y12298 = ~n31898 ;
  assign y12299 = n31901 ;
  assign y12300 = ~n31902 ;
  assign y12301 = n31903 ;
  assign y12302 = ~n31906 ;
  assign y12303 = ~1'b0 ;
  assign y12304 = ~n31909 ;
  assign y12305 = ~1'b0 ;
  assign y12306 = n31910 ;
  assign y12307 = ~n31911 ;
  assign y12308 = n31914 ;
  assign y12309 = n31917 ;
  assign y12310 = n31920 ;
  assign y12311 = ~n31921 ;
  assign y12312 = ~1'b0 ;
  assign y12313 = n31931 ;
  assign y12314 = n31933 ;
  assign y12315 = n31934 ;
  assign y12316 = ~n3810 ;
  assign y12317 = ~1'b0 ;
  assign y12318 = n31935 ;
  assign y12319 = 1'b0 ;
  assign y12320 = ~1'b0 ;
  assign y12321 = ~n31938 ;
  assign y12322 = n31942 ;
  assign y12323 = n31943 ;
  assign y12324 = ~n31945 ;
  assign y12325 = n15086 ;
  assign y12326 = ~1'b0 ;
  assign y12327 = n31948 ;
  assign y12328 = ~n31952 ;
  assign y12329 = n31954 ;
  assign y12330 = n31959 ;
  assign y12331 = n31960 ;
  assign y12332 = ~1'b0 ;
  assign y12333 = ~n31963 ;
  assign y12334 = ~n31964 ;
  assign y12335 = n31969 ;
  assign y12336 = ~n31971 ;
  assign y12337 = n31976 ;
  assign y12338 = n31978 ;
  assign y12339 = ~1'b0 ;
  assign y12340 = ~n6062 ;
  assign y12341 = n31981 ;
  assign y12342 = ~n31984 ;
  assign y12343 = n31986 ;
  assign y12344 = ~1'b0 ;
  assign y12345 = ~n31987 ;
  assign y12346 = ~n31990 ;
  assign y12347 = n7124 ;
  assign y12348 = n31996 ;
  assign y12349 = n31997 ;
  assign y12350 = ~n31998 ;
  assign y12351 = n32001 ;
  assign y12352 = ~n32002 ;
  assign y12353 = ~n32011 ;
  assign y12354 = ~n32013 ;
  assign y12355 = ~1'b0 ;
  assign y12356 = ~n32014 ;
  assign y12357 = ~n32016 ;
  assign y12358 = ~1'b0 ;
  assign y12359 = n32021 ;
  assign y12360 = ~n32026 ;
  assign y12361 = n32033 ;
  assign y12362 = ~n32034 ;
  assign y12363 = ~n32035 ;
  assign y12364 = ~n32039 ;
  assign y12365 = n32042 ;
  assign y12366 = n32045 ;
  assign y12367 = n32047 ;
  assign y12368 = ~1'b0 ;
  assign y12369 = ~n32051 ;
  assign y12370 = n32052 ;
  assign y12371 = ~n32053 ;
  assign y12372 = n32054 ;
  assign y12373 = ~1'b0 ;
  assign y12374 = n32056 ;
  assign y12375 = ~n32057 ;
  assign y12376 = n32058 ;
  assign y12377 = ~1'b0 ;
  assign y12378 = ~1'b0 ;
  assign y12379 = ~n32059 ;
  assign y12380 = n32060 ;
  assign y12381 = n32065 ;
  assign y12382 = ~1'b0 ;
  assign y12383 = ~n32066 ;
  assign y12384 = n32069 ;
  assign y12385 = ~n32072 ;
  assign y12386 = ~n32074 ;
  assign y12387 = ~n32075 ;
  assign y12388 = ~1'b0 ;
  assign y12389 = ~n32076 ;
  assign y12390 = n32082 ;
  assign y12391 = ~n32086 ;
  assign y12392 = ~1'b0 ;
  assign y12393 = ~1'b0 ;
  assign y12394 = ~1'b0 ;
  assign y12395 = ~1'b0 ;
  assign y12396 = ~n32087 ;
  assign y12397 = n32090 ;
  assign y12398 = ~n32098 ;
  assign y12399 = ~n32101 ;
  assign y12400 = ~1'b0 ;
  assign y12401 = n32103 ;
  assign y12402 = ~n32106 ;
  assign y12403 = ~n32108 ;
  assign y12404 = n32109 ;
  assign y12405 = ~n32110 ;
  assign y12406 = ~1'b0 ;
  assign y12407 = n32113 ;
  assign y12408 = ~1'b0 ;
  assign y12409 = n32114 ;
  assign y12410 = ~n32115 ;
  assign y12411 = 1'b0 ;
  assign y12412 = ~n32118 ;
  assign y12413 = ~n32124 ;
  assign y12414 = ~n32127 ;
  assign y12415 = n32130 ;
  assign y12416 = ~n32136 ;
  assign y12417 = ~1'b0 ;
  assign y12418 = n32144 ;
  assign y12419 = n5793 ;
  assign y12420 = n32146 ;
  assign y12421 = n32147 ;
  assign y12422 = ~n32148 ;
  assign y12423 = ~n32152 ;
  assign y12424 = ~n19042 ;
  assign y12425 = n32153 ;
  assign y12426 = ~1'b0 ;
  assign y12427 = n32156 ;
  assign y12428 = ~n32157 ;
  assign y12429 = ~n32159 ;
  assign y12430 = ~n32160 ;
  assign y12431 = n32162 ;
  assign y12432 = ~n32164 ;
  assign y12433 = ~n32165 ;
  assign y12434 = ~n32172 ;
  assign y12435 = n32173 ;
  assign y12436 = ~n32174 ;
  assign y12437 = n32178 ;
  assign y12438 = ~1'b0 ;
  assign y12439 = ~1'b0 ;
  assign y12440 = ~1'b0 ;
  assign y12441 = ~n32179 ;
  assign y12442 = ~n32180 ;
  assign y12443 = n32181 ;
  assign y12444 = n32184 ;
  assign y12445 = ~n32185 ;
  assign y12446 = ~n32186 ;
  assign y12447 = ~n32189 ;
  assign y12448 = ~1'b0 ;
  assign y12449 = ~n32192 ;
  assign y12450 = n32027 ;
  assign y12451 = ~n32195 ;
  assign y12452 = ~1'b0 ;
  assign y12453 = n32197 ;
  assign y12454 = ~1'b0 ;
  assign y12455 = ~1'b0 ;
  assign y12456 = ~n32201 ;
  assign y12457 = ~n32202 ;
  assign y12458 = ~n32205 ;
  assign y12459 = ~1'b0 ;
  assign y12460 = n32206 ;
  assign y12461 = n32208 ;
  assign y12462 = ~1'b0 ;
  assign y12463 = ~1'b0 ;
  assign y12464 = ~n32211 ;
  assign y12465 = ~n32214 ;
  assign y12466 = ~n32215 ;
  assign y12467 = ~n32220 ;
  assign y12468 = ~1'b0 ;
  assign y12469 = n32224 ;
  assign y12470 = ~n32225 ;
  assign y12471 = ~n32228 ;
  assign y12472 = ~n32229 ;
  assign y12473 = ~n32231 ;
  assign y12474 = ~n32232 ;
  assign y12475 = n32241 ;
  assign y12476 = ~1'b0 ;
  assign y12477 = n32242 ;
  assign y12478 = ~n32244 ;
  assign y12479 = ~n32247 ;
  assign y12480 = n32250 ;
  assign y12481 = n32252 ;
  assign y12482 = ~n32255 ;
  assign y12483 = ~n32256 ;
  assign y12484 = ~1'b0 ;
  assign y12485 = ~n32257 ;
  assign y12486 = ~1'b0 ;
  assign y12487 = ~1'b0 ;
  assign y12488 = n32262 ;
  assign y12489 = ~n32264 ;
  assign y12490 = n32268 ;
  assign y12491 = ~n32272 ;
  assign y12492 = n32278 ;
  assign y12493 = ~n32280 ;
  assign y12494 = ~1'b0 ;
  assign y12495 = ~n8236 ;
  assign y12496 = n32284 ;
  assign y12497 = n32285 ;
  assign y12498 = ~1'b0 ;
  assign y12499 = ~1'b0 ;
  assign y12500 = ~n32286 ;
  assign y12501 = n32287 ;
  assign y12502 = ~n31199 ;
  assign y12503 = ~n32289 ;
  assign y12504 = n32294 ;
  assign y12505 = ~n32305 ;
  assign y12506 = n32306 ;
  assign y12507 = n32310 ;
  assign y12508 = n32311 ;
  assign y12509 = ~n32312 ;
  assign y12510 = ~1'b0 ;
  assign y12511 = ~1'b0 ;
  assign y12512 = n32315 ;
  assign y12513 = ~1'b0 ;
  assign y12514 = n32316 ;
  assign y12515 = n32317 ;
  assign y12516 = n32318 ;
  assign y12517 = n32320 ;
  assign y12518 = n32324 ;
  assign y12519 = ~1'b0 ;
  assign y12520 = ~1'b0 ;
  assign y12521 = n32331 ;
  assign y12522 = ~1'b0 ;
  assign y12523 = ~1'b0 ;
  assign y12524 = n32333 ;
  assign y12525 = n32335 ;
  assign y12526 = ~n32337 ;
  assign y12527 = ~n20501 ;
  assign y12528 = n32339 ;
  assign y12529 = ~n32341 ;
  assign y12530 = ~1'b0 ;
  assign y12531 = ~n32343 ;
  assign y12532 = ~n32348 ;
  assign y12533 = n32352 ;
  assign y12534 = n32353 ;
  assign y12535 = ~n32357 ;
  assign y12536 = ~n32362 ;
  assign y12537 = ~1'b0 ;
  assign y12538 = ~n32363 ;
  assign y12539 = n32365 ;
  assign y12540 = ~n32366 ;
  assign y12541 = ~1'b0 ;
  assign y12542 = ~n32369 ;
  assign y12543 = ~1'b0 ;
  assign y12544 = ~1'b0 ;
  assign y12545 = n32371 ;
  assign y12546 = ~1'b0 ;
  assign y12547 = n32374 ;
  assign y12548 = n32379 ;
  assign y12549 = n32387 ;
  assign y12550 = ~1'b0 ;
  assign y12551 = n32389 ;
  assign y12552 = n32395 ;
  assign y12553 = ~n32400 ;
  assign y12554 = ~n32402 ;
  assign y12555 = n32405 ;
  assign y12556 = ~n32411 ;
  assign y12557 = ~1'b0 ;
  assign y12558 = n32414 ;
  assign y12559 = ~1'b0 ;
  assign y12560 = n32415 ;
  assign y12561 = 1'b0 ;
  assign y12562 = n32416 ;
  assign y12563 = n32418 ;
  assign y12564 = n32419 ;
  assign y12565 = n32420 ;
  assign y12566 = n32422 ;
  assign y12567 = ~1'b0 ;
  assign y12568 = n32424 ;
  assign y12569 = n32427 ;
  assign y12570 = ~n32429 ;
  assign y12571 = ~n32430 ;
  assign y12572 = ~n32432 ;
  assign y12573 = n32435 ;
  assign y12574 = ~n32436 ;
  assign y12575 = n32444 ;
  assign y12576 = ~n32447 ;
  assign y12577 = n32448 ;
  assign y12578 = n32449 ;
  assign y12579 = n32451 ;
  assign y12580 = n32455 ;
  assign y12581 = ~1'b0 ;
  assign y12582 = n32458 ;
  assign y12583 = ~n32461 ;
  assign y12584 = n15961 ;
  assign y12585 = ~n32464 ;
  assign y12586 = ~1'b0 ;
  assign y12587 = ~n32467 ;
  assign y12588 = ~1'b0 ;
  assign y12589 = ~n32471 ;
  assign y12590 = ~n32474 ;
  assign y12591 = n32475 ;
  assign y12592 = ~1'b0 ;
  assign y12593 = n31794 ;
  assign y12594 = n32478 ;
  assign y12595 = ~n32481 ;
  assign y12596 = ~1'b0 ;
  assign y12597 = 1'b0 ;
  assign y12598 = n3515 ;
  assign y12599 = n32485 ;
  assign y12600 = ~n32486 ;
  assign y12601 = ~n32489 ;
  assign y12602 = n15741 ;
  assign y12603 = ~n32490 ;
  assign y12604 = ~n32492 ;
  assign y12605 = n32494 ;
  assign y12606 = n26797 ;
  assign y12607 = n2394 ;
  assign y12608 = ~n32495 ;
  assign y12609 = n32501 ;
  assign y12610 = n32502 ;
  assign y12611 = n32505 ;
  assign y12612 = n32507 ;
  assign y12613 = ~n32511 ;
  assign y12614 = ~n32513 ;
  assign y12615 = ~n32515 ;
  assign y12616 = n32517 ;
  assign y12617 = ~n32521 ;
  assign y12618 = ~1'b0 ;
  assign y12619 = n32524 ;
  assign y12620 = n32526 ;
  assign y12621 = ~n32528 ;
  assign y12622 = ~n32531 ;
  assign y12623 = ~n32533 ;
  assign y12624 = n32535 ;
  assign y12625 = ~n32538 ;
  assign y12626 = ~n32539 ;
  assign y12627 = ~n32540 ;
  assign y12628 = ~1'b0 ;
  assign y12629 = ~1'b0 ;
  assign y12630 = n32542 ;
  assign y12631 = ~n32546 ;
  assign y12632 = n32547 ;
  assign y12633 = n32548 ;
  assign y12634 = ~1'b0 ;
  assign y12635 = n32550 ;
  assign y12636 = ~n32556 ;
  assign y12637 = ~n13495 ;
  assign y12638 = ~n32558 ;
  assign y12639 = ~1'b0 ;
  assign y12640 = n32563 ;
  assign y12641 = ~n32565 ;
  assign y12642 = ~n32567 ;
  assign y12643 = ~n32571 ;
  assign y12644 = n32579 ;
  assign y12645 = ~n32581 ;
  assign y12646 = ~n32583 ;
  assign y12647 = ~1'b0 ;
  assign y12648 = ~1'b0 ;
  assign y12649 = n32592 ;
  assign y12650 = n4310 ;
  assign y12651 = n32595 ;
  assign y12652 = ~n32597 ;
  assign y12653 = ~n32601 ;
  assign y12654 = ~1'b0 ;
  assign y12655 = ~1'b0 ;
  assign y12656 = n32602 ;
  assign y12657 = n32603 ;
  assign y12658 = ~1'b0 ;
  assign y12659 = n32606 ;
  assign y12660 = ~n32607 ;
  assign y12661 = ~n32609 ;
  assign y12662 = ~n32611 ;
  assign y12663 = ~n32615 ;
  assign y12664 = ~n32618 ;
  assign y12665 = ~n17769 ;
  assign y12666 = ~1'b0 ;
  assign y12667 = ~n32619 ;
  assign y12668 = n32624 ;
  assign y12669 = ~n32631 ;
  assign y12670 = n32632 ;
  assign y12671 = n32636 ;
  assign y12672 = n32637 ;
  assign y12673 = n32640 ;
  assign y12674 = ~1'b0 ;
  assign y12675 = ~1'b0 ;
  assign y12676 = n32644 ;
  assign y12677 = n32645 ;
  assign y12678 = n32646 ;
  assign y12679 = n5146 ;
  assign y12680 = n32647 ;
  assign y12681 = ~1'b0 ;
  assign y12682 = n32651 ;
  assign y12683 = n32652 ;
  assign y12684 = ~n32653 ;
  assign y12685 = ~n32656 ;
  assign y12686 = ~n32661 ;
  assign y12687 = ~1'b0 ;
  assign y12688 = ~n32662 ;
  assign y12689 = n32664 ;
  assign y12690 = n32668 ;
  assign y12691 = n32669 ;
  assign y12692 = n32670 ;
  assign y12693 = ~n32675 ;
  assign y12694 = n32678 ;
  assign y12695 = ~n32680 ;
  assign y12696 = n32684 ;
  assign y12697 = ~1'b0 ;
  assign y12698 = ~n32687 ;
  assign y12699 = ~n32694 ;
  assign y12700 = ~1'b0 ;
  assign y12701 = n32697 ;
  assign y12702 = ~1'b0 ;
  assign y12703 = n32702 ;
  assign y12704 = ~1'b0 ;
  assign y12705 = n32703 ;
  assign y12706 = ~n13102 ;
  assign y12707 = ~1'b0 ;
  assign y12708 = ~1'b0 ;
  assign y12709 = ~1'b0 ;
  assign y12710 = n32704 ;
  assign y12711 = ~1'b0 ;
  assign y12712 = ~n32708 ;
  assign y12713 = ~n32712 ;
  assign y12714 = ~n32716 ;
  assign y12715 = n32717 ;
  assign y12716 = n32719 ;
  assign y12717 = n32720 ;
  assign y12718 = n32721 ;
  assign y12719 = ~n14914 ;
  assign y12720 = ~n32726 ;
  assign y12721 = ~n32730 ;
  assign y12722 = n32734 ;
  assign y12723 = ~1'b0 ;
  assign y12724 = n32738 ;
  assign y12725 = ~n32739 ;
  assign y12726 = ~1'b0 ;
  assign y12727 = ~1'b0 ;
  assign y12728 = n32740 ;
  assign y12729 = n32750 ;
  assign y12730 = ~1'b0 ;
  assign y12731 = ~1'b0 ;
  assign y12732 = n32751 ;
  assign y12733 = ~n32758 ;
  assign y12734 = ~n32759 ;
  assign y12735 = ~n32760 ;
  assign y12736 = ~n32761 ;
  assign y12737 = ~n32764 ;
  assign y12738 = n32770 ;
  assign y12739 = ~n32772 ;
  assign y12740 = ~n32774 ;
  assign y12741 = ~1'b0 ;
  assign y12742 = ~1'b0 ;
  assign y12743 = n32777 ;
  assign y12744 = n32778 ;
  assign y12745 = ~n24153 ;
  assign y12746 = ~1'b0 ;
  assign y12747 = ~n32783 ;
  assign y12748 = ~n32789 ;
  assign y12749 = ~n32793 ;
  assign y12750 = n32794 ;
  assign y12751 = n32796 ;
  assign y12752 = ~n32798 ;
  assign y12753 = ~n32800 ;
  assign y12754 = n32801 ;
  assign y12755 = n32803 ;
  assign y12756 = n32804 ;
  assign y12757 = n32807 ;
  assign y12758 = ~n32808 ;
  assign y12759 = ~1'b0 ;
  assign y12760 = n32810 ;
  assign y12761 = ~n32812 ;
  assign y12762 = ~1'b0 ;
  assign y12763 = ~n32814 ;
  assign y12764 = n32816 ;
  assign y12765 = n32823 ;
  assign y12766 = ~n32824 ;
  assign y12767 = ~n32826 ;
  assign y12768 = ~1'b0 ;
  assign y12769 = ~n32830 ;
  assign y12770 = ~n32832 ;
  assign y12771 = n32833 ;
  assign y12772 = ~n32835 ;
  assign y12773 = ~n32837 ;
  assign y12774 = ~n12226 ;
  assign y12775 = n32841 ;
  assign y12776 = ~n32844 ;
  assign y12777 = n32845 ;
  assign y12778 = n32849 ;
  assign y12779 = ~1'b0 ;
  assign y12780 = ~1'b0 ;
  assign y12781 = ~1'b0 ;
  assign y12782 = n32857 ;
  assign y12783 = ~n32858 ;
  assign y12784 = ~n32860 ;
  assign y12785 = ~n32865 ;
  assign y12786 = n32866 ;
  assign y12787 = ~n32867 ;
  assign y12788 = ~n32870 ;
  assign y12789 = ~n32871 ;
  assign y12790 = ~n32878 ;
  assign y12791 = n32879 ;
  assign y12792 = ~1'b0 ;
  assign y12793 = n32883 ;
  assign y12794 = n32884 ;
  assign y12795 = ~1'b0 ;
  assign y12796 = n32887 ;
  assign y12797 = n32888 ;
  assign y12798 = n32890 ;
  assign y12799 = n32894 ;
  assign y12800 = ~n32896 ;
  assign y12801 = n32900 ;
  assign y12802 = ~1'b0 ;
  assign y12803 = n32909 ;
  assign y12804 = ~n32912 ;
  assign y12805 = ~n32914 ;
  assign y12806 = ~n32915 ;
  assign y12807 = ~n32916 ;
  assign y12808 = ~1'b0 ;
  assign y12809 = ~1'b0 ;
  assign y12810 = ~n32917 ;
  assign y12811 = n32919 ;
  assign y12812 = ~1'b0 ;
  assign y12813 = ~n32920 ;
  assign y12814 = n32924 ;
  assign y12815 = ~n32929 ;
  assign y12816 = ~1'b0 ;
  assign y12817 = n32933 ;
  assign y12818 = ~n32936 ;
  assign y12819 = ~n32942 ;
  assign y12820 = n32944 ;
  assign y12821 = ~n9837 ;
  assign y12822 = n32946 ;
  assign y12823 = ~n32952 ;
  assign y12824 = n32953 ;
  assign y12825 = ~1'b0 ;
  assign y12826 = n32955 ;
  assign y12827 = ~n32956 ;
  assign y12828 = ~n32965 ;
  assign y12829 = n32967 ;
  assign y12830 = ~n32969 ;
  assign y12831 = n32970 ;
  assign y12832 = n32977 ;
  assign y12833 = ~n32982 ;
  assign y12834 = ~1'b0 ;
  assign y12835 = ~n32983 ;
  assign y12836 = n32984 ;
  assign y12837 = 1'b0 ;
  assign y12838 = ~1'b0 ;
  assign y12839 = ~n32986 ;
  assign y12840 = n32992 ;
  assign y12841 = n32998 ;
  assign y12842 = n33001 ;
  assign y12843 = ~n33005 ;
  assign y12844 = ~n33006 ;
  assign y12845 = n33011 ;
  assign y12846 = ~1'b0 ;
  assign y12847 = ~n33015 ;
  assign y12848 = ~n33016 ;
  assign y12849 = ~n33018 ;
  assign y12850 = ~n18833 ;
  assign y12851 = n33020 ;
  assign y12852 = ~n33022 ;
  assign y12853 = ~1'b0 ;
  assign y12854 = ~n33025 ;
  assign y12855 = n33028 ;
  assign y12856 = ~n8025 ;
  assign y12857 = ~1'b0 ;
  assign y12858 = n33030 ;
  assign y12859 = ~n33034 ;
  assign y12860 = n33038 ;
  assign y12861 = ~1'b0 ;
  assign y12862 = ~n33043 ;
  assign y12863 = n33045 ;
  assign y12864 = n33046 ;
  assign y12865 = ~1'b0 ;
  assign y12866 = n31071 ;
  assign y12867 = ~n33049 ;
  assign y12868 = n33052 ;
  assign y12869 = n33054 ;
  assign y12870 = n33056 ;
  assign y12871 = ~n33059 ;
  assign y12872 = n33063 ;
  assign y12873 = ~n33065 ;
  assign y12874 = ~1'b0 ;
  assign y12875 = ~n33067 ;
  assign y12876 = n33068 ;
  assign y12877 = n33069 ;
  assign y12878 = n33071 ;
  assign y12879 = ~1'b0 ;
  assign y12880 = ~1'b0 ;
  assign y12881 = ~1'b0 ;
  assign y12882 = 1'b0 ;
  assign y12883 = n33073 ;
  assign y12884 = n33076 ;
  assign y12885 = n33078 ;
  assign y12886 = ~n33080 ;
  assign y12887 = ~1'b0 ;
  assign y12888 = n33082 ;
  assign y12889 = n33083 ;
  assign y12890 = ~n33086 ;
  assign y12891 = n33087 ;
  assign y12892 = ~n33089 ;
  assign y12893 = ~n33096 ;
  assign y12894 = ~1'b0 ;
  assign y12895 = ~n33100 ;
  assign y12896 = ~1'b0 ;
  assign y12897 = n33103 ;
  assign y12898 = ~n33104 ;
  assign y12899 = ~n33105 ;
  assign y12900 = ~n33107 ;
  assign y12901 = ~n33108 ;
  assign y12902 = n33111 ;
  assign y12903 = ~n33114 ;
  assign y12904 = ~n33119 ;
  assign y12905 = ~1'b0 ;
  assign y12906 = ~n33122 ;
  assign y12907 = n33123 ;
  assign y12908 = ~n33125 ;
  assign y12909 = ~n33127 ;
  assign y12910 = ~n33128 ;
  assign y12911 = ~1'b0 ;
  assign y12912 = ~n33129 ;
  assign y12913 = n33133 ;
  assign y12914 = n33136 ;
  assign y12915 = ~1'b0 ;
  assign y12916 = ~n33138 ;
  assign y12917 = n33140 ;
  assign y12918 = ~1'b0 ;
  assign y12919 = ~1'b0 ;
  assign y12920 = n33141 ;
  assign y12921 = x178 ;
  assign y12922 = ~n33144 ;
  assign y12923 = ~n33148 ;
  assign y12924 = n33154 ;
  assign y12925 = ~1'b0 ;
  assign y12926 = ~1'b0 ;
  assign y12927 = ~n33155 ;
  assign y12928 = ~n33156 ;
  assign y12929 = ~n33160 ;
  assign y12930 = ~n33162 ;
  assign y12931 = ~1'b0 ;
  assign y12932 = ~n33167 ;
  assign y12933 = ~n33168 ;
  assign y12934 = ~1'b0 ;
  assign y12935 = n33170 ;
  assign y12936 = ~n33171 ;
  assign y12937 = n33172 ;
  assign y12938 = n33174 ;
  assign y12939 = n33176 ;
  assign y12940 = n33182 ;
  assign y12941 = n33184 ;
  assign y12942 = n33190 ;
  assign y12943 = n33195 ;
  assign y12944 = ~n33201 ;
  assign y12945 = ~n33203 ;
  assign y12946 = ~n33205 ;
  assign y12947 = ~1'b0 ;
  assign y12948 = ~n33206 ;
  assign y12949 = ~n33207 ;
  assign y12950 = ~n33212 ;
  assign y12951 = ~n15296 ;
  assign y12952 = ~1'b0 ;
  assign y12953 = n33215 ;
  assign y12954 = n33216 ;
  assign y12955 = n33218 ;
  assign y12956 = n33219 ;
  assign y12957 = n33221 ;
  assign y12958 = n33222 ;
  assign y12959 = ~n33223 ;
  assign y12960 = ~n33225 ;
  assign y12961 = n33228 ;
  assign y12962 = n33230 ;
  assign y12963 = ~n33232 ;
  assign y12964 = n9680 ;
  assign y12965 = ~n33233 ;
  assign y12966 = ~n33237 ;
  assign y12967 = ~n33238 ;
  assign y12968 = ~1'b0 ;
  assign y12969 = ~n33241 ;
  assign y12970 = n33246 ;
  assign y12971 = ~n33248 ;
  assign y12972 = ~1'b0 ;
  assign y12973 = n33251 ;
  assign y12974 = n33258 ;
  assign y12975 = ~1'b0 ;
  assign y12976 = ~1'b0 ;
  assign y12977 = n33261 ;
  assign y12978 = ~1'b0 ;
  assign y12979 = ~1'b0 ;
  assign y12980 = ~1'b0 ;
  assign y12981 = ~n33267 ;
  assign y12982 = ~n33268 ;
  assign y12983 = ~n33270 ;
  assign y12984 = n33273 ;
  assign y12985 = n33274 ;
  assign y12986 = ~1'b0 ;
  assign y12987 = n33276 ;
  assign y12988 = n33283 ;
  assign y12989 = ~n14224 ;
  assign y12990 = n33284 ;
  assign y12991 = ~n33285 ;
  assign y12992 = ~n33286 ;
  assign y12993 = n33291 ;
  assign y12994 = n33293 ;
  assign y12995 = n33299 ;
  assign y12996 = ~n33301 ;
  assign y12997 = ~n33302 ;
  assign y12998 = ~n33304 ;
  assign y12999 = ~n33311 ;
  assign y13000 = ~n33312 ;
  assign y13001 = ~n33316 ;
  assign y13002 = ~n33318 ;
  assign y13003 = n33321 ;
  assign y13004 = n33323 ;
  assign y13005 = ~n33328 ;
  assign y13006 = n33331 ;
  assign y13007 = n33334 ;
  assign y13008 = ~1'b0 ;
  assign y13009 = ~n33336 ;
  assign y13010 = n33340 ;
  assign y13011 = ~1'b0 ;
  assign y13012 = ~n33344 ;
  assign y13013 = ~1'b0 ;
  assign y13014 = ~n33349 ;
  assign y13015 = n33352 ;
  assign y13016 = n3452 ;
  assign y13017 = ~1'b0 ;
  assign y13018 = n33354 ;
  assign y13019 = ~n14063 ;
  assign y13020 = ~n33355 ;
  assign y13021 = n4326 ;
  assign y13022 = ~n33356 ;
  assign y13023 = n33358 ;
  assign y13024 = n33360 ;
  assign y13025 = ~1'b0 ;
  assign y13026 = ~1'b0 ;
  assign y13027 = ~1'b0 ;
  assign y13028 = n33364 ;
  assign y13029 = ~n33366 ;
  assign y13030 = ~n33367 ;
  assign y13031 = ~n33369 ;
  assign y13032 = ~1'b0 ;
  assign y13033 = ~1'b0 ;
  assign y13034 = ~1'b0 ;
  assign y13035 = n33373 ;
  assign y13036 = n33374 ;
  assign y13037 = n33376 ;
  assign y13038 = ~n33377 ;
  assign y13039 = ~n33379 ;
  assign y13040 = ~n33380 ;
  assign y13041 = n33385 ;
  assign y13042 = ~n33387 ;
  assign y13043 = ~n33389 ;
  assign y13044 = ~n33393 ;
  assign y13045 = n33395 ;
  assign y13046 = n33397 ;
  assign y13047 = ~n33400 ;
  assign y13048 = ~n33403 ;
  assign y13049 = ~n33405 ;
  assign y13050 = ~n33410 ;
  assign y13051 = n33411 ;
  assign y13052 = ~1'b0 ;
  assign y13053 = ~1'b0 ;
  assign y13054 = n33416 ;
  assign y13055 = ~n32659 ;
  assign y13056 = ~n33422 ;
  assign y13057 = n33425 ;
  assign y13058 = ~1'b0 ;
  assign y13059 = n33427 ;
  assign y13060 = ~n33432 ;
  assign y13061 = ~n33435 ;
  assign y13062 = ~n33436 ;
  assign y13063 = n33437 ;
  assign y13064 = ~n33439 ;
  assign y13065 = ~n33440 ;
  assign y13066 = ~n33443 ;
  assign y13067 = ~1'b0 ;
  assign y13068 = 1'b0 ;
  assign y13069 = n33452 ;
  assign y13070 = n33454 ;
  assign y13071 = n33457 ;
  assign y13072 = ~1'b0 ;
  assign y13073 = ~1'b0 ;
  assign y13074 = n33458 ;
  assign y13075 = ~n33459 ;
  assign y13076 = n33463 ;
  assign y13077 = n33465 ;
  assign y13078 = ~n33466 ;
  assign y13079 = n33471 ;
  assign y13080 = ~n33475 ;
  assign y13081 = n33477 ;
  assign y13082 = ~1'b0 ;
  assign y13083 = ~1'b0 ;
  assign y13084 = ~n33479 ;
  assign y13085 = ~n33480 ;
  assign y13086 = ~1'b0 ;
  assign y13087 = ~n33482 ;
  assign y13088 = ~n33507 ;
  assign y13089 = ~n33509 ;
  assign y13090 = n28096 ;
  assign y13091 = n33511 ;
  assign y13092 = n33515 ;
  assign y13093 = ~1'b0 ;
  assign y13094 = ~n33521 ;
  assign y13095 = ~1'b0 ;
  assign y13096 = ~n33523 ;
  assign y13097 = n33525 ;
  assign y13098 = n33526 ;
  assign y13099 = ~n33527 ;
  assign y13100 = ~n33528 ;
  assign y13101 = n33535 ;
  assign y13102 = n33537 ;
  assign y13103 = ~n29364 ;
  assign y13104 = ~n33539 ;
  assign y13105 = ~n33540 ;
  assign y13106 = n33544 ;
  assign y13107 = ~n33547 ;
  assign y13108 = ~1'b0 ;
  assign y13109 = ~n33548 ;
  assign y13110 = ~1'b0 ;
  assign y13111 = ~n33550 ;
  assign y13112 = ~1'b0 ;
  assign y13113 = ~n33554 ;
  assign y13114 = ~n33557 ;
  assign y13115 = n33558 ;
  assign y13116 = ~1'b0 ;
  assign y13117 = ~1'b0 ;
  assign y13118 = n33560 ;
  assign y13119 = n33567 ;
  assign y13120 = ~n33570 ;
  assign y13121 = n33571 ;
  assign y13122 = ~n33575 ;
  assign y13123 = ~n33576 ;
  assign y13124 = n28086 ;
  assign y13125 = ~n5047 ;
  assign y13126 = ~n33578 ;
  assign y13127 = ~1'b0 ;
  assign y13128 = ~n7382 ;
  assign y13129 = n33580 ;
  assign y13130 = ~1'b0 ;
  assign y13131 = ~n33583 ;
  assign y13132 = ~1'b0 ;
  assign y13133 = ~n33589 ;
  assign y13134 = n33595 ;
  assign y13135 = n33596 ;
  assign y13136 = ~n33604 ;
  assign y13137 = n33605 ;
  assign y13138 = ~n33607 ;
  assign y13139 = ~1'b0 ;
  assign y13140 = n33613 ;
  assign y13141 = ~n33616 ;
  assign y13142 = ~1'b0 ;
  assign y13143 = ~n33620 ;
  assign y13144 = ~n33621 ;
  assign y13145 = n33626 ;
  assign y13146 = n33630 ;
  assign y13147 = ~n33632 ;
  assign y13148 = ~1'b0 ;
  assign y13149 = n33634 ;
  assign y13150 = n33638 ;
  assign y13151 = n33639 ;
  assign y13152 = ~n33642 ;
  assign y13153 = n33645 ;
  assign y13154 = ~1'b0 ;
  assign y13155 = ~n33648 ;
  assign y13156 = n33649 ;
  assign y13157 = ~1'b0 ;
  assign y13158 = ~n31682 ;
  assign y13159 = ~n2993 ;
  assign y13160 = ~n33652 ;
  assign y13161 = n33656 ;
  assign y13162 = n33657 ;
  assign y13163 = n33658 ;
  assign y13164 = ~n33659 ;
  assign y13165 = ~n33665 ;
  assign y13166 = n33668 ;
  assign y13167 = ~n33672 ;
  assign y13168 = n33673 ;
  assign y13169 = ~n33675 ;
  assign y13170 = ~1'b0 ;
  assign y13171 = n33680 ;
  assign y13172 = n33682 ;
  assign y13173 = ~n33683 ;
  assign y13174 = n33684 ;
  assign y13175 = ~n33686 ;
  assign y13176 = ~n33687 ;
  assign y13177 = n33689 ;
  assign y13178 = ~1'b0 ;
  assign y13179 = ~n33692 ;
  assign y13180 = ~n33697 ;
  assign y13181 = ~1'b0 ;
  assign y13182 = n33699 ;
  assign y13183 = n33700 ;
  assign y13184 = ~1'b0 ;
  assign y13185 = ~n33702 ;
  assign y13186 = ~1'b0 ;
  assign y13187 = ~n33706 ;
  assign y13188 = ~1'b0 ;
  assign y13189 = ~n33708 ;
  assign y13190 = n33709 ;
  assign y13191 = n18597 ;
  assign y13192 = ~n33712 ;
  assign y13193 = ~1'b0 ;
  assign y13194 = ~n33718 ;
  assign y13195 = n33721 ;
  assign y13196 = n33722 ;
  assign y13197 = ~n33725 ;
  assign y13198 = ~n33733 ;
  assign y13199 = ~1'b0 ;
  assign y13200 = n33743 ;
  assign y13201 = ~n33747 ;
  assign y13202 = ~1'b0 ;
  assign y13203 = n33749 ;
  assign y13204 = n14465 ;
  assign y13205 = ~n33750 ;
  assign y13206 = ~n33752 ;
  assign y13207 = ~1'b0 ;
  assign y13208 = ~1'b0 ;
  assign y13209 = n33755 ;
  assign y13210 = ~1'b0 ;
  assign y13211 = ~1'b0 ;
  assign y13212 = ~1'b0 ;
  assign y13213 = ~n33757 ;
  assign y13214 = n19204 ;
  assign y13215 = n23929 ;
  assign y13216 = ~n33758 ;
  assign y13217 = ~n33760 ;
  assign y13218 = ~n33761 ;
  assign y13219 = ~n33764 ;
  assign y13220 = ~1'b0 ;
  assign y13221 = ~n33766 ;
  assign y13222 = n33769 ;
  assign y13223 = n33770 ;
  assign y13224 = n33772 ;
  assign y13225 = ~n33775 ;
  assign y13226 = ~n33782 ;
  assign y13227 = n33789 ;
  assign y13228 = ~n33791 ;
  assign y13229 = n33796 ;
  assign y13230 = n33798 ;
  assign y13231 = n33801 ;
  assign y13232 = n33802 ;
  assign y13233 = n33803 ;
  assign y13234 = ~n33808 ;
  assign y13235 = ~n21288 ;
  assign y13236 = n33815 ;
  assign y13237 = ~1'b0 ;
  assign y13238 = n33817 ;
  assign y13239 = ~n33819 ;
  assign y13240 = n33821 ;
  assign y13241 = ~n33823 ;
  assign y13242 = ~n33825 ;
  assign y13243 = ~n33827 ;
  assign y13244 = ~1'b0 ;
  assign y13245 = n33831 ;
  assign y13246 = n33832 ;
  assign y13247 = ~n33833 ;
  assign y13248 = ~n33836 ;
  assign y13249 = ~1'b0 ;
  assign y13250 = ~1'b0 ;
  assign y13251 = n33839 ;
  assign y13252 = ~1'b0 ;
  assign y13253 = ~1'b0 ;
  assign y13254 = ~n33841 ;
  assign y13255 = ~n33842 ;
  assign y13256 = ~n33851 ;
  assign y13257 = ~n33853 ;
  assign y13258 = ~n33858 ;
  assign y13259 = n586 ;
  assign y13260 = ~n33860 ;
  assign y13261 = ~n33863 ;
  assign y13262 = n33865 ;
  assign y13263 = ~n33867 ;
  assign y13264 = ~n33868 ;
  assign y13265 = ~n2841 ;
  assign y13266 = ~1'b0 ;
  assign y13267 = ~1'b0 ;
  assign y13268 = ~1'b0 ;
  assign y13269 = n33870 ;
  assign y13270 = n33871 ;
  assign y13271 = n33873 ;
  assign y13272 = ~n33874 ;
  assign y13273 = ~n33878 ;
  assign y13274 = ~n33879 ;
  assign y13275 = n33881 ;
  assign y13276 = n33882 ;
  assign y13277 = n33885 ;
  assign y13278 = 1'b0 ;
  assign y13279 = n33886 ;
  assign y13280 = ~1'b0 ;
  assign y13281 = ~1'b0 ;
  assign y13282 = ~n33888 ;
  assign y13283 = ~1'b0 ;
  assign y13284 = n33895 ;
  assign y13285 = n33899 ;
  assign y13286 = ~n33900 ;
  assign y13287 = ~n33902 ;
  assign y13288 = ~n33906 ;
  assign y13289 = n33908 ;
  assign y13290 = ~1'b0 ;
  assign y13291 = n33910 ;
  assign y13292 = ~n33913 ;
  assign y13293 = ~n33918 ;
  assign y13294 = ~n33920 ;
  assign y13295 = ~n33922 ;
  assign y13296 = ~1'b0 ;
  assign y13297 = ~1'b0 ;
  assign y13298 = ~1'b0 ;
  assign y13299 = ~n33923 ;
  assign y13300 = n33924 ;
  assign y13301 = n33930 ;
  assign y13302 = ~n33933 ;
  assign y13303 = ~n33936 ;
  assign y13304 = n33937 ;
  assign y13305 = ~n33939 ;
  assign y13306 = ~n22251 ;
  assign y13307 = ~1'b0 ;
  assign y13308 = n33940 ;
  assign y13309 = ~n33944 ;
  assign y13310 = ~1'b0 ;
  assign y13311 = n33948 ;
  assign y13312 = n33950 ;
  assign y13313 = n33953 ;
  assign y13314 = n33959 ;
  assign y13315 = n33961 ;
  assign y13316 = n33968 ;
  assign y13317 = n33970 ;
  assign y13318 = n33971 ;
  assign y13319 = n33973 ;
  assign y13320 = ~n33974 ;
  assign y13321 = n33975 ;
  assign y13322 = n33978 ;
  assign y13323 = n33979 ;
  assign y13324 = n33980 ;
  assign y13325 = n33981 ;
  assign y13326 = ~n33985 ;
  assign y13327 = n33988 ;
  assign y13328 = n33989 ;
  assign y13329 = ~n30201 ;
  assign y13330 = ~n33995 ;
  assign y13331 = 1'b0 ;
  assign y13332 = n33998 ;
  assign y13333 = ~n34001 ;
  assign y13334 = ~1'b0 ;
  assign y13335 = n34004 ;
  assign y13336 = n34006 ;
  assign y13337 = ~1'b0 ;
  assign y13338 = ~1'b0 ;
  assign y13339 = ~n34010 ;
  assign y13340 = ~1'b0 ;
  assign y13341 = ~n34012 ;
  assign y13342 = ~n34013 ;
  assign y13343 = ~n34015 ;
  assign y13344 = n34016 ;
  assign y13345 = n34026 ;
  assign y13346 = ~n34028 ;
  assign y13347 = ~n34029 ;
  assign y13348 = n34030 ;
  assign y13349 = n34033 ;
  assign y13350 = n34034 ;
  assign y13351 = ~n34036 ;
  assign y13352 = ~1'b0 ;
  assign y13353 = ~n34039 ;
  assign y13354 = n34040 ;
  assign y13355 = ~n34041 ;
  assign y13356 = ~1'b0 ;
  assign y13357 = ~n34042 ;
  assign y13358 = ~n34044 ;
  assign y13359 = ~n34045 ;
  assign y13360 = ~n34046 ;
  assign y13361 = ~n34048 ;
  assign y13362 = n34050 ;
  assign y13363 = ~1'b0 ;
  assign y13364 = n34059 ;
  assign y13365 = ~n34061 ;
  assign y13366 = n34064 ;
  assign y13367 = ~n34065 ;
  assign y13368 = n34066 ;
  assign y13369 = ~1'b0 ;
  assign y13370 = n34072 ;
  assign y13371 = n34079 ;
  assign y13372 = n34085 ;
  assign y13373 = ~n34092 ;
  assign y13374 = ~n34093 ;
  assign y13375 = ~n34098 ;
  assign y13376 = n34100 ;
  assign y13377 = n34104 ;
  assign y13378 = ~n34106 ;
  assign y13379 = ~n34111 ;
  assign y13380 = n34113 ;
  assign y13381 = n34116 ;
  assign y13382 = ~n34117 ;
  assign y13383 = ~n34121 ;
  assign y13384 = ~n34123 ;
  assign y13385 = n34125 ;
  assign y13386 = ~n34126 ;
  assign y13387 = ~n34133 ;
  assign y13388 = ~n34135 ;
  assign y13389 = ~n34138 ;
  assign y13390 = ~n34139 ;
  assign y13391 = ~1'b0 ;
  assign y13392 = n34140 ;
  assign y13393 = ~n34144 ;
  assign y13394 = ~n34148 ;
  assign y13395 = ~n34151 ;
  assign y13396 = ~n28439 ;
  assign y13397 = ~1'b0 ;
  assign y13398 = n34152 ;
  assign y13399 = n34155 ;
  assign y13400 = ~n34162 ;
  assign y13401 = n34165 ;
  assign y13402 = n34166 ;
  assign y13403 = ~n34178 ;
  assign y13404 = ~n34180 ;
  assign y13405 = ~1'b0 ;
  assign y13406 = ~1'b0 ;
  assign y13407 = ~1'b0 ;
  assign y13408 = ~1'b0 ;
  assign y13409 = n34181 ;
  assign y13410 = ~n34183 ;
  assign y13411 = ~n34188 ;
  assign y13412 = n34193 ;
  assign y13413 = ~n34203 ;
  assign y13414 = ~n34204 ;
  assign y13415 = ~1'b0 ;
  assign y13416 = n34208 ;
  assign y13417 = n34210 ;
  assign y13418 = ~n34215 ;
  assign y13419 = ~n4851 ;
  assign y13420 = ~n34221 ;
  assign y13421 = ~n34224 ;
  assign y13422 = n34226 ;
  assign y13423 = n34227 ;
  assign y13424 = ~n34230 ;
  assign y13425 = n15462 ;
  assign y13426 = ~n34231 ;
  assign y13427 = n34232 ;
  assign y13428 = ~n34233 ;
  assign y13429 = ~n34234 ;
  assign y13430 = n34242 ;
  assign y13431 = ~1'b0 ;
  assign y13432 = ~n34243 ;
  assign y13433 = ~1'b0 ;
  assign y13434 = n34244 ;
  assign y13435 = ~n34246 ;
  assign y13436 = ~1'b0 ;
  assign y13437 = n34249 ;
  assign y13438 = n34250 ;
  assign y13439 = ~n34256 ;
  assign y13440 = n34258 ;
  assign y13441 = ~n34261 ;
  assign y13442 = ~n34267 ;
  assign y13443 = n34274 ;
  assign y13444 = n34275 ;
  assign y13445 = ~n34276 ;
  assign y13446 = 1'b0 ;
  assign y13447 = n29073 ;
  assign y13448 = n34278 ;
  assign y13449 = n34280 ;
  assign y13450 = ~1'b0 ;
  assign y13451 = n34285 ;
  assign y13452 = ~n34288 ;
  assign y13453 = n34289 ;
  assign y13454 = 1'b0 ;
  assign y13455 = ~1'b0 ;
  assign y13456 = ~1'b0 ;
  assign y13457 = ~n34291 ;
  assign y13458 = n34294 ;
  assign y13459 = n34297 ;
  assign y13460 = ~1'b0 ;
  assign y13461 = ~n34304 ;
  assign y13462 = n34314 ;
  assign y13463 = n34316 ;
  assign y13464 = n34319 ;
  assign y13465 = ~1'b0 ;
  assign y13466 = ~n34324 ;
  assign y13467 = ~n34327 ;
  assign y13468 = ~1'b0 ;
  assign y13469 = n34329 ;
  assign y13470 = ~n34333 ;
  assign y13471 = n34340 ;
  assign y13472 = ~n34343 ;
  assign y13473 = ~n34347 ;
  assign y13474 = ~n34348 ;
  assign y13475 = ~1'b0 ;
  assign y13476 = ~n34350 ;
  assign y13477 = ~n34351 ;
  assign y13478 = n34353 ;
  assign y13479 = n34358 ;
  assign y13480 = ~n34359 ;
  assign y13481 = n34363 ;
  assign y13482 = n34367 ;
  assign y13483 = n34369 ;
  assign y13484 = n34370 ;
  assign y13485 = n19204 ;
  assign y13486 = ~n34372 ;
  assign y13487 = ~1'b0 ;
  assign y13488 = ~n34376 ;
  assign y13489 = ~n34377 ;
  assign y13490 = ~n34379 ;
  assign y13491 = n34380 ;
  assign y13492 = ~1'b0 ;
  assign y13493 = ~n34384 ;
  assign y13494 = n34386 ;
  assign y13495 = n34389 ;
  assign y13496 = ~1'b0 ;
  assign y13497 = ~n34392 ;
  assign y13498 = ~1'b0 ;
  assign y13499 = n34395 ;
  assign y13500 = ~n34399 ;
  assign y13501 = ~n34400 ;
  assign y13502 = ~n34401 ;
  assign y13503 = n34403 ;
  assign y13504 = ~1'b0 ;
  assign y13505 = n34409 ;
  assign y13506 = n22678 ;
  assign y13507 = n34412 ;
  assign y13508 = n34413 ;
  assign y13509 = n34415 ;
  assign y13510 = n34417 ;
  assign y13511 = n34418 ;
  assign y13512 = ~n34419 ;
  assign y13513 = ~n34421 ;
  assign y13514 = ~1'b0 ;
  assign y13515 = n34422 ;
  assign y13516 = n34427 ;
  assign y13517 = ~n34430 ;
  assign y13518 = ~1'b0 ;
  assign y13519 = ~n34431 ;
  assign y13520 = ~n34432 ;
  assign y13521 = ~n34434 ;
  assign y13522 = ~1'b0 ;
  assign y13523 = n34436 ;
  assign y13524 = ~1'b0 ;
  assign y13525 = ~1'b0 ;
  assign y13526 = n34440 ;
  assign y13527 = ~n34444 ;
  assign y13528 = ~n34445 ;
  assign y13529 = ~n34446 ;
  assign y13530 = n34448 ;
  assign y13531 = n34450 ;
  assign y13532 = 1'b0 ;
  assign y13533 = 1'b0 ;
  assign y13534 = ~n17301 ;
  assign y13535 = n34451 ;
  assign y13536 = ~n34453 ;
  assign y13537 = ~n34456 ;
  assign y13538 = ~1'b0 ;
  assign y13539 = n34457 ;
  assign y13540 = ~n34460 ;
  assign y13541 = n34463 ;
  assign y13542 = n34464 ;
  assign y13543 = n34467 ;
  assign y13544 = ~1'b0 ;
  assign y13545 = ~n34471 ;
  assign y13546 = ~n34472 ;
  assign y13547 = n34482 ;
  assign y13548 = ~n34483 ;
  assign y13549 = n34485 ;
  assign y13550 = ~1'b0 ;
  assign y13551 = n34486 ;
  assign y13552 = n34490 ;
  assign y13553 = ~1'b0 ;
  assign y13554 = ~1'b0 ;
  assign y13555 = n34492 ;
  assign y13556 = n34497 ;
  assign y13557 = ~n6627 ;
  assign y13558 = n34498 ;
  assign y13559 = ~n34501 ;
  assign y13560 = ~1'b0 ;
  assign y13561 = ~n34504 ;
  assign y13562 = n34505 ;
  assign y13563 = n34506 ;
  assign y13564 = ~n34509 ;
  assign y13565 = ~n34511 ;
  assign y13566 = ~1'b0 ;
  assign y13567 = n34513 ;
  assign y13568 = n4993 ;
  assign y13569 = ~n34514 ;
  assign y13570 = ~n34516 ;
  assign y13571 = ~n34518 ;
  assign y13572 = ~1'b0 ;
  assign y13573 = ~1'b0 ;
  assign y13574 = ~1'b0 ;
  assign y13575 = ~n34522 ;
  assign y13576 = n34526 ;
  assign y13577 = ~n34531 ;
  assign y13578 = n34532 ;
  assign y13579 = n34534 ;
  assign y13580 = ~n34535 ;
  assign y13581 = n34537 ;
  assign y13582 = n34541 ;
  assign y13583 = ~n34551 ;
  assign y13584 = ~n34554 ;
  assign y13585 = ~n34556 ;
  assign y13586 = 1'b0 ;
  assign y13587 = ~n34557 ;
  assign y13588 = n34561 ;
  assign y13589 = ~n34564 ;
  assign y13590 = ~n34567 ;
  assign y13591 = n34568 ;
  assign y13592 = ~n34572 ;
  assign y13593 = ~1'b0 ;
  assign y13594 = ~1'b0 ;
  assign y13595 = ~1'b0 ;
  assign y13596 = ~n34573 ;
  assign y13597 = n34576 ;
  assign y13598 = n34579 ;
  assign y13599 = ~n34580 ;
  assign y13600 = ~1'b0 ;
  assign y13601 = ~1'b0 ;
  assign y13602 = ~1'b0 ;
  assign y13603 = ~n34581 ;
  assign y13604 = n34582 ;
  assign y13605 = ~n34583 ;
  assign y13606 = ~n34584 ;
  assign y13607 = ~n34585 ;
  assign y13608 = ~n34587 ;
  assign y13609 = n34591 ;
  assign y13610 = n34593 ;
  assign y13611 = ~n34595 ;
  assign y13612 = ~n34600 ;
  assign y13613 = ~n34608 ;
  assign y13614 = ~1'b0 ;
  assign y13615 = ~1'b0 ;
  assign y13616 = n34609 ;
  assign y13617 = ~1'b0 ;
  assign y13618 = n34610 ;
  assign y13619 = ~n34614 ;
  assign y13620 = ~n34620 ;
  assign y13621 = ~n34622 ;
  assign y13622 = 1'b0 ;
  assign y13623 = ~1'b0 ;
  assign y13624 = n34625 ;
  assign y13625 = ~n34626 ;
  assign y13626 = n34627 ;
  assign y13627 = n34630 ;
  assign y13628 = ~1'b0 ;
  assign y13629 = n34631 ;
  assign y13630 = ~n12458 ;
  assign y13631 = n34633 ;
  assign y13632 = n34634 ;
  assign y13633 = ~1'b0 ;
  assign y13634 = ~1'b0 ;
  assign y13635 = ~n34636 ;
  assign y13636 = ~n34638 ;
  assign y13637 = 1'b0 ;
  assign y13638 = ~1'b0 ;
  assign y13639 = ~n34647 ;
  assign y13640 = ~n34651 ;
  assign y13641 = ~n34653 ;
  assign y13642 = ~1'b0 ;
  assign y13643 = ~n34656 ;
  assign y13644 = n34664 ;
  assign y13645 = ~n34668 ;
  assign y13646 = n34669 ;
  assign y13647 = n34670 ;
  assign y13648 = n34673 ;
  assign y13649 = n34674 ;
  assign y13650 = ~1'b0 ;
  assign y13651 = ~n34676 ;
  assign y13652 = n34677 ;
  assign y13653 = ~1'b0 ;
  assign y13654 = 1'b0 ;
  assign y13655 = n34683 ;
  assign y13656 = n34684 ;
  assign y13657 = 1'b0 ;
  assign y13658 = ~1'b0 ;
  assign y13659 = n34686 ;
  assign y13660 = ~n34689 ;
  assign y13661 = n34691 ;
  assign y13662 = n34694 ;
  assign y13663 = ~n34696 ;
  assign y13664 = ~1'b0 ;
  assign y13665 = n34697 ;
  assign y13666 = ~1'b0 ;
  assign y13667 = ~n34698 ;
  assign y13668 = n34699 ;
  assign y13669 = ~n24862 ;
  assign y13670 = ~n34702 ;
  assign y13671 = n34703 ;
  assign y13672 = ~n34707 ;
  assign y13673 = ~n34710 ;
  assign y13674 = n34712 ;
  assign y13675 = ~n34713 ;
  assign y13676 = n34715 ;
  assign y13677 = n34717 ;
  assign y13678 = ~n34718 ;
  assign y13679 = n34721 ;
  assign y13680 = ~n34724 ;
  assign y13681 = ~1'b0 ;
  assign y13682 = ~1'b0 ;
  assign y13683 = ~1'b0 ;
  assign y13684 = n34725 ;
  assign y13685 = ~n34726 ;
  assign y13686 = ~1'b0 ;
  assign y13687 = n34727 ;
  assign y13688 = n15721 ;
  assign y13689 = ~n34728 ;
  assign y13690 = n34733 ;
  assign y13691 = ~n24506 ;
  assign y13692 = ~1'b0 ;
  assign y13693 = n34737 ;
  assign y13694 = ~n26134 ;
  assign y13695 = n34740 ;
  assign y13696 = ~n34741 ;
  assign y13697 = ~n33242 ;
  assign y13698 = n34745 ;
  assign y13699 = n34749 ;
  assign y13700 = n34756 ;
  assign y13701 = ~1'b0 ;
  assign y13702 = n34758 ;
  assign y13703 = ~n34760 ;
  assign y13704 = ~n34761 ;
  assign y13705 = ~n34763 ;
  assign y13706 = n34765 ;
  assign y13707 = ~1'b0 ;
  assign y13708 = ~1'b0 ;
  assign y13709 = n34769 ;
  assign y13710 = n34770 ;
  assign y13711 = ~n34771 ;
  assign y13712 = ~1'b0 ;
  assign y13713 = ~n34772 ;
  assign y13714 = ~1'b0 ;
  assign y13715 = ~1'b0 ;
  assign y13716 = ~n34775 ;
  assign y13717 = ~n34778 ;
  assign y13718 = ~n34779 ;
  assign y13719 = ~n34780 ;
  assign y13720 = n34781 ;
  assign y13721 = n34787 ;
  assign y13722 = n34789 ;
  assign y13723 = n34793 ;
  assign y13724 = ~1'b0 ;
  assign y13725 = n34797 ;
  assign y13726 = n34801 ;
  assign y13727 = n34804 ;
  assign y13728 = ~n34805 ;
  assign y13729 = ~1'b0 ;
  assign y13730 = n34807 ;
  assign y13731 = ~1'b0 ;
  assign y13732 = ~n34808 ;
  assign y13733 = ~n34810 ;
  assign y13734 = n34812 ;
  assign y13735 = ~n34815 ;
  assign y13736 = ~n34816 ;
  assign y13737 = n34817 ;
  assign y13738 = n34819 ;
  assign y13739 = n34820 ;
  assign y13740 = ~1'b0 ;
  assign y13741 = n34822 ;
  assign y13742 = ~1'b0 ;
  assign y13743 = ~n34823 ;
  assign y13744 = ~n34824 ;
  assign y13745 = ~1'b0 ;
  assign y13746 = ~n34825 ;
  assign y13747 = ~n34826 ;
  assign y13748 = ~1'b0 ;
  assign y13749 = ~n34828 ;
  assign y13750 = ~n34829 ;
  assign y13751 = ~n34839 ;
  assign y13752 = ~n34840 ;
  assign y13753 = n34842 ;
  assign y13754 = ~n34845 ;
  assign y13755 = n34846 ;
  assign y13756 = ~1'b0 ;
  assign y13757 = n34848 ;
  assign y13758 = ~1'b0 ;
  assign y13759 = ~1'b0 ;
  assign y13760 = n4220 ;
  assign y13761 = ~n34849 ;
  assign y13762 = ~n34850 ;
  assign y13763 = ~n34855 ;
  assign y13764 = ~1'b0 ;
  assign y13765 = ~1'b0 ;
  assign y13766 = 1'b0 ;
  assign y13767 = ~n34857 ;
  assign y13768 = n34860 ;
  assign y13769 = n34865 ;
  assign y13770 = n34871 ;
  assign y13771 = n34872 ;
  assign y13772 = ~1'b0 ;
  assign y13773 = ~n34874 ;
  assign y13774 = ~1'b0 ;
  assign y13775 = ~1'b0 ;
  assign y13776 = ~n34878 ;
  assign y13777 = n34880 ;
  assign y13778 = n34884 ;
  assign y13779 = ~n34888 ;
  assign y13780 = ~n34897 ;
  assign y13781 = ~1'b0 ;
  assign y13782 = ~n34898 ;
  assign y13783 = ~n32593 ;
  assign y13784 = n34899 ;
  assign y13785 = ~n34902 ;
  assign y13786 = ~1'b0 ;
  assign y13787 = n34904 ;
  assign y13788 = ~n5095 ;
  assign y13789 = n7450 ;
  assign y13790 = n34917 ;
  assign y13791 = ~n34918 ;
  assign y13792 = 1'b0 ;
  assign y13793 = ~n34919 ;
  assign y13794 = ~1'b0 ;
  assign y13795 = ~n34921 ;
  assign y13796 = ~n34924 ;
  assign y13797 = ~n34927 ;
  assign y13798 = ~n34928 ;
  assign y13799 = ~n34931 ;
  assign y13800 = ~n34933 ;
  assign y13801 = ~n34934 ;
  assign y13802 = ~n34936 ;
  assign y13803 = n34938 ;
  assign y13804 = n34940 ;
  assign y13805 = ~n34946 ;
  assign y13806 = ~1'b0 ;
  assign y13807 = ~1'b0 ;
  assign y13808 = ~n34950 ;
  assign y13809 = n34951 ;
  assign y13810 = ~n34956 ;
  assign y13811 = ~n34957 ;
  assign y13812 = ~1'b0 ;
  assign y13813 = ~1'b0 ;
  assign y13814 = n34959 ;
  assign y13815 = 1'b0 ;
  assign y13816 = ~n34964 ;
  assign y13817 = n34966 ;
  assign y13818 = n34969 ;
  assign y13819 = ~n34970 ;
  assign y13820 = ~n34972 ;
  assign y13821 = ~n34974 ;
  assign y13822 = ~n34980 ;
  assign y13823 = n34984 ;
  assign y13824 = ~n34985 ;
  assign y13825 = ~n12779 ;
  assign y13826 = ~n34986 ;
  assign y13827 = ~n34987 ;
  assign y13828 = ~n21122 ;
  assign y13829 = 1'b0 ;
  assign y13830 = ~n34990 ;
  assign y13831 = ~1'b0 ;
  assign y13832 = n34992 ;
  assign y13833 = n34994 ;
  assign y13834 = ~n35002 ;
  assign y13835 = n35004 ;
  assign y13836 = ~n2009 ;
  assign y13837 = n35007 ;
  assign y13838 = ~1'b0 ;
  assign y13839 = n35009 ;
  assign y13840 = ~n35020 ;
  assign y13841 = ~n35022 ;
  assign y13842 = ~1'b0 ;
  assign y13843 = ~n35029 ;
  assign y13844 = ~n35031 ;
  assign y13845 = ~n35032 ;
  assign y13846 = n35033 ;
  assign y13847 = ~n35039 ;
  assign y13848 = n35043 ;
  assign y13849 = ~n35044 ;
  assign y13850 = n35050 ;
  assign y13851 = n35052 ;
  assign y13852 = n35055 ;
  assign y13853 = n35057 ;
  assign y13854 = n35060 ;
  assign y13855 = ~n13348 ;
  assign y13856 = ~n35062 ;
  assign y13857 = ~n35063 ;
  assign y13858 = ~1'b0 ;
  assign y13859 = n35067 ;
  assign y13860 = ~n35068 ;
  assign y13861 = n35071 ;
  assign y13862 = n35078 ;
  assign y13863 = n35080 ;
  assign y13864 = ~n35082 ;
  assign y13865 = n35084 ;
  assign y13866 = ~1'b0 ;
  assign y13867 = ~n35086 ;
  assign y13868 = ~1'b0 ;
  assign y13869 = n35088 ;
  assign y13870 = n35089 ;
  assign y13871 = ~n35090 ;
  assign y13872 = n35094 ;
  assign y13873 = n35098 ;
  assign y13874 = n35100 ;
  assign y13875 = ~1'b0 ;
  assign y13876 = n35102 ;
  assign y13877 = n35105 ;
  assign y13878 = ~n35107 ;
  assign y13879 = n35108 ;
  assign y13880 = n35109 ;
  assign y13881 = ~n35111 ;
  assign y13882 = ~1'b0 ;
  assign y13883 = ~n35120 ;
  assign y13884 = ~1'b0 ;
  assign y13885 = ~n35122 ;
  assign y13886 = ~n35123 ;
  assign y13887 = ~n35125 ;
  assign y13888 = ~n35128 ;
  assign y13889 = ~1'b0 ;
  assign y13890 = ~n35132 ;
  assign y13891 = n35133 ;
  assign y13892 = ~1'b0 ;
  assign y13893 = ~n35137 ;
  assign y13894 = ~n35140 ;
  assign y13895 = ~n35143 ;
  assign y13896 = ~n35146 ;
  assign y13897 = ~1'b0 ;
  assign y13898 = ~n35153 ;
  assign y13899 = ~n35156 ;
  assign y13900 = n35159 ;
  assign y13901 = n35161 ;
  assign y13902 = ~n35162 ;
  assign y13903 = n35168 ;
  assign y13904 = n22186 ;
  assign y13905 = n35172 ;
  assign y13906 = ~n35178 ;
  assign y13907 = ~n35183 ;
  assign y13908 = ~1'b0 ;
  assign y13909 = n35189 ;
  assign y13910 = n35193 ;
  assign y13911 = ~n35195 ;
  assign y13912 = ~1'b0 ;
  assign y13913 = n35198 ;
  assign y13914 = n35203 ;
  assign y13915 = ~n35213 ;
  assign y13916 = n35214 ;
  assign y13917 = n35217 ;
  assign y13918 = ~1'b0 ;
  assign y13919 = ~n35220 ;
  assign y13920 = n35224 ;
  assign y13921 = n35226 ;
  assign y13922 = n35227 ;
  assign y13923 = ~n35228 ;
  assign y13924 = ~1'b0 ;
  assign y13925 = n35232 ;
  assign y13926 = n28502 ;
  assign y13927 = ~n35235 ;
  assign y13928 = n35236 ;
  assign y13929 = ~n26614 ;
  assign y13930 = ~1'b0 ;
  assign y13931 = n35238 ;
  assign y13932 = ~1'b0 ;
  assign y13933 = n35241 ;
  assign y13934 = ~n35242 ;
  assign y13935 = n35244 ;
  assign y13936 = ~n35247 ;
  assign y13937 = ~n35251 ;
  assign y13938 = n35258 ;
  assign y13939 = n35259 ;
  assign y13940 = ~1'b0 ;
  assign y13941 = ~1'b0 ;
  assign y13942 = n35262 ;
  assign y13943 = n35267 ;
  assign y13944 = n35268 ;
  assign y13945 = n35275 ;
  assign y13946 = ~n35277 ;
  assign y13947 = ~n35279 ;
  assign y13948 = ~1'b0 ;
  assign y13949 = ~n35283 ;
  assign y13950 = ~n35285 ;
  assign y13951 = ~n35289 ;
  assign y13952 = n35291 ;
  assign y13953 = n35292 ;
  assign y13954 = ~n35293 ;
  assign y13955 = ~1'b0 ;
  assign y13956 = ~1'b0 ;
  assign y13957 = n35296 ;
  assign y13958 = ~1'b0 ;
  assign y13959 = ~1'b0 ;
  assign y13960 = 1'b0 ;
  assign y13961 = ~n35302 ;
  assign y13962 = ~n35303 ;
  assign y13963 = ~n35304 ;
  assign y13964 = ~n35306 ;
  assign y13965 = n35308 ;
  assign y13966 = n35313 ;
  assign y13967 = ~n8839 ;
  assign y13968 = ~1'b0 ;
  assign y13969 = 1'b0 ;
  assign y13970 = ~n35315 ;
  assign y13971 = n35321 ;
  assign y13972 = n35322 ;
  assign y13973 = n35325 ;
  assign y13974 = n35332 ;
  assign y13975 = n35336 ;
  assign y13976 = n35344 ;
  assign y13977 = n35346 ;
  assign y13978 = ~n35350 ;
  assign y13979 = n35351 ;
  assign y13980 = ~1'b0 ;
  assign y13981 = ~n35355 ;
  assign y13982 = ~n35357 ;
  assign y13983 = ~n35361 ;
  assign y13984 = ~n35363 ;
  assign y13985 = n35364 ;
  assign y13986 = n35367 ;
  assign y13987 = n35373 ;
  assign y13988 = n35378 ;
  assign y13989 = n35380 ;
  assign y13990 = ~n35381 ;
  assign y13991 = n35383 ;
  assign y13992 = ~n35385 ;
  assign y13993 = ~n35387 ;
  assign y13994 = ~n35388 ;
  assign y13995 = n35390 ;
  assign y13996 = n35391 ;
  assign y13997 = ~n35397 ;
  assign y13998 = ~1'b0 ;
  assign y13999 = n35398 ;
  assign y14000 = ~n35399 ;
  assign y14001 = ~n35401 ;
  assign y14002 = ~n35402 ;
  assign y14003 = n35404 ;
  assign y14004 = ~n35407 ;
  assign y14005 = ~1'b0 ;
  assign y14006 = n35408 ;
  assign y14007 = ~n35412 ;
  assign y14008 = n35413 ;
  assign y14009 = ~1'b0 ;
  assign y14010 = n35414 ;
  assign y14011 = ~n35417 ;
  assign y14012 = ~n35419 ;
  assign y14013 = ~1'b0 ;
  assign y14014 = n35420 ;
  assign y14015 = n35422 ;
  assign y14016 = n35428 ;
  assign y14017 = n35430 ;
  assign y14018 = n35432 ;
  assign y14019 = ~1'b0 ;
  assign y14020 = n35436 ;
  assign y14021 = ~1'b0 ;
  assign y14022 = n35438 ;
  assign y14023 = n35439 ;
  assign y14024 = n35441 ;
  assign y14025 = n35445 ;
  assign y14026 = ~1'b0 ;
  assign y14027 = n35448 ;
  assign y14028 = n35449 ;
  assign y14029 = ~n35452 ;
  assign y14030 = n35456 ;
  assign y14031 = ~n35461 ;
  assign y14032 = n35463 ;
  assign y14033 = n35465 ;
  assign y14034 = n35471 ;
  assign y14035 = n35475 ;
  assign y14036 = ~1'b0 ;
  assign y14037 = n35480 ;
  assign y14038 = n35482 ;
  assign y14039 = ~n35484 ;
  assign y14040 = ~1'b0 ;
  assign y14041 = ~n35486 ;
  assign y14042 = ~n35487 ;
  assign y14043 = n35488 ;
  assign y14044 = n35492 ;
  assign y14045 = n35495 ;
  assign y14046 = n11167 ;
  assign y14047 = ~1'b0 ;
  assign y14048 = n35500 ;
  assign y14049 = ~n35505 ;
  assign y14050 = ~n35509 ;
  assign y14051 = n35511 ;
  assign y14052 = n35518 ;
  assign y14053 = ~n35520 ;
  assign y14054 = ~1'b0 ;
  assign y14055 = n35523 ;
  assign y14056 = ~n35528 ;
  assign y14057 = ~n35531 ;
  assign y14058 = ~n35532 ;
  assign y14059 = ~n35534 ;
  assign y14060 = n35535 ;
  assign y14061 = n35537 ;
  assign y14062 = ~n35539 ;
  assign y14063 = n35541 ;
  assign y14064 = ~n35545 ;
  assign y14065 = ~1'b0 ;
  assign y14066 = n35546 ;
  assign y14067 = n35550 ;
  assign y14068 = n35551 ;
  assign y14069 = n35552 ;
  assign y14070 = ~n35554 ;
  assign y14071 = ~n35564 ;
  assign y14072 = n35565 ;
  assign y14073 = n35566 ;
  assign y14074 = 1'b0 ;
  assign y14075 = ~n35567 ;
  assign y14076 = n35569 ;
  assign y14077 = ~1'b0 ;
  assign y14078 = ~n35572 ;
  assign y14079 = ~n35574 ;
  assign y14080 = n35578 ;
  assign y14081 = ~1'b0 ;
  assign y14082 = n35581 ;
  assign y14083 = ~n35583 ;
  assign y14084 = ~n35584 ;
  assign y14085 = ~n35586 ;
  assign y14086 = ~n35590 ;
  assign y14087 = ~n35592 ;
  assign y14088 = n35596 ;
  assign y14089 = ~1'b0 ;
  assign y14090 = ~n35597 ;
  assign y14091 = n35599 ;
  assign y14092 = ~n35601 ;
  assign y14093 = ~n35602 ;
  assign y14094 = n35603 ;
  assign y14095 = ~1'b0 ;
  assign y14096 = ~n35606 ;
  assign y14097 = ~n35608 ;
  assign y14098 = n35609 ;
  assign y14099 = n35611 ;
  assign y14100 = n35613 ;
  assign y14101 = ~n35614 ;
  assign y14102 = n35615 ;
  assign y14103 = ~n35618 ;
  assign y14104 = n35620 ;
  assign y14105 = ~1'b0 ;
  assign y14106 = n35623 ;
  assign y14107 = ~n35628 ;
  assign y14108 = ~1'b0 ;
  assign y14109 = ~n35630 ;
  assign y14110 = n35631 ;
  assign y14111 = ~n35635 ;
  assign y14112 = n35638 ;
  assign y14113 = ~n35639 ;
  assign y14114 = ~1'b0 ;
  assign y14115 = n35640 ;
  assign y14116 = ~n35643 ;
  assign y14117 = ~n35652 ;
  assign y14118 = n35653 ;
  assign y14119 = ~n35656 ;
  assign y14120 = ~n35659 ;
  assign y14121 = n35660 ;
  assign y14122 = ~n35664 ;
  assign y14123 = ~1'b0 ;
  assign y14124 = ~n35666 ;
  assign y14125 = ~n35671 ;
  assign y14126 = n35673 ;
  assign y14127 = ~n35675 ;
  assign y14128 = n35677 ;
  assign y14129 = n35679 ;
  assign y14130 = n35682 ;
  assign y14131 = ~n35684 ;
  assign y14132 = n35686 ;
  assign y14133 = ~1'b0 ;
  assign y14134 = n35687 ;
  assign y14135 = n35692 ;
  assign y14136 = ~1'b0 ;
  assign y14137 = n35694 ;
  assign y14138 = n35697 ;
  assign y14139 = ~n35698 ;
  assign y14140 = n35702 ;
  assign y14141 = n903 ;
  assign y14142 = ~n35704 ;
  assign y14143 = ~1'b0 ;
  assign y14144 = ~n35706 ;
  assign y14145 = ~1'b0 ;
  assign y14146 = ~n35711 ;
  assign y14147 = n35712 ;
  assign y14148 = n35717 ;
  assign y14149 = ~n35720 ;
  assign y14150 = ~1'b0 ;
  assign y14151 = n35728 ;
  assign y14152 = ~1'b0 ;
  assign y14153 = ~n35730 ;
  assign y14154 = ~n35731 ;
  assign y14155 = ~n35733 ;
  assign y14156 = ~1'b0 ;
  assign y14157 = n35737 ;
  assign y14158 = ~1'b0 ;
  assign y14159 = n35738 ;
  assign y14160 = ~n35739 ;
  assign y14161 = n6719 ;
  assign y14162 = ~1'b0 ;
  assign y14163 = n35740 ;
  assign y14164 = n35741 ;
  assign y14165 = n11510 ;
  assign y14166 = n35743 ;
  assign y14167 = ~n35745 ;
  assign y14168 = ~n35749 ;
  assign y14169 = ~n35750 ;
  assign y14170 = ~n35752 ;
  assign y14171 = ~n35753 ;
  assign y14172 = ~1'b0 ;
  assign y14173 = n35759 ;
  assign y14174 = ~n35760 ;
  assign y14175 = ~n35761 ;
  assign y14176 = ~n35762 ;
  assign y14177 = ~1'b0 ;
  assign y14178 = n35765 ;
  assign y14179 = 1'b0 ;
  assign y14180 = n35768 ;
  assign y14181 = n35773 ;
  assign y14182 = n35779 ;
  assign y14183 = ~n35780 ;
  assign y14184 = ~n35784 ;
  assign y14185 = n35786 ;
  assign y14186 = ~n35787 ;
  assign y14187 = ~n35789 ;
  assign y14188 = n35790 ;
  assign y14189 = ~1'b0 ;
  assign y14190 = n35792 ;
  assign y14191 = n35793 ;
  assign y14192 = ~1'b0 ;
  assign y14193 = n35795 ;
  assign y14194 = ~n35798 ;
  assign y14195 = ~n35803 ;
  assign y14196 = n35805 ;
  assign y14197 = ~1'b0 ;
  assign y14198 = ~1'b0 ;
  assign y14199 = n35806 ;
  assign y14200 = n35810 ;
  assign y14201 = n35814 ;
  assign y14202 = ~n35815 ;
  assign y14203 = ~n35817 ;
  assign y14204 = ~1'b0 ;
  assign y14205 = n35820 ;
  assign y14206 = ~n35822 ;
  assign y14207 = n35826 ;
  assign y14208 = ~n35828 ;
  assign y14209 = ~n35833 ;
  assign y14210 = ~n35835 ;
  assign y14211 = ~n35836 ;
  assign y14212 = ~n27776 ;
  assign y14213 = ~n35838 ;
  assign y14214 = ~n35840 ;
  assign y14215 = ~n35843 ;
  assign y14216 = ~n35844 ;
  assign y14217 = ~n35845 ;
  assign y14218 = ~1'b0 ;
  assign y14219 = ~1'b0 ;
  assign y14220 = ~1'b0 ;
  assign y14221 = ~n35851 ;
  assign y14222 = n35856 ;
  assign y14223 = n35861 ;
  assign y14224 = ~n35862 ;
  assign y14225 = ~n35868 ;
  assign y14226 = ~1'b0 ;
  assign y14227 = ~1'b0 ;
  assign y14228 = ~1'b0 ;
  assign y14229 = n35869 ;
  assign y14230 = n14836 ;
  assign y14231 = ~1'b0 ;
  assign y14232 = n35870 ;
  assign y14233 = ~n35873 ;
  assign y14234 = n35876 ;
  assign y14235 = n35881 ;
  assign y14236 = ~n35888 ;
  assign y14237 = n35889 ;
  assign y14238 = ~n35897 ;
  assign y14239 = n35902 ;
  assign y14240 = ~n35904 ;
  assign y14241 = n35907 ;
  assign y14242 = ~1'b0 ;
  assign y14243 = ~1'b0 ;
  assign y14244 = ~1'b0 ;
  assign y14245 = ~n35911 ;
  assign y14246 = n35913 ;
  assign y14247 = ~n35914 ;
  assign y14248 = n35916 ;
  assign y14249 = n35921 ;
  assign y14250 = ~n35925 ;
  assign y14251 = ~1'b0 ;
  assign y14252 = ~1'b0 ;
  assign y14253 = n35926 ;
  assign y14254 = n35927 ;
  assign y14255 = ~n35929 ;
  assign y14256 = n30022 ;
  assign y14257 = ~n35931 ;
  assign y14258 = n35937 ;
  assign y14259 = ~n35940 ;
  assign y14260 = n35942 ;
  assign y14261 = n35943 ;
  assign y14262 = n35945 ;
  assign y14263 = ~1'b0 ;
  assign y14264 = 1'b0 ;
  assign y14265 = ~1'b0 ;
  assign y14266 = n35947 ;
  assign y14267 = n35948 ;
  assign y14268 = ~n35949 ;
  assign y14269 = n35952 ;
  assign y14270 = n35955 ;
  assign y14271 = n35958 ;
  assign y14272 = n35963 ;
  assign y14273 = ~n35968 ;
  assign y14274 = ~n35969 ;
  assign y14275 = ~n35974 ;
  assign y14276 = n35981 ;
  assign y14277 = n35983 ;
  assign y14278 = ~n35985 ;
  assign y14279 = ~1'b0 ;
  assign y14280 = ~n35992 ;
  assign y14281 = ~1'b0 ;
  assign y14282 = ~n35997 ;
  assign y14283 = ~n35998 ;
  assign y14284 = ~n35999 ;
  assign y14285 = n36001 ;
  assign y14286 = n36009 ;
  assign y14287 = ~n36010 ;
  assign y14288 = ~1'b0 ;
  assign y14289 = ~n36014 ;
  assign y14290 = n31456 ;
  assign y14291 = ~n36016 ;
  assign y14292 = ~1'b0 ;
  assign y14293 = ~n36022 ;
  assign y14294 = ~n36026 ;
  assign y14295 = ~n36027 ;
  assign y14296 = ~n36029 ;
  assign y14297 = ~n36043 ;
  assign y14298 = ~n36044 ;
  assign y14299 = ~1'b0 ;
  assign y14300 = ~1'b0 ;
  assign y14301 = ~n36046 ;
  assign y14302 = n36049 ;
  assign y14303 = ~n36050 ;
  assign y14304 = n36053 ;
  assign y14305 = ~n11013 ;
  assign y14306 = n36054 ;
  assign y14307 = ~1'b0 ;
  assign y14308 = ~1'b0 ;
  assign y14309 = ~n36055 ;
  assign y14310 = ~n36059 ;
  assign y14311 = ~n36060 ;
  assign y14312 = ~n36063 ;
  assign y14313 = ~n36065 ;
  assign y14314 = ~n36068 ;
  assign y14315 = ~n36072 ;
  assign y14316 = n36073 ;
  assign y14317 = ~1'b0 ;
  assign y14318 = n36075 ;
  assign y14319 = ~n36078 ;
  assign y14320 = ~1'b0 ;
  assign y14321 = n36080 ;
  assign y14322 = ~n36081 ;
  assign y14323 = ~n36083 ;
  assign y14324 = ~1'b0 ;
  assign y14325 = ~1'b0 ;
  assign y14326 = ~1'b0 ;
  assign y14327 = ~n36084 ;
  assign y14328 = ~n36086 ;
  assign y14329 = ~1'b0 ;
  assign y14330 = ~n36090 ;
  assign y14331 = n36094 ;
  assign y14332 = n36095 ;
  assign y14333 = ~n36098 ;
  assign y14334 = n36100 ;
  assign y14335 = ~n36104 ;
  assign y14336 = ~n36106 ;
  assign y14337 = n36107 ;
  assign y14338 = ~n36108 ;
  assign y14339 = ~n36109 ;
  assign y14340 = ~n36110 ;
  assign y14341 = n36112 ;
  assign y14342 = n36118 ;
  assign y14343 = ~1'b0 ;
  assign y14344 = ~n36121 ;
  assign y14345 = n36123 ;
  assign y14346 = ~n36131 ;
  assign y14347 = ~n36133 ;
  assign y14348 = n36137 ;
  assign y14349 = ~1'b0 ;
  assign y14350 = ~n36138 ;
  assign y14351 = ~n36144 ;
  assign y14352 = ~1'b0 ;
  assign y14353 = ~n36146 ;
  assign y14354 = ~n36148 ;
  assign y14355 = n36149 ;
  assign y14356 = n36156 ;
  assign y14357 = ~n33256 ;
  assign y14358 = ~n36161 ;
  assign y14359 = n36163 ;
  assign y14360 = n36166 ;
  assign y14361 = ~n22346 ;
  assign y14362 = ~n36171 ;
  assign y14363 = n36173 ;
  assign y14364 = ~n36176 ;
  assign y14365 = ~n36177 ;
  assign y14366 = ~1'b0 ;
  assign y14367 = ~n36180 ;
  assign y14368 = ~n36184 ;
  assign y14369 = ~n36193 ;
  assign y14370 = n36197 ;
  assign y14371 = ~1'b0 ;
  assign y14372 = n36201 ;
  assign y14373 = n36205 ;
  assign y14374 = n36207 ;
  assign y14375 = ~n36209 ;
  assign y14376 = ~n36210 ;
  assign y14377 = n36212 ;
  assign y14378 = n36216 ;
  assign y14379 = 1'b0 ;
  assign y14380 = 1'b0 ;
  assign y14381 = n36217 ;
  assign y14382 = ~n36219 ;
  assign y14383 = ~n1134 ;
  assign y14384 = n36221 ;
  assign y14385 = ~1'b0 ;
  assign y14386 = ~n36226 ;
  assign y14387 = ~1'b0 ;
  assign y14388 = ~n36229 ;
  assign y14389 = ~n36233 ;
  assign y14390 = ~n36238 ;
  assign y14391 = n36239 ;
  assign y14392 = n36241 ;
  assign y14393 = ~1'b0 ;
  assign y14394 = ~n2849 ;
  assign y14395 = ~n36244 ;
  assign y14396 = n36251 ;
  assign y14397 = n36253 ;
  assign y14398 = ~n36255 ;
  assign y14399 = ~1'b0 ;
  assign y14400 = ~n26410 ;
  assign y14401 = n36263 ;
  assign y14402 = n36268 ;
  assign y14403 = ~n36269 ;
  assign y14404 = ~1'b0 ;
  assign y14405 = ~1'b0 ;
  assign y14406 = n36270 ;
  assign y14407 = n36273 ;
  assign y14408 = ~n36275 ;
  assign y14409 = n3475 ;
  assign y14410 = n36276 ;
  assign y14411 = ~1'b0 ;
  assign y14412 = n36278 ;
  assign y14413 = ~1'b0 ;
  assign y14414 = ~n36286 ;
  assign y14415 = n5432 ;
  assign y14416 = ~1'b0 ;
  assign y14417 = n36287 ;
  assign y14418 = ~n36292 ;
  assign y14419 = n36295 ;
  assign y14420 = ~1'b0 ;
  assign y14421 = n11871 ;
  assign y14422 = n36297 ;
  assign y14423 = ~1'b0 ;
  assign y14424 = n36298 ;
  assign y14425 = ~1'b0 ;
  assign y14426 = ~n36301 ;
  assign y14427 = n36302 ;
  assign y14428 = ~n36305 ;
  assign y14429 = n36307 ;
  assign y14430 = ~1'b0 ;
  assign y14431 = ~n36309 ;
  assign y14432 = n36310 ;
  assign y14433 = ~1'b0 ;
  assign y14434 = ~n36322 ;
  assign y14435 = ~n36326 ;
  assign y14436 = n36332 ;
  assign y14437 = n36333 ;
  assign y14438 = ~n36334 ;
  assign y14439 = ~n36337 ;
  assign y14440 = 1'b0 ;
  assign y14441 = ~1'b0 ;
  assign y14442 = ~1'b0 ;
  assign y14443 = n36338 ;
  assign y14444 = ~n36342 ;
  assign y14445 = ~n36344 ;
  assign y14446 = ~n36346 ;
  assign y14447 = ~n36349 ;
  assign y14448 = ~n36355 ;
  assign y14449 = ~n36357 ;
  assign y14450 = ~1'b0 ;
  assign y14451 = ~n36359 ;
  assign y14452 = n36360 ;
  assign y14453 = n36363 ;
  assign y14454 = n36364 ;
  assign y14455 = n36365 ;
  assign y14456 = ~n36366 ;
  assign y14457 = 1'b0 ;
  assign y14458 = n36369 ;
  assign y14459 = ~n36373 ;
  assign y14460 = n36376 ;
  assign y14461 = ~n36377 ;
  assign y14462 = n36382 ;
  assign y14463 = ~n36387 ;
  assign y14464 = n36390 ;
  assign y14465 = ~n36392 ;
  assign y14466 = ~1'b0 ;
  assign y14467 = ~n36396 ;
  assign y14468 = ~n36403 ;
  assign y14469 = ~n32574 ;
  assign y14470 = n36407 ;
  assign y14471 = ~n36409 ;
  assign y14472 = n36416 ;
  assign y14473 = ~1'b0 ;
  assign y14474 = n36418 ;
  assign y14475 = ~1'b0 ;
  assign y14476 = n36419 ;
  assign y14477 = ~1'b0 ;
  assign y14478 = n36422 ;
  assign y14479 = n36425 ;
  assign y14480 = ~n36426 ;
  assign y14481 = n4434 ;
  assign y14482 = ~n36427 ;
  assign y14483 = ~1'b0 ;
  assign y14484 = ~n36430 ;
  assign y14485 = ~n36432 ;
  assign y14486 = n36437 ;
  assign y14487 = ~1'b0 ;
  assign y14488 = ~1'b0 ;
  assign y14489 = n36439 ;
  assign y14490 = ~1'b0 ;
  assign y14491 = ~n36444 ;
  assign y14492 = ~n36450 ;
  assign y14493 = ~n30699 ;
  assign y14494 = n36452 ;
  assign y14495 = n36453 ;
  assign y14496 = ~n36454 ;
  assign y14497 = ~n36455 ;
  assign y14498 = n36456 ;
  assign y14499 = ~n36460 ;
  assign y14500 = n36462 ;
  assign y14501 = ~n36467 ;
  assign y14502 = n36469 ;
  assign y14503 = n36470 ;
  assign y14504 = ~n36476 ;
  assign y14505 = n36479 ;
  assign y14506 = ~n36480 ;
  assign y14507 = ~1'b0 ;
  assign y14508 = n36481 ;
  assign y14509 = ~n36482 ;
  assign y14510 = ~1'b0 ;
  assign y14511 = n36486 ;
  assign y14512 = ~n36489 ;
  assign y14513 = n36492 ;
  assign y14514 = n36493 ;
  assign y14515 = ~n36495 ;
  assign y14516 = ~n36500 ;
  assign y14517 = n36503 ;
  assign y14518 = ~n36505 ;
  assign y14519 = ~n36509 ;
  assign y14520 = n36510 ;
  assign y14521 = ~n36513 ;
  assign y14522 = n36514 ;
  assign y14523 = n9376 ;
  assign y14524 = ~n36516 ;
  assign y14525 = ~n36517 ;
  assign y14526 = ~n36518 ;
  assign y14527 = n36520 ;
  assign y14528 = n36525 ;
  assign y14529 = ~n36527 ;
  assign y14530 = ~n36529 ;
  assign y14531 = ~n36535 ;
  assign y14532 = ~n36537 ;
  assign y14533 = n36540 ;
  assign y14534 = ~1'b0 ;
  assign y14535 = ~1'b0 ;
  assign y14536 = ~n36545 ;
  assign y14537 = n36548 ;
  assign y14538 = n36549 ;
  assign y14539 = ~n36554 ;
  assign y14540 = ~n36555 ;
  assign y14541 = ~1'b0 ;
  assign y14542 = ~n7416 ;
  assign y14543 = ~1'b0 ;
  assign y14544 = ~1'b0 ;
  assign y14545 = ~n36558 ;
  assign y14546 = n36561 ;
  assign y14547 = ~n36564 ;
  assign y14548 = ~1'b0 ;
  assign y14549 = ~1'b0 ;
  assign y14550 = n36567 ;
  assign y14551 = ~1'b0 ;
  assign y14552 = ~1'b0 ;
  assign y14553 = ~1'b0 ;
  assign y14554 = n36568 ;
  assign y14555 = n36570 ;
  assign y14556 = n36571 ;
  assign y14557 = ~n36573 ;
  assign y14558 = ~n36576 ;
  assign y14559 = ~1'b0 ;
  assign y14560 = ~n36582 ;
  assign y14561 = ~1'b0 ;
  assign y14562 = n36583 ;
  assign y14563 = n36584 ;
  assign y14564 = n36594 ;
  assign y14565 = n36599 ;
  assign y14566 = n36600 ;
  assign y14567 = ~n36601 ;
  assign y14568 = ~1'b0 ;
  assign y14569 = ~1'b0 ;
  assign y14570 = 1'b0 ;
  assign y14571 = n36602 ;
  assign y14572 = ~1'b0 ;
  assign y14573 = n36603 ;
  assign y14574 = ~n36605 ;
  assign y14575 = ~n36607 ;
  assign y14576 = ~1'b0 ;
  assign y14577 = ~n36609 ;
  assign y14578 = ~n36611 ;
  assign y14579 = n11620 ;
  assign y14580 = n36617 ;
  assign y14581 = n36620 ;
  assign y14582 = n36624 ;
  assign y14583 = n36629 ;
  assign y14584 = ~1'b0 ;
  assign y14585 = n36630 ;
  assign y14586 = ~n36632 ;
  assign y14587 = ~1'b0 ;
  assign y14588 = ~n36634 ;
  assign y14589 = ~n36636 ;
  assign y14590 = ~n36640 ;
  assign y14591 = n36645 ;
  assign y14592 = n36650 ;
  assign y14593 = ~1'b0 ;
  assign y14594 = ~1'b0 ;
  assign y14595 = 1'b0 ;
  assign y14596 = ~1'b0 ;
  assign y14597 = ~n36652 ;
  assign y14598 = n36653 ;
  assign y14599 = ~n36654 ;
  assign y14600 = n36656 ;
  assign y14601 = n36661 ;
  assign y14602 = n36663 ;
  assign y14603 = n36665 ;
  assign y14604 = ~1'b0 ;
  assign y14605 = ~n36667 ;
  assign y14606 = n36669 ;
  assign y14607 = ~1'b0 ;
  assign y14608 = ~n36670 ;
  assign y14609 = n36671 ;
  assign y14610 = n8556 ;
  assign y14611 = n36674 ;
  assign y14612 = ~1'b0 ;
  assign y14613 = ~n1339 ;
  assign y14614 = ~1'b0 ;
  assign y14615 = n36678 ;
  assign y14616 = n36681 ;
  assign y14617 = n36684 ;
  assign y14618 = n18479 ;
  assign y14619 = ~n36690 ;
  assign y14620 = n36692 ;
  assign y14621 = ~n36695 ;
  assign y14622 = ~1'b0 ;
  assign y14623 = ~n36698 ;
  assign y14624 = ~n36700 ;
  assign y14625 = ~1'b0 ;
  assign y14626 = ~n36701 ;
  assign y14627 = ~n36702 ;
  assign y14628 = n36703 ;
  assign y14629 = n36704 ;
  assign y14630 = n36705 ;
  assign y14631 = ~1'b0 ;
  assign y14632 = ~1'b0 ;
  assign y14633 = ~n36707 ;
  assign y14634 = ~1'b0 ;
  assign y14635 = ~n36712 ;
  assign y14636 = n36716 ;
  assign y14637 = ~n36717 ;
  assign y14638 = n36718 ;
  assign y14639 = ~1'b0 ;
  assign y14640 = ~n36720 ;
  assign y14641 = ~1'b0 ;
  assign y14642 = ~1'b0 ;
  assign y14643 = ~1'b0 ;
  assign y14644 = ~n36726 ;
  assign y14645 = n36730 ;
  assign y14646 = n36732 ;
  assign y14647 = ~n36734 ;
  assign y14648 = ~n36742 ;
  assign y14649 = ~1'b0 ;
  assign y14650 = ~n36743 ;
  assign y14651 = n25059 ;
  assign y14652 = n36745 ;
  assign y14653 = ~n36749 ;
  assign y14654 = ~n36750 ;
  assign y14655 = n36753 ;
  assign y14656 = ~1'b0 ;
  assign y14657 = n36755 ;
  assign y14658 = ~n36757 ;
  assign y14659 = ~n36761 ;
  assign y14660 = ~1'b0 ;
  assign y14661 = n36763 ;
  assign y14662 = n36767 ;
  assign y14663 = ~n36768 ;
  assign y14664 = ~n36770 ;
  assign y14665 = ~n36775 ;
  assign y14666 = ~1'b0 ;
  assign y14667 = ~1'b0 ;
  assign y14668 = n22297 ;
  assign y14669 = ~n36776 ;
  assign y14670 = ~n36780 ;
  assign y14671 = ~n36784 ;
  assign y14672 = ~1'b0 ;
  assign y14673 = ~1'b0 ;
  assign y14674 = ~1'b0 ;
  assign y14675 = n36788 ;
  assign y14676 = ~n36791 ;
  assign y14677 = n36792 ;
  assign y14678 = ~n36797 ;
  assign y14679 = 1'b0 ;
  assign y14680 = n36800 ;
  assign y14681 = n36803 ;
  assign y14682 = ~n36806 ;
  assign y14683 = n36807 ;
  assign y14684 = n36816 ;
  assign y14685 = ~n36821 ;
  assign y14686 = ~n36823 ;
  assign y14687 = ~n36827 ;
  assign y14688 = ~1'b0 ;
  assign y14689 = ~n36829 ;
  assign y14690 = n36831 ;
  assign y14691 = n36839 ;
  assign y14692 = n36841 ;
  assign y14693 = ~n36847 ;
  assign y14694 = ~n36850 ;
  assign y14695 = ~n36854 ;
  assign y14696 = ~1'b0 ;
  assign y14697 = ~1'b0 ;
  assign y14698 = ~1'b0 ;
  assign y14699 = ~n36858 ;
  assign y14700 = n36860 ;
  assign y14701 = n36861 ;
  assign y14702 = ~n36868 ;
  assign y14703 = n36873 ;
  assign y14704 = n36874 ;
  assign y14705 = n36875 ;
  assign y14706 = ~n36879 ;
  assign y14707 = ~1'b0 ;
  assign y14708 = n36880 ;
  assign y14709 = ~n36882 ;
  assign y14710 = ~1'b0 ;
  assign y14711 = ~n36885 ;
  assign y14712 = n36886 ;
  assign y14713 = ~1'b0 ;
  assign y14714 = ~1'b0 ;
  assign y14715 = ~1'b0 ;
  assign y14716 = ~n36893 ;
  assign y14717 = ~n36899 ;
  assign y14718 = ~n36901 ;
  assign y14719 = ~n36903 ;
  assign y14720 = ~n36904 ;
  assign y14721 = n36906 ;
  assign y14722 = n36907 ;
  assign y14723 = n36910 ;
  assign y14724 = ~n36912 ;
  assign y14725 = ~1'b0 ;
  assign y14726 = ~1'b0 ;
  assign y14727 = ~n36913 ;
  assign y14728 = ~n36914 ;
  assign y14729 = ~n36915 ;
  assign y14730 = ~1'b0 ;
  assign y14731 = n36917 ;
  assign y14732 = ~1'b0 ;
  assign y14733 = ~n3736 ;
  assign y14734 = ~n36918 ;
  assign y14735 = n36921 ;
  assign y14736 = n36927 ;
  assign y14737 = ~1'b0 ;
  assign y14738 = ~n36930 ;
  assign y14739 = 1'b0 ;
  assign y14740 = ~n36933 ;
  assign y14741 = n36935 ;
  assign y14742 = n36936 ;
  assign y14743 = ~n36937 ;
  assign y14744 = n36939 ;
  assign y14745 = ~n36943 ;
  assign y14746 = ~n36945 ;
  assign y14747 = ~1'b0 ;
  assign y14748 = n36947 ;
  assign y14749 = n36948 ;
  assign y14750 = ~n36954 ;
  assign y14751 = ~1'b0 ;
  assign y14752 = ~1'b0 ;
  assign y14753 = ~n36958 ;
  assign y14754 = ~n36961 ;
  assign y14755 = ~1'b0 ;
  assign y14756 = ~n36968 ;
  assign y14757 = ~n36972 ;
  assign y14758 = n6341 ;
  assign y14759 = ~n36975 ;
  assign y14760 = n36977 ;
  assign y14761 = ~n17270 ;
  assign y14762 = ~n36985 ;
  assign y14763 = ~n36990 ;
  assign y14764 = ~n36991 ;
  assign y14765 = n36993 ;
  assign y14766 = n36999 ;
  assign y14767 = n37002 ;
  assign y14768 = ~n37004 ;
  assign y14769 = ~1'b0 ;
  assign y14770 = ~1'b0 ;
  assign y14771 = ~n37005 ;
  assign y14772 = ~n37008 ;
  assign y14773 = 1'b0 ;
  assign y14774 = n37010 ;
  assign y14775 = ~1'b0 ;
  assign y14776 = n37013 ;
  assign y14777 = n37018 ;
  assign y14778 = ~n37020 ;
  assign y14779 = ~n37021 ;
  assign y14780 = ~n37024 ;
  assign y14781 = n37025 ;
  assign y14782 = n37032 ;
  assign y14783 = ~n37035 ;
  assign y14784 = ~n37043 ;
  assign y14785 = n37045 ;
  assign y14786 = ~1'b0 ;
  assign y14787 = ~1'b0 ;
  assign y14788 = ~n37047 ;
  assign y14789 = n37050 ;
  assign y14790 = n37052 ;
  assign y14791 = ~n37056 ;
  assign y14792 = ~n37057 ;
  assign y14793 = ~n37063 ;
  assign y14794 = n37064 ;
  assign y14795 = ~1'b0 ;
  assign y14796 = n37066 ;
  assign y14797 = ~1'b0 ;
  assign y14798 = n37069 ;
  assign y14799 = n37076 ;
  assign y14800 = n37078 ;
  assign y14801 = n37079 ;
  assign y14802 = ~n37083 ;
  assign y14803 = n37087 ;
  assign y14804 = n37088 ;
  assign y14805 = n37091 ;
  assign y14806 = n37092 ;
  assign y14807 = n37095 ;
  assign y14808 = ~n37097 ;
  assign y14809 = ~n37099 ;
  assign y14810 = ~n37104 ;
  assign y14811 = ~1'b0 ;
  assign y14812 = ~n37105 ;
  assign y14813 = ~n37111 ;
  assign y14814 = n37124 ;
  assign y14815 = ~n37125 ;
  assign y14816 = ~1'b0 ;
  assign y14817 = ~n37127 ;
  assign y14818 = ~n37131 ;
  assign y14819 = n37134 ;
  assign y14820 = ~n37135 ;
  assign y14821 = ~n37136 ;
  assign y14822 = n37142 ;
  assign y14823 = ~n4404 ;
  assign y14824 = n37143 ;
  assign y14825 = n37145 ;
  assign y14826 = ~1'b0 ;
  assign y14827 = ~n37149 ;
  assign y14828 = ~n37150 ;
  assign y14829 = ~1'b0 ;
  assign y14830 = ~n37156 ;
  assign y14831 = ~1'b0 ;
  assign y14832 = n37158 ;
  assign y14833 = n37159 ;
  assign y14834 = n36343 ;
  assign y14835 = ~n37164 ;
  assign y14836 = n37168 ;
  assign y14837 = ~n37169 ;
  assign y14838 = n37171 ;
  assign y14839 = n37172 ;
  assign y14840 = ~n37175 ;
  assign y14841 = n37181 ;
  assign y14842 = ~n37183 ;
  assign y14843 = n37184 ;
  assign y14844 = ~n37187 ;
  assign y14845 = ~1'b0 ;
  assign y14846 = ~1'b0 ;
  assign y14847 = ~n37188 ;
  assign y14848 = n37189 ;
  assign y14849 = ~1'b0 ;
  assign y14850 = ~n37191 ;
  assign y14851 = n37192 ;
  assign y14852 = n37194 ;
  assign y14853 = ~1'b0 ;
  assign y14854 = n37198 ;
  assign y14855 = ~1'b0 ;
  assign y14856 = ~n37200 ;
  assign y14857 = n37202 ;
  assign y14858 = n37203 ;
  assign y14859 = n37204 ;
  assign y14860 = ~1'b0 ;
  assign y14861 = n37206 ;
  assign y14862 = n37214 ;
  assign y14863 = ~n37215 ;
  assign y14864 = ~n37219 ;
  assign y14865 = n37222 ;
  assign y14866 = n37223 ;
  assign y14867 = ~n37226 ;
  assign y14868 = n37227 ;
  assign y14869 = ~n37228 ;
  assign y14870 = ~1'b0 ;
  assign y14871 = ~1'b0 ;
  assign y14872 = n37230 ;
  assign y14873 = ~n37239 ;
  assign y14874 = ~n37240 ;
  assign y14875 = ~n37242 ;
  assign y14876 = ~n37247 ;
  assign y14877 = ~n37257 ;
  assign y14878 = 1'b0 ;
  assign y14879 = 1'b0 ;
  assign y14880 = ~n37259 ;
  assign y14881 = ~n37261 ;
  assign y14882 = ~n37262 ;
  assign y14883 = ~1'b0 ;
  assign y14884 = ~n37265 ;
  assign y14885 = ~n37266 ;
  assign y14886 = n37269 ;
  assign y14887 = n37273 ;
  assign y14888 = n37276 ;
  assign y14889 = ~n37278 ;
  assign y14890 = n37280 ;
  assign y14891 = ~1'b0 ;
  assign y14892 = n37281 ;
  assign y14893 = ~n37288 ;
  assign y14894 = n37292 ;
  assign y14895 = ~n37293 ;
  assign y14896 = ~n37296 ;
  assign y14897 = ~1'b0 ;
  assign y14898 = ~n37298 ;
  assign y14899 = ~1'b0 ;
  assign y14900 = n37302 ;
  assign y14901 = n37304 ;
  assign y14902 = n37307 ;
  assign y14903 = n37313 ;
  assign y14904 = n37314 ;
  assign y14905 = ~n37315 ;
  assign y14906 = ~1'b0 ;
  assign y14907 = ~n37317 ;
  assign y14908 = ~n37322 ;
  assign y14909 = ~1'b0 ;
  assign y14910 = n37326 ;
  assign y14911 = n37329 ;
  assign y14912 = ~n37330 ;
  assign y14913 = n37334 ;
  assign y14914 = n37335 ;
  assign y14915 = ~n37343 ;
  assign y14916 = ~n37344 ;
  assign y14917 = n37345 ;
  assign y14918 = ~n37349 ;
  assign y14919 = ~n37350 ;
  assign y14920 = ~n37353 ;
  assign y14921 = ~n37354 ;
  assign y14922 = ~n37355 ;
  assign y14923 = ~n37358 ;
  assign y14924 = n37361 ;
  assign y14925 = ~1'b0 ;
  assign y14926 = ~n23253 ;
  assign y14927 = ~n37362 ;
  assign y14928 = ~1'b0 ;
  assign y14929 = ~1'b0 ;
  assign y14930 = n37364 ;
  assign y14931 = n37368 ;
  assign y14932 = ~1'b0 ;
  assign y14933 = ~n37372 ;
  assign y14934 = n37375 ;
  assign y14935 = ~n37376 ;
  assign y14936 = ~n37377 ;
  assign y14937 = ~1'b0 ;
  assign y14938 = ~1'b0 ;
  assign y14939 = n37379 ;
  assign y14940 = ~1'b0 ;
  assign y14941 = ~1'b0 ;
  assign y14942 = n37383 ;
  assign y14943 = n37385 ;
  assign y14944 = ~n37394 ;
  assign y14945 = ~n37395 ;
  assign y14946 = ~n37396 ;
  assign y14947 = ~n37400 ;
  assign y14948 = ~n37402 ;
  assign y14949 = ~n37407 ;
  assign y14950 = ~n37408 ;
  assign y14951 = ~n37412 ;
  assign y14952 = n37415 ;
  assign y14953 = ~n37416 ;
  assign y14954 = ~n37418 ;
  assign y14955 = ~1'b0 ;
  assign y14956 = n37421 ;
  assign y14957 = ~1'b0 ;
  assign y14958 = n37422 ;
  assign y14959 = n37425 ;
  assign y14960 = ~n37430 ;
  assign y14961 = n37434 ;
  assign y14962 = ~n37437 ;
  assign y14963 = ~1'b0 ;
  assign y14964 = ~1'b0 ;
  assign y14965 = ~1'b0 ;
  assign y14966 = ~1'b0 ;
  assign y14967 = ~n37441 ;
  assign y14968 = n37442 ;
  assign y14969 = n37454 ;
  assign y14970 = ~n37458 ;
  assign y14971 = ~1'b0 ;
  assign y14972 = ~n37461 ;
  assign y14973 = ~n37464 ;
  assign y14974 = ~n37467 ;
  assign y14975 = ~n37475 ;
  assign y14976 = n37477 ;
  assign y14977 = ~n37478 ;
  assign y14978 = ~n37479 ;
  assign y14979 = ~n37481 ;
  assign y14980 = n37484 ;
  assign y14981 = n37485 ;
  assign y14982 = ~n37488 ;
  assign y14983 = n37494 ;
  assign y14984 = ~n37498 ;
  assign y14985 = ~n37507 ;
  assign y14986 = ~1'b0 ;
  assign y14987 = ~1'b0 ;
  assign y14988 = ~1'b0 ;
  assign y14989 = ~n37509 ;
  assign y14990 = n37512 ;
  assign y14991 = ~n37519 ;
  assign y14992 = n37521 ;
  assign y14993 = ~n37526 ;
  assign y14994 = ~n37527 ;
  assign y14995 = ~n37531 ;
  assign y14996 = n32573 ;
  assign y14997 = n37538 ;
  assign y14998 = n37540 ;
  assign y14999 = ~n37544 ;
  assign y15000 = ~1'b0 ;
  assign y15001 = ~1'b0 ;
  assign y15002 = ~1'b0 ;
  assign y15003 = ~1'b0 ;
  assign y15004 = ~1'b0 ;
  assign y15005 = ~n37545 ;
  assign y15006 = n37546 ;
  assign y15007 = n37547 ;
  assign y15008 = n37551 ;
  assign y15009 = ~1'b0 ;
  assign y15010 = ~1'b0 ;
  assign y15011 = n21486 ;
  assign y15012 = ~1'b0 ;
  assign y15013 = n37557 ;
  assign y15014 = x252 ;
  assign y15015 = ~n37558 ;
  assign y15016 = n37563 ;
  assign y15017 = n37566 ;
  assign y15018 = ~1'b0 ;
  assign y15019 = ~1'b0 ;
  assign y15020 = n15950 ;
  assign y15021 = ~1'b0 ;
  assign y15022 = ~n37569 ;
  assign y15023 = n37570 ;
  assign y15024 = ~1'b0 ;
  assign y15025 = ~n37571 ;
  assign y15026 = ~1'b0 ;
  assign y15027 = n37573 ;
  assign y15028 = ~1'b0 ;
  assign y15029 = n21291 ;
  assign y15030 = n37574 ;
  assign y15031 = n37575 ;
  assign y15032 = ~n37579 ;
  assign y15033 = ~n37581 ;
  assign y15034 = ~1'b0 ;
  assign y15035 = ~1'b0 ;
  assign y15036 = n37582 ;
  assign y15037 = n37583 ;
  assign y15038 = ~n37585 ;
  assign y15039 = n37588 ;
  assign y15040 = ~1'b0 ;
  assign y15041 = ~1'b0 ;
  assign y15042 = ~n37591 ;
  assign y15043 = ~n37595 ;
  assign y15044 = ~n37598 ;
  assign y15045 = n37599 ;
  assign y15046 = n37602 ;
  assign y15047 = ~n37605 ;
  assign y15048 = ~n37611 ;
  assign y15049 = n37615 ;
  assign y15050 = ~n37617 ;
  assign y15051 = ~n37618 ;
  assign y15052 = ~1'b0 ;
  assign y15053 = ~n37621 ;
  assign y15054 = n37622 ;
  assign y15055 = ~n37631 ;
  assign y15056 = ~n37633 ;
  assign y15057 = n7653 ;
  assign y15058 = n37634 ;
  assign y15059 = ~1'b0 ;
  assign y15060 = ~n37635 ;
  assign y15061 = ~1'b0 ;
  assign y15062 = n37637 ;
  assign y15063 = ~1'b0 ;
  assign y15064 = n37643 ;
  assign y15065 = ~n37644 ;
  assign y15066 = ~n37647 ;
  assign y15067 = n37650 ;
  assign y15068 = ~n37654 ;
  assign y15069 = ~1'b0 ;
  assign y15070 = ~n37655 ;
  assign y15071 = ~1'b0 ;
  assign y15072 = ~n37658 ;
  assign y15073 = ~n37659 ;
  assign y15074 = ~n37662 ;
  assign y15075 = ~1'b0 ;
  assign y15076 = n37664 ;
  assign y15077 = ~n37669 ;
  assign y15078 = 1'b0 ;
  assign y15079 = n37670 ;
  assign y15080 = ~1'b0 ;
  assign y15081 = n37671 ;
  assign y15082 = n37674 ;
  assign y15083 = n37676 ;
  assign y15084 = ~n37678 ;
  assign y15085 = ~n37681 ;
  assign y15086 = n37683 ;
  assign y15087 = ~1'b0 ;
  assign y15088 = ~1'b0 ;
  assign y15089 = n37686 ;
  assign y15090 = ~n37687 ;
  assign y15091 = n37690 ;
  assign y15092 = ~n37691 ;
  assign y15093 = 1'b0 ;
  assign y15094 = ~1'b0 ;
  assign y15095 = ~1'b0 ;
  assign y15096 = ~1'b0 ;
  assign y15097 = ~n37696 ;
  assign y15098 = n37697 ;
  assign y15099 = ~n37702 ;
  assign y15100 = n37703 ;
  assign y15101 = n37705 ;
  assign y15102 = n37707 ;
  assign y15103 = ~1'b0 ;
  assign y15104 = ~1'b0 ;
  assign y15105 = ~1'b0 ;
  assign y15106 = ~1'b0 ;
  assign y15107 = ~n37708 ;
  assign y15108 = ~n37709 ;
  assign y15109 = ~1'b0 ;
  assign y15110 = ~1'b0 ;
  assign y15111 = n37710 ;
  assign y15112 = n37711 ;
  assign y15113 = ~1'b0 ;
  assign y15114 = n37713 ;
  assign y15115 = ~n37715 ;
  assign y15116 = n37723 ;
  assign y15117 = ~n37724 ;
  assign y15118 = n37725 ;
  assign y15119 = ~n37731 ;
  assign y15120 = ~n37733 ;
  assign y15121 = n37735 ;
  assign y15122 = n5899 ;
  assign y15123 = ~n37736 ;
  assign y15124 = ~1'b0 ;
  assign y15125 = n37738 ;
  assign y15126 = n37741 ;
  assign y15127 = n37743 ;
  assign y15128 = n37752 ;
  assign y15129 = n37754 ;
  assign y15130 = n37755 ;
  assign y15131 = ~n37756 ;
  assign y15132 = ~n37759 ;
  assign y15133 = n37760 ;
  assign y15134 = n37765 ;
  assign y15135 = ~n37769 ;
  assign y15136 = ~n37771 ;
  assign y15137 = ~1'b0 ;
  assign y15138 = n37773 ;
  assign y15139 = n37774 ;
  assign y15140 = ~n37777 ;
  assign y15141 = ~n37779 ;
  assign y15142 = ~n37784 ;
  assign y15143 = n37786 ;
  assign y15144 = n37788 ;
  assign y15145 = ~n37791 ;
  assign y15146 = ~n37792 ;
  assign y15147 = ~1'b0 ;
  assign y15148 = ~n37799 ;
  assign y15149 = ~n37802 ;
  assign y15150 = ~n37803 ;
  assign y15151 = ~n37804 ;
  assign y15152 = ~1'b0 ;
  assign y15153 = ~1'b0 ;
  assign y15154 = n37808 ;
  assign y15155 = ~1'b0 ;
  assign y15156 = ~n37812 ;
  assign y15157 = n37813 ;
  assign y15158 = ~n6647 ;
  assign y15159 = n37822 ;
  assign y15160 = ~n37826 ;
  assign y15161 = ~1'b0 ;
  assign y15162 = ~n37832 ;
  assign y15163 = n37834 ;
  assign y15164 = n37835 ;
  assign y15165 = ~n37838 ;
  assign y15166 = ~1'b0 ;
  assign y15167 = ~1'b0 ;
  assign y15168 = ~n37841 ;
  assign y15169 = n37844 ;
  assign y15170 = n37846 ;
  assign y15171 = ~1'b0 ;
  assign y15172 = ~n37848 ;
  assign y15173 = ~1'b0 ;
  assign y15174 = ~n32642 ;
  assign y15175 = n37849 ;
  assign y15176 = n37851 ;
  assign y15177 = n37854 ;
  assign y15178 = ~1'b0 ;
  assign y15179 = ~n37858 ;
  assign y15180 = ~n37859 ;
  assign y15181 = n37863 ;
  assign y15182 = ~n25580 ;
  assign y15183 = n37865 ;
  assign y15184 = n37866 ;
  assign y15185 = n37871 ;
  assign y15186 = n37877 ;
  assign y15187 = n37879 ;
  assign y15188 = n37886 ;
  assign y15189 = ~1'b0 ;
  assign y15190 = n37887 ;
  assign y15191 = ~n37890 ;
  assign y15192 = n37892 ;
  assign y15193 = ~n37894 ;
  assign y15194 = ~n37897 ;
  assign y15195 = n37898 ;
  assign y15196 = ~n37899 ;
  assign y15197 = n37902 ;
  assign y15198 = n37906 ;
  assign y15199 = ~n37911 ;
  assign y15200 = n37917 ;
  assign y15201 = ~n37918 ;
  assign y15202 = ~n37923 ;
  assign y15203 = 1'b0 ;
  assign y15204 = ~1'b0 ;
  assign y15205 = ~n37924 ;
  assign y15206 = ~n37930 ;
  assign y15207 = n37934 ;
  assign y15208 = ~1'b0 ;
  assign y15209 = ~1'b0 ;
  assign y15210 = n37937 ;
  assign y15211 = ~1'b0 ;
  assign y15212 = ~n37939 ;
  assign y15213 = n37940 ;
  assign y15214 = ~n37941 ;
  assign y15215 = n37945 ;
  assign y15216 = n37947 ;
  assign y15217 = n37949 ;
  assign y15218 = ~1'b0 ;
  assign y15219 = ~n17721 ;
  assign y15220 = ~1'b0 ;
  assign y15221 = n37951 ;
  assign y15222 = n37953 ;
  assign y15223 = ~n37954 ;
  assign y15224 = ~1'b0 ;
  assign y15225 = ~1'b0 ;
  assign y15226 = ~n37958 ;
  assign y15227 = n37962 ;
  assign y15228 = ~1'b0 ;
  assign y15229 = n37965 ;
  assign y15230 = ~n37966 ;
  assign y15231 = ~n37967 ;
  assign y15232 = ~n37972 ;
  assign y15233 = ~n37979 ;
  assign y15234 = n37980 ;
  assign y15235 = ~n37982 ;
  assign y15236 = n37987 ;
  assign y15237 = n37989 ;
  assign y15238 = ~n37990 ;
  assign y15239 = n37992 ;
  assign y15240 = ~n38001 ;
  assign y15241 = ~1'b0 ;
  assign y15242 = ~n38002 ;
  assign y15243 = 1'b0 ;
  assign y15244 = ~1'b0 ;
  assign y15245 = n38004 ;
  assign y15246 = n38005 ;
  assign y15247 = ~n38008 ;
  assign y15248 = ~n38013 ;
  assign y15249 = n38016 ;
  assign y15250 = ~n38017 ;
  assign y15251 = n38018 ;
  assign y15252 = n38021 ;
  assign y15253 = ~1'b0 ;
  assign y15254 = ~1'b0 ;
  assign y15255 = 1'b0 ;
  assign y15256 = ~n38024 ;
  assign y15257 = n38025 ;
  assign y15258 = n3633 ;
  assign y15259 = n38028 ;
  assign y15260 = n38035 ;
  assign y15261 = n38039 ;
  assign y15262 = ~1'b0 ;
  assign y15263 = ~n38040 ;
  assign y15264 = ~n38044 ;
  assign y15265 = n38045 ;
  assign y15266 = n38052 ;
  assign y15267 = ~n38053 ;
  assign y15268 = ~1'b0 ;
  assign y15269 = ~1'b0 ;
  assign y15270 = ~n38054 ;
  assign y15271 = n38055 ;
  assign y15272 = ~n38059 ;
  assign y15273 = n38061 ;
  assign y15274 = ~n38062 ;
  assign y15275 = n38065 ;
  assign y15276 = ~n38068 ;
  assign y15277 = n38069 ;
  assign y15278 = ~n38072 ;
  assign y15279 = ~n38074 ;
  assign y15280 = ~1'b0 ;
  assign y15281 = n38076 ;
  assign y15282 = ~n38079 ;
  assign y15283 = n38084 ;
  assign y15284 = n38086 ;
  assign y15285 = ~n38091 ;
  assign y15286 = ~n38095 ;
  assign y15287 = ~n38098 ;
  assign y15288 = ~n38103 ;
  assign y15289 = n38105 ;
  assign y15290 = ~n38111 ;
  assign y15291 = ~n38113 ;
  assign y15292 = n38116 ;
  assign y15293 = ~n38123 ;
  assign y15294 = ~1'b0 ;
  assign y15295 = ~n38126 ;
  assign y15296 = ~1'b0 ;
  assign y15297 = n38129 ;
  assign y15298 = ~n38132 ;
  assign y15299 = ~n38137 ;
  assign y15300 = ~1'b0 ;
  assign y15301 = ~1'b0 ;
  assign y15302 = ~1'b0 ;
  assign y15303 = 1'b0 ;
  assign y15304 = ~n13554 ;
  assign y15305 = ~n38141 ;
  assign y15306 = n38148 ;
  assign y15307 = ~1'b0 ;
  assign y15308 = ~1'b0 ;
  assign y15309 = ~1'b0 ;
  assign y15310 = n38152 ;
  assign y15311 = n38154 ;
  assign y15312 = ~1'b0 ;
  assign y15313 = n38155 ;
  assign y15314 = ~n38158 ;
  assign y15315 = ~n38160 ;
  assign y15316 = ~n38162 ;
  assign y15317 = ~1'b0 ;
  assign y15318 = ~1'b0 ;
  assign y15319 = n38163 ;
  assign y15320 = ~1'b0 ;
  assign y15321 = ~n38166 ;
  assign y15322 = n38167 ;
  assign y15323 = ~1'b0 ;
  assign y15324 = n38168 ;
  assign y15325 = ~1'b0 ;
  assign y15326 = ~n38170 ;
  assign y15327 = ~1'b0 ;
  assign y15328 = ~1'b0 ;
  assign y15329 = n38172 ;
  assign y15330 = ~n38181 ;
  assign y15331 = n38184 ;
  assign y15332 = ~n38185 ;
  assign y15333 = ~n38194 ;
  assign y15334 = n38197 ;
  assign y15335 = n38200 ;
  assign y15336 = n38202 ;
  assign y15337 = n38203 ;
  assign y15338 = ~1'b0 ;
  assign y15339 = ~n38205 ;
  assign y15340 = n38208 ;
  assign y15341 = ~n38210 ;
  assign y15342 = n38213 ;
  assign y15343 = ~n38217 ;
  assign y15344 = ~n38219 ;
  assign y15345 = n13583 ;
  assign y15346 = ~1'b0 ;
  assign y15347 = ~n38221 ;
  assign y15348 = ~n38223 ;
  assign y15349 = ~n38224 ;
  assign y15350 = ~n38225 ;
  assign y15351 = n38227 ;
  assign y15352 = ~n38228 ;
  assign y15353 = n38229 ;
  assign y15354 = n38235 ;
  assign y15355 = ~n38238 ;
  assign y15356 = n22044 ;
  assign y15357 = n38241 ;
  assign y15358 = ~1'b0 ;
  assign y15359 = ~n38245 ;
  assign y15360 = n38248 ;
  assign y15361 = n38250 ;
  assign y15362 = ~n38251 ;
  assign y15363 = ~n38255 ;
  assign y15364 = ~n38258 ;
  assign y15365 = ~1'b0 ;
  assign y15366 = ~n38260 ;
  assign y15367 = ~n38266 ;
  assign y15368 = ~1'b0 ;
  assign y15369 = ~1'b0 ;
  assign y15370 = n38267 ;
  assign y15371 = n38271 ;
  assign y15372 = ~1'b0 ;
  assign y15373 = ~1'b0 ;
  assign y15374 = ~n38273 ;
  assign y15375 = ~1'b0 ;
  assign y15376 = n38280 ;
  assign y15377 = ~n38281 ;
  assign y15378 = ~n38282 ;
  assign y15379 = n38283 ;
  assign y15380 = ~n38287 ;
  assign y15381 = ~1'b0 ;
  assign y15382 = n38290 ;
  assign y15383 = ~n38296 ;
  assign y15384 = ~n38297 ;
  assign y15385 = n38299 ;
  assign y15386 = ~1'b0 ;
  assign y15387 = n38306 ;
  assign y15388 = ~n38308 ;
  assign y15389 = ~n38318 ;
  assign y15390 = n38319 ;
  assign y15391 = ~n38320 ;
  assign y15392 = ~n38321 ;
  assign y15393 = n38328 ;
  assign y15394 = ~n38331 ;
  assign y15395 = n38333 ;
  assign y15396 = ~n38337 ;
  assign y15397 = n38340 ;
  assign y15398 = ~n38342 ;
  assign y15399 = ~1'b0 ;
  assign y15400 = n38345 ;
  assign y15401 = ~n38346 ;
  assign y15402 = n38349 ;
  assign y15403 = ~n38355 ;
  assign y15404 = ~n38357 ;
  assign y15405 = n38362 ;
  assign y15406 = ~1'b0 ;
  assign y15407 = ~1'b0 ;
  assign y15408 = ~n38364 ;
  assign y15409 = ~1'b0 ;
  assign y15410 = ~1'b0 ;
  assign y15411 = ~n38367 ;
  assign y15412 = n38369 ;
  assign y15413 = n38370 ;
  assign y15414 = n38372 ;
  assign y15415 = ~1'b0 ;
  assign y15416 = ~n38373 ;
  assign y15417 = ~1'b0 ;
  assign y15418 = ~1'b0 ;
  assign y15419 = n38381 ;
  assign y15420 = n38389 ;
  assign y15421 = ~n38392 ;
  assign y15422 = ~n38394 ;
  assign y15423 = ~n38396 ;
  assign y15424 = n38399 ;
  assign y15425 = ~n38401 ;
  assign y15426 = n38403 ;
  assign y15427 = ~n38405 ;
  assign y15428 = ~1'b0 ;
  assign y15429 = ~n38410 ;
  assign y15430 = n38412 ;
  assign y15431 = ~n38424 ;
  assign y15432 = ~1'b0 ;
  assign y15433 = n38425 ;
  assign y15434 = n38426 ;
  assign y15435 = ~n38427 ;
  assign y15436 = ~1'b0 ;
  assign y15437 = n38428 ;
  assign y15438 = ~n38429 ;
  assign y15439 = ~n38430 ;
  assign y15440 = n38431 ;
  assign y15441 = ~1'b0 ;
  assign y15442 = n38433 ;
  assign y15443 = n38437 ;
  assign y15444 = ~1'b0 ;
  assign y15445 = ~n38446 ;
  assign y15446 = n38448 ;
  assign y15447 = ~n38449 ;
  assign y15448 = n38451 ;
  assign y15449 = ~1'b0 ;
  assign y15450 = ~n38454 ;
  assign y15451 = n38457 ;
  assign y15452 = ~1'b0 ;
  assign y15453 = n38458 ;
  assign y15454 = ~n38461 ;
  assign y15455 = ~n38462 ;
  assign y15456 = n38464 ;
  assign y15457 = n38465 ;
  assign y15458 = ~1'b0 ;
  assign y15459 = n38466 ;
  assign y15460 = n38467 ;
  assign y15461 = n38469 ;
  assign y15462 = n38470 ;
  assign y15463 = n38478 ;
  assign y15464 = ~n38479 ;
  assign y15465 = ~1'b0 ;
  assign y15466 = n38481 ;
  assign y15467 = ~n38489 ;
  assign y15468 = ~1'b0 ;
  assign y15469 = n38497 ;
  assign y15470 = ~1'b0 ;
  assign y15471 = n32573 ;
  assign y15472 = n38500 ;
  assign y15473 = ~1'b0 ;
  assign y15474 = n38501 ;
  assign y15475 = ~n38502 ;
  assign y15476 = n38504 ;
  assign y15477 = ~n38505 ;
  assign y15478 = n38507 ;
  assign y15479 = n38511 ;
  assign y15480 = ~1'b0 ;
  assign y15481 = ~1'b0 ;
  assign y15482 = n38513 ;
  assign y15483 = ~1'b0 ;
  assign y15484 = ~1'b0 ;
  assign y15485 = ~n38517 ;
  assign y15486 = n38518 ;
  assign y15487 = ~n38519 ;
  assign y15488 = n38520 ;
  assign y15489 = n38522 ;
  assign y15490 = ~1'b0 ;
  assign y15491 = ~1'b0 ;
  assign y15492 = n38525 ;
  assign y15493 = n38526 ;
  assign y15494 = ~n38527 ;
  assign y15495 = ~1'b0 ;
  assign y15496 = ~n38529 ;
  assign y15497 = ~1'b0 ;
  assign y15498 = ~n38536 ;
  assign y15499 = n38537 ;
  assign y15500 = ~n38538 ;
  assign y15501 = ~n38540 ;
  assign y15502 = ~1'b0 ;
  assign y15503 = n38548 ;
  assign y15504 = ~n38551 ;
  assign y15505 = ~1'b0 ;
  assign y15506 = n7535 ;
  assign y15507 = n38552 ;
  assign y15508 = ~n38553 ;
  assign y15509 = ~n38560 ;
  assign y15510 = ~n38562 ;
  assign y15511 = ~n38564 ;
  assign y15512 = n38567 ;
  assign y15513 = n38570 ;
  assign y15514 = n38572 ;
  assign y15515 = ~1'b0 ;
  assign y15516 = ~n38573 ;
  assign y15517 = ~1'b0 ;
  assign y15518 = n38576 ;
  assign y15519 = n38578 ;
  assign y15520 = ~n38582 ;
  assign y15521 = ~n38584 ;
  assign y15522 = ~n38586 ;
  assign y15523 = ~1'b0 ;
  assign y15524 = n38588 ;
  assign y15525 = n38590 ;
  assign y15526 = ~n38593 ;
  assign y15527 = n38594 ;
  assign y15528 = n38598 ;
  assign y15529 = ~n38601 ;
  assign y15530 = ~n38604 ;
  assign y15531 = ~n38605 ;
  assign y15532 = n38608 ;
  assign y15533 = ~1'b0 ;
  assign y15534 = ~1'b0 ;
  assign y15535 = n38612 ;
  assign y15536 = n38616 ;
  assign y15537 = ~n38618 ;
  assign y15538 = ~1'b0 ;
  assign y15539 = n38620 ;
  assign y15540 = n38623 ;
  assign y15541 = ~n38625 ;
  assign y15542 = n38626 ;
  assign y15543 = ~n38629 ;
  assign y15544 = ~n38630 ;
  assign y15545 = n38631 ;
  assign y15546 = ~n38632 ;
  assign y15547 = n38636 ;
  assign y15548 = ~1'b0 ;
  assign y15549 = ~n38637 ;
  assign y15550 = ~n3813 ;
  assign y15551 = ~n38641 ;
  assign y15552 = ~n38642 ;
  assign y15553 = ~n38643 ;
  assign y15554 = n38647 ;
  assign y15555 = n38650 ;
  assign y15556 = ~n38651 ;
  assign y15557 = n38653 ;
  assign y15558 = ~1'b0 ;
  assign y15559 = n38654 ;
  assign y15560 = ~n38656 ;
  assign y15561 = ~n38657 ;
  assign y15562 = n38658 ;
  assign y15563 = n38659 ;
  assign y15564 = ~n38660 ;
  assign y15565 = ~1'b0 ;
  assign y15566 = ~n38665 ;
  assign y15567 = n38669 ;
  assign y15568 = n38675 ;
  assign y15569 = n38677 ;
  assign y15570 = n38678 ;
  assign y15571 = ~1'b0 ;
  assign y15572 = ~1'b0 ;
  assign y15573 = ~n7599 ;
  assign y15574 = n38681 ;
  assign y15575 = ~1'b0 ;
  assign y15576 = n38685 ;
  assign y15577 = ~n38686 ;
  assign y15578 = ~n38687 ;
  assign y15579 = ~n38689 ;
  assign y15580 = n38691 ;
  assign y15581 = ~n38694 ;
  assign y15582 = ~1'b0 ;
  assign y15583 = ~1'b0 ;
  assign y15584 = ~1'b0 ;
  assign y15585 = n38698 ;
  assign y15586 = ~n38702 ;
  assign y15587 = ~n38706 ;
  assign y15588 = ~n38710 ;
  assign y15589 = ~n38714 ;
  assign y15590 = n38715 ;
  assign y15591 = ~n38717 ;
  assign y15592 = ~1'b0 ;
  assign y15593 = n38719 ;
  assign y15594 = ~1'b0 ;
  assign y15595 = n38726 ;
  assign y15596 = n38729 ;
  assign y15597 = n38734 ;
  assign y15598 = n38735 ;
  assign y15599 = ~n38736 ;
  assign y15600 = n38738 ;
  assign y15601 = n38740 ;
  assign y15602 = n38743 ;
  assign y15603 = ~n38746 ;
  assign y15604 = n38750 ;
  assign y15605 = n38751 ;
  assign y15606 = ~n38757 ;
  assign y15607 = ~1'b0 ;
  assign y15608 = ~n38758 ;
  assign y15609 = n38759 ;
  assign y15610 = n38765 ;
  assign y15611 = ~n38772 ;
  assign y15612 = n38779 ;
  assign y15613 = ~1'b0 ;
  assign y15614 = ~n38782 ;
  assign y15615 = n38785 ;
  assign y15616 = n38787 ;
  assign y15617 = n38792 ;
  assign y15618 = n38793 ;
  assign y15619 = ~n38795 ;
  assign y15620 = ~1'b0 ;
  assign y15621 = ~n38798 ;
  assign y15622 = ~n38799 ;
  assign y15623 = ~1'b0 ;
  assign y15624 = ~n38801 ;
  assign y15625 = n38804 ;
  assign y15626 = n38807 ;
  assign y15627 = n38814 ;
  assign y15628 = n38818 ;
  assign y15629 = ~1'b0 ;
  assign y15630 = ~n19413 ;
  assign y15631 = ~1'b0 ;
  assign y15632 = n38821 ;
  assign y15633 = n2756 ;
  assign y15634 = n38822 ;
  assign y15635 = n511 ;
  assign y15636 = ~n38826 ;
  assign y15637 = ~1'b0 ;
  assign y15638 = ~1'b0 ;
  assign y15639 = ~1'b0 ;
  assign y15640 = n38827 ;
  assign y15641 = ~n38828 ;
  assign y15642 = n38829 ;
  assign y15643 = ~n38830 ;
  assign y15644 = ~n38835 ;
  assign y15645 = n38836 ;
  assign y15646 = ~n38838 ;
  assign y15647 = ~n38839 ;
  assign y15648 = n38842 ;
  assign y15649 = ~n38843 ;
  assign y15650 = n38844 ;
  assign y15651 = ~n38849 ;
  assign y15652 = n38852 ;
  assign y15653 = n38853 ;
  assign y15654 = ~n38856 ;
  assign y15655 = n38857 ;
  assign y15656 = ~n38859 ;
  assign y15657 = n38860 ;
  assign y15658 = ~n38862 ;
  assign y15659 = n38865 ;
  assign y15660 = ~1'b0 ;
  assign y15661 = ~n38869 ;
  assign y15662 = n38871 ;
  assign y15663 = n38873 ;
  assign y15664 = n38882 ;
  assign y15665 = n38883 ;
  assign y15666 = n38885 ;
  assign y15667 = ~n38890 ;
  assign y15668 = n38892 ;
  assign y15669 = ~n38895 ;
  assign y15670 = n38896 ;
  assign y15671 = ~1'b0 ;
  assign y15672 = n38900 ;
  assign y15673 = n38902 ;
  assign y15674 = n38905 ;
  assign y15675 = ~n38913 ;
  assign y15676 = ~1'b0 ;
  assign y15677 = n38916 ;
  assign y15678 = ~1'b0 ;
  assign y15679 = ~1'b0 ;
  assign y15680 = ~n38919 ;
  assign y15681 = ~n38920 ;
  assign y15682 = n38929 ;
  assign y15683 = n38930 ;
  assign y15684 = n38933 ;
  assign y15685 = ~n38936 ;
  assign y15686 = ~n38938 ;
  assign y15687 = n38939 ;
  assign y15688 = n38945 ;
  assign y15689 = n38946 ;
  assign y15690 = ~n38947 ;
  assign y15691 = ~n38948 ;
  assign y15692 = n38950 ;
  assign y15693 = ~n38951 ;
  assign y15694 = n38954 ;
  assign y15695 = n38959 ;
  assign y15696 = n38960 ;
  assign y15697 = ~n38961 ;
  assign y15698 = n38968 ;
  assign y15699 = n38969 ;
  assign y15700 = n38970 ;
  assign y15701 = ~n38972 ;
  assign y15702 = ~n38982 ;
  assign y15703 = ~1'b0 ;
  assign y15704 = ~n38986 ;
  assign y15705 = n1496 ;
  assign y15706 = ~n38988 ;
  assign y15707 = ~1'b0 ;
  assign y15708 = ~1'b0 ;
  assign y15709 = ~1'b0 ;
  assign y15710 = ~1'b0 ;
  assign y15711 = ~n38989 ;
  assign y15712 = ~n38990 ;
  assign y15713 = n38991 ;
  assign y15714 = ~1'b0 ;
  assign y15715 = ~1'b0 ;
  assign y15716 = n38995 ;
  assign y15717 = ~n38999 ;
  assign y15718 = ~n39006 ;
  assign y15719 = ~1'b0 ;
  assign y15720 = n39009 ;
  assign y15721 = n39012 ;
  assign y15722 = ~n3156 ;
  assign y15723 = n39015 ;
  assign y15724 = ~n39018 ;
  assign y15725 = ~1'b0 ;
  assign y15726 = n39019 ;
  assign y15727 = n39025 ;
  assign y15728 = n39026 ;
  assign y15729 = n39027 ;
  assign y15730 = ~1'b0 ;
  assign y15731 = ~n39028 ;
  assign y15732 = ~n39029 ;
  assign y15733 = ~n4266 ;
  assign y15734 = ~1'b0 ;
  assign y15735 = ~1'b0 ;
  assign y15736 = ~n39030 ;
  assign y15737 = ~n39034 ;
  assign y15738 = n39035 ;
  assign y15739 = ~n39038 ;
  assign y15740 = ~1'b0 ;
  assign y15741 = n39043 ;
  assign y15742 = n39047 ;
  assign y15743 = n39052 ;
  assign y15744 = n39054 ;
  assign y15745 = ~n39057 ;
  assign y15746 = ~n39066 ;
  assign y15747 = ~n39067 ;
  assign y15748 = ~n39070 ;
  assign y15749 = n39071 ;
  assign y15750 = n39073 ;
  assign y15751 = ~n39076 ;
  assign y15752 = ~n39078 ;
  assign y15753 = n39079 ;
  assign y15754 = ~n14634 ;
  assign y15755 = n39083 ;
  assign y15756 = ~1'b0 ;
  assign y15757 = ~1'b0 ;
  assign y15758 = ~n39084 ;
  assign y15759 = ~n39085 ;
  assign y15760 = n39090 ;
  assign y15761 = n39091 ;
  assign y15762 = ~1'b0 ;
  assign y15763 = ~1'b0 ;
  assign y15764 = ~n39093 ;
  assign y15765 = n39098 ;
  assign y15766 = ~1'b0 ;
  assign y15767 = n39099 ;
  assign y15768 = ~n14859 ;
  assign y15769 = ~n39106 ;
  assign y15770 = ~1'b0 ;
  assign y15771 = ~1'b0 ;
  assign y15772 = ~n39112 ;
  assign y15773 = ~1'b0 ;
  assign y15774 = ~n39113 ;
  assign y15775 = n39115 ;
  assign y15776 = n39116 ;
  assign y15777 = ~1'b0 ;
  assign y15778 = ~n39118 ;
  assign y15779 = n39120 ;
  assign y15780 = ~n39125 ;
  assign y15781 = ~n39132 ;
  assign y15782 = ~n39133 ;
  assign y15783 = ~n1869 ;
  assign y15784 = ~1'b0 ;
  assign y15785 = ~1'b0 ;
  assign y15786 = ~n39138 ;
  assign y15787 = n39140 ;
  assign y15788 = n39141 ;
  assign y15789 = ~n39143 ;
  assign y15790 = ~n39146 ;
  assign y15791 = ~n39147 ;
  assign y15792 = ~n39148 ;
  assign y15793 = ~n39150 ;
  assign y15794 = ~1'b0 ;
  assign y15795 = n39151 ;
  assign y15796 = ~n39155 ;
  assign y15797 = ~1'b0 ;
  assign y15798 = ~n4882 ;
  assign y15799 = ~n39157 ;
  assign y15800 = ~1'b0 ;
  assign y15801 = ~1'b0 ;
  assign y15802 = ~1'b0 ;
  assign y15803 = n39159 ;
  assign y15804 = ~n39160 ;
  assign y15805 = ~n21612 ;
  assign y15806 = n39163 ;
  assign y15807 = n39165 ;
  assign y15808 = ~n39168 ;
  assign y15809 = ~n39171 ;
  assign y15810 = ~n39172 ;
  assign y15811 = ~1'b0 ;
  assign y15812 = ~n39174 ;
  assign y15813 = ~n39175 ;
  assign y15814 = n39179 ;
  assign y15815 = n39181 ;
  assign y15816 = n39184 ;
  assign y15817 = ~n39188 ;
  assign y15818 = 1'b0 ;
  assign y15819 = ~1'b0 ;
  assign y15820 = n39189 ;
  assign y15821 = ~n39192 ;
  assign y15822 = n39203 ;
  assign y15823 = ~n39209 ;
  assign y15824 = ~n39210 ;
  assign y15825 = n39212 ;
  assign y15826 = n39213 ;
  assign y15827 = ~1'b0 ;
  assign y15828 = n39214 ;
  assign y15829 = n39216 ;
  assign y15830 = n39218 ;
  assign y15831 = ~n39220 ;
  assign y15832 = n39230 ;
  assign y15833 = ~n39231 ;
  assign y15834 = n39232 ;
  assign y15835 = ~1'b0 ;
  assign y15836 = ~1'b0 ;
  assign y15837 = ~n39237 ;
  assign y15838 = ~1'b0 ;
  assign y15839 = ~1'b0 ;
  assign y15840 = n39242 ;
  assign y15841 = ~n39243 ;
  assign y15842 = ~n39250 ;
  assign y15843 = ~n39257 ;
  assign y15844 = ~1'b0 ;
  assign y15845 = ~1'b0 ;
  assign y15846 = ~1'b0 ;
  assign y15847 = n39259 ;
  assign y15848 = ~n39263 ;
  assign y15849 = ~1'b0 ;
  assign y15850 = n39267 ;
  assign y15851 = n39276 ;
  assign y15852 = ~n39278 ;
  assign y15853 = ~n39280 ;
  assign y15854 = n39285 ;
  assign y15855 = ~n39287 ;
  assign y15856 = ~n39289 ;
  assign y15857 = n39295 ;
  assign y15858 = ~1'b0 ;
  assign y15859 = ~n39296 ;
  assign y15860 = ~n39301 ;
  assign y15861 = n39302 ;
  assign y15862 = n39304 ;
  assign y15863 = ~1'b0 ;
  assign y15864 = ~1'b0 ;
  assign y15865 = n39307 ;
  assign y15866 = ~1'b0 ;
  assign y15867 = ~n39312 ;
  assign y15868 = n39316 ;
  assign y15869 = n39318 ;
  assign y15870 = ~n39319 ;
  assign y15871 = n39323 ;
  assign y15872 = n39327 ;
  assign y15873 = n39330 ;
  assign y15874 = ~1'b0 ;
  assign y15875 = ~n39332 ;
  assign y15876 = ~n39335 ;
  assign y15877 = ~n39341 ;
  assign y15878 = ~n8658 ;
  assign y15879 = n37021 ;
  assign y15880 = n39343 ;
  assign y15881 = n39346 ;
  assign y15882 = ~1'b0 ;
  assign y15883 = n39347 ;
  assign y15884 = ~n39350 ;
  assign y15885 = ~n39351 ;
  assign y15886 = ~n39356 ;
  assign y15887 = n39360 ;
  assign y15888 = ~n39361 ;
  assign y15889 = ~n39362 ;
  assign y15890 = ~1'b0 ;
  assign y15891 = ~1'b0 ;
  assign y15892 = ~n39367 ;
  assign y15893 = ~n39371 ;
  assign y15894 = ~n24464 ;
  assign y15895 = ~n39374 ;
  assign y15896 = ~n39375 ;
  assign y15897 = n39377 ;
  assign y15898 = ~n39379 ;
  assign y15899 = ~1'b0 ;
  assign y15900 = ~n39380 ;
  assign y15901 = ~1'b0 ;
  assign y15902 = n39383 ;
  assign y15903 = ~n39386 ;
  assign y15904 = ~n39387 ;
  assign y15905 = n39390 ;
  assign y15906 = n3107 ;
  assign y15907 = ~1'b0 ;
  assign y15908 = ~n39392 ;
  assign y15909 = n39395 ;
  assign y15910 = ~n39396 ;
  assign y15911 = ~1'b0 ;
  assign y15912 = ~n39401 ;
  assign y15913 = ~1'b0 ;
  assign y15914 = n39403 ;
  assign y15915 = ~n39404 ;
  assign y15916 = ~n39407 ;
  assign y15917 = n39408 ;
  assign y15918 = ~n39409 ;
  assign y15919 = ~n39411 ;
  assign y15920 = ~1'b0 ;
  assign y15921 = ~1'b0 ;
  assign y15922 = n39413 ;
  assign y15923 = n39416 ;
  assign y15924 = n39419 ;
  assign y15925 = n39421 ;
  assign y15926 = ~n39425 ;
  assign y15927 = n39427 ;
  assign y15928 = n39431 ;
  assign y15929 = ~n39434 ;
  assign y15930 = n39435 ;
  assign y15931 = ~n39437 ;
  assign y15932 = ~n39438 ;
  assign y15933 = ~n39440 ;
  assign y15934 = ~n39441 ;
  assign y15935 = ~1'b0 ;
  assign y15936 = n39442 ;
  assign y15937 = ~n39445 ;
  assign y15938 = n39446 ;
  assign y15939 = ~n39448 ;
  assign y15940 = ~n39450 ;
  assign y15941 = ~n39451 ;
  assign y15942 = ~n39456 ;
  assign y15943 = n39462 ;
  assign y15944 = ~n39464 ;
  assign y15945 = ~1'b0 ;
  assign y15946 = ~1'b0 ;
  assign y15947 = ~n39467 ;
  assign y15948 = n39468 ;
  assign y15949 = n39469 ;
  assign y15950 = ~n39470 ;
  assign y15951 = n7873 ;
  assign y15952 = ~1'b0 ;
  assign y15953 = ~1'b0 ;
  assign y15954 = n39471 ;
  assign y15955 = ~1'b0 ;
  assign y15956 = ~n39474 ;
  assign y15957 = n39475 ;
  assign y15958 = ~n39476 ;
  assign y15959 = n39478 ;
  assign y15960 = ~n39481 ;
  assign y15961 = ~n39483 ;
  assign y15962 = n39484 ;
  assign y15963 = n39489 ;
  assign y15964 = ~n39492 ;
  assign y15965 = 1'b0 ;
  assign y15966 = n39496 ;
  assign y15967 = n37095 ;
  assign y15968 = ~n39497 ;
  assign y15969 = n39498 ;
  assign y15970 = ~n39501 ;
  assign y15971 = ~1'b0 ;
  assign y15972 = ~n39503 ;
  assign y15973 = ~1'b0 ;
  assign y15974 = n39505 ;
  assign y15975 = ~n39507 ;
  assign y15976 = ~n39508 ;
  assign y15977 = n39514 ;
  assign y15978 = ~1'b0 ;
  assign y15979 = ~1'b0 ;
  assign y15980 = n39516 ;
  assign y15981 = ~n39519 ;
  assign y15982 = n39525 ;
  assign y15983 = ~1'b0 ;
  assign y15984 = ~n39532 ;
  assign y15985 = ~1'b0 ;
  assign y15986 = ~n39533 ;
  assign y15987 = n39535 ;
  assign y15988 = n39537 ;
  assign y15989 = ~n39540 ;
  assign y15990 = ~1'b0 ;
  assign y15991 = n39544 ;
  assign y15992 = ~n39545 ;
  assign y15993 = ~1'b0 ;
  assign y15994 = ~1'b0 ;
  assign y15995 = n39549 ;
  assign y15996 = ~n39552 ;
  assign y15997 = ~n39554 ;
  assign y15998 = n39555 ;
  assign y15999 = n39557 ;
  assign y16000 = n34525 ;
  assign y16001 = ~n39559 ;
  assign y16002 = n39560 ;
  assign y16003 = n39565 ;
  assign y16004 = ~n39569 ;
  assign y16005 = n39575 ;
  assign y16006 = ~1'b0 ;
  assign y16007 = ~n39580 ;
  assign y16008 = n39582 ;
  assign y16009 = n39584 ;
  assign y16010 = n39585 ;
  assign y16011 = n6321 ;
  assign y16012 = ~1'b0 ;
  assign y16013 = ~1'b0 ;
  assign y16014 = ~1'b0 ;
  assign y16015 = n39587 ;
  assign y16016 = ~1'b0 ;
  assign y16017 = ~n39589 ;
  assign y16018 = n39590 ;
  assign y16019 = n39591 ;
  assign y16020 = ~1'b0 ;
  assign y16021 = n39594 ;
  assign y16022 = ~1'b0 ;
  assign y16023 = ~1'b0 ;
  assign y16024 = ~1'b0 ;
  assign y16025 = n39602 ;
  assign y16026 = ~1'b0 ;
  assign y16027 = n39605 ;
  assign y16028 = ~n39606 ;
  assign y16029 = ~n39611 ;
  assign y16030 = n39614 ;
  assign y16031 = ~n39616 ;
  assign y16032 = n39617 ;
  assign y16033 = ~1'b0 ;
  assign y16034 = ~n9000 ;
  assign y16035 = n39622 ;
  assign y16036 = 1'b0 ;
  assign y16037 = ~n39623 ;
  assign y16038 = ~n39625 ;
  assign y16039 = n39626 ;
  assign y16040 = ~1'b0 ;
  assign y16041 = n39631 ;
  assign y16042 = ~1'b0 ;
  assign y16043 = n39633 ;
  assign y16044 = ~n39635 ;
  assign y16045 = ~n39643 ;
  assign y16046 = ~1'b0 ;
  assign y16047 = ~1'b0 ;
  assign y16048 = ~n39644 ;
  assign y16049 = ~1'b0 ;
  assign y16050 = ~n39646 ;
  assign y16051 = n39647 ;
  assign y16052 = n39650 ;
  assign y16053 = ~n39654 ;
  assign y16054 = ~n39655 ;
  assign y16055 = ~1'b0 ;
  assign y16056 = ~1'b0 ;
  assign y16057 = ~1'b0 ;
  assign y16058 = ~n39656 ;
  assign y16059 = n39658 ;
  assign y16060 = ~n39660 ;
  assign y16061 = n39661 ;
  assign y16062 = ~1'b0 ;
  assign y16063 = ~1'b0 ;
  assign y16064 = n39663 ;
  assign y16065 = n39670 ;
  assign y16066 = n39672 ;
  assign y16067 = ~1'b0 ;
  assign y16068 = ~1'b0 ;
  assign y16069 = n39677 ;
  assign y16070 = n39678 ;
  assign y16071 = ~n39682 ;
  assign y16072 = n39685 ;
  assign y16073 = n39695 ;
  assign y16074 = ~1'b0 ;
  assign y16075 = ~n39698 ;
  assign y16076 = n39699 ;
  assign y16077 = n39700 ;
  assign y16078 = n39701 ;
  assign y16079 = ~n36710 ;
  assign y16080 = ~n39703 ;
  assign y16081 = n39704 ;
  assign y16082 = ~n39706 ;
  assign y16083 = 1'b0 ;
  assign y16084 = n39708 ;
  assign y16085 = ~n39711 ;
  assign y16086 = ~1'b0 ;
  assign y16087 = ~n39713 ;
  assign y16088 = ~n39714 ;
  assign y16089 = ~n39722 ;
  assign y16090 = ~n39723 ;
  assign y16091 = ~n39728 ;
  assign y16092 = n39729 ;
  assign y16093 = ~1'b0 ;
  assign y16094 = n39730 ;
  assign y16095 = n39736 ;
  assign y16096 = ~n39739 ;
  assign y16097 = ~n39740 ;
  assign y16098 = n39741 ;
  assign y16099 = ~n39748 ;
  assign y16100 = ~n39749 ;
  assign y16101 = n39755 ;
  assign y16102 = ~1'b0 ;
  assign y16103 = n5199 ;
  assign y16104 = n39757 ;
  assign y16105 = ~n39763 ;
  assign y16106 = n39767 ;
  assign y16107 = ~n39771 ;
  assign y16108 = ~n39773 ;
  assign y16109 = ~n39775 ;
  assign y16110 = n39780 ;
  assign y16111 = ~n39783 ;
  assign y16112 = n39785 ;
  assign y16113 = n39786 ;
  assign y16114 = ~n39788 ;
  assign y16115 = n39790 ;
  assign y16116 = ~n39791 ;
  assign y16117 = ~n39794 ;
  assign y16118 = ~n39797 ;
  assign y16119 = ~n39801 ;
  assign y16120 = ~1'b0 ;
  assign y16121 = ~n39806 ;
  assign y16122 = n39808 ;
  assign y16123 = n39811 ;
  assign y16124 = n39813 ;
  assign y16125 = ~1'b0 ;
  assign y16126 = n39814 ;
  assign y16127 = n39815 ;
  assign y16128 = n16661 ;
  assign y16129 = n39816 ;
  assign y16130 = n39819 ;
  assign y16131 = ~n39821 ;
  assign y16132 = ~n39822 ;
  assign y16133 = ~n39829 ;
  assign y16134 = ~1'b0 ;
  assign y16135 = ~n39831 ;
  assign y16136 = n39834 ;
  assign y16137 = ~n39838 ;
  assign y16138 = ~n39844 ;
  assign y16139 = ~1'b0 ;
  assign y16140 = ~n39852 ;
  assign y16141 = 1'b0 ;
  assign y16142 = n39854 ;
  assign y16143 = ~1'b0 ;
  assign y16144 = ~n39856 ;
  assign y16145 = ~1'b0 ;
  assign y16146 = n39857 ;
  assign y16147 = ~n39867 ;
  assign y16148 = ~1'b0 ;
  assign y16149 = n39870 ;
  assign y16150 = ~n39872 ;
  assign y16151 = ~1'b0 ;
  assign y16152 = ~1'b0 ;
  assign y16153 = ~n39876 ;
  assign y16154 = ~n39877 ;
  assign y16155 = ~n39878 ;
  assign y16156 = 1'b0 ;
  assign y16157 = n39882 ;
  assign y16158 = ~n39885 ;
  assign y16159 = n39887 ;
  assign y16160 = n39889 ;
  assign y16161 = 1'b0 ;
  assign y16162 = n39890 ;
  assign y16163 = n39892 ;
  assign y16164 = n39893 ;
  assign y16165 = ~n39894 ;
  assign y16166 = ~n39897 ;
  assign y16167 = n39899 ;
  assign y16168 = ~1'b0 ;
  assign y16169 = ~1'b0 ;
  assign y16170 = n39906 ;
  assign y16171 = n39909 ;
  assign y16172 = n39911 ;
  assign y16173 = ~1'b0 ;
  assign y16174 = ~n39913 ;
  assign y16175 = n39915 ;
  assign y16176 = n39921 ;
  assign y16177 = ~1'b0 ;
  assign y16178 = n39926 ;
  assign y16179 = n39927 ;
  assign y16180 = ~n39930 ;
  assign y16181 = ~n39931 ;
  assign y16182 = ~n39932 ;
  assign y16183 = ~n39933 ;
  assign y16184 = ~n39937 ;
  assign y16185 = ~1'b0 ;
  assign y16186 = n39942 ;
  assign y16187 = n39944 ;
  assign y16188 = n39946 ;
  assign y16189 = ~n39947 ;
  assign y16190 = ~n39948 ;
  assign y16191 = n39950 ;
  assign y16192 = ~n39953 ;
  assign y16193 = ~1'b0 ;
  assign y16194 = ~1'b0 ;
  assign y16195 = ~n39956 ;
  assign y16196 = ~n4202 ;
  assign y16197 = n39957 ;
  assign y16198 = n39960 ;
  assign y16199 = ~1'b0 ;
  assign y16200 = ~1'b0 ;
  assign y16201 = n39961 ;
  assign y16202 = ~1'b0 ;
  assign y16203 = ~n39962 ;
  assign y16204 = 1'b0 ;
  assign y16205 = n39964 ;
  assign y16206 = ~n39966 ;
  assign y16207 = ~1'b0 ;
  assign y16208 = ~n39967 ;
  assign y16209 = ~1'b0 ;
  assign y16210 = ~n39968 ;
  assign y16211 = ~n39970 ;
  assign y16212 = ~n39972 ;
  assign y16213 = ~n39975 ;
  assign y16214 = n39976 ;
  assign y16215 = ~n39977 ;
  assign y16216 = ~1'b0 ;
  assign y16217 = n39978 ;
  assign y16218 = n39980 ;
  assign y16219 = ~n39982 ;
  assign y16220 = n39985 ;
  assign y16221 = ~n39986 ;
  assign y16222 = n39987 ;
  assign y16223 = ~n39993 ;
  assign y16224 = ~n39994 ;
  assign y16225 = ~n39995 ;
  assign y16226 = n32763 ;
  assign y16227 = ~1'b0 ;
  assign y16228 = n39996 ;
  assign y16229 = n39997 ;
  assign y16230 = ~n39999 ;
  assign y16231 = ~1'b0 ;
  assign y16232 = ~1'b0 ;
  assign y16233 = ~n40001 ;
  assign y16234 = n40002 ;
  assign y16235 = n40003 ;
  assign y16236 = n40004 ;
  assign y16237 = n1725 ;
  assign y16238 = ~n40006 ;
  assign y16239 = ~n40007 ;
  assign y16240 = ~n40010 ;
  assign y16241 = ~n40011 ;
  assign y16242 = ~n40018 ;
  assign y16243 = n40020 ;
  assign y16244 = n40021 ;
  assign y16245 = ~n40025 ;
  assign y16246 = n40026 ;
  assign y16247 = n40028 ;
  assign y16248 = ~n40029 ;
  assign y16249 = n40031 ;
  assign y16250 = ~1'b0 ;
  assign y16251 = ~1'b0 ;
  assign y16252 = ~n40033 ;
  assign y16253 = n6179 ;
  assign y16254 = ~1'b0 ;
  assign y16255 = ~n40036 ;
  assign y16256 = ~n40037 ;
  assign y16257 = n40038 ;
  assign y16258 = ~1'b0 ;
  assign y16259 = ~n40047 ;
  assign y16260 = n40048 ;
  assign y16261 = n40049 ;
  assign y16262 = n40054 ;
  assign y16263 = ~1'b0 ;
  assign y16264 = n40055 ;
  assign y16265 = ~n40056 ;
  assign y16266 = n40057 ;
  assign y16267 = ~n40059 ;
  assign y16268 = ~n40061 ;
  assign y16269 = ~1'b0 ;
  assign y16270 = n40064 ;
  assign y16271 = n40068 ;
  assign y16272 = ~n40072 ;
  assign y16273 = n40075 ;
  assign y16274 = ~n40077 ;
  assign y16275 = ~1'b0 ;
  assign y16276 = n40078 ;
  assign y16277 = n40085 ;
  assign y16278 = ~1'b0 ;
  assign y16279 = n40091 ;
  assign y16280 = n40092 ;
  assign y16281 = ~n40093 ;
  assign y16282 = ~1'b0 ;
  assign y16283 = ~n40094 ;
  assign y16284 = n40096 ;
  assign y16285 = ~n40098 ;
  assign y16286 = n40101 ;
  assign y16287 = ~n40104 ;
  assign y16288 = ~n40109 ;
  assign y16289 = ~n40110 ;
  assign y16290 = ~1'b0 ;
  assign y16291 = n40113 ;
  assign y16292 = n40115 ;
  assign y16293 = n40117 ;
  assign y16294 = ~n40119 ;
  assign y16295 = ~n40130 ;
  assign y16296 = n40135 ;
  assign y16297 = n40139 ;
  assign y16298 = ~1'b0 ;
  assign y16299 = n40144 ;
  assign y16300 = ~1'b0 ;
  assign y16301 = n40150 ;
  assign y16302 = ~1'b0 ;
  assign y16303 = ~n40152 ;
  assign y16304 = ~n40153 ;
  assign y16305 = ~n40159 ;
  assign y16306 = ~1'b0 ;
  assign y16307 = n40161 ;
  assign y16308 = n40162 ;
  assign y16309 = n40163 ;
  assign y16310 = ~1'b0 ;
  assign y16311 = n40167 ;
  assign y16312 = ~n40168 ;
  assign y16313 = ~n40169 ;
  assign y16314 = n40170 ;
  assign y16315 = n40172 ;
  assign y16316 = n40175 ;
  assign y16317 = n40178 ;
  assign y16318 = ~n40180 ;
  assign y16319 = n40185 ;
  assign y16320 = n1367 ;
  assign y16321 = ~1'b0 ;
  assign y16322 = n40187 ;
  assign y16323 = ~n40190 ;
  assign y16324 = ~n31995 ;
  assign y16325 = ~n40192 ;
  assign y16326 = n40195 ;
  assign y16327 = ~n40198 ;
  assign y16328 = ~n40200 ;
  assign y16329 = n40201 ;
  assign y16330 = ~1'b0 ;
  assign y16331 = ~n40202 ;
  assign y16332 = ~n40205 ;
  assign y16333 = ~1'b0 ;
  assign y16334 = n40206 ;
  assign y16335 = ~1'b0 ;
  assign y16336 = ~n40207 ;
  assign y16337 = ~n40209 ;
  assign y16338 = ~1'b0 ;
  assign y16339 = n40211 ;
  assign y16340 = n21339 ;
  assign y16341 = ~n40213 ;
  assign y16342 = n40216 ;
  assign y16343 = ~1'b0 ;
  assign y16344 = n40217 ;
  assign y16345 = ~n40218 ;
  assign y16346 = ~n40226 ;
  assign y16347 = n40227 ;
  assign y16348 = ~n40228 ;
  assign y16349 = n40230 ;
  assign y16350 = ~1'b0 ;
  assign y16351 = ~n40232 ;
  assign y16352 = n40233 ;
  assign y16353 = ~1'b0 ;
  assign y16354 = ~n40234 ;
  assign y16355 = ~n11909 ;
  assign y16356 = n40237 ;
  assign y16357 = ~1'b0 ;
  assign y16358 = ~1'b0 ;
  assign y16359 = ~n40241 ;
  assign y16360 = ~1'b0 ;
  assign y16361 = ~1'b0 ;
  assign y16362 = n40244 ;
  assign y16363 = n40245 ;
  assign y16364 = ~n40246 ;
  assign y16365 = ~n40247 ;
  assign y16366 = ~1'b0 ;
  assign y16367 = n40252 ;
  assign y16368 = ~1'b0 ;
  assign y16369 = n40255 ;
  assign y16370 = n33651 ;
  assign y16371 = n40257 ;
  assign y16372 = ~n40260 ;
  assign y16373 = n30355 ;
  assign y16374 = ~1'b0 ;
  assign y16375 = ~n40262 ;
  assign y16376 = ~1'b0 ;
  assign y16377 = ~n40265 ;
  assign y16378 = n40271 ;
  assign y16379 = ~1'b0 ;
  assign y16380 = ~1'b0 ;
  assign y16381 = n40272 ;
  assign y16382 = ~1'b0 ;
  assign y16383 = n40273 ;
  assign y16384 = n40275 ;
  assign y16385 = n40278 ;
  assign y16386 = ~n40282 ;
  assign y16387 = ~n40285 ;
  assign y16388 = ~n40287 ;
  assign y16389 = n40289 ;
  assign y16390 = ~n40291 ;
  assign y16391 = n40296 ;
  assign y16392 = ~n40297 ;
  assign y16393 = ~n40299 ;
  assign y16394 = n40300 ;
  assign y16395 = n40301 ;
  assign y16396 = n40302 ;
  assign y16397 = ~n40306 ;
  assign y16398 = ~n40308 ;
  assign y16399 = n40309 ;
  assign y16400 = n40311 ;
  assign y16401 = ~n40313 ;
  assign y16402 = n40316 ;
  assign y16403 = n40317 ;
  assign y16404 = ~n40318 ;
  assign y16405 = ~1'b0 ;
  assign y16406 = ~n40323 ;
  assign y16407 = ~1'b0 ;
  assign y16408 = n40327 ;
  assign y16409 = ~n27268 ;
  assign y16410 = n23581 ;
  assign y16411 = n40330 ;
  assign y16412 = n40333 ;
  assign y16413 = ~n40334 ;
  assign y16414 = ~1'b0 ;
  assign y16415 = ~1'b0 ;
  assign y16416 = n40338 ;
  assign y16417 = ~n40340 ;
  assign y16418 = n40341 ;
  assign y16419 = ~n40342 ;
  assign y16420 = ~n40343 ;
  assign y16421 = ~n40345 ;
  assign y16422 = ~n30307 ;
  assign y16423 = n40351 ;
  assign y16424 = n40353 ;
  assign y16425 = ~n40354 ;
  assign y16426 = ~n16325 ;
  assign y16427 = ~n34605 ;
  assign y16428 = n40357 ;
  assign y16429 = ~n40358 ;
  assign y16430 = n40359 ;
  assign y16431 = n40360 ;
  assign y16432 = n40361 ;
  assign y16433 = n1925 ;
  assign y16434 = n1579 ;
  assign y16435 = ~n40362 ;
  assign y16436 = ~n40367 ;
  assign y16437 = ~n40371 ;
  assign y16438 = ~1'b0 ;
  assign y16439 = ~n40373 ;
  assign y16440 = ~1'b0 ;
  assign y16441 = ~1'b0 ;
  assign y16442 = n40374 ;
  assign y16443 = ~n40376 ;
  assign y16444 = ~n40377 ;
  assign y16445 = n40380 ;
  assign y16446 = n40381 ;
  assign y16447 = ~n40388 ;
  assign y16448 = ~n40391 ;
  assign y16449 = ~1'b0 ;
  assign y16450 = ~1'b0 ;
  assign y16451 = n40401 ;
  assign y16452 = ~n40402 ;
  assign y16453 = ~n40403 ;
  assign y16454 = ~n40407 ;
  assign y16455 = n40410 ;
  assign y16456 = ~n40413 ;
  assign y16457 = ~n40414 ;
  assign y16458 = n40416 ;
  assign y16459 = n40417 ;
  assign y16460 = 1'b0 ;
  assign y16461 = ~n40420 ;
  assign y16462 = ~n40422 ;
  assign y16463 = ~n40426 ;
  assign y16464 = ~n40428 ;
  assign y16465 = n40431 ;
  assign y16466 = ~1'b0 ;
  assign y16467 = ~1'b0 ;
  assign y16468 = n40432 ;
  assign y16469 = n40433 ;
  assign y16470 = ~n40437 ;
  assign y16471 = n40441 ;
  assign y16472 = n40448 ;
  assign y16473 = ~1'b0 ;
  assign y16474 = ~1'b0 ;
  assign y16475 = ~1'b0 ;
  assign y16476 = n40450 ;
  assign y16477 = n40451 ;
  assign y16478 = ~n40452 ;
  assign y16479 = ~n40453 ;
  assign y16480 = ~n40457 ;
  assign y16481 = ~1'b0 ;
  assign y16482 = n40463 ;
  assign y16483 = ~1'b0 ;
  assign y16484 = n40465 ;
  assign y16485 = ~1'b0 ;
  assign y16486 = ~n28991 ;
  assign y16487 = ~n40468 ;
  assign y16488 = n40472 ;
  assign y16489 = ~n40477 ;
  assign y16490 = ~n40478 ;
  assign y16491 = ~n40480 ;
  assign y16492 = n40484 ;
  assign y16493 = n40486 ;
  assign y16494 = ~n40493 ;
  assign y16495 = n40494 ;
  assign y16496 = n26696 ;
  assign y16497 = ~n40495 ;
  assign y16498 = ~n40497 ;
  assign y16499 = ~1'b0 ;
  assign y16500 = n40502 ;
  assign y16501 = ~1'b0 ;
  assign y16502 = n40503 ;
  assign y16503 = ~n40505 ;
  assign y16504 = n31769 ;
  assign y16505 = ~1'b0 ;
  assign y16506 = ~1'b0 ;
  assign y16507 = n40507 ;
  assign y16508 = n32898 ;
  assign y16509 = ~n40509 ;
  assign y16510 = ~1'b0 ;
  assign y16511 = ~n40513 ;
  assign y16512 = ~n40517 ;
  assign y16513 = ~n40518 ;
  assign y16514 = ~1'b0 ;
  assign y16515 = ~n40520 ;
  assign y16516 = ~1'b0 ;
  assign y16517 = ~n40522 ;
  assign y16518 = ~n40526 ;
  assign y16519 = n40529 ;
  assign y16520 = n40536 ;
  assign y16521 = ~n40538 ;
  assign y16522 = ~n40541 ;
  assign y16523 = n40543 ;
  assign y16524 = ~1'b0 ;
  assign y16525 = ~n40545 ;
  assign y16526 = ~n40552 ;
  assign y16527 = ~n40557 ;
  assign y16528 = n40558 ;
  assign y16529 = n40559 ;
  assign y16530 = n40563 ;
  assign y16531 = n40565 ;
  assign y16532 = n40567 ;
  assign y16533 = n18600 ;
  assign y16534 = ~1'b0 ;
  assign y16535 = n40568 ;
  assign y16536 = ~n40570 ;
  assign y16537 = ~n40574 ;
  assign y16538 = ~n40575 ;
  assign y16539 = 1'b0 ;
  assign y16540 = n40576 ;
  assign y16541 = ~n40578 ;
  assign y16542 = n40582 ;
  assign y16543 = n40584 ;
  assign y16544 = n40586 ;
  assign y16545 = n40590 ;
  assign y16546 = ~n40591 ;
  assign y16547 = ~n21692 ;
  assign y16548 = ~n40592 ;
  assign y16549 = n40594 ;
  assign y16550 = n40598 ;
  assign y16551 = ~n40599 ;
  assign y16552 = ~1'b0 ;
  assign y16553 = n2992 ;
  assign y16554 = ~n40600 ;
  assign y16555 = ~n40601 ;
  assign y16556 = ~n40602 ;
  assign y16557 = n2094 ;
  assign y16558 = ~1'b0 ;
  assign y16559 = n40607 ;
  assign y16560 = ~1'b0 ;
  assign y16561 = ~n40608 ;
  assign y16562 = ~n40610 ;
  assign y16563 = ~n40611 ;
  assign y16564 = ~n40612 ;
  assign y16565 = ~n40614 ;
  assign y16566 = n40617 ;
  assign y16567 = ~n40618 ;
  assign y16568 = ~1'b0 ;
  assign y16569 = ~1'b0 ;
  assign y16570 = ~n40620 ;
  assign y16571 = ~n40625 ;
  assign y16572 = n40627 ;
  assign y16573 = ~n40629 ;
  assign y16574 = ~1'b0 ;
  assign y16575 = n40630 ;
  assign y16576 = ~n40631 ;
  assign y16577 = ~n40632 ;
  assign y16578 = ~n40635 ;
  assign y16579 = ~n40637 ;
  assign y16580 = n40640 ;
  assign y16581 = ~1'b0 ;
  assign y16582 = ~n40643 ;
  assign y16583 = n40646 ;
  assign y16584 = n40647 ;
  assign y16585 = ~n40654 ;
  assign y16586 = ~n40657 ;
  assign y16587 = ~n40658 ;
  assign y16588 = n40661 ;
  assign y16589 = n40663 ;
  assign y16590 = ~1'b0 ;
  assign y16591 = ~n40665 ;
  assign y16592 = ~n40672 ;
  assign y16593 = ~1'b0 ;
  assign y16594 = n40675 ;
  assign y16595 = ~n40676 ;
  assign y16596 = n40679 ;
  assign y16597 = ~n40681 ;
  assign y16598 = ~1'b0 ;
  assign y16599 = n40683 ;
  assign y16600 = n40687 ;
  assign y16601 = ~1'b0 ;
  assign y16602 = ~n40691 ;
  assign y16603 = n40698 ;
  assign y16604 = ~n40700 ;
  assign y16605 = ~n40701 ;
  assign y16606 = n40702 ;
  assign y16607 = ~1'b0 ;
  assign y16608 = ~n40704 ;
  assign y16609 = n40706 ;
  assign y16610 = ~n40711 ;
  assign y16611 = n40712 ;
  assign y16612 = ~n40715 ;
  assign y16613 = n40718 ;
  assign y16614 = ~n40719 ;
  assign y16615 = ~1'b0 ;
  assign y16616 = ~1'b0 ;
  assign y16617 = ~n40720 ;
  assign y16618 = ~n40722 ;
  assign y16619 = n40723 ;
  assign y16620 = ~1'b0 ;
  assign y16621 = ~1'b0 ;
  assign y16622 = ~1'b0 ;
  assign y16623 = 1'b0 ;
  assign y16624 = ~n40725 ;
  assign y16625 = ~1'b0 ;
  assign y16626 = n40726 ;
  assign y16627 = ~n40730 ;
  assign y16628 = ~1'b0 ;
  assign y16629 = ~n40732 ;
  assign y16630 = ~n40733 ;
  assign y16631 = ~1'b0 ;
  assign y16632 = n40734 ;
  assign y16633 = n40739 ;
  assign y16634 = n40741 ;
  assign y16635 = ~n40744 ;
  assign y16636 = ~1'b0 ;
  assign y16637 = ~1'b0 ;
  assign y16638 = ~1'b0 ;
  assign y16639 = n40745 ;
  assign y16640 = ~1'b0 ;
  assign y16641 = ~1'b0 ;
  assign y16642 = n40746 ;
  assign y16643 = ~n40748 ;
  assign y16644 = ~n40750 ;
  assign y16645 = n40752 ;
  assign y16646 = ~n40755 ;
  assign y16647 = ~1'b0 ;
  assign y16648 = ~n40757 ;
  assign y16649 = n40760 ;
  assign y16650 = ~n40763 ;
  assign y16651 = ~n40769 ;
  assign y16652 = ~1'b0 ;
  assign y16653 = n40771 ;
  assign y16654 = ~n40775 ;
  assign y16655 = n40776 ;
  assign y16656 = ~1'b0 ;
  assign y16657 = ~n40777 ;
  assign y16658 = n40778 ;
  assign y16659 = ~n40779 ;
  assign y16660 = ~n40781 ;
  assign y16661 = ~n40785 ;
  assign y16662 = n40787 ;
  assign y16663 = ~1'b0 ;
  assign y16664 = n40788 ;
  assign y16665 = n40791 ;
  assign y16666 = ~1'b0 ;
  assign y16667 = n40792 ;
  assign y16668 = n40793 ;
  assign y16669 = ~n40794 ;
  assign y16670 = n40795 ;
  assign y16671 = ~1'b0 ;
  assign y16672 = ~1'b0 ;
  assign y16673 = ~n40797 ;
  assign y16674 = n40801 ;
  assign y16675 = n40802 ;
  assign y16676 = n40804 ;
  assign y16677 = n40807 ;
  assign y16678 = n6644 ;
  assign y16679 = n40808 ;
  assign y16680 = ~n40815 ;
  assign y16681 = n38629 ;
  assign y16682 = ~n40818 ;
  assign y16683 = ~1'b0 ;
  assign y16684 = ~1'b0 ;
  assign y16685 = ~n12541 ;
  assign y16686 = ~n40819 ;
  assign y16687 = ~n40820 ;
  assign y16688 = ~n40823 ;
  assign y16689 = ~n40825 ;
  assign y16690 = ~1'b0 ;
  assign y16691 = n40829 ;
  assign y16692 = n40837 ;
  assign y16693 = ~n40840 ;
  assign y16694 = n40848 ;
  assign y16695 = ~n40854 ;
  assign y16696 = ~n40858 ;
  assign y16697 = ~n40860 ;
  assign y16698 = ~1'b0 ;
  assign y16699 = ~1'b0 ;
  assign y16700 = n40867 ;
  assign y16701 = ~1'b0 ;
  assign y16702 = ~n40872 ;
  assign y16703 = ~1'b0 ;
  assign y16704 = n40873 ;
  assign y16705 = ~n40879 ;
  assign y16706 = ~1'b0 ;
  assign y16707 = ~1'b0 ;
  assign y16708 = ~1'b0 ;
  assign y16709 = n40881 ;
  assign y16710 = ~n40883 ;
  assign y16711 = n40884 ;
  assign y16712 = n40886 ;
  assign y16713 = n40889 ;
  assign y16714 = ~1'b0 ;
  assign y16715 = ~1'b0 ;
  assign y16716 = n40891 ;
  assign y16717 = n40894 ;
  assign y16718 = ~1'b0 ;
  assign y16719 = n40897 ;
  assign y16720 = n40901 ;
  assign y16721 = n40904 ;
  assign y16722 = ~n40905 ;
  assign y16723 = n40907 ;
  assign y16724 = n40911 ;
  assign y16725 = ~n40916 ;
  assign y16726 = n40917 ;
  assign y16727 = n40921 ;
  assign y16728 = n40922 ;
  assign y16729 = ~n40923 ;
  assign y16730 = n40927 ;
  assign y16731 = ~n40931 ;
  assign y16732 = n40933 ;
  assign y16733 = ~1'b0 ;
  assign y16734 = n40935 ;
  assign y16735 = n40936 ;
  assign y16736 = ~n40939 ;
  assign y16737 = n40941 ;
  assign y16738 = n40942 ;
  assign y16739 = n40944 ;
  assign y16740 = n33200 ;
  assign y16741 = ~n40946 ;
  assign y16742 = n40948 ;
  assign y16743 = n40956 ;
  assign y16744 = ~1'b0 ;
  assign y16745 = ~n40960 ;
  assign y16746 = ~1'b0 ;
  assign y16747 = n40961 ;
  assign y16748 = ~n40966 ;
  assign y16749 = ~1'b0 ;
  assign y16750 = n7842 ;
  assign y16751 = n40967 ;
  assign y16752 = ~n40971 ;
  assign y16753 = ~n25040 ;
  assign y16754 = ~n40975 ;
  assign y16755 = n40976 ;
  assign y16756 = ~1'b0 ;
  assign y16757 = ~1'b0 ;
  assign y16758 = ~1'b0 ;
  assign y16759 = ~1'b0 ;
  assign y16760 = n40979 ;
  assign y16761 = ~n40981 ;
  assign y16762 = ~n40982 ;
  assign y16763 = ~n40984 ;
  assign y16764 = ~n40985 ;
  assign y16765 = ~n40986 ;
  assign y16766 = ~n40987 ;
  assign y16767 = ~n40989 ;
  assign y16768 = ~1'b0 ;
  assign y16769 = ~n40990 ;
  assign y16770 = ~n40991 ;
  assign y16771 = n40995 ;
  assign y16772 = ~1'b0 ;
  assign y16773 = ~n40998 ;
  assign y16774 = ~n40999 ;
  assign y16775 = ~1'b0 ;
  assign y16776 = ~n41000 ;
  assign y16777 = ~n41007 ;
  assign y16778 = ~n41008 ;
  assign y16779 = ~n41016 ;
  assign y16780 = n41018 ;
  assign y16781 = ~1'b0 ;
  assign y16782 = n41020 ;
  assign y16783 = ~1'b0 ;
  assign y16784 = ~n41023 ;
  assign y16785 = n41025 ;
  assign y16786 = n41029 ;
  assign y16787 = ~1'b0 ;
  assign y16788 = ~1'b0 ;
  assign y16789 = ~1'b0 ;
  assign y16790 = ~n41031 ;
  assign y16791 = ~n41032 ;
  assign y16792 = n41033 ;
  assign y16793 = ~n41035 ;
  assign y16794 = ~n41036 ;
  assign y16795 = n41039 ;
  assign y16796 = ~n41041 ;
  assign y16797 = n41044 ;
  assign y16798 = ~n41047 ;
  assign y16799 = n41049 ;
  assign y16800 = ~n41052 ;
  assign y16801 = n41054 ;
  assign y16802 = n41058 ;
  assign y16803 = n41060 ;
  assign y16804 = ~1'b0 ;
  assign y16805 = ~n41069 ;
  assign y16806 = ~n41070 ;
  assign y16807 = ~n41075 ;
  assign y16808 = n41077 ;
  assign y16809 = n41078 ;
  assign y16810 = ~1'b0 ;
  assign y16811 = n41079 ;
  assign y16812 = n41084 ;
  assign y16813 = ~1'b0 ;
  assign y16814 = ~1'b0 ;
  assign y16815 = n41085 ;
  assign y16816 = ~n41095 ;
  assign y16817 = n41096 ;
  assign y16818 = ~n41098 ;
  assign y16819 = ~1'b0 ;
  assign y16820 = n41100 ;
  assign y16821 = n41102 ;
  assign y16822 = ~n41107 ;
  assign y16823 = ~n41109 ;
  assign y16824 = n41111 ;
  assign y16825 = ~1'b0 ;
  assign y16826 = ~1'b0 ;
  assign y16827 = ~n41115 ;
  assign y16828 = ~n41116 ;
  assign y16829 = ~n41118 ;
  assign y16830 = ~1'b0 ;
  assign y16831 = n41119 ;
  assign y16832 = ~n41122 ;
  assign y16833 = ~n41125 ;
  assign y16834 = ~n41128 ;
  assign y16835 = ~1'b0 ;
  assign y16836 = n41129 ;
  assign y16837 = ~n41131 ;
  assign y16838 = ~n41134 ;
  assign y16839 = n41135 ;
  assign y16840 = ~1'b0 ;
  assign y16841 = ~n19488 ;
  assign y16842 = n41137 ;
  assign y16843 = ~n41138 ;
  assign y16844 = n41141 ;
  assign y16845 = n41144 ;
  assign y16846 = ~n41152 ;
  assign y16847 = n41153 ;
  assign y16848 = ~n41163 ;
  assign y16849 = n41165 ;
  assign y16850 = n41166 ;
  assign y16851 = ~1'b0 ;
  assign y16852 = ~1'b0 ;
  assign y16853 = ~n41167 ;
  assign y16854 = ~n41173 ;
  assign y16855 = n41174 ;
  assign y16856 = n41178 ;
  assign y16857 = n41179 ;
  assign y16858 = n41180 ;
  assign y16859 = 1'b0 ;
  assign y16860 = n41182 ;
  assign y16861 = ~1'b0 ;
  assign y16862 = ~n41184 ;
  assign y16863 = ~n41186 ;
  assign y16864 = n41188 ;
  assign y16865 = ~n41190 ;
  assign y16866 = n41191 ;
  assign y16867 = ~1'b0 ;
  assign y16868 = ~1'b0 ;
  assign y16869 = ~n41193 ;
  assign y16870 = ~n19821 ;
  assign y16871 = n41199 ;
  assign y16872 = n41202 ;
  assign y16873 = ~n41203 ;
  assign y16874 = n41205 ;
  assign y16875 = ~n41206 ;
  assign y16876 = ~n41214 ;
  assign y16877 = ~n41216 ;
  assign y16878 = ~n41223 ;
  assign y16879 = ~1'b0 ;
  assign y16880 = ~1'b0 ;
  assign y16881 = n41231 ;
  assign y16882 = n41233 ;
  assign y16883 = n41235 ;
  assign y16884 = ~n41237 ;
  assign y16885 = ~n41240 ;
  assign y16886 = ~n24098 ;
  assign y16887 = ~1'b0 ;
  assign y16888 = ~1'b0 ;
  assign y16889 = n41248 ;
  assign y16890 = n41250 ;
  assign y16891 = ~1'b0 ;
  assign y16892 = ~n6184 ;
  assign y16893 = n41252 ;
  assign y16894 = ~1'b0 ;
  assign y16895 = n41254 ;
  assign y16896 = ~1'b0 ;
  assign y16897 = ~n41259 ;
  assign y16898 = n41261 ;
  assign y16899 = ~n41264 ;
  assign y16900 = 1'b0 ;
  assign y16901 = n41267 ;
  assign y16902 = ~n41270 ;
  assign y16903 = ~1'b0 ;
  assign y16904 = n41271 ;
  assign y16905 = ~n41274 ;
  assign y16906 = ~n41275 ;
  assign y16907 = n41276 ;
  assign y16908 = n41277 ;
  assign y16909 = n41280 ;
  assign y16910 = ~n41281 ;
  assign y16911 = ~1'b0 ;
  assign y16912 = ~n41283 ;
  assign y16913 = ~n41289 ;
  assign y16914 = n35462 ;
  assign y16915 = n41293 ;
  assign y16916 = ~n41294 ;
  assign y16917 = ~1'b0 ;
  assign y16918 = ~1'b0 ;
  assign y16919 = n41295 ;
  assign y16920 = ~n41296 ;
  assign y16921 = ~n41297 ;
  assign y16922 = n41299 ;
  assign y16923 = n41301 ;
  assign y16924 = ~n41303 ;
  assign y16925 = n41307 ;
  assign y16926 = n41309 ;
  assign y16927 = 1'b0 ;
  assign y16928 = 1'b0 ;
  assign y16929 = ~1'b0 ;
  assign y16930 = n41310 ;
  assign y16931 = n7235 ;
  assign y16932 = ~n41311 ;
  assign y16933 = n41319 ;
  assign y16934 = ~1'b0 ;
  assign y16935 = ~n41323 ;
  assign y16936 = ~n41325 ;
  assign y16937 = ~1'b0 ;
  assign y16938 = ~1'b0 ;
  assign y16939 = n41326 ;
  assign y16940 = ~n41330 ;
  assign y16941 = ~n41331 ;
  assign y16942 = ~n41335 ;
  assign y16943 = ~1'b0 ;
  assign y16944 = ~1'b0 ;
  assign y16945 = ~1'b0 ;
  assign y16946 = ~n41342 ;
  assign y16947 = ~1'b0 ;
  assign y16948 = n41346 ;
  assign y16949 = n41347 ;
  assign y16950 = n41348 ;
  assign y16951 = n41351 ;
  assign y16952 = n41355 ;
  assign y16953 = ~1'b0 ;
  assign y16954 = ~n41358 ;
  assign y16955 = ~n41360 ;
  assign y16956 = ~n41362 ;
  assign y16957 = ~1'b0 ;
  assign y16958 = ~n41364 ;
  assign y16959 = n41365 ;
  assign y16960 = n41367 ;
  assign y16961 = n41373 ;
  assign y16962 = ~n41377 ;
  assign y16963 = n41378 ;
  assign y16964 = ~n41382 ;
  assign y16965 = ~n41383 ;
  assign y16966 = ~1'b0 ;
  assign y16967 = n41384 ;
  assign y16968 = n41387 ;
  assign y16969 = ~n41390 ;
  assign y16970 = ~n41393 ;
  assign y16971 = ~n41399 ;
  assign y16972 = ~n41410 ;
  assign y16973 = ~1'b0 ;
  assign y16974 = ~1'b0 ;
  assign y16975 = n41414 ;
  assign y16976 = ~n41416 ;
  assign y16977 = n41417 ;
  assign y16978 = ~1'b0 ;
  assign y16979 = ~n41419 ;
  assign y16980 = n41421 ;
  assign y16981 = n41429 ;
  assign y16982 = n41431 ;
  assign y16983 = ~n41432 ;
  assign y16984 = ~n41433 ;
  assign y16985 = ~n41435 ;
  assign y16986 = n37176 ;
  assign y16987 = ~1'b0 ;
  assign y16988 = ~n41438 ;
  assign y16989 = n41442 ;
  assign y16990 = ~n41443 ;
  assign y16991 = n41444 ;
  assign y16992 = n41446 ;
  assign y16993 = n41452 ;
  assign y16994 = ~n9644 ;
  assign y16995 = ~n41454 ;
  assign y16996 = n41456 ;
  assign y16997 = ~n41458 ;
  assign y16998 = ~n41459 ;
  assign y16999 = n41460 ;
  assign y17000 = ~n41461 ;
  assign y17001 = n41463 ;
  assign y17002 = n41468 ;
  assign y17003 = n41469 ;
  assign y17004 = n41472 ;
  assign y17005 = ~n41473 ;
  assign y17006 = n41474 ;
  assign y17007 = n41475 ;
  assign y17008 = ~n41476 ;
  assign y17009 = ~n41485 ;
  assign y17010 = ~n41486 ;
  assign y17011 = ~n41488 ;
  assign y17012 = ~1'b0 ;
  assign y17013 = ~n41490 ;
  assign y17014 = ~n41491 ;
  assign y17015 = ~n41493 ;
  assign y17016 = ~n41496 ;
  assign y17017 = n41501 ;
  assign y17018 = n41504 ;
  assign y17019 = ~1'b0 ;
  assign y17020 = n41506 ;
  assign y17021 = ~n41508 ;
  assign y17022 = ~1'b0 ;
  assign y17023 = ~1'b0 ;
  assign y17024 = ~n41512 ;
  assign y17025 = n41513 ;
  assign y17026 = ~n41516 ;
  assign y17027 = n41526 ;
  assign y17028 = ~n41529 ;
  assign y17029 = ~1'b0 ;
  assign y17030 = ~n16837 ;
  assign y17031 = ~n41531 ;
  assign y17032 = ~n41534 ;
  assign y17033 = ~1'b0 ;
  assign y17034 = n41535 ;
  assign y17035 = n41541 ;
  assign y17036 = ~n41545 ;
  assign y17037 = ~1'b0 ;
  assign y17038 = n41547 ;
  assign y17039 = n20450 ;
  assign y17040 = ~n41548 ;
  assign y17041 = n41549 ;
  assign y17042 = n10732 ;
  assign y17043 = ~n41553 ;
  assign y17044 = n41556 ;
  assign y17045 = n41561 ;
  assign y17046 = n41563 ;
  assign y17047 = ~n41565 ;
  assign y17048 = ~n41568 ;
  assign y17049 = n41569 ;
  assign y17050 = ~n41570 ;
  assign y17051 = ~n41576 ;
  assign y17052 = n41578 ;
  assign y17053 = n41582 ;
  assign y17054 = n41583 ;
  assign y17055 = ~n41590 ;
  assign y17056 = 1'b0 ;
  assign y17057 = ~n41591 ;
  assign y17058 = ~n41593 ;
  assign y17059 = n41595 ;
  assign y17060 = ~n41598 ;
  assign y17061 = n41599 ;
  assign y17062 = ~n41601 ;
  assign y17063 = ~n41603 ;
  assign y17064 = ~n41605 ;
  assign y17065 = ~n41607 ;
  assign y17066 = n41610 ;
  assign y17067 = n41612 ;
  assign y17068 = ~n41613 ;
  assign y17069 = ~1'b0 ;
  assign y17070 = ~n41617 ;
  assign y17071 = ~n41618 ;
  assign y17072 = ~n41622 ;
  assign y17073 = ~n41626 ;
  assign y17074 = ~n41629 ;
  assign y17075 = ~n41630 ;
  assign y17076 = ~n41631 ;
  assign y17077 = n41632 ;
  assign y17078 = n41634 ;
  assign y17079 = n41637 ;
  assign y17080 = n41638 ;
  assign y17081 = ~n41644 ;
  assign y17082 = ~n41647 ;
  assign y17083 = ~n41648 ;
  assign y17084 = ~n41649 ;
  assign y17085 = ~n41650 ;
  assign y17086 = n41654 ;
  assign y17087 = ~n41663 ;
  assign y17088 = ~1'b0 ;
  assign y17089 = n41664 ;
  assign y17090 = ~n41665 ;
  assign y17091 = n41669 ;
  assign y17092 = ~n41670 ;
  assign y17093 = ~n41678 ;
  assign y17094 = ~1'b0 ;
  assign y17095 = n41682 ;
  assign y17096 = ~n41684 ;
  assign y17097 = ~1'b0 ;
  assign y17098 = n41685 ;
  assign y17099 = ~n41687 ;
  assign y17100 = ~n41690 ;
  assign y17101 = ~n41693 ;
  assign y17102 = ~n41694 ;
  assign y17103 = n41701 ;
  assign y17104 = ~1'b0 ;
  assign y17105 = ~n41704 ;
  assign y17106 = n41707 ;
  assign y17107 = n41709 ;
  assign y17108 = n41716 ;
  assign y17109 = ~n41720 ;
  assign y17110 = ~1'b0 ;
  assign y17111 = ~1'b0 ;
  assign y17112 = n41722 ;
  assign y17113 = n14262 ;
  assign y17114 = ~1'b0 ;
  assign y17115 = ~n41725 ;
  assign y17116 = ~n41726 ;
  assign y17117 = ~n41727 ;
  assign y17118 = ~n41729 ;
  assign y17119 = ~1'b0 ;
  assign y17120 = ~n41730 ;
  assign y17121 = n41733 ;
  assign y17122 = n41735 ;
  assign y17123 = ~n41736 ;
  assign y17124 = ~n41739 ;
  assign y17125 = n41743 ;
  assign y17126 = n41747 ;
  assign y17127 = n41748 ;
  assign y17128 = n41753 ;
  assign y17129 = ~n41755 ;
  assign y17130 = ~n41760 ;
  assign y17131 = n41762 ;
  assign y17132 = ~1'b0 ;
  assign y17133 = ~n41765 ;
  assign y17134 = n41766 ;
  assign y17135 = n41768 ;
  assign y17136 = ~n41772 ;
  assign y17137 = ~n34796 ;
  assign y17138 = n41776 ;
  assign y17139 = ~1'b0 ;
  assign y17140 = ~n41781 ;
  assign y17141 = n41782 ;
  assign y17142 = ~n27190 ;
  assign y17143 = n41788 ;
  assign y17144 = ~n41790 ;
  assign y17145 = n41791 ;
  assign y17146 = ~n41792 ;
  assign y17147 = ~n41794 ;
  assign y17148 = n41798 ;
  assign y17149 = ~n41799 ;
  assign y17150 = ~1'b0 ;
  assign y17151 = ~n41800 ;
  assign y17152 = n41806 ;
  assign y17153 = ~n41807 ;
  assign y17154 = ~1'b0 ;
  assign y17155 = ~n41810 ;
  assign y17156 = ~1'b0 ;
  assign y17157 = n41812 ;
  assign y17158 = ~n41814 ;
  assign y17159 = ~n41816 ;
  assign y17160 = ~n9863 ;
  assign y17161 = ~n41818 ;
  assign y17162 = n41822 ;
  assign y17163 = ~n41823 ;
  assign y17164 = ~n41825 ;
  assign y17165 = ~n41827 ;
  assign y17166 = n41828 ;
  assign y17167 = n41831 ;
  assign y17168 = ~n41834 ;
  assign y17169 = ~n41838 ;
  assign y17170 = 1'b0 ;
  assign y17171 = n41839 ;
  assign y17172 = ~n41842 ;
  assign y17173 = n41848 ;
  assign y17174 = ~n41849 ;
  assign y17175 = n41850 ;
  assign y17176 = ~n41854 ;
  assign y17177 = ~1'b0 ;
  assign y17178 = n41856 ;
  assign y17179 = ~n41858 ;
  assign y17180 = ~n41864 ;
  assign y17181 = n41867 ;
  assign y17182 = n41868 ;
  assign y17183 = n41869 ;
  assign y17184 = ~n41874 ;
  assign y17185 = n41881 ;
  assign y17186 = ~n41882 ;
  assign y17187 = ~n41884 ;
  assign y17188 = ~1'b0 ;
  assign y17189 = ~n41886 ;
  assign y17190 = ~n41888 ;
  assign y17191 = n41889 ;
  assign y17192 = n41891 ;
  assign y17193 = ~n41899 ;
  assign y17194 = n9566 ;
  assign y17195 = ~1'b0 ;
  assign y17196 = ~n3644 ;
  assign y17197 = n41900 ;
  assign y17198 = ~n41902 ;
  assign y17199 = ~n41903 ;
  assign y17200 = n41909 ;
  assign y17201 = n41914 ;
  assign y17202 = ~n41917 ;
  assign y17203 = ~n41921 ;
  assign y17204 = n41922 ;
  assign y17205 = n41925 ;
  assign y17206 = ~n41930 ;
  assign y17207 = n41932 ;
  assign y17208 = ~1'b0 ;
  assign y17209 = n41933 ;
  assign y17210 = n41936 ;
  assign y17211 = ~n41937 ;
  assign y17212 = ~n41943 ;
  assign y17213 = ~n41944 ;
  assign y17214 = ~n41949 ;
  assign y17215 = n41951 ;
  assign y17216 = ~n41953 ;
  assign y17217 = n41961 ;
  assign y17218 = ~n41964 ;
  assign y17219 = n41966 ;
  assign y17220 = ~n41968 ;
  assign y17221 = ~1'b0 ;
  assign y17222 = ~n665 ;
  assign y17223 = ~1'b0 ;
  assign y17224 = ~n41969 ;
  assign y17225 = ~n41973 ;
  assign y17226 = ~n41974 ;
  assign y17227 = n41977 ;
  assign y17228 = ~1'b0 ;
  assign y17229 = ~1'b0 ;
  assign y17230 = ~n41982 ;
  assign y17231 = ~1'b0 ;
  assign y17232 = n41984 ;
  assign y17233 = ~1'b0 ;
  assign y17234 = n41985 ;
  assign y17235 = ~n41986 ;
  assign y17236 = ~n41987 ;
  assign y17237 = ~1'b0 ;
  assign y17238 = ~n41989 ;
  assign y17239 = n41994 ;
  assign y17240 = n41996 ;
  assign y17241 = ~n41997 ;
  assign y17242 = ~n42003 ;
  assign y17243 = ~n42005 ;
  assign y17244 = n42006 ;
  assign y17245 = ~n42008 ;
  assign y17246 = ~n42012 ;
  assign y17247 = ~n42013 ;
  assign y17248 = n42015 ;
  assign y17249 = n42016 ;
  assign y17250 = ~n42019 ;
  assign y17251 = ~n6045 ;
  assign y17252 = n42021 ;
  assign y17253 = n42023 ;
  assign y17254 = ~n42031 ;
  assign y17255 = n19113 ;
  assign y17256 = ~n42032 ;
  assign y17257 = ~1'b0 ;
  assign y17258 = n42037 ;
  assign y17259 = ~n42038 ;
  assign y17260 = ~n42040 ;
  assign y17261 = n42046 ;
  assign y17262 = n15366 ;
  assign y17263 = n42047 ;
  assign y17264 = n42048 ;
  assign y17265 = ~n42051 ;
  assign y17266 = ~1'b0 ;
  assign y17267 = ~1'b0 ;
  assign y17268 = ~1'b0 ;
  assign y17269 = n42053 ;
  assign y17270 = ~1'b0 ;
  assign y17271 = n42058 ;
  assign y17272 = n42061 ;
  assign y17273 = n42065 ;
  assign y17274 = ~n42067 ;
  assign y17275 = ~n42068 ;
  assign y17276 = n42069 ;
  assign y17277 = ~1'b0 ;
  assign y17278 = ~n42073 ;
  assign y17279 = ~n42077 ;
  assign y17280 = n42079 ;
  assign y17281 = n42083 ;
  assign y17282 = ~n42085 ;
  assign y17283 = ~1'b0 ;
  assign y17284 = ~n42089 ;
  assign y17285 = ~1'b0 ;
  assign y17286 = ~1'b0 ;
  assign y17287 = n42092 ;
  assign y17288 = ~n42093 ;
  assign y17289 = n42101 ;
  assign y17290 = ~n42102 ;
  assign y17291 = ~n42107 ;
  assign y17292 = n42110 ;
  assign y17293 = ~1'b0 ;
  assign y17294 = n42111 ;
  assign y17295 = ~1'b0 ;
  assign y17296 = ~1'b0 ;
  assign y17297 = n42114 ;
  assign y17298 = ~n42117 ;
  assign y17299 = ~1'b0 ;
  assign y17300 = n42119 ;
  assign y17301 = ~n42123 ;
  assign y17302 = ~1'b0 ;
  assign y17303 = ~1'b0 ;
  assign y17304 = n42125 ;
  assign y17305 = n42135 ;
  assign y17306 = n42139 ;
  assign y17307 = n42141 ;
  assign y17308 = ~n42142 ;
  assign y17309 = ~n42146 ;
  assign y17310 = ~n42147 ;
  assign y17311 = n42151 ;
  assign y17312 = ~1'b0 ;
  assign y17313 = ~n42155 ;
  assign y17314 = ~n42156 ;
  assign y17315 = n42157 ;
  assign y17316 = ~n42162 ;
  assign y17317 = ~n42169 ;
  assign y17318 = ~1'b0 ;
  assign y17319 = ~n42171 ;
  assign y17320 = ~1'b0 ;
  assign y17321 = ~n42173 ;
  assign y17322 = ~n42174 ;
  assign y17323 = n42175 ;
  assign y17324 = n42179 ;
  assign y17325 = n42183 ;
  assign y17326 = x253 ;
  assign y17327 = ~n42184 ;
  assign y17328 = ~n42187 ;
  assign y17329 = ~n36689 ;
  assign y17330 = n42188 ;
  assign y17331 = ~n42193 ;
  assign y17332 = ~n42198 ;
  assign y17333 = n42201 ;
  assign y17334 = n42202 ;
  assign y17335 = ~n42203 ;
  assign y17336 = ~1'b0 ;
  assign y17337 = n42205 ;
  assign y17338 = n42206 ;
  assign y17339 = n12167 ;
  assign y17340 = ~n42212 ;
  assign y17341 = n42213 ;
  assign y17342 = ~n42217 ;
  assign y17343 = n42218 ;
  assign y17344 = ~n42221 ;
  assign y17345 = ~1'b0 ;
  assign y17346 = ~1'b0 ;
  assign y17347 = ~n42223 ;
  assign y17348 = n42227 ;
  assign y17349 = ~n42231 ;
  assign y17350 = ~1'b0 ;
  assign y17351 = n42234 ;
  assign y17352 = ~n42235 ;
  assign y17353 = ~1'b0 ;
  assign y17354 = ~1'b0 ;
  assign y17355 = n42237 ;
  assign y17356 = n30201 ;
  assign y17357 = ~n42240 ;
  assign y17358 = ~n42241 ;
  assign y17359 = ~n42243 ;
  assign y17360 = n42244 ;
  assign y17361 = ~1'b0 ;
  assign y17362 = ~n42245 ;
  assign y17363 = ~1'b0 ;
  assign y17364 = ~1'b0 ;
  assign y17365 = n42248 ;
  assign y17366 = n42252 ;
  assign y17367 = n42254 ;
  assign y17368 = n42255 ;
  assign y17369 = n42256 ;
  assign y17370 = ~1'b0 ;
  assign y17371 = ~n12679 ;
  assign y17372 = n42263 ;
  assign y17373 = ~n42265 ;
  assign y17374 = n42268 ;
  assign y17375 = ~n42271 ;
  assign y17376 = ~n42272 ;
  assign y17377 = ~n42278 ;
  assign y17378 = ~n42290 ;
  assign y17379 = ~n42291 ;
  assign y17380 = ~1'b0 ;
  assign y17381 = ~1'b0 ;
  assign y17382 = ~1'b0 ;
  assign y17383 = ~1'b0 ;
  assign y17384 = ~n42294 ;
  assign y17385 = n42295 ;
  assign y17386 = n42301 ;
  assign y17387 = n42302 ;
  assign y17388 = ~1'b0 ;
  assign y17389 = ~n42303 ;
  assign y17390 = n42304 ;
  assign y17391 = n42308 ;
  assign y17392 = ~n42311 ;
  assign y17393 = n42313 ;
  assign y17394 = n42315 ;
  assign y17395 = ~1'b0 ;
  assign y17396 = ~n42319 ;
  assign y17397 = n42320 ;
  assign y17398 = ~1'b0 ;
  assign y17399 = ~1'b0 ;
  assign y17400 = ~n42325 ;
  assign y17401 = ~n42326 ;
  assign y17402 = n42327 ;
  assign y17403 = ~n42328 ;
  assign y17404 = n42329 ;
  assign y17405 = ~1'b0 ;
  assign y17406 = ~n42331 ;
  assign y17407 = ~1'b0 ;
  assign y17408 = ~1'b0 ;
  assign y17409 = n42334 ;
  assign y17410 = n42336 ;
  assign y17411 = ~n9847 ;
  assign y17412 = ~1'b0 ;
  assign y17413 = n42340 ;
  assign y17414 = ~1'b0 ;
  assign y17415 = ~n42341 ;
  assign y17416 = ~1'b0 ;
  assign y17417 = ~n42343 ;
  assign y17418 = n42346 ;
  assign y17419 = ~n42351 ;
  assign y17420 = n42355 ;
  assign y17421 = n42359 ;
  assign y17422 = n42360 ;
  assign y17423 = n42362 ;
  assign y17424 = ~1'b0 ;
  assign y17425 = n42364 ;
  assign y17426 = ~n42371 ;
  assign y17427 = ~n31965 ;
  assign y17428 = n42372 ;
  assign y17429 = ~n42373 ;
  assign y17430 = n42374 ;
  assign y17431 = n42377 ;
  assign y17432 = n42381 ;
  assign y17433 = ~1'b0 ;
  assign y17434 = n42382 ;
  assign y17435 = ~1'b0 ;
  assign y17436 = ~n42386 ;
  assign y17437 = n42387 ;
  assign y17438 = ~n42390 ;
  assign y17439 = n42391 ;
  assign y17440 = ~1'b0 ;
  assign y17441 = n42393 ;
  assign y17442 = ~n42401 ;
  assign y17443 = ~1'b0 ;
  assign y17444 = ~n42403 ;
  assign y17445 = ~n42404 ;
  assign y17446 = ~n42405 ;
  assign y17447 = ~n42407 ;
  assign y17448 = n42408 ;
  assign y17449 = ~1'b0 ;
  assign y17450 = ~n42414 ;
  assign y17451 = n42416 ;
  assign y17452 = n42418 ;
  assign y17453 = ~n42422 ;
  assign y17454 = n42426 ;
  assign y17455 = n42429 ;
  assign y17456 = ~n42432 ;
  assign y17457 = ~1'b0 ;
  assign y17458 = ~1'b0 ;
  assign y17459 = n42436 ;
  assign y17460 = n42438 ;
  assign y17461 = ~1'b0 ;
  assign y17462 = n42439 ;
  assign y17463 = n42440 ;
  assign y17464 = ~n42442 ;
  assign y17465 = n9564 ;
  assign y17466 = ~n42444 ;
  assign y17467 = n42446 ;
  assign y17468 = n42447 ;
  assign y17469 = ~n42448 ;
  assign y17470 = n11334 ;
  assign y17471 = n42449 ;
  assign y17472 = ~n42451 ;
  assign y17473 = ~n42455 ;
  assign y17474 = ~n42459 ;
  assign y17475 = ~n42462 ;
  assign y17476 = n42463 ;
  assign y17477 = ~1'b0 ;
  assign y17478 = ~n42464 ;
  assign y17479 = ~1'b0 ;
  assign y17480 = n42466 ;
  assign y17481 = ~n42468 ;
  assign y17482 = n42476 ;
  assign y17483 = n42478 ;
  assign y17484 = n42481 ;
  assign y17485 = n42485 ;
  assign y17486 = ~n42491 ;
  assign y17487 = n42492 ;
  assign y17488 = n42494 ;
  assign y17489 = ~n42495 ;
  assign y17490 = ~n42496 ;
  assign y17491 = ~n42498 ;
  assign y17492 = n42499 ;
  assign y17493 = n42501 ;
  assign y17494 = n42505 ;
  assign y17495 = ~1'b0 ;
  assign y17496 = ~n42509 ;
  assign y17497 = ~1'b0 ;
  assign y17498 = ~n42510 ;
  assign y17499 = ~n42511 ;
  assign y17500 = n42518 ;
  assign y17501 = ~n42519 ;
  assign y17502 = n42521 ;
  assign y17503 = n42522 ;
  assign y17504 = ~n42528 ;
  assign y17505 = ~n42529 ;
  assign y17506 = ~n42533 ;
  assign y17507 = ~n42537 ;
  assign y17508 = n42538 ;
  assign y17509 = n42539 ;
  assign y17510 = ~1'b0 ;
  assign y17511 = ~n42546 ;
  assign y17512 = n42550 ;
  assign y17513 = ~n42552 ;
  assign y17514 = ~n42554 ;
  assign y17515 = ~1'b0 ;
  assign y17516 = ~n2296 ;
  assign y17517 = n14789 ;
  assign y17518 = ~n42555 ;
  assign y17519 = n42558 ;
  assign y17520 = ~1'b0 ;
  assign y17521 = n42561 ;
  assign y17522 = n42565 ;
  assign y17523 = ~n42570 ;
  assign y17524 = ~1'b0 ;
  assign y17525 = n42571 ;
  assign y17526 = ~n42572 ;
  assign y17527 = n42573 ;
  assign y17528 = n42574 ;
  assign y17529 = n42576 ;
  assign y17530 = n42579 ;
  assign y17531 = ~1'b0 ;
  assign y17532 = ~n42582 ;
  assign y17533 = ~n42585 ;
  assign y17534 = ~n42591 ;
  assign y17535 = n42592 ;
  assign y17536 = ~1'b0 ;
  assign y17537 = ~1'b0 ;
  assign y17538 = ~n42593 ;
  assign y17539 = ~n42595 ;
  assign y17540 = n42597 ;
  assign y17541 = ~1'b0 ;
  assign y17542 = n42598 ;
  assign y17543 = n42600 ;
  assign y17544 = ~1'b0 ;
  assign y17545 = n42602 ;
  assign y17546 = n42603 ;
  assign y17547 = ~1'b0 ;
  assign y17548 = ~n42605 ;
  assign y17549 = ~1'b0 ;
  assign y17550 = ~n42606 ;
  assign y17551 = n42607 ;
  assign y17552 = n42610 ;
  assign y17553 = n42615 ;
  assign y17554 = n42617 ;
  assign y17555 = n42620 ;
  assign y17556 = ~1'b0 ;
  assign y17557 = 1'b0 ;
  assign y17558 = ~1'b0 ;
  assign y17559 = n42622 ;
  assign y17560 = n42625 ;
  assign y17561 = ~1'b0 ;
  assign y17562 = ~n42627 ;
  assign y17563 = ~n42630 ;
  assign y17564 = n42632 ;
  assign y17565 = ~n42635 ;
  assign y17566 = ~1'b0 ;
  assign y17567 = n2444 ;
  assign y17568 = ~n42637 ;
  assign y17569 = n42638 ;
  assign y17570 = n42639 ;
  assign y17571 = n42640 ;
  assign y17572 = ~n42641 ;
  assign y17573 = ~n42642 ;
  assign y17574 = ~n42645 ;
  assign y17575 = ~n42646 ;
  assign y17576 = ~1'b0 ;
  assign y17577 = n42653 ;
  assign y17578 = ~n42656 ;
  assign y17579 = ~n42658 ;
  assign y17580 = n42661 ;
  assign y17581 = n42663 ;
  assign y17582 = ~n42664 ;
  assign y17583 = ~n42671 ;
  assign y17584 = n42674 ;
  assign y17585 = ~1'b0 ;
  assign y17586 = ~n42678 ;
  assign y17587 = ~1'b0 ;
  assign y17588 = ~n42683 ;
  assign y17589 = n42684 ;
  assign y17590 = n42688 ;
  assign y17591 = n42692 ;
  assign y17592 = n42699 ;
  assign y17593 = n42700 ;
  assign y17594 = ~1'b0 ;
  assign y17595 = ~1'b0 ;
  assign y17596 = ~n42706 ;
  assign y17597 = n42708 ;
  assign y17598 = n42711 ;
  assign y17599 = ~n42712 ;
  assign y17600 = ~1'b0 ;
  assign y17601 = n42714 ;
  assign y17602 = ~1'b0 ;
  assign y17603 = ~1'b0 ;
  assign y17604 = ~n42715 ;
  assign y17605 = ~1'b0 ;
  assign y17606 = n42717 ;
  assign y17607 = n42719 ;
  assign y17608 = n3596 ;
  assign y17609 = ~n42721 ;
  assign y17610 = n42723 ;
  assign y17611 = ~1'b0 ;
  assign y17612 = ~n42725 ;
  assign y17613 = n4868 ;
  assign y17614 = ~1'b0 ;
  assign y17615 = ~n42726 ;
  assign y17616 = ~n42728 ;
  assign y17617 = ~n14929 ;
  assign y17618 = n42730 ;
  assign y17619 = ~1'b0 ;
  assign y17620 = n42732 ;
  assign y17621 = ~n42735 ;
  assign y17622 = ~n42738 ;
  assign y17623 = n42740 ;
  assign y17624 = n42745 ;
  assign y17625 = n42746 ;
  assign y17626 = n42747 ;
  assign y17627 = ~n42750 ;
  assign y17628 = n42751 ;
  assign y17629 = ~n42752 ;
  assign y17630 = ~n42754 ;
  assign y17631 = ~n42755 ;
  assign y17632 = n42761 ;
  assign y17633 = ~n42765 ;
  assign y17634 = ~n16358 ;
  assign y17635 = ~n42766 ;
  assign y17636 = n42767 ;
  assign y17637 = ~n42770 ;
  assign y17638 = n42772 ;
  assign y17639 = ~n42773 ;
  assign y17640 = n42774 ;
  assign y17641 = ~1'b0 ;
  assign y17642 = n42777 ;
  assign y17643 = ~n42778 ;
  assign y17644 = n13710 ;
  assign y17645 = n42780 ;
  assign y17646 = n1629 ;
  assign y17647 = n42782 ;
  assign y17648 = ~n42786 ;
  assign y17649 = ~1'b0 ;
  assign y17650 = ~n42787 ;
  assign y17651 = n42791 ;
  assign y17652 = ~n42793 ;
  assign y17653 = n42794 ;
  assign y17654 = ~n42796 ;
  assign y17655 = ~1'b0 ;
  assign y17656 = ~1'b0 ;
  assign y17657 = ~n42799 ;
  assign y17658 = ~1'b0 ;
  assign y17659 = n42807 ;
  assign y17660 = n42808 ;
  assign y17661 = n42809 ;
  assign y17662 = ~n42811 ;
  assign y17663 = ~n42813 ;
  assign y17664 = 1'b0 ;
  assign y17665 = ~n9109 ;
  assign y17666 = 1'b0 ;
  assign y17667 = n42815 ;
  assign y17668 = ~n42817 ;
  assign y17669 = 1'b0 ;
  assign y17670 = n424 ;
  assign y17671 = n42822 ;
  assign y17672 = ~1'b0 ;
  assign y17673 = n42823 ;
  assign y17674 = ~1'b0 ;
  assign y17675 = n42827 ;
  assign y17676 = ~1'b0 ;
  assign y17677 = ~1'b0 ;
  assign y17678 = ~n42829 ;
  assign y17679 = ~1'b0 ;
  assign y17680 = n42830 ;
  assign y17681 = n1711 ;
  assign y17682 = n42832 ;
  assign y17683 = ~n42834 ;
  assign y17684 = ~1'b0 ;
  assign y17685 = ~1'b0 ;
  assign y17686 = ~1'b0 ;
  assign y17687 = n42838 ;
  assign y17688 = ~1'b0 ;
  assign y17689 = ~1'b0 ;
  assign y17690 = ~n42839 ;
  assign y17691 = ~n42840 ;
  assign y17692 = ~n42845 ;
  assign y17693 = ~n42849 ;
  assign y17694 = ~n42853 ;
  assign y17695 = ~1'b0 ;
  assign y17696 = n42854 ;
  assign y17697 = ~1'b0 ;
  assign y17698 = ~n42855 ;
  assign y17699 = n42856 ;
  assign y17700 = ~n42857 ;
  assign y17701 = n42860 ;
  assign y17702 = ~n42862 ;
  assign y17703 = ~n42865 ;
  assign y17704 = ~1'b0 ;
  assign y17705 = n42871 ;
  assign y17706 = n42872 ;
  assign y17707 = ~1'b0 ;
  assign y17708 = n42873 ;
  assign y17709 = n42876 ;
  assign y17710 = n42878 ;
  assign y17711 = ~n4827 ;
  assign y17712 = n1197 ;
  assign y17713 = n42879 ;
  assign y17714 = n21192 ;
  assign y17715 = ~n42883 ;
  assign y17716 = ~1'b0 ;
  assign y17717 = n35596 ;
  assign y17718 = ~n42888 ;
  assign y17719 = ~n42892 ;
  assign y17720 = ~n42894 ;
  assign y17721 = n42895 ;
  assign y17722 = ~1'b0 ;
  assign y17723 = n42897 ;
  assign y17724 = ~1'b0 ;
  assign y17725 = n42901 ;
  assign y17726 = n42902 ;
  assign y17727 = n31152 ;
  assign y17728 = n42907 ;
  assign y17729 = ~n42912 ;
  assign y17730 = ~n42913 ;
  assign y17731 = ~n42917 ;
  assign y17732 = n42922 ;
  assign y17733 = ~1'b0 ;
  assign y17734 = ~1'b0 ;
  assign y17735 = n42923 ;
  assign y17736 = n42925 ;
  assign y17737 = ~n42928 ;
  assign y17738 = ~n42929 ;
  assign y17739 = ~n42931 ;
  assign y17740 = ~n42932 ;
  assign y17741 = n42940 ;
  assign y17742 = n12269 ;
  assign y17743 = ~n42941 ;
  assign y17744 = ~1'b0 ;
  assign y17745 = n42942 ;
  assign y17746 = ~1'b0 ;
  assign y17747 = ~1'b0 ;
  assign y17748 = n42945 ;
  assign y17749 = ~n42947 ;
  assign y17750 = n42948 ;
  assign y17751 = ~1'b0 ;
  assign y17752 = n42950 ;
  assign y17753 = n42952 ;
  assign y17754 = ~n42954 ;
  assign y17755 = ~n42958 ;
  assign y17756 = ~n42966 ;
  assign y17757 = n42970 ;
  assign y17758 = ~n42975 ;
  assign y17759 = n7638 ;
  assign y17760 = n42976 ;
  assign y17761 = n42978 ;
  assign y17762 = ~1'b0 ;
  assign y17763 = ~n42980 ;
  assign y17764 = ~1'b0 ;
  assign y17765 = ~1'b0 ;
  assign y17766 = 1'b0 ;
  assign y17767 = ~n42982 ;
  assign y17768 = ~1'b0 ;
  assign y17769 = ~n42987 ;
  assign y17770 = n42988 ;
  assign y17771 = ~n42989 ;
  assign y17772 = ~1'b0 ;
  assign y17773 = ~n42990 ;
  assign y17774 = n42994 ;
  assign y17775 = ~1'b0 ;
  assign y17776 = ~n42995 ;
  assign y17777 = ~1'b0 ;
  assign y17778 = n42996 ;
  assign y17779 = n42999 ;
  assign y17780 = n43002 ;
  assign y17781 = n43004 ;
  assign y17782 = n43007 ;
  assign y17783 = ~n43009 ;
  assign y17784 = ~1'b0 ;
  assign y17785 = ~1'b0 ;
  assign y17786 = ~1'b0 ;
  assign y17787 = ~n43013 ;
  assign y17788 = ~1'b0 ;
  assign y17789 = ~n21084 ;
  assign y17790 = ~n43016 ;
  assign y17791 = ~n43023 ;
  assign y17792 = ~n43026 ;
  assign y17793 = n43029 ;
  assign y17794 = n43030 ;
  assign y17795 = ~n43034 ;
  assign y17796 = n43037 ;
  assign y17797 = n43039 ;
  assign y17798 = ~n43042 ;
  assign y17799 = n4619 ;
  assign y17800 = n43044 ;
  assign y17801 = n43046 ;
  assign y17802 = ~1'b0 ;
  assign y17803 = n43047 ;
  assign y17804 = ~n43049 ;
  assign y17805 = n43053 ;
  assign y17806 = ~n43054 ;
  assign y17807 = ~n43056 ;
  assign y17808 = ~n43059 ;
  assign y17809 = ~n43061 ;
  assign y17810 = n22088 ;
  assign y17811 = ~1'b0 ;
  assign y17812 = ~n43063 ;
  assign y17813 = ~n43064 ;
  assign y17814 = ~1'b0 ;
  assign y17815 = ~n14274 ;
  assign y17816 = n43068 ;
  assign y17817 = ~n43070 ;
  assign y17818 = ~n43072 ;
  assign y17819 = n43073 ;
  assign y17820 = ~n43074 ;
  assign y17821 = ~n43076 ;
  assign y17822 = n43078 ;
  assign y17823 = n43081 ;
  assign y17824 = ~1'b0 ;
  assign y17825 = n43089 ;
  assign y17826 = n43091 ;
  assign y17827 = ~n43092 ;
  assign y17828 = ~n43093 ;
  assign y17829 = n43097 ;
  assign y17830 = n40879 ;
  assign y17831 = ~1'b0 ;
  assign y17832 = n43101 ;
  assign y17833 = n43104 ;
  assign y17834 = n43111 ;
  assign y17835 = n43112 ;
  assign y17836 = n43114 ;
  assign y17837 = n43119 ;
  assign y17838 = n43120 ;
  assign y17839 = ~1'b0 ;
  assign y17840 = n43122 ;
  assign y17841 = ~1'b0 ;
  assign y17842 = n43125 ;
  assign y17843 = ~n43129 ;
  assign y17844 = 1'b0 ;
  assign y17845 = ~n43132 ;
  assign y17846 = ~1'b0 ;
  assign y17847 = ~n43135 ;
  assign y17848 = ~n43138 ;
  assign y17849 = n43140 ;
  assign y17850 = ~n43141 ;
  assign y17851 = n43144 ;
  assign y17852 = ~n43145 ;
  assign y17853 = n18289 ;
  assign y17854 = ~n43147 ;
  assign y17855 = ~n43148 ;
  assign y17856 = ~n43149 ;
  assign y17857 = n43150 ;
  assign y17858 = ~n43152 ;
  assign y17859 = n43154 ;
  assign y17860 = n43155 ;
  assign y17861 = n28283 ;
  assign y17862 = n43157 ;
  assign y17863 = n43159 ;
  assign y17864 = ~1'b0 ;
  assign y17865 = n43161 ;
  assign y17866 = n43164 ;
  assign y17867 = ~n43166 ;
  assign y17868 = ~n43169 ;
  assign y17869 = n43171 ;
  assign y17870 = n43172 ;
  assign y17871 = n43175 ;
  assign y17872 = n43176 ;
  assign y17873 = ~n43180 ;
  assign y17874 = n43181 ;
  assign y17875 = n43182 ;
  assign y17876 = ~1'b0 ;
  assign y17877 = ~1'b0 ;
  assign y17878 = ~1'b0 ;
  assign y17879 = ~n43183 ;
  assign y17880 = n43186 ;
  assign y17881 = n26618 ;
  assign y17882 = n43187 ;
  assign y17883 = ~n43190 ;
  assign y17884 = ~n43195 ;
  assign y17885 = n43198 ;
  assign y17886 = ~n43206 ;
  assign y17887 = n43211 ;
  assign y17888 = ~n43214 ;
  assign y17889 = n43217 ;
  assign y17890 = ~n43221 ;
  assign y17891 = n43224 ;
  assign y17892 = n43227 ;
  assign y17893 = n43230 ;
  assign y17894 = ~1'b0 ;
  assign y17895 = ~n43237 ;
  assign y17896 = ~1'b0 ;
  assign y17897 = ~1'b0 ;
  assign y17898 = ~n43239 ;
  assign y17899 = n43240 ;
  assign y17900 = ~n43246 ;
  assign y17901 = ~n43250 ;
  assign y17902 = n43251 ;
  assign y17903 = n43255 ;
  assign y17904 = ~n43257 ;
  assign y17905 = n43258 ;
  assign y17906 = ~1'b0 ;
  assign y17907 = ~1'b0 ;
  assign y17908 = ~n43259 ;
  assign y17909 = n43260 ;
  assign y17910 = n43263 ;
  assign y17911 = ~n43265 ;
  assign y17912 = ~n43269 ;
  assign y17913 = ~n43274 ;
  assign y17914 = ~n43275 ;
  assign y17915 = ~1'b0 ;
  assign y17916 = n43280 ;
  assign y17917 = ~n43282 ;
  assign y17918 = n43284 ;
  assign y17919 = n43285 ;
  assign y17920 = n43290 ;
  assign y17921 = n43291 ;
  assign y17922 = n43292 ;
  assign y17923 = n43298 ;
  assign y17924 = ~n43300 ;
  assign y17925 = n43306 ;
  assign y17926 = ~n26429 ;
  assign y17927 = n43307 ;
  assign y17928 = ~1'b0 ;
  assign y17929 = ~1'b0 ;
  assign y17930 = ~n43311 ;
  assign y17931 = ~n20925 ;
  assign y17932 = ~n43313 ;
  assign y17933 = n43315 ;
  assign y17934 = n43316 ;
  assign y17935 = ~n31751 ;
  assign y17936 = ~n43319 ;
  assign y17937 = ~n43322 ;
  assign y17938 = ~1'b0 ;
  assign y17939 = n43323 ;
  assign y17940 = ~n43325 ;
  assign y17941 = ~n43326 ;
  assign y17942 = ~n43328 ;
  assign y17943 = n43330 ;
  assign y17944 = ~n43333 ;
  assign y17945 = n43335 ;
  assign y17946 = n43337 ;
  assign y17947 = ~1'b0 ;
  assign y17948 = ~n43342 ;
  assign y17949 = n43345 ;
  assign y17950 = n43347 ;
  assign y17951 = n43349 ;
  assign y17952 = ~n43350 ;
  assign y17953 = ~n43353 ;
  assign y17954 = ~n43357 ;
  assign y17955 = n43360 ;
  assign y17956 = ~n9071 ;
  assign y17957 = ~1'b0 ;
  assign y17958 = n43361 ;
  assign y17959 = ~n43364 ;
  assign y17960 = ~1'b0 ;
  assign y17961 = n43366 ;
  assign y17962 = n43375 ;
  assign y17963 = ~n21466 ;
  assign y17964 = ~n43378 ;
  assign y17965 = n43381 ;
  assign y17966 = ~n43383 ;
  assign y17967 = ~1'b0 ;
  assign y17968 = n43388 ;
  assign y17969 = ~n43391 ;
  assign y17970 = ~n40634 ;
  assign y17971 = ~n43392 ;
  assign y17972 = ~n43393 ;
  assign y17973 = n6435 ;
  assign y17974 = ~n43399 ;
  assign y17975 = ~1'b0 ;
  assign y17976 = ~n43400 ;
  assign y17977 = n43401 ;
  assign y17978 = n43402 ;
  assign y17979 = ~n43403 ;
  assign y17980 = ~n43404 ;
  assign y17981 = ~1'b0 ;
  assign y17982 = ~n43411 ;
  assign y17983 = ~n43415 ;
  assign y17984 = ~1'b0 ;
  assign y17985 = ~1'b0 ;
  assign y17986 = n43416 ;
  assign y17987 = ~n43417 ;
  assign y17988 = ~n43418 ;
  assign y17989 = ~1'b0 ;
  assign y17990 = ~1'b0 ;
  assign y17991 = ~1'b0 ;
  assign y17992 = ~n20319 ;
  assign y17993 = n43419 ;
  assign y17994 = ~1'b0 ;
  assign y17995 = ~n43423 ;
  assign y17996 = ~n43424 ;
  assign y17997 = ~n43425 ;
  assign y17998 = n40845 ;
  assign y17999 = ~n43428 ;
  assign y18000 = n43432 ;
  assign y18001 = ~1'b0 ;
  assign y18002 = n43433 ;
  assign y18003 = n14262 ;
  assign y18004 = ~1'b0 ;
  assign y18005 = ~1'b0 ;
  assign y18006 = ~n43434 ;
  assign y18007 = ~n43436 ;
  assign y18008 = ~n43439 ;
  assign y18009 = ~1'b0 ;
  assign y18010 = ~1'b0 ;
  assign y18011 = ~n43445 ;
  assign y18012 = n43449 ;
  assign y18013 = ~n43452 ;
  assign y18014 = ~n43457 ;
  assign y18015 = n43458 ;
  assign y18016 = n43459 ;
  assign y18017 = n43464 ;
  assign y18018 = ~n43468 ;
  assign y18019 = ~n43470 ;
  assign y18020 = ~1'b0 ;
  assign y18021 = ~n43471 ;
  assign y18022 = ~1'b0 ;
  assign y18023 = n43476 ;
  assign y18024 = ~n43478 ;
  assign y18025 = ~n43481 ;
  assign y18026 = n43485 ;
  assign y18027 = n43487 ;
  assign y18028 = n43496 ;
  assign y18029 = ~1'b0 ;
  assign y18030 = ~1'b0 ;
  assign y18031 = n43498 ;
  assign y18032 = ~n43500 ;
  assign y18033 = n4558 ;
  assign y18034 = n43502 ;
  assign y18035 = ~n43505 ;
  assign y18036 = ~n43507 ;
  assign y18037 = n43510 ;
  assign y18038 = ~1'b0 ;
  assign y18039 = ~1'b0 ;
  assign y18040 = n43513 ;
  assign y18041 = ~1'b0 ;
  assign y18042 = ~n15632 ;
  assign y18043 = ~n7684 ;
  assign y18044 = ~n43517 ;
  assign y18045 = ~n43521 ;
  assign y18046 = ~n43524 ;
  assign y18047 = ~n43525 ;
  assign y18048 = n43529 ;
  assign y18049 = ~1'b0 ;
  assign y18050 = ~n43530 ;
  assign y18051 = n43532 ;
  assign y18052 = n43534 ;
  assign y18053 = ~n43536 ;
  assign y18054 = ~n43539 ;
  assign y18055 = ~n43540 ;
  assign y18056 = n43541 ;
  assign y18057 = ~n43542 ;
  assign y18058 = n43543 ;
  assign y18059 = ~1'b0 ;
  assign y18060 = n43544 ;
  assign y18061 = ~n43545 ;
  assign y18062 = ~1'b0 ;
  assign y18063 = ~n43546 ;
  assign y18064 = ~n43548 ;
  assign y18065 = ~n43550 ;
  assign y18066 = n43552 ;
  assign y18067 = ~n43553 ;
  assign y18068 = ~n43557 ;
  assign y18069 = ~1'b0 ;
  assign y18070 = ~1'b0 ;
  assign y18071 = ~1'b0 ;
  assign y18072 = ~1'b0 ;
  assign y18073 = ~n43559 ;
  assign y18074 = n43561 ;
  assign y18075 = ~n43563 ;
  assign y18076 = ~1'b0 ;
  assign y18077 = ~n43564 ;
  assign y18078 = n697 ;
  assign y18079 = n43567 ;
  assign y18080 = n43571 ;
  assign y18081 = n43572 ;
  assign y18082 = ~n35371 ;
  assign y18083 = ~n43575 ;
  assign y18084 = 1'b0 ;
  assign y18085 = n43577 ;
  assign y18086 = ~n43579 ;
  assign y18087 = ~1'b0 ;
  assign y18088 = n43580 ;
  assign y18089 = ~n43588 ;
  assign y18090 = n43589 ;
  assign y18091 = ~n43591 ;
  assign y18092 = ~1'b0 ;
  assign y18093 = ~n43592 ;
  assign y18094 = ~1'b0 ;
  assign y18095 = ~1'b0 ;
  assign y18096 = ~n43596 ;
  assign y18097 = n43600 ;
  assign y18098 = n43602 ;
  assign y18099 = ~n43603 ;
  assign y18100 = ~n43606 ;
  assign y18101 = n43607 ;
  assign y18102 = n43611 ;
  assign y18103 = n43612 ;
  assign y18104 = ~n43616 ;
  assign y18105 = n43618 ;
  assign y18106 = ~n43619 ;
  assign y18107 = n43621 ;
  assign y18108 = ~1'b0 ;
  assign y18109 = ~n43622 ;
  assign y18110 = ~n43623 ;
  assign y18111 = n43626 ;
  assign y18112 = n43627 ;
  assign y18113 = n43628 ;
  assign y18114 = ~n43630 ;
  assign y18115 = ~n43632 ;
  assign y18116 = ~n43633 ;
  assign y18117 = ~n43644 ;
  assign y18118 = n43645 ;
  assign y18119 = ~n43648 ;
  assign y18120 = n43649 ;
  assign y18121 = ~n43653 ;
  assign y18122 = ~n43654 ;
  assign y18123 = n43655 ;
  assign y18124 = n43657 ;
  assign y18125 = n43658 ;
  assign y18126 = ~n43661 ;
  assign y18127 = ~1'b0 ;
  assign y18128 = n43664 ;
  assign y18129 = ~n43666 ;
  assign y18130 = n43667 ;
  assign y18131 = n43669 ;
  assign y18132 = n43670 ;
  assign y18133 = ~n43672 ;
  assign y18134 = ~1'b0 ;
  assign y18135 = n43673 ;
  assign y18136 = ~n43675 ;
  assign y18137 = ~n43676 ;
  assign y18138 = n43162 ;
  assign y18139 = ~n43679 ;
  assign y18140 = n43680 ;
  assign y18141 = n43682 ;
  assign y18142 = n43684 ;
  assign y18143 = n43688 ;
  assign y18144 = ~n43690 ;
  assign y18145 = ~n43692 ;
  assign y18146 = ~n43700 ;
  assign y18147 = ~n43701 ;
  assign y18148 = ~1'b0 ;
  assign y18149 = ~1'b0 ;
  assign y18150 = ~n43704 ;
  assign y18151 = ~n43705 ;
  assign y18152 = ~n43708 ;
  assign y18153 = n43711 ;
  assign y18154 = n43717 ;
  assign y18155 = ~n43720 ;
  assign y18156 = ~1'b0 ;
  assign y18157 = n43723 ;
  assign y18158 = n43727 ;
  assign y18159 = n43730 ;
  assign y18160 = n28248 ;
  assign y18161 = n43732 ;
  assign y18162 = ~n43733 ;
  assign y18163 = ~n43734 ;
  assign y18164 = ~n43739 ;
  assign y18165 = ~1'b0 ;
  assign y18166 = ~1'b0 ;
  assign y18167 = n43741 ;
  assign y18168 = n43745 ;
  assign y18169 = ~n43750 ;
  assign y18170 = ~n43752 ;
  assign y18171 = n43754 ;
  assign y18172 = ~n43757 ;
  assign y18173 = n43758 ;
  assign y18174 = n43759 ;
  assign y18175 = ~1'b0 ;
  assign y18176 = ~n43761 ;
  assign y18177 = ~n43763 ;
  assign y18178 = n43765 ;
  assign y18179 = ~1'b0 ;
  assign y18180 = ~1'b0 ;
  assign y18181 = n43772 ;
  assign y18182 = ~n43773 ;
  assign y18183 = n43774 ;
  assign y18184 = n43779 ;
  assign y18185 = ~n43782 ;
  assign y18186 = n43786 ;
  assign y18187 = 1'b0 ;
  assign y18188 = ~n43790 ;
  assign y18189 = ~1'b0 ;
  assign y18190 = ~1'b0 ;
  assign y18191 = n9596 ;
  assign y18192 = ~n43792 ;
  assign y18193 = n43794 ;
  assign y18194 = ~1'b0 ;
  assign y18195 = ~1'b0 ;
  assign y18196 = n43799 ;
  assign y18197 = ~n43800 ;
  assign y18198 = ~n43801 ;
  assign y18199 = n6418 ;
  assign y18200 = ~n43804 ;
  assign y18201 = ~n33938 ;
  assign y18202 = ~n43811 ;
  assign y18203 = n29828 ;
  assign y18204 = ~n43815 ;
  assign y18205 = ~n43816 ;
  assign y18206 = n43818 ;
  assign y18207 = n43820 ;
  assign y18208 = n43821 ;
  assign y18209 = ~1'b0 ;
  assign y18210 = ~n43823 ;
  assign y18211 = n43824 ;
  assign y18212 = n43826 ;
  assign y18213 = ~n43829 ;
  assign y18214 = n43831 ;
  assign y18215 = n43833 ;
  assign y18216 = ~n43834 ;
  assign y18217 = ~1'b0 ;
  assign y18218 = ~n43837 ;
  assign y18219 = n43842 ;
  assign y18220 = 1'b0 ;
  assign y18221 = n43844 ;
  assign y18222 = n43851 ;
  assign y18223 = ~1'b0 ;
  assign y18224 = n43853 ;
  assign y18225 = n43858 ;
  assign y18226 = n19503 ;
  assign y18227 = ~1'b0 ;
  assign y18228 = ~n43859 ;
  assign y18229 = n43862 ;
  assign y18230 = ~n43863 ;
  assign y18231 = ~1'b0 ;
  assign y18232 = n43866 ;
  assign y18233 = ~1'b0 ;
  assign y18234 = ~1'b0 ;
  assign y18235 = ~n43867 ;
  assign y18236 = n43871 ;
  assign y18237 = n43872 ;
  assign y18238 = ~n43873 ;
  assign y18239 = ~1'b0 ;
  assign y18240 = ~n43876 ;
  assign y18241 = ~1'b0 ;
  assign y18242 = ~n43878 ;
  assign y18243 = ~1'b0 ;
  assign y18244 = ~1'b0 ;
  assign y18245 = n43885 ;
  assign y18246 = n43886 ;
  assign y18247 = ~n43887 ;
  assign y18248 = ~n43888 ;
  assign y18249 = n43890 ;
  assign y18250 = ~n43892 ;
  assign y18251 = ~1'b0 ;
  assign y18252 = ~n43896 ;
  assign y18253 = ~1'b0 ;
  assign y18254 = ~n43897 ;
  assign y18255 = n43899 ;
  assign y18256 = ~n43900 ;
  assign y18257 = n43904 ;
  assign y18258 = ~1'b0 ;
  assign y18259 = ~1'b0 ;
  assign y18260 = n43908 ;
  assign y18261 = ~1'b0 ;
  assign y18262 = ~n43913 ;
  assign y18263 = ~1'b0 ;
  assign y18264 = ~n43914 ;
  assign y18265 = ~n43917 ;
  assign y18266 = n43920 ;
  assign y18267 = ~1'b0 ;
  assign y18268 = ~n43923 ;
  assign y18269 = n43924 ;
  assign y18270 = ~1'b0 ;
  assign y18271 = ~1'b0 ;
  assign y18272 = ~n43929 ;
  assign y18273 = ~n43935 ;
  assign y18274 = ~n43936 ;
  assign y18275 = n43937 ;
  assign y18276 = n37567 ;
  assign y18277 = ~1'b0 ;
  assign y18278 = n43938 ;
  assign y18279 = n43939 ;
  assign y18280 = ~1'b0 ;
  assign y18281 = ~n785 ;
  assign y18282 = n43942 ;
  assign y18283 = ~n43945 ;
  assign y18284 = n43946 ;
  assign y18285 = ~1'b0 ;
  assign y18286 = ~n43947 ;
  assign y18287 = n43948 ;
  assign y18288 = ~n43950 ;
  assign y18289 = ~1'b0 ;
  assign y18290 = n43952 ;
  assign y18291 = n43956 ;
  assign y18292 = ~1'b0 ;
  assign y18293 = ~1'b0 ;
  assign y18294 = n43958 ;
  assign y18295 = n43960 ;
  assign y18296 = n43965 ;
  assign y18297 = ~1'b0 ;
  assign y18298 = ~n43967 ;
  assign y18299 = ~n43968 ;
  assign y18300 = ~n43971 ;
  assign y18301 = ~1'b0 ;
  assign y18302 = ~n3715 ;
  assign y18303 = ~n43972 ;
  assign y18304 = ~n43974 ;
  assign y18305 = n43975 ;
  assign y18306 = ~n43977 ;
  assign y18307 = ~n43981 ;
  assign y18308 = ~n43985 ;
  assign y18309 = n43988 ;
  assign y18310 = n43991 ;
  assign y18311 = ~n38014 ;
  assign y18312 = ~n43992 ;
  assign y18313 = ~n43994 ;
  assign y18314 = ~n43995 ;
  assign y18315 = ~n43998 ;
  assign y18316 = ~1'b0 ;
  assign y18317 = ~1'b0 ;
  assign y18318 = n44001 ;
  assign y18319 = n44003 ;
  assign y18320 = n44008 ;
  assign y18321 = ~n44009 ;
  assign y18322 = ~n44010 ;
  assign y18323 = n44011 ;
  assign y18324 = n44015 ;
  assign y18325 = n44017 ;
  assign y18326 = ~1'b0 ;
  assign y18327 = ~1'b0 ;
  assign y18328 = ~n44019 ;
  assign y18329 = n44020 ;
  assign y18330 = n44022 ;
  assign y18331 = n44030 ;
  assign y18332 = ~n44032 ;
  assign y18333 = ~n44033 ;
  assign y18334 = n44037 ;
  assign y18335 = n44038 ;
  assign y18336 = n44039 ;
  assign y18337 = ~n44040 ;
  assign y18338 = ~1'b0 ;
  assign y18339 = ~n44042 ;
  assign y18340 = ~n44045 ;
  assign y18341 = n44048 ;
  assign y18342 = n44049 ;
  assign y18343 = ~n44053 ;
  assign y18344 = ~1'b0 ;
  assign y18345 = n44054 ;
  assign y18346 = ~n44055 ;
  assign y18347 = x157 ;
  assign y18348 = ~n44056 ;
  assign y18349 = n44060 ;
  assign y18350 = ~n44061 ;
  assign y18351 = ~n44063 ;
  assign y18352 = n1481 ;
  assign y18353 = n44064 ;
  assign y18354 = n44065 ;
  assign y18355 = n44066 ;
  assign y18356 = 1'b0 ;
  assign y18357 = n44071 ;
  assign y18358 = n44072 ;
  assign y18359 = ~1'b0 ;
  assign y18360 = ~1'b0 ;
  assign y18361 = ~n44073 ;
  assign y18362 = ~n44075 ;
  assign y18363 = ~1'b0 ;
  assign y18364 = ~1'b0 ;
  assign y18365 = n44076 ;
  assign y18366 = ~n44078 ;
  assign y18367 = n44082 ;
  assign y18368 = n44085 ;
  assign y18369 = n44091 ;
  assign y18370 = ~n44093 ;
  assign y18371 = n44096 ;
  assign y18372 = ~n44097 ;
  assign y18373 = ~1'b0 ;
  assign y18374 = n44098 ;
  assign y18375 = n44099 ;
  assign y18376 = n44100 ;
  assign y18377 = ~n21563 ;
  assign y18378 = ~1'b0 ;
  assign y18379 = n24129 ;
  assign y18380 = n44102 ;
  assign y18381 = ~1'b0 ;
  assign y18382 = n44104 ;
  assign y18383 = ~n44106 ;
  assign y18384 = ~n44107 ;
  assign y18385 = ~n44109 ;
  assign y18386 = n44112 ;
  assign y18387 = n44113 ;
  assign y18388 = ~n44115 ;
  assign y18389 = ~n44118 ;
  assign y18390 = n44121 ;
  assign y18391 = n44123 ;
  assign y18392 = ~1'b0 ;
  assign y18393 = n4514 ;
  assign y18394 = n44128 ;
  assign y18395 = ~n44129 ;
  assign y18396 = ~1'b0 ;
  assign y18397 = ~1'b0 ;
  assign y18398 = ~n44131 ;
  assign y18399 = n44135 ;
  assign y18400 = n44136 ;
  assign y18401 = ~1'b0 ;
  assign y18402 = ~1'b0 ;
  assign y18403 = ~n44139 ;
  assign y18404 = n44140 ;
  assign y18405 = ~1'b0 ;
  assign y18406 = ~n44142 ;
  assign y18407 = 1'b0 ;
  assign y18408 = ~n44144 ;
  assign y18409 = ~n44146 ;
  assign y18410 = ~1'b0 ;
  assign y18411 = ~n44147 ;
  assign y18412 = ~n44150 ;
  assign y18413 = ~n44153 ;
  assign y18414 = ~n44154 ;
  assign y18415 = ~n44156 ;
  assign y18416 = ~n44160 ;
  assign y18417 = ~1'b0 ;
  assign y18418 = n44165 ;
  assign y18419 = ~1'b0 ;
  assign y18420 = ~n44169 ;
  assign y18421 = ~n44176 ;
  assign y18422 = n44179 ;
  assign y18423 = ~n44180 ;
  assign y18424 = ~n44181 ;
  assign y18425 = ~n44182 ;
  assign y18426 = n44184 ;
  assign y18427 = ~1'b0 ;
  assign y18428 = ~n44187 ;
  assign y18429 = ~1'b0 ;
  assign y18430 = ~1'b0 ;
  assign y18431 = ~n44189 ;
  assign y18432 = ~n44191 ;
  assign y18433 = n44197 ;
  assign y18434 = n44198 ;
  assign y18435 = ~n44199 ;
  assign y18436 = ~n44201 ;
  assign y18437 = ~1'b0 ;
  assign y18438 = ~n44204 ;
  assign y18439 = n44206 ;
  assign y18440 = n44208 ;
  assign y18441 = n44212 ;
  assign y18442 = n44219 ;
  assign y18443 = n44220 ;
  assign y18444 = ~n44221 ;
  assign y18445 = ~n44224 ;
  assign y18446 = n44227 ;
  assign y18447 = ~1'b0 ;
  assign y18448 = ~n44229 ;
  assign y18449 = ~n2590 ;
  assign y18450 = ~1'b0 ;
  assign y18451 = ~1'b0 ;
  assign y18452 = ~1'b0 ;
  assign y18453 = n44231 ;
  assign y18454 = 1'b0 ;
  assign y18455 = ~n44239 ;
  assign y18456 = ~n44242 ;
  assign y18457 = ~1'b0 ;
  assign y18458 = ~n44245 ;
  assign y18459 = n44249 ;
  assign y18460 = n44250 ;
  assign y18461 = n44252 ;
  assign y18462 = n44255 ;
  assign y18463 = n44256 ;
  assign y18464 = n44257 ;
  assign y18465 = ~n44260 ;
  assign y18466 = n44261 ;
  assign y18467 = n44267 ;
  assign y18468 = ~1'b0 ;
  assign y18469 = ~1'b0 ;
  assign y18470 = ~n44272 ;
  assign y18471 = ~1'b0 ;
  assign y18472 = ~n31187 ;
  assign y18473 = ~n44276 ;
  assign y18474 = ~n44277 ;
  assign y18475 = n44278 ;
  assign y18476 = n44283 ;
  assign y18477 = ~1'b0 ;
  assign y18478 = ~1'b0 ;
  assign y18479 = ~n44287 ;
  assign y18480 = n44288 ;
  assign y18481 = ~n44292 ;
  assign y18482 = n44301 ;
  assign y18483 = ~n44303 ;
  assign y18484 = n44304 ;
  assign y18485 = ~n44306 ;
  assign y18486 = ~1'b0 ;
  assign y18487 = ~n44310 ;
  assign y18488 = ~n44312 ;
  assign y18489 = n3007 ;
  assign y18490 = n44314 ;
  assign y18491 = n44316 ;
  assign y18492 = n44320 ;
  assign y18493 = n44323 ;
  assign y18494 = ~n44326 ;
  assign y18495 = ~n44327 ;
  assign y18496 = n44328 ;
  assign y18497 = ~1'b0 ;
  assign y18498 = ~n44329 ;
  assign y18499 = n44333 ;
  assign y18500 = ~1'b0 ;
  assign y18501 = n44337 ;
  assign y18502 = ~n44341 ;
  assign y18503 = n44344 ;
  assign y18504 = n44349 ;
  assign y18505 = ~n44352 ;
  assign y18506 = ~n44355 ;
  assign y18507 = ~1'b0 ;
  assign y18508 = n44356 ;
  assign y18509 = n44357 ;
  assign y18510 = ~n44360 ;
  assign y18511 = ~n44361 ;
  assign y18512 = ~n44363 ;
  assign y18513 = n44367 ;
  assign y18514 = ~n44368 ;
  assign y18515 = n44369 ;
  assign y18516 = n44373 ;
  assign y18517 = ~n44375 ;
  assign y18518 = n44376 ;
  assign y18519 = ~1'b0 ;
  assign y18520 = ~n44380 ;
  assign y18521 = ~1'b0 ;
  assign y18522 = ~n44383 ;
  assign y18523 = ~n44387 ;
  assign y18524 = n44390 ;
  assign y18525 = ~n44391 ;
  assign y18526 = ~n44393 ;
  assign y18527 = ~n44394 ;
  assign y18528 = n44395 ;
  assign y18529 = n44398 ;
  assign y18530 = n44401 ;
  assign y18531 = n44403 ;
  assign y18532 = n44404 ;
  assign y18533 = n44407 ;
  assign y18534 = ~n44408 ;
  assign y18535 = n44410 ;
  assign y18536 = 1'b0 ;
  assign y18537 = n44411 ;
  assign y18538 = ~1'b0 ;
  assign y18539 = n44413 ;
  assign y18540 = ~1'b0 ;
  assign y18541 = ~n44414 ;
  assign y18542 = ~1'b0 ;
  assign y18543 = ~1'b0 ;
  assign y18544 = n44417 ;
  assign y18545 = ~n44420 ;
  assign y18546 = ~1'b0 ;
  assign y18547 = n44422 ;
  assign y18548 = ~n44423 ;
  assign y18549 = ~1'b0 ;
  assign y18550 = ~n44428 ;
  assign y18551 = ~1'b0 ;
  assign y18552 = n44431 ;
  assign y18553 = ~n44432 ;
  assign y18554 = ~n44436 ;
  assign y18555 = ~n44441 ;
  assign y18556 = ~n44445 ;
  assign y18557 = ~n44448 ;
  assign y18558 = n44451 ;
  assign y18559 = ~1'b0 ;
  assign y18560 = n44452 ;
  assign y18561 = n44453 ;
  assign y18562 = n44456 ;
  assign y18563 = n44460 ;
  assign y18564 = ~n44462 ;
  assign y18565 = ~n39398 ;
  assign y18566 = ~1'b0 ;
  assign y18567 = ~n44466 ;
  assign y18568 = ~1'b0 ;
  assign y18569 = n44468 ;
  assign y18570 = n44471 ;
  assign y18571 = ~n44473 ;
  assign y18572 = ~n44474 ;
  assign y18573 = ~n44476 ;
  assign y18574 = ~1'b0 ;
  assign y18575 = n44480 ;
  assign y18576 = ~1'b0 ;
  assign y18577 = n44481 ;
  assign y18578 = ~n44484 ;
  assign y18579 = n44485 ;
  assign y18580 = ~n44488 ;
  assign y18581 = ~n44491 ;
  assign y18582 = n44492 ;
  assign y18583 = ~1'b0 ;
  assign y18584 = ~n44493 ;
  assign y18585 = ~n44494 ;
  assign y18586 = n44496 ;
  assign y18587 = ~1'b0 ;
  assign y18588 = ~n44497 ;
  assign y18589 = ~n44499 ;
  assign y18590 = n44500 ;
  assign y18591 = ~1'b0 ;
  assign y18592 = n13554 ;
  assign y18593 = n44505 ;
  assign y18594 = n44506 ;
  assign y18595 = n44508 ;
  assign y18596 = ~n44509 ;
  assign y18597 = n44510 ;
  assign y18598 = ~n44511 ;
  assign y18599 = n44514 ;
  assign y18600 = ~n44516 ;
  assign y18601 = n44517 ;
  assign y18602 = ~1'b0 ;
  assign y18603 = ~1'b0 ;
  assign y18604 = ~n44518 ;
  assign y18605 = ~n44519 ;
  assign y18606 = n44520 ;
  assign y18607 = ~n44521 ;
  assign y18608 = ~n44524 ;
  assign y18609 = ~n44525 ;
  assign y18610 = n44536 ;
  assign y18611 = ~1'b0 ;
  assign y18612 = 1'b0 ;
  assign y18613 = n44538 ;
  assign y18614 = ~n44539 ;
  assign y18615 = n44547 ;
  assign y18616 = ~n44550 ;
  assign y18617 = ~1'b0 ;
  assign y18618 = ~n44551 ;
  assign y18619 = ~n44553 ;
  assign y18620 = ~n2754 ;
  assign y18621 = ~1'b0 ;
  assign y18622 = n44555 ;
  assign y18623 = ~1'b0 ;
  assign y18624 = ~n44559 ;
  assign y18625 = ~n44566 ;
  assign y18626 = n44567 ;
  assign y18627 = ~n26175 ;
  assign y18628 = n44569 ;
  assign y18629 = n44577 ;
  assign y18630 = n44578 ;
  assign y18631 = n44584 ;
  assign y18632 = ~n44586 ;
  assign y18633 = ~1'b0 ;
  assign y18634 = ~n44588 ;
  assign y18635 = n44590 ;
  assign y18636 = n44592 ;
  assign y18637 = ~n44598 ;
  assign y18638 = ~1'b0 ;
  assign y18639 = ~n44601 ;
  assign y18640 = n44602 ;
  assign y18641 = n44607 ;
  assign y18642 = n44609 ;
  assign y18643 = ~1'b0 ;
  assign y18644 = ~n44610 ;
  assign y18645 = ~1'b0 ;
  assign y18646 = ~1'b0 ;
  assign y18647 = ~n44612 ;
  assign y18648 = ~n44613 ;
  assign y18649 = ~n44616 ;
  assign y18650 = n44617 ;
  assign y18651 = ~n44621 ;
  assign y18652 = n44623 ;
  assign y18653 = n44625 ;
  assign y18654 = ~1'b0 ;
  assign y18655 = n44626 ;
  assign y18656 = n44627 ;
  assign y18657 = ~n44629 ;
  assign y18658 = n44632 ;
  assign y18659 = ~n44637 ;
  assign y18660 = n44643 ;
  assign y18661 = ~1'b0 ;
  assign y18662 = ~n44645 ;
  assign y18663 = ~1'b0 ;
  assign y18664 = ~n44646 ;
  assign y18665 = ~n44647 ;
  assign y18666 = ~n44648 ;
  assign y18667 = ~n44655 ;
  assign y18668 = n44656 ;
  assign y18669 = ~1'b0 ;
  assign y18670 = ~n44657 ;
  assign y18671 = ~n44660 ;
  assign y18672 = n44664 ;
  assign y18673 = ~1'b0 ;
  assign y18674 = ~1'b0 ;
  assign y18675 = ~1'b0 ;
  assign y18676 = n44666 ;
  assign y18677 = ~n44667 ;
  assign y18678 = 1'b0 ;
  assign y18679 = n44668 ;
  assign y18680 = ~n44669 ;
  assign y18681 = n44672 ;
  assign y18682 = ~n44676 ;
  assign y18683 = n44678 ;
  assign y18684 = ~n44680 ;
  assign y18685 = n44683 ;
  assign y18686 = ~n44684 ;
  assign y18687 = ~1'b0 ;
  assign y18688 = n44685 ;
  assign y18689 = ~n44687 ;
  assign y18690 = ~n44690 ;
  assign y18691 = ~1'b0 ;
  assign y18692 = n44694 ;
  assign y18693 = ~1'b0 ;
  assign y18694 = n44696 ;
  assign y18695 = ~1'b0 ;
  assign y18696 = ~n44697 ;
  assign y18697 = n44699 ;
  assign y18698 = n44701 ;
  assign y18699 = ~n44702 ;
  assign y18700 = ~n44706 ;
  assign y18701 = n44711 ;
  assign y18702 = ~n44713 ;
  assign y18703 = ~1'b0 ;
  assign y18704 = ~n44715 ;
  assign y18705 = ~1'b0 ;
  assign y18706 = ~n44722 ;
  assign y18707 = ~n44724 ;
  assign y18708 = n44731 ;
  assign y18709 = n44732 ;
  assign y18710 = n44734 ;
  assign y18711 = ~n44735 ;
  assign y18712 = n44736 ;
  assign y18713 = ~1'b0 ;
  assign y18714 = ~1'b0 ;
  assign y18715 = n44738 ;
  assign y18716 = ~1'b0 ;
  assign y18717 = n44739 ;
  assign y18718 = ~n44742 ;
  assign y18719 = ~n5492 ;
  assign y18720 = n44743 ;
  assign y18721 = n44744 ;
  assign y18722 = ~n44746 ;
  assign y18723 = ~1'b0 ;
  assign y18724 = ~n44753 ;
  assign y18725 = n44755 ;
  assign y18726 = n44758 ;
  assign y18727 = n44760 ;
  assign y18728 = ~n44768 ;
  assign y18729 = n44773 ;
  assign y18730 = ~n44774 ;
  assign y18731 = ~n44775 ;
  assign y18732 = 1'b0 ;
  assign y18733 = n44776 ;
  assign y18734 = ~n44777 ;
  assign y18735 = ~1'b0 ;
  assign y18736 = n44780 ;
  assign y18737 = ~n44781 ;
  assign y18738 = ~n44786 ;
  assign y18739 = ~n44789 ;
  assign y18740 = ~n44793 ;
  assign y18741 = n44794 ;
  assign y18742 = ~n44797 ;
  assign y18743 = ~n44801 ;
  assign y18744 = n44802 ;
  assign y18745 = ~1'b0 ;
  assign y18746 = n44803 ;
  assign y18747 = n44804 ;
  assign y18748 = n44807 ;
  assign y18749 = n44817 ;
  assign y18750 = n23967 ;
  assign y18751 = ~n44820 ;
  assign y18752 = n44821 ;
  assign y18753 = n44822 ;
  assign y18754 = n44825 ;
  assign y18755 = 1'b0 ;
  assign y18756 = ~1'b0 ;
  assign y18757 = n44827 ;
  assign y18758 = n44829 ;
  assign y18759 = n44831 ;
  assign y18760 = ~1'b0 ;
  assign y18761 = ~1'b0 ;
  assign y18762 = n44833 ;
  assign y18763 = n44835 ;
  assign y18764 = ~1'b0 ;
  assign y18765 = n33336 ;
  assign y18766 = ~1'b0 ;
  assign y18767 = n44837 ;
  assign y18768 = ~n44838 ;
  assign y18769 = ~n44839 ;
  assign y18770 = n44845 ;
  assign y18771 = n44847 ;
  assign y18772 = n37209 ;
  assign y18773 = n44849 ;
  assign y18774 = ~n44851 ;
  assign y18775 = ~n44852 ;
  assign y18776 = ~1'b0 ;
  assign y18777 = n44855 ;
  assign y18778 = ~n44861 ;
  assign y18779 = n44862 ;
  assign y18780 = n44866 ;
  assign y18781 = ~n44868 ;
  assign y18782 = ~1'b0 ;
  assign y18783 = 1'b0 ;
  assign y18784 = ~n44871 ;
  assign y18785 = n44873 ;
  assign y18786 = ~1'b0 ;
  assign y18787 = ~1'b0 ;
  assign y18788 = 1'b0 ;
  assign y18789 = n44877 ;
  assign y18790 = ~n44878 ;
  assign y18791 = n44880 ;
  assign y18792 = ~1'b0 ;
  assign y18793 = ~n44882 ;
  assign y18794 = ~n44883 ;
  assign y18795 = ~n44885 ;
  assign y18796 = n44888 ;
  assign y18797 = ~n44891 ;
  assign y18798 = ~n44892 ;
  assign y18799 = ~n5011 ;
  assign y18800 = ~1'b0 ;
  assign y18801 = ~n44894 ;
  assign y18802 = ~n44895 ;
  assign y18803 = ~1'b0 ;
  assign y18804 = ~1'b0 ;
  assign y18805 = n44896 ;
  assign y18806 = ~n44897 ;
  assign y18807 = n44900 ;
  assign y18808 = n44902 ;
  assign y18809 = n44904 ;
  assign y18810 = ~n44906 ;
  assign y18811 = ~n44908 ;
  assign y18812 = ~n44914 ;
  assign y18813 = ~n44917 ;
  assign y18814 = ~1'b0 ;
  assign y18815 = n44918 ;
  assign y18816 = ~n44919 ;
  assign y18817 = ~1'b0 ;
  assign y18818 = ~n44921 ;
  assign y18819 = n44923 ;
  assign y18820 = n44924 ;
  assign y18821 = ~n44925 ;
  assign y18822 = ~n44926 ;
  assign y18823 = n43903 ;
  assign y18824 = ~n44928 ;
  assign y18825 = n44931 ;
  assign y18826 = n44935 ;
  assign y18827 = n44937 ;
  assign y18828 = ~1'b0 ;
  assign y18829 = n44940 ;
  assign y18830 = ~n44943 ;
  assign y18831 = ~1'b0 ;
  assign y18832 = n44944 ;
  assign y18833 = n44946 ;
  assign y18834 = ~n44947 ;
  assign y18835 = ~n44951 ;
  assign y18836 = n44953 ;
  assign y18837 = n44955 ;
  assign y18838 = ~n44962 ;
  assign y18839 = ~1'b0 ;
  assign y18840 = ~1'b0 ;
  assign y18841 = ~1'b0 ;
  assign y18842 = ~1'b0 ;
  assign y18843 = n44964 ;
  assign y18844 = ~n44971 ;
  assign y18845 = ~n44973 ;
  assign y18846 = n44974 ;
  assign y18847 = n44977 ;
  assign y18848 = n44978 ;
  assign y18849 = n44979 ;
  assign y18850 = n44981 ;
  assign y18851 = ~n44984 ;
  assign y18852 = n44988 ;
  assign y18853 = n44989 ;
  assign y18854 = ~n37251 ;
  assign y18855 = n44992 ;
  assign y18856 = n44995 ;
  assign y18857 = ~1'b0 ;
  assign y18858 = ~n44996 ;
  assign y18859 = ~n45000 ;
  assign y18860 = ~n45003 ;
  assign y18861 = ~n45004 ;
  assign y18862 = n45008 ;
  assign y18863 = ~1'b0 ;
  assign y18864 = ~n45010 ;
  assign y18865 = ~n45014 ;
  assign y18866 = n45016 ;
  assign y18867 = ~n45022 ;
  assign y18868 = ~n45026 ;
  assign y18869 = ~n3344 ;
  assign y18870 = n45027 ;
  assign y18871 = n45028 ;
  assign y18872 = ~n45029 ;
  assign y18873 = 1'b0 ;
  assign y18874 = ~n45034 ;
  assign y18875 = n45035 ;
  assign y18876 = ~n40590 ;
  assign y18877 = n45037 ;
  assign y18878 = 1'b0 ;
  assign y18879 = ~1'b0 ;
  assign y18880 = n45038 ;
  assign y18881 = n39255 ;
  assign y18882 = n45042 ;
  assign y18883 = n45046 ;
  assign y18884 = ~n45048 ;
  assign y18885 = n8836 ;
  assign y18886 = ~n35019 ;
  assign y18887 = ~n45050 ;
  assign y18888 = ~1'b0 ;
  assign y18889 = ~n45054 ;
  assign y18890 = ~n45055 ;
  assign y18891 = ~n45056 ;
  assign y18892 = n45059 ;
  assign y18893 = ~n45060 ;
  assign y18894 = ~1'b0 ;
  assign y18895 = n45061 ;
  assign y18896 = ~n45062 ;
  assign y18897 = ~1'b0 ;
  assign y18898 = n45064 ;
  assign y18899 = ~1'b0 ;
  assign y18900 = n45065 ;
  assign y18901 = ~n45066 ;
  assign y18902 = ~1'b0 ;
  assign y18903 = ~n45069 ;
  assign y18904 = ~1'b0 ;
  assign y18905 = n45078 ;
  assign y18906 = n45081 ;
  assign y18907 = ~1'b0 ;
  assign y18908 = ~n45082 ;
  assign y18909 = ~n45083 ;
  assign y18910 = n45084 ;
  assign y18911 = ~n45087 ;
  assign y18912 = ~1'b0 ;
  assign y18913 = ~1'b0 ;
  assign y18914 = n45091 ;
  assign y18915 = ~1'b0 ;
  assign y18916 = n45094 ;
  assign y18917 = ~1'b0 ;
  assign y18918 = n45096 ;
  assign y18919 = ~n45100 ;
  assign y18920 = ~n45101 ;
  assign y18921 = ~n45105 ;
  assign y18922 = ~1'b0 ;
  assign y18923 = n45106 ;
  assign y18924 = ~1'b0 ;
  assign y18925 = n45110 ;
  assign y18926 = n45112 ;
  assign y18927 = n45113 ;
  assign y18928 = ~n45114 ;
  assign y18929 = n45115 ;
  assign y18930 = n45120 ;
  assign y18931 = ~n45125 ;
  assign y18932 = n45128 ;
  assign y18933 = ~n45130 ;
  assign y18934 = ~n45133 ;
  assign y18935 = n45135 ;
  assign y18936 = n45138 ;
  assign y18937 = ~1'b0 ;
  assign y18938 = n45139 ;
  assign y18939 = ~n45143 ;
  assign y18940 = n45145 ;
  assign y18941 = n45166 ;
  assign y18942 = ~n45168 ;
  assign y18943 = ~n45170 ;
  assign y18944 = ~n45172 ;
  assign y18945 = ~n45173 ;
  assign y18946 = n23037 ;
  assign y18947 = ~1'b0 ;
  assign y18948 = n45174 ;
  assign y18949 = ~n45176 ;
  assign y18950 = n45179 ;
  assign y18951 = n45181 ;
  assign y18952 = ~1'b0 ;
  assign y18953 = n45185 ;
  assign y18954 = n45186 ;
  assign y18955 = n45189 ;
  assign y18956 = ~n45190 ;
  assign y18957 = ~1'b0 ;
  assign y18958 = n45194 ;
  assign y18959 = n45199 ;
  assign y18960 = ~n45200 ;
  assign y18961 = ~n45201 ;
  assign y18962 = n45204 ;
  assign y18963 = ~1'b0 ;
  assign y18964 = ~n45209 ;
  assign y18965 = ~n45211 ;
  assign y18966 = ~1'b0 ;
  assign y18967 = ~1'b0 ;
  assign y18968 = ~1'b0 ;
  assign y18969 = ~n45213 ;
  assign y18970 = n45215 ;
  assign y18971 = ~n45217 ;
  assign y18972 = n45220 ;
  assign y18973 = n45223 ;
  assign y18974 = ~n45225 ;
  assign y18975 = ~n45227 ;
  assign y18976 = n45229 ;
  assign y18977 = ~n45231 ;
  assign y18978 = ~n45233 ;
  assign y18979 = ~n45235 ;
  assign y18980 = ~1'b0 ;
  assign y18981 = n32786 ;
  assign y18982 = ~n45238 ;
  assign y18983 = ~n45239 ;
  assign y18984 = n45241 ;
  assign y18985 = n45243 ;
  assign y18986 = ~n45246 ;
  assign y18987 = n45247 ;
  assign y18988 = n45252 ;
  assign y18989 = ~1'b0 ;
  assign y18990 = ~n45253 ;
  assign y18991 = n45254 ;
  assign y18992 = ~n45259 ;
  assign y18993 = ~n45260 ;
  assign y18994 = ~n45265 ;
  assign y18995 = ~1'b0 ;
  assign y18996 = n35561 ;
  assign y18997 = ~1'b0 ;
  assign y18998 = ~n45267 ;
  assign y18999 = ~n45269 ;
  assign y19000 = ~n45271 ;
  assign y19001 = n45276 ;
  assign y19002 = n45277 ;
  assign y19003 = n45278 ;
  assign y19004 = n45280 ;
  assign y19005 = ~n11251 ;
  assign y19006 = n45285 ;
  assign y19007 = ~1'b0 ;
  assign y19008 = 1'b0 ;
  assign y19009 = ~n45286 ;
  assign y19010 = ~n45287 ;
  assign y19011 = ~n45288 ;
  assign y19012 = n45290 ;
  assign y19013 = n45293 ;
  assign y19014 = n45303 ;
  assign y19015 = ~n45304 ;
  assign y19016 = ~n45305 ;
  assign y19017 = ~n3649 ;
  assign y19018 = ~1'b0 ;
  assign y19019 = n5478 ;
  assign y19020 = ~n45306 ;
  assign y19021 = ~n45311 ;
  assign y19022 = ~n45312 ;
  assign y19023 = n45319 ;
  assign y19024 = ~1'b0 ;
  assign y19025 = ~n45321 ;
  assign y19026 = ~1'b0 ;
  assign y19027 = ~1'b0 ;
  assign y19028 = ~n45323 ;
  assign y19029 = 1'b0 ;
  assign y19030 = ~n45324 ;
  assign y19031 = n45326 ;
  assign y19032 = ~n45331 ;
  assign y19033 = 1'b0 ;
  assign y19034 = ~n45333 ;
  assign y19035 = ~n45340 ;
  assign y19036 = ~n45341 ;
  assign y19037 = ~n45344 ;
  assign y19038 = n45345 ;
  assign y19039 = ~n45349 ;
  assign y19040 = ~n45351 ;
  assign y19041 = ~n45352 ;
  assign y19042 = n45353 ;
  assign y19043 = n45361 ;
  assign y19044 = n45368 ;
  assign y19045 = ~1'b0 ;
  assign y19046 = ~n45369 ;
  assign y19047 = ~1'b0 ;
  assign y19048 = n45371 ;
  assign y19049 = n45373 ;
  assign y19050 = n45375 ;
  assign y19051 = ~n45380 ;
  assign y19052 = n45381 ;
  assign y19053 = ~n45384 ;
  assign y19054 = n45387 ;
  assign y19055 = ~n45393 ;
  assign y19056 = n45397 ;
  assign y19057 = ~n45398 ;
  assign y19058 = ~1'b0 ;
  assign y19059 = n45399 ;
  assign y19060 = n45400 ;
  assign y19061 = n45403 ;
  assign y19062 = ~n45409 ;
  assign y19063 = ~n45410 ;
  assign y19064 = n45413 ;
  assign y19065 = n45415 ;
  assign y19066 = ~n45416 ;
  assign y19067 = ~n45419 ;
  assign y19068 = ~n45420 ;
  assign y19069 = n45421 ;
  assign y19070 = n45425 ;
  assign y19071 = n45427 ;
  assign y19072 = ~1'b0 ;
  assign y19073 = n45431 ;
  assign y19074 = n45433 ;
  assign y19075 = ~n45437 ;
  assign y19076 = ~n45440 ;
  assign y19077 = ~n45444 ;
  assign y19078 = ~n45449 ;
  assign y19079 = ~n45450 ;
  assign y19080 = ~1'b0 ;
  assign y19081 = ~1'b0 ;
  assign y19082 = ~1'b0 ;
  assign y19083 = ~1'b0 ;
  assign y19084 = ~1'b0 ;
  assign y19085 = ~1'b0 ;
  assign y19086 = ~1'b0 ;
  assign y19087 = ~n45451 ;
  assign y19088 = n45452 ;
  assign y19089 = n45455 ;
  assign y19090 = ~n45456 ;
  assign y19091 = ~n3302 ;
  assign y19092 = ~n45457 ;
  assign y19093 = ~n45459 ;
  assign y19094 = n45460 ;
  assign y19095 = n45462 ;
  assign y19096 = n45467 ;
  assign y19097 = n45471 ;
  assign y19098 = n45473 ;
  assign y19099 = ~n45477 ;
  assign y19100 = ~1'b0 ;
  assign y19101 = n45485 ;
  assign y19102 = n45487 ;
  assign y19103 = ~n45490 ;
  assign y19104 = ~1'b0 ;
  assign y19105 = n45493 ;
  assign y19106 = n45497 ;
  assign y19107 = ~n45501 ;
  assign y19108 = n45506 ;
  assign y19109 = n45507 ;
  assign y19110 = n45508 ;
  assign y19111 = n45510 ;
  assign y19112 = ~n45513 ;
  assign y19113 = ~n45515 ;
  assign y19114 = n45517 ;
  assign y19115 = n45518 ;
  assign y19116 = n45524 ;
  assign y19117 = ~1'b0 ;
  assign y19118 = n45526 ;
  assign y19119 = ~n45528 ;
  assign y19120 = n45533 ;
  assign y19121 = n45538 ;
  assign y19122 = ~1'b0 ;
  assign y19123 = ~n45542 ;
  assign y19124 = ~n45545 ;
  assign y19125 = ~1'b0 ;
  assign y19126 = ~n45547 ;
  assign y19127 = ~1'b0 ;
  assign y19128 = ~n45548 ;
  assign y19129 = ~n45549 ;
  assign y19130 = ~n45551 ;
  assign y19131 = ~n45553 ;
  assign y19132 = ~1'b0 ;
  assign y19133 = ~n38211 ;
  assign y19134 = n45555 ;
  assign y19135 = ~n45559 ;
  assign y19136 = n45562 ;
  assign y19137 = n45563 ;
  assign y19138 = ~1'b0 ;
  assign y19139 = n45564 ;
  assign y19140 = n45565 ;
  assign y19141 = ~n45566 ;
  assign y19142 = ~n8647 ;
  assign y19143 = ~n45567 ;
  assign y19144 = ~1'b0 ;
  assign y19145 = ~n45569 ;
  assign y19146 = ~1'b0 ;
  assign y19147 = ~1'b0 ;
  assign y19148 = n45572 ;
  assign y19149 = ~n45574 ;
  assign y19150 = ~n45575 ;
  assign y19151 = ~n45576 ;
  assign y19152 = ~1'b0 ;
  assign y19153 = n45577 ;
  assign y19154 = ~1'b0 ;
  assign y19155 = n45579 ;
  assign y19156 = n45581 ;
  assign y19157 = n45583 ;
  assign y19158 = n45586 ;
  assign y19159 = 1'b0 ;
  assign y19160 = ~1'b0 ;
  assign y19161 = ~n45588 ;
  assign y19162 = n45589 ;
  assign y19163 = n45596 ;
  assign y19164 = ~1'b0 ;
  assign y19165 = n45597 ;
  assign y19166 = ~n45599 ;
  assign y19167 = ~n45601 ;
  assign y19168 = ~1'b0 ;
  assign y19169 = ~n45603 ;
  assign y19170 = ~n45604 ;
  assign y19171 = ~n45606 ;
  assign y19172 = n45608 ;
  assign y19173 = n45609 ;
  assign y19174 = ~n45611 ;
  assign y19175 = n18191 ;
  assign y19176 = ~n45613 ;
  assign y19177 = ~1'b0 ;
  assign y19178 = ~1'b0 ;
  assign y19179 = ~n45616 ;
  assign y19180 = ~n45617 ;
  assign y19181 = ~n45620 ;
  assign y19182 = n45621 ;
  assign y19183 = ~1'b0 ;
  assign y19184 = n45624 ;
  assign y19185 = ~1'b0 ;
  assign y19186 = ~n45626 ;
  assign y19187 = ~n45627 ;
  assign y19188 = ~n45628 ;
  assign y19189 = ~n45642 ;
  assign y19190 = n45643 ;
  assign y19191 = ~n45645 ;
  assign y19192 = n45647 ;
  assign y19193 = ~n45648 ;
  assign y19194 = ~n45654 ;
  assign y19195 = ~1'b0 ;
  assign y19196 = ~n45659 ;
  assign y19197 = ~n45664 ;
  assign y19198 = ~1'b0 ;
  assign y19199 = n45665 ;
  assign y19200 = ~n45667 ;
  assign y19201 = ~n45669 ;
  assign y19202 = n45672 ;
  assign y19203 = ~1'b0 ;
  assign y19204 = n45674 ;
  assign y19205 = ~1'b0 ;
  assign y19206 = n45678 ;
  assign y19207 = n45680 ;
  assign y19208 = ~n45684 ;
  assign y19209 = n45687 ;
  assign y19210 = ~n45689 ;
  assign y19211 = ~n45697 ;
  assign y19212 = ~n45698 ;
  assign y19213 = n45702 ;
  assign y19214 = ~n45707 ;
  assign y19215 = ~n45709 ;
  assign y19216 = ~1'b0 ;
  assign y19217 = ~n28872 ;
  assign y19218 = n45711 ;
  assign y19219 = n45718 ;
  assign y19220 = ~n45726 ;
  assign y19221 = ~n45728 ;
  assign y19222 = ~n45738 ;
  assign y19223 = n45739 ;
  assign y19224 = ~1'b0 ;
  assign y19225 = n45744 ;
  assign y19226 = ~1'b0 ;
  assign y19227 = ~1'b0 ;
  assign y19228 = ~1'b0 ;
  assign y19229 = n45746 ;
  assign y19230 = ~n45747 ;
  assign y19231 = ~n45748 ;
  assign y19232 = ~n45750 ;
  assign y19233 = n44534 ;
  assign y19234 = ~1'b0 ;
  assign y19235 = ~n45753 ;
  assign y19236 = n45758 ;
  assign y19237 = ~1'b0 ;
  assign y19238 = ~1'b0 ;
  assign y19239 = n45759 ;
  assign y19240 = ~n45760 ;
  assign y19241 = n45761 ;
  assign y19242 = n45764 ;
  assign y19243 = ~n45769 ;
  assign y19244 = n45771 ;
  assign y19245 = ~1'b0 ;
  assign y19246 = ~n45773 ;
  assign y19247 = ~1'b0 ;
  assign y19248 = ~1'b0 ;
  assign y19249 = ~1'b0 ;
  assign y19250 = n45776 ;
  assign y19251 = ~n45779 ;
  assign y19252 = ~n45780 ;
  assign y19253 = n45781 ;
  assign y19254 = ~n45784 ;
  assign y19255 = n45785 ;
  assign y19256 = ~n45788 ;
  assign y19257 = n45791 ;
  assign y19258 = n45792 ;
  assign y19259 = ~n45794 ;
  assign y19260 = ~1'b0 ;
  assign y19261 = n42985 ;
  assign y19262 = n45796 ;
  assign y19263 = n45799 ;
  assign y19264 = ~1'b0 ;
  assign y19265 = n45801 ;
  assign y19266 = ~n45805 ;
  assign y19267 = ~n45807 ;
  assign y19268 = n45809 ;
  assign y19269 = ~1'b0 ;
  assign y19270 = n45810 ;
  assign y19271 = n45817 ;
  assign y19272 = ~n45820 ;
  assign y19273 = ~1'b0 ;
  assign y19274 = ~1'b0 ;
  assign y19275 = n45822 ;
  assign y19276 = ~n45824 ;
  assign y19277 = ~n45826 ;
  assign y19278 = ~1'b0 ;
  assign y19279 = n23867 ;
  assign y19280 = n45827 ;
  assign y19281 = n45831 ;
  assign y19282 = n45832 ;
  assign y19283 = ~n45834 ;
  assign y19284 = ~1'b0 ;
  assign y19285 = ~n45835 ;
  assign y19286 = n45836 ;
  assign y19287 = n45840 ;
  assign y19288 = ~n45841 ;
  assign y19289 = ~n45845 ;
  assign y19290 = ~n45850 ;
  assign y19291 = ~n45851 ;
  assign y19292 = ~n45852 ;
  assign y19293 = ~n45854 ;
  assign y19294 = 1'b0 ;
  assign y19295 = n45855 ;
  assign y19296 = n45856 ;
  assign y19297 = ~n45858 ;
  assign y19298 = n45859 ;
  assign y19299 = ~n7468 ;
  assign y19300 = ~n45860 ;
  assign y19301 = ~n45865 ;
  assign y19302 = ~n45869 ;
  assign y19303 = ~1'b0 ;
  assign y19304 = ~1'b0 ;
  assign y19305 = n45873 ;
  assign y19306 = ~n45879 ;
  assign y19307 = n45881 ;
  assign y19308 = ~1'b0 ;
  assign y19309 = ~n45882 ;
  assign y19310 = ~n45883 ;
  assign y19311 = ~n45884 ;
  assign y19312 = ~n45885 ;
  assign y19313 = n45887 ;
  assign y19314 = ~1'b0 ;
  assign y19315 = ~n45889 ;
  assign y19316 = ~n45891 ;
  assign y19317 = ~n45895 ;
  assign y19318 = n45896 ;
  assign y19319 = n45897 ;
  assign y19320 = ~n45902 ;
  assign y19321 = ~1'b0 ;
  assign y19322 = ~n19770 ;
  assign y19323 = 1'b0 ;
  assign y19324 = ~1'b0 ;
  assign y19325 = n45906 ;
  assign y19326 = ~1'b0 ;
  assign y19327 = ~n45908 ;
  assign y19328 = ~n45910 ;
  assign y19329 = n19737 ;
  assign y19330 = n45911 ;
  assign y19331 = ~1'b0 ;
  assign y19332 = n45912 ;
  assign y19333 = ~1'b0 ;
  assign y19334 = ~n45914 ;
  assign y19335 = ~n45915 ;
  assign y19336 = ~1'b0 ;
  assign y19337 = 1'b0 ;
  assign y19338 = n45918 ;
  assign y19339 = ~n45919 ;
  assign y19340 = n45920 ;
  assign y19341 = n45923 ;
  assign y19342 = ~n45925 ;
  assign y19343 = n45928 ;
  assign y19344 = ~n45929 ;
  assign y19345 = ~n45931 ;
  assign y19346 = ~n45934 ;
  assign y19347 = n45935 ;
  assign y19348 = ~n45939 ;
  assign y19349 = ~n45945 ;
  assign y19350 = ~n45947 ;
  assign y19351 = ~n45948 ;
  assign y19352 = ~n45949 ;
  assign y19353 = n45953 ;
  assign y19354 = ~1'b0 ;
  assign y19355 = ~n45955 ;
  assign y19356 = ~1'b0 ;
  assign y19357 = ~n45957 ;
  assign y19358 = ~n45961 ;
  assign y19359 = ~n45964 ;
  assign y19360 = ~n45967 ;
  assign y19361 = n45973 ;
  assign y19362 = ~n45979 ;
  assign y19363 = ~n45981 ;
  assign y19364 = ~1'b0 ;
  assign y19365 = n45983 ;
  assign y19366 = n36164 ;
  assign y19367 = n45984 ;
  assign y19368 = n45988 ;
  assign y19369 = n45990 ;
  assign y19370 = ~1'b0 ;
  assign y19371 = n45991 ;
  assign y19372 = ~n45997 ;
  assign y19373 = ~n46000 ;
  assign y19374 = ~n46002 ;
  assign y19375 = ~1'b0 ;
  assign y19376 = n46003 ;
  assign y19377 = n46004 ;
  assign y19378 = n46007 ;
  assign y19379 = ~n46011 ;
  assign y19380 = ~n46017 ;
  assign y19381 = ~n46019 ;
  assign y19382 = ~n46020 ;
  assign y19383 = 1'b0 ;
  assign y19384 = n46021 ;
  assign y19385 = n46023 ;
  assign y19386 = ~1'b0 ;
  assign y19387 = n46025 ;
  assign y19388 = ~1'b0 ;
  assign y19389 = ~n46027 ;
  assign y19390 = ~1'b0 ;
  assign y19391 = ~1'b0 ;
  assign y19392 = ~1'b0 ;
  assign y19393 = ~n46028 ;
  assign y19394 = ~n46033 ;
  assign y19395 = ~n46035 ;
  assign y19396 = n46037 ;
  assign y19397 = ~n46040 ;
  assign y19398 = ~n46042 ;
  assign y19399 = n46043 ;
  assign y19400 = ~n17078 ;
  assign y19401 = n46048 ;
  assign y19402 = n46051 ;
  assign y19403 = ~n46054 ;
  assign y19404 = ~n46056 ;
  assign y19405 = n46060 ;
  assign y19406 = n46061 ;
  assign y19407 = ~1'b0 ;
  assign y19408 = ~n46062 ;
  assign y19409 = ~1'b0 ;
  assign y19410 = n32218 ;
  assign y19411 = n46064 ;
  assign y19412 = ~n46068 ;
  assign y19413 = ~n46069 ;
  assign y19414 = ~n46070 ;
  assign y19415 = ~n46072 ;
  assign y19416 = ~1'b0 ;
  assign y19417 = n46074 ;
  assign y19418 = ~1'b0 ;
  assign y19419 = n46079 ;
  assign y19420 = ~n46081 ;
  assign y19421 = ~n33773 ;
  assign y19422 = ~n46083 ;
  assign y19423 = n46089 ;
  assign y19424 = n46092 ;
  assign y19425 = ~n46094 ;
  assign y19426 = ~1'b0 ;
  assign y19427 = ~1'b0 ;
  assign y19428 = ~1'b0 ;
  assign y19429 = n46100 ;
  assign y19430 = ~n46103 ;
  assign y19431 = n46105 ;
  assign y19432 = n46106 ;
  assign y19433 = n21695 ;
  assign y19434 = 1'b0 ;
  assign y19435 = n46108 ;
  assign y19436 = ~n46109 ;
  assign y19437 = ~n46110 ;
  assign y19438 = ~n46113 ;
  assign y19439 = n46115 ;
  assign y19440 = n46117 ;
  assign y19441 = n43296 ;
  assign y19442 = ~n46119 ;
  assign y19443 = n9478 ;
  assign y19444 = ~1'b0 ;
  assign y19445 = ~1'b0 ;
  assign y19446 = n29984 ;
  assign y19447 = n46123 ;
  assign y19448 = ~n46124 ;
  assign y19449 = ~n46128 ;
  assign y19450 = 1'b0 ;
  assign y19451 = ~n46129 ;
  assign y19452 = ~n46134 ;
  assign y19453 = ~n46136 ;
  assign y19454 = ~n46138 ;
  assign y19455 = ~1'b0 ;
  assign y19456 = ~1'b0 ;
  assign y19457 = n46142 ;
  assign y19458 = n46144 ;
  assign y19459 = ~1'b0 ;
  assign y19460 = n46146 ;
  assign y19461 = ~1'b0 ;
  assign y19462 = n46151 ;
  assign y19463 = ~n18365 ;
  assign y19464 = ~n46152 ;
  assign y19465 = ~n46154 ;
  assign y19466 = ~1'b0 ;
  assign y19467 = n46156 ;
  assign y19468 = n46160 ;
  assign y19469 = 1'b0 ;
  assign y19470 = n46162 ;
  assign y19471 = n46163 ;
  assign y19472 = n46164 ;
  assign y19473 = n46169 ;
  assign y19474 = n46172 ;
  assign y19475 = n46173 ;
  assign y19476 = n46175 ;
  assign y19477 = ~n46179 ;
  assign y19478 = ~n46180 ;
  assign y19479 = ~n46185 ;
  assign y19480 = ~n46187 ;
  assign y19481 = n46189 ;
  assign y19482 = n46190 ;
  assign y19483 = n46194 ;
  assign y19484 = n46195 ;
  assign y19485 = n46196 ;
  assign y19486 = n46197 ;
  assign y19487 = ~n46200 ;
  assign y19488 = n46202 ;
  assign y19489 = ~1'b0 ;
  assign y19490 = n46204 ;
  assign y19491 = ~1'b0 ;
  assign y19492 = ~n46213 ;
  assign y19493 = ~1'b0 ;
  assign y19494 = ~n46214 ;
  assign y19495 = n46217 ;
  assign y19496 = n46218 ;
  assign y19497 = ~1'b0 ;
  assign y19498 = ~1'b0 ;
  assign y19499 = ~1'b0 ;
  assign y19500 = ~n46224 ;
  assign y19501 = n46228 ;
  assign y19502 = ~n46235 ;
  assign y19503 = ~n46236 ;
  assign y19504 = ~n8198 ;
  assign y19505 = ~1'b0 ;
  assign y19506 = ~1'b0 ;
  assign y19507 = ~n12671 ;
  assign y19508 = ~n46238 ;
  assign y19509 = n46239 ;
  assign y19510 = ~1'b0 ;
  assign y19511 = ~1'b0 ;
  assign y19512 = ~n46246 ;
  assign y19513 = n46251 ;
  assign y19514 = n46252 ;
  assign y19515 = ~n46253 ;
  assign y19516 = ~n46255 ;
  assign y19517 = ~1'b0 ;
  assign y19518 = ~n46257 ;
  assign y19519 = n46259 ;
  assign y19520 = ~1'b0 ;
  assign y19521 = ~n46264 ;
  assign y19522 = n46266 ;
  assign y19523 = n46272 ;
  assign y19524 = n46273 ;
  assign y19525 = ~n46276 ;
  assign y19526 = ~n46278 ;
  assign y19527 = ~n27832 ;
  assign y19528 = ~1'b0 ;
  assign y19529 = ~n46280 ;
  assign y19530 = n14690 ;
  assign y19531 = ~1'b0 ;
  assign y19532 = n39973 ;
  assign y19533 = n46281 ;
  assign y19534 = n46283 ;
  assign y19535 = n46284 ;
  assign y19536 = ~n46285 ;
  assign y19537 = ~1'b0 ;
  assign y19538 = ~1'b0 ;
  assign y19539 = ~n46292 ;
  assign y19540 = ~1'b0 ;
  assign y19541 = ~1'b0 ;
  assign y19542 = ~1'b0 ;
  assign y19543 = ~n46297 ;
  assign y19544 = n46299 ;
  assign y19545 = n46301 ;
  assign y19546 = n46307 ;
  assign y19547 = ~n46310 ;
  assign y19548 = ~n46312 ;
  assign y19549 = ~n46313 ;
  assign y19550 = ~n46316 ;
  assign y19551 = ~1'b0 ;
  assign y19552 = n46322 ;
  assign y19553 = ~n46323 ;
  assign y19554 = ~n46325 ;
  assign y19555 = n46327 ;
  assign y19556 = ~n46329 ;
  assign y19557 = n46331 ;
  assign y19558 = ~1'b0 ;
  assign y19559 = n46335 ;
  assign y19560 = n28021 ;
  assign y19561 = ~1'b0 ;
  assign y19562 = n46337 ;
  assign y19563 = n46338 ;
  assign y19564 = ~1'b0 ;
  assign y19565 = ~n46339 ;
  assign y19566 = n46340 ;
  assign y19567 = ~n46344 ;
  assign y19568 = ~n46349 ;
  assign y19569 = ~1'b0 ;
  assign y19570 = n46351 ;
  assign y19571 = ~1'b0 ;
  assign y19572 = ~n46356 ;
  assign y19573 = n46358 ;
  assign y19574 = ~1'b0 ;
  assign y19575 = ~1'b0 ;
  assign y19576 = n46362 ;
  assign y19577 = n46364 ;
  assign y19578 = n46365 ;
  assign y19579 = n17555 ;
  assign y19580 = ~n46368 ;
  assign y19581 = n46371 ;
  assign y19582 = n46374 ;
  assign y19583 = ~n46377 ;
  assign y19584 = ~n46379 ;
  assign y19585 = ~n46382 ;
  assign y19586 = ~n46383 ;
  assign y19587 = ~n46384 ;
  assign y19588 = n46387 ;
  assign y19589 = n46388 ;
  assign y19590 = ~n46390 ;
  assign y19591 = ~n46391 ;
  assign y19592 = ~1'b0 ;
  assign y19593 = n46393 ;
  assign y19594 = ~1'b0 ;
  assign y19595 = n46395 ;
  assign y19596 = ~n46402 ;
  assign y19597 = ~n46403 ;
  assign y19598 = ~n46404 ;
  assign y19599 = ~n46405 ;
  assign y19600 = ~1'b0 ;
  assign y19601 = ~1'b0 ;
  assign y19602 = ~n46406 ;
  assign y19603 = ~n19580 ;
  assign y19604 = ~n46408 ;
  assign y19605 = ~1'b0 ;
  assign y19606 = ~n46409 ;
  assign y19607 = ~n46410 ;
  assign y19608 = ~1'b0 ;
  assign y19609 = ~1'b0 ;
  assign y19610 = ~1'b0 ;
  assign y19611 = ~n46413 ;
  assign y19612 = ~n46418 ;
  assign y19613 = 1'b0 ;
  assign y19614 = ~n46420 ;
  assign y19615 = ~n46425 ;
  assign y19616 = ~n46426 ;
  assign y19617 = ~n46428 ;
  assign y19618 = n46429 ;
  assign y19619 = n46431 ;
  assign y19620 = n46434 ;
  assign y19621 = ~1'b0 ;
  assign y19622 = ~1'b0 ;
  assign y19623 = n46435 ;
  assign y19624 = n46439 ;
  assign y19625 = ~n46441 ;
  assign y19626 = ~n33347 ;
  assign y19627 = n46444 ;
  assign y19628 = ~n46453 ;
  assign y19629 = n46455 ;
  assign y19630 = ~1'b0 ;
  assign y19631 = ~n46459 ;
  assign y19632 = ~n46464 ;
  assign y19633 = ~1'b0 ;
  assign y19634 = ~n46465 ;
  assign y19635 = n46467 ;
  assign y19636 = n46468 ;
  assign y19637 = n46469 ;
  assign y19638 = n29585 ;
  assign y19639 = ~n46470 ;
  assign y19640 = n46473 ;
  assign y19641 = ~1'b0 ;
  assign y19642 = ~1'b0 ;
  assign y19643 = ~1'b0 ;
  assign y19644 = n46477 ;
  assign y19645 = ~n46479 ;
  assign y19646 = n46481 ;
  assign y19647 = n46482 ;
  assign y19648 = ~n46483 ;
  assign y19649 = ~n46484 ;
  assign y19650 = n46488 ;
  assign y19651 = ~n46490 ;
  assign y19652 = ~1'b0 ;
  assign y19653 = ~1'b0 ;
  assign y19654 = ~n46492 ;
  assign y19655 = 1'b0 ;
  assign y19656 = ~1'b0 ;
  assign y19657 = ~n46494 ;
  assign y19658 = ~n46496 ;
  assign y19659 = n46497 ;
  assign y19660 = ~n46498 ;
  assign y19661 = ~n46502 ;
  assign y19662 = n46504 ;
  assign y19663 = ~1'b0 ;
  assign y19664 = ~1'b0 ;
  assign y19665 = ~n46506 ;
  assign y19666 = ~1'b0 ;
  assign y19667 = ~1'b0 ;
  assign y19668 = ~n46508 ;
  assign y19669 = n46509 ;
  assign y19670 = ~n46510 ;
  assign y19671 = n46512 ;
  assign y19672 = ~n46514 ;
  assign y19673 = n46516 ;
  assign y19674 = ~1'b0 ;
  assign y19675 = ~1'b0 ;
  assign y19676 = n46519 ;
  assign y19677 = ~n46520 ;
  assign y19678 = n46521 ;
  assign y19679 = n46523 ;
  assign y19680 = ~n46524 ;
  assign y19681 = n46525 ;
  assign y19682 = n27843 ;
  assign y19683 = ~1'b0 ;
  assign y19684 = ~1'b0 ;
  assign y19685 = ~n46528 ;
  assign y19686 = ~n46529 ;
  assign y19687 = ~1'b0 ;
  assign y19688 = ~n46532 ;
  assign y19689 = n46533 ;
  assign y19690 = n46534 ;
  assign y19691 = n46535 ;
  assign y19692 = ~1'b0 ;
  assign y19693 = ~1'b0 ;
  assign y19694 = ~1'b0 ;
  assign y19695 = n46544 ;
  assign y19696 = ~n46545 ;
  assign y19697 = n46546 ;
  assign y19698 = ~n46548 ;
  assign y19699 = ~1'b0 ;
  assign y19700 = ~n46549 ;
  assign y19701 = ~n46550 ;
  assign y19702 = ~n46551 ;
  assign y19703 = ~n46554 ;
  assign y19704 = n46556 ;
  assign y19705 = n46566 ;
  assign y19706 = ~n46569 ;
  assign y19707 = ~n46571 ;
  assign y19708 = n46573 ;
  assign y19709 = n46574 ;
  assign y19710 = ~n46575 ;
  assign y19711 = ~n46578 ;
  assign y19712 = n46583 ;
  assign y19713 = ~n46584 ;
  assign y19714 = ~1'b0 ;
  assign y19715 = n46588 ;
  assign y19716 = ~1'b0 ;
  assign y19717 = n46589 ;
  assign y19718 = ~n46590 ;
  assign y19719 = ~n46591 ;
  assign y19720 = n46592 ;
  assign y19721 = ~n46593 ;
  assign y19722 = n46595 ;
  assign y19723 = ~n46602 ;
  assign y19724 = ~1'b0 ;
  assign y19725 = ~n46605 ;
  assign y19726 = ~n46607 ;
  assign y19727 = n46613 ;
  assign y19728 = ~n46619 ;
  assign y19729 = ~1'b0 ;
  assign y19730 = n46620 ;
  assign y19731 = n46621 ;
  assign y19732 = ~n46625 ;
  assign y19733 = ~n46627 ;
  assign y19734 = ~n46632 ;
  assign y19735 = n46634 ;
  assign y19736 = ~n46635 ;
  assign y19737 = n46639 ;
  assign y19738 = ~1'b0 ;
  assign y19739 = ~n46644 ;
  assign y19740 = n46645 ;
  assign y19741 = ~n46646 ;
  assign y19742 = ~n46651 ;
  assign y19743 = ~1'b0 ;
  assign y19744 = 1'b0 ;
  assign y19745 = ~n46655 ;
  assign y19746 = ~1'b0 ;
  assign y19747 = ~n46656 ;
  assign y19748 = ~n46661 ;
  assign y19749 = ~1'b0 ;
  assign y19750 = n46662 ;
  assign y19751 = n46665 ;
  assign y19752 = ~n46666 ;
  assign y19753 = ~n46667 ;
  assign y19754 = ~1'b0 ;
  assign y19755 = n46671 ;
  assign y19756 = ~n46672 ;
  assign y19757 = ~1'b0 ;
  assign y19758 = ~n46674 ;
  assign y19759 = n46679 ;
  assign y19760 = ~n46685 ;
  assign y19761 = n46686 ;
  assign y19762 = ~n46687 ;
  assign y19763 = n46688 ;
  assign y19764 = ~n46689 ;
  assign y19765 = ~1'b0 ;
  assign y19766 = ~1'b0 ;
  assign y19767 = n46691 ;
  assign y19768 = ~n46693 ;
  assign y19769 = ~n46695 ;
  assign y19770 = n46698 ;
  assign y19771 = n46702 ;
  assign y19772 = ~n46707 ;
  assign y19773 = n46708 ;
  assign y19774 = ~n46710 ;
  assign y19775 = ~n46713 ;
  assign y19776 = n46714 ;
  assign y19777 = ~1'b0 ;
  assign y19778 = ~n46715 ;
  assign y19779 = ~1'b0 ;
  assign y19780 = n46717 ;
  assign y19781 = n16466 ;
  assign y19782 = ~1'b0 ;
  assign y19783 = ~n46718 ;
  assign y19784 = ~n46719 ;
  assign y19785 = ~n46722 ;
  assign y19786 = ~n46723 ;
  assign y19787 = n46724 ;
  assign y19788 = ~1'b0 ;
  assign y19789 = ~n46726 ;
  assign y19790 = ~1'b0 ;
  assign y19791 = ~1'b0 ;
  assign y19792 = ~n46728 ;
  assign y19793 = n46729 ;
  assign y19794 = n46730 ;
  assign y19795 = n46733 ;
  assign y19796 = n46735 ;
  assign y19797 = n46737 ;
  assign y19798 = ~n46742 ;
  assign y19799 = ~1'b0 ;
  assign y19800 = ~n46743 ;
  assign y19801 = n46745 ;
  assign y19802 = ~n46749 ;
  assign y19803 = n46753 ;
  assign y19804 = n46754 ;
  assign y19805 = ~n46757 ;
  assign y19806 = n46761 ;
  assign y19807 = ~n46762 ;
  assign y19808 = ~1'b0 ;
  assign y19809 = ~n46768 ;
  assign y19810 = ~n46771 ;
  assign y19811 = n46772 ;
  assign y19812 = ~1'b0 ;
  assign y19813 = n46774 ;
  assign y19814 = ~1'b0 ;
  assign y19815 = ~n46783 ;
  assign y19816 = n46790 ;
  assign y19817 = ~1'b0 ;
  assign y19818 = ~n46791 ;
  assign y19819 = ~n46793 ;
  assign y19820 = ~n46794 ;
  assign y19821 = ~n46796 ;
  assign y19822 = ~n46798 ;
  assign y19823 = ~1'b0 ;
  assign y19824 = n46801 ;
  assign y19825 = ~1'b0 ;
  assign y19826 = ~n46804 ;
  assign y19827 = n46810 ;
  assign y19828 = ~n46812 ;
  assign y19829 = ~1'b0 ;
  assign y19830 = ~n46813 ;
  assign y19831 = n46814 ;
  assign y19832 = ~1'b0 ;
  assign y19833 = ~n46815 ;
  assign y19834 = ~n46817 ;
  assign y19835 = ~n46819 ;
  assign y19836 = n46823 ;
  assign y19837 = ~n46824 ;
  assign y19838 = ~n46825 ;
  assign y19839 = ~1'b0 ;
  assign y19840 = n46827 ;
  assign y19841 = n46828 ;
  assign y19842 = ~n46831 ;
  assign y19843 = ~n46834 ;
  assign y19844 = ~1'b0 ;
  assign y19845 = ~n46835 ;
  assign y19846 = ~n30859 ;
  assign y19847 = n46836 ;
  assign y19848 = n46838 ;
  assign y19849 = ~n46840 ;
  assign y19850 = 1'b0 ;
  assign y19851 = n38149 ;
  assign y19852 = n46841 ;
  assign y19853 = ~n46843 ;
  assign y19854 = ~n46845 ;
  assign y19855 = n46846 ;
  assign y19856 = ~n46847 ;
  assign y19857 = n46848 ;
  assign y19858 = ~n28788 ;
  assign y19859 = ~n46851 ;
  assign y19860 = ~n46853 ;
  assign y19861 = n46857 ;
  assign y19862 = ~1'b0 ;
  assign y19863 = ~n46860 ;
  assign y19864 = ~1'b0 ;
  assign y19865 = ~n46862 ;
  assign y19866 = n46865 ;
  assign y19867 = n46868 ;
  assign y19868 = ~n46869 ;
  assign y19869 = ~n22879 ;
  assign y19870 = ~1'b0 ;
  assign y19871 = ~n46872 ;
  assign y19872 = ~n27142 ;
  assign y19873 = n46876 ;
  assign y19874 = n46878 ;
  assign y19875 = n46880 ;
  assign y19876 = n46881 ;
  assign y19877 = n46882 ;
  assign y19878 = ~1'b0 ;
  assign y19879 = n46883 ;
  assign y19880 = n46884 ;
  assign y19881 = ~n46889 ;
  assign y19882 = ~n6891 ;
  assign y19883 = ~1'b0 ;
  assign y19884 = n46892 ;
  assign y19885 = n46897 ;
  assign y19886 = ~1'b0 ;
  assign y19887 = n46898 ;
  assign y19888 = n46900 ;
  assign y19889 = n46901 ;
  assign y19890 = ~n46908 ;
  assign y19891 = ~n46910 ;
  assign y19892 = n46911 ;
  assign y19893 = ~n46912 ;
  assign y19894 = ~n46916 ;
  assign y19895 = n46920 ;
  assign y19896 = ~n46929 ;
  assign y19897 = n46932 ;
  assign y19898 = n46936 ;
  assign y19899 = ~n46937 ;
  assign y19900 = n43698 ;
  assign y19901 = n46939 ;
  assign y19902 = n46941 ;
  assign y19903 = ~1'b0 ;
  assign y19904 = ~1'b0 ;
  assign y19905 = ~n46942 ;
  assign y19906 = ~n46944 ;
  assign y19907 = ~n16656 ;
  assign y19908 = n46946 ;
  assign y19909 = n46948 ;
  assign y19910 = ~n46950 ;
  assign y19911 = n46952 ;
  assign y19912 = ~1'b0 ;
  assign y19913 = ~1'b0 ;
  assign y19914 = ~n46954 ;
  assign y19915 = ~n46958 ;
  assign y19916 = n46961 ;
  assign y19917 = n46962 ;
  assign y19918 = ~n46968 ;
  assign y19919 = n46969 ;
  assign y19920 = n46971 ;
  assign y19921 = ~n46980 ;
  assign y19922 = n46982 ;
  assign y19923 = ~n46986 ;
  assign y19924 = n46989 ;
  assign y19925 = ~n46992 ;
  assign y19926 = ~n46995 ;
  assign y19927 = n46997 ;
  assign y19928 = ~n47000 ;
  assign y19929 = ~n47002 ;
  assign y19930 = ~1'b0 ;
  assign y19931 = ~1'b0 ;
  assign y19932 = n47004 ;
  assign y19933 = ~n47005 ;
  assign y19934 = ~n47006 ;
  assign y19935 = ~n47009 ;
  assign y19936 = ~n47012 ;
  assign y19937 = 1'b0 ;
  assign y19938 = ~1'b0 ;
  assign y19939 = 1'b0 ;
  assign y19940 = ~1'b0 ;
  assign y19941 = n47015 ;
  assign y19942 = ~n47019 ;
  assign y19943 = ~n47020 ;
  assign y19944 = n47023 ;
  assign y19945 = ~1'b0 ;
  assign y19946 = n47024 ;
  assign y19947 = ~n47026 ;
  assign y19948 = n47028 ;
  assign y19949 = ~n47030 ;
  assign y19950 = ~1'b0 ;
  assign y19951 = ~n47031 ;
  assign y19952 = ~n7910 ;
  assign y19953 = n47036 ;
  assign y19954 = ~1'b0 ;
  assign y19955 = n47037 ;
  assign y19956 = ~1'b0 ;
  assign y19957 = ~1'b0 ;
  assign y19958 = ~1'b0 ;
  assign y19959 = n47038 ;
  assign y19960 = n47041 ;
  assign y19961 = ~n47042 ;
  assign y19962 = ~n47045 ;
  assign y19963 = ~n47046 ;
  assign y19964 = 1'b0 ;
  assign y19965 = n44927 ;
  assign y19966 = n47048 ;
  assign y19967 = ~1'b0 ;
  assign y19968 = ~n24780 ;
  assign y19969 = ~n47051 ;
  assign y19970 = ~n47053 ;
  assign y19971 = ~n47056 ;
  assign y19972 = ~n47059 ;
  assign y19973 = n47063 ;
  assign y19974 = 1'b0 ;
  assign y19975 = n47064 ;
  assign y19976 = ~n47066 ;
  assign y19977 = ~1'b0 ;
  assign y19978 = ~1'b0 ;
  assign y19979 = ~n47067 ;
  assign y19980 = n47068 ;
  assign y19981 = ~n47070 ;
  assign y19982 = ~n47071 ;
  assign y19983 = ~n47072 ;
  assign y19984 = n47076 ;
  assign y19985 = n47077 ;
  assign y19986 = ~n47084 ;
  assign y19987 = ~1'b0 ;
  assign y19988 = ~n47086 ;
  assign y19989 = n47090 ;
  assign y19990 = n47095 ;
  assign y19991 = ~1'b0 ;
  assign y19992 = n47096 ;
  assign y19993 = ~n47097 ;
  assign y19994 = n47098 ;
  assign y19995 = ~n47099 ;
  assign y19996 = ~n47101 ;
  assign y19997 = ~n14634 ;
  assign y19998 = n47104 ;
  assign y19999 = ~1'b0 ;
  assign y20000 = n47106 ;
  assign y20001 = ~1'b0 ;
  assign y20002 = n47109 ;
  assign y20003 = n47110 ;
  assign y20004 = n47111 ;
  assign y20005 = n47112 ;
  assign y20006 = ~1'b0 ;
  assign y20007 = ~n47117 ;
  assign y20008 = ~n47118 ;
  assign y20009 = ~n47120 ;
  assign y20010 = ~1'b0 ;
  assign y20011 = ~1'b0 ;
  assign y20012 = ~n47125 ;
  assign y20013 = ~n47127 ;
  assign y20014 = ~n47128 ;
  assign y20015 = ~n47129 ;
  assign y20016 = ~n47131 ;
  assign y20017 = ~n47133 ;
  assign y20018 = ~n47135 ;
  assign y20019 = ~1'b0 ;
  assign y20020 = ~1'b0 ;
  assign y20021 = ~n47136 ;
  assign y20022 = n47137 ;
  assign y20023 = ~n47140 ;
  assign y20024 = n47141 ;
  assign y20025 = n4454 ;
  assign y20026 = ~n47142 ;
  assign y20027 = ~n47143 ;
  assign y20028 = ~n47144 ;
  assign y20029 = ~n47149 ;
  assign y20030 = n3763 ;
  assign y20031 = n47153 ;
  assign y20032 = ~1'b0 ;
  assign y20033 = n47156 ;
  assign y20034 = n47157 ;
  assign y20035 = n47161 ;
  assign y20036 = n47162 ;
  assign y20037 = n47163 ;
  assign y20038 = n47167 ;
  assign y20039 = ~n47168 ;
  assign y20040 = ~n13268 ;
  assign y20041 = ~1'b0 ;
  assign y20042 = ~1'b0 ;
  assign y20043 = ~1'b0 ;
  assign y20044 = n47174 ;
  assign y20045 = ~n47175 ;
  assign y20046 = ~n47176 ;
  assign y20047 = n47177 ;
  assign y20048 = ~n47181 ;
  assign y20049 = ~1'b0 ;
  assign y20050 = ~1'b0 ;
  assign y20051 = ~n47184 ;
  assign y20052 = n47186 ;
  assign y20053 = ~n47189 ;
  assign y20054 = n47194 ;
  assign y20055 = ~1'b0 ;
  assign y20056 = ~n47199 ;
  assign y20057 = n47200 ;
  assign y20058 = ~n47203 ;
  assign y20059 = n47204 ;
  assign y20060 = n23213 ;
  assign y20061 = ~1'b0 ;
  assign y20062 = ~1'b0 ;
  assign y20063 = ~1'b0 ;
  assign y20064 = ~n47206 ;
  assign y20065 = n47209 ;
  assign y20066 = ~n47215 ;
  assign y20067 = ~n47219 ;
  assign y20068 = n47220 ;
  assign y20069 = n47221 ;
  assign y20070 = n47222 ;
  assign y20071 = ~n47224 ;
  assign y20072 = ~n47226 ;
  assign y20073 = ~n47228 ;
  assign y20074 = ~1'b0 ;
  assign y20075 = ~n47230 ;
  assign y20076 = ~n47231 ;
  assign y20077 = ~1'b0 ;
  assign y20078 = n47233 ;
  assign y20079 = ~n47236 ;
  assign y20080 = ~n47241 ;
  assign y20081 = ~1'b0 ;
  assign y20082 = n47243 ;
  assign y20083 = ~1'b0 ;
  assign y20084 = n47244 ;
  assign y20085 = ~n47248 ;
  assign y20086 = n661 ;
  assign y20087 = ~n47252 ;
  assign y20088 = n32776 ;
  assign y20089 = ~n47257 ;
  assign y20090 = ~n47258 ;
  assign y20091 = n47262 ;
  assign y20092 = n47264 ;
  assign y20093 = ~1'b0 ;
  assign y20094 = n47265 ;
  assign y20095 = n47269 ;
  assign y20096 = ~n25448 ;
  assign y20097 = n47271 ;
  assign y20098 = n47273 ;
  assign y20099 = n47274 ;
  assign y20100 = n47276 ;
  assign y20101 = ~n47278 ;
  assign y20102 = ~1'b0 ;
  assign y20103 = ~1'b0 ;
  assign y20104 = ~n47280 ;
  assign y20105 = ~n47283 ;
  assign y20106 = ~n47285 ;
  assign y20107 = ~n47286 ;
  assign y20108 = ~n47287 ;
  assign y20109 = n47292 ;
  assign y20110 = n47295 ;
  assign y20111 = ~1'b0 ;
  assign y20112 = ~n47296 ;
  assign y20113 = n47297 ;
  assign y20114 = ~1'b0 ;
  assign y20115 = ~n47299 ;
  assign y20116 = ~1'b0 ;
  assign y20117 = n47309 ;
  assign y20118 = n47310 ;
  assign y20119 = ~n47311 ;
  assign y20120 = ~n47312 ;
  assign y20121 = n47313 ;
  assign y20122 = ~n47314 ;
  assign y20123 = n47316 ;
  assign y20124 = n47317 ;
  assign y20125 = ~n47319 ;
  assign y20126 = ~1'b0 ;
  assign y20127 = n47328 ;
  assign y20128 = n47330 ;
  assign y20129 = ~n47333 ;
  assign y20130 = ~n47334 ;
  assign y20131 = ~1'b0 ;
  assign y20132 = ~1'b0 ;
  assign y20133 = ~1'b0 ;
  assign y20134 = n47335 ;
  assign y20135 = ~n47338 ;
  assign y20136 = ~n47341 ;
  assign y20137 = ~n47345 ;
  assign y20138 = ~n47347 ;
  assign y20139 = n47353 ;
  assign y20140 = n47356 ;
  assign y20141 = n47357 ;
  assign y20142 = n47363 ;
  assign y20143 = n47365 ;
  assign y20144 = ~1'b0 ;
  assign y20145 = n47367 ;
  assign y20146 = ~1'b0 ;
  assign y20147 = n47368 ;
  assign y20148 = ~n47369 ;
  assign y20149 = ~n47370 ;
  assign y20150 = n47374 ;
  assign y20151 = ~n47376 ;
  assign y20152 = ~n47377 ;
  assign y20153 = ~1'b0 ;
  assign y20154 = ~1'b0 ;
  assign y20155 = n47380 ;
  assign y20156 = n47384 ;
  assign y20157 = n47385 ;
  assign y20158 = n47386 ;
  assign y20159 = ~n47391 ;
  assign y20160 = n47395 ;
  assign y20161 = ~1'b0 ;
  assign y20162 = ~1'b0 ;
  assign y20163 = ~n47398 ;
  assign y20164 = ~n47399 ;
  assign y20165 = ~n47402 ;
  assign y20166 = n47404 ;
  assign y20167 = ~n47406 ;
  assign y20168 = ~n47414 ;
  assign y20169 = ~1'b0 ;
  assign y20170 = n47418 ;
  assign y20171 = ~1'b0 ;
  assign y20172 = ~n47420 ;
  assign y20173 = n47421 ;
  assign y20174 = n47422 ;
  assign y20175 = ~n47423 ;
  assign y20176 = ~n47425 ;
  assign y20177 = ~n47426 ;
  assign y20178 = ~n47427 ;
  assign y20179 = ~n47430 ;
  assign y20180 = ~1'b0 ;
  assign y20181 = ~n47432 ;
  assign y20182 = n47435 ;
  assign y20183 = ~n47438 ;
  assign y20184 = ~n16559 ;
  assign y20185 = n47441 ;
  assign y20186 = n47443 ;
  assign y20187 = ~n47445 ;
  assign y20188 = ~1'b0 ;
  assign y20189 = ~n47447 ;
  assign y20190 = ~1'b0 ;
  assign y20191 = ~n47449 ;
  assign y20192 = ~n47451 ;
  assign y20193 = ~1'b0 ;
  assign y20194 = ~n47452 ;
  assign y20195 = n47457 ;
  assign y20196 = ~n47459 ;
  assign y20197 = ~n47462 ;
  assign y20198 = n11548 ;
  assign y20199 = ~1'b0 ;
  assign y20200 = ~n47466 ;
  assign y20201 = ~n47478 ;
  assign y20202 = n47479 ;
  assign y20203 = ~1'b0 ;
  assign y20204 = ~n47481 ;
  assign y20205 = ~n47484 ;
  assign y20206 = ~n47485 ;
  assign y20207 = ~n47487 ;
  assign y20208 = ~1'b0 ;
  assign y20209 = n47488 ;
  assign y20210 = ~1'b0 ;
  assign y20211 = ~n7745 ;
  assign y20212 = ~n47490 ;
  assign y20213 = ~n47493 ;
  assign y20214 = ~1'b0 ;
  assign y20215 = n47494 ;
  assign y20216 = n47495 ;
  assign y20217 = ~n47496 ;
  assign y20218 = ~1'b0 ;
  assign y20219 = ~1'b0 ;
  assign y20220 = n38948 ;
  assign y20221 = n47498 ;
  assign y20222 = ~n47500 ;
  assign y20223 = ~n47501 ;
  assign y20224 = ~n47502 ;
  assign y20225 = ~n47503 ;
  assign y20226 = n47505 ;
  assign y20227 = n47509 ;
  assign y20228 = ~n47511 ;
  assign y20229 = 1'b0 ;
  assign y20230 = ~1'b0 ;
  assign y20231 = n44613 ;
  assign y20232 = ~n47512 ;
  assign y20233 = n47513 ;
  assign y20234 = ~n47515 ;
  assign y20235 = ~n47517 ;
  assign y20236 = n47520 ;
  assign y20237 = ~n47521 ;
  assign y20238 = n47522 ;
  assign y20239 = n47525 ;
  assign y20240 = n28528 ;
  assign y20241 = ~1'b0 ;
  assign y20242 = ~1'b0 ;
  assign y20243 = n47531 ;
  assign y20244 = ~n47533 ;
  assign y20245 = ~n47538 ;
  assign y20246 = n47539 ;
  assign y20247 = ~n47541 ;
  assign y20248 = n47542 ;
  assign y20249 = n27034 ;
  assign y20250 = ~n47543 ;
  assign y20251 = n47544 ;
  assign y20252 = ~n47550 ;
  assign y20253 = ~1'b0 ;
  assign y20254 = n47553 ;
  assign y20255 = ~1'b0 ;
  assign y20256 = n47556 ;
  assign y20257 = ~n47557 ;
  assign y20258 = ~n47560 ;
  assign y20259 = ~n33500 ;
  assign y20260 = n47566 ;
  assign y20261 = n47567 ;
  assign y20262 = ~1'b0 ;
  assign y20263 = ~1'b0 ;
  assign y20264 = ~n47569 ;
  assign y20265 = n47570 ;
  assign y20266 = ~1'b0 ;
  assign y20267 = n47573 ;
  assign y20268 = n47576 ;
  assign y20269 = n47577 ;
  assign y20270 = n47581 ;
  assign y20271 = ~n47582 ;
  assign y20272 = ~n47585 ;
  assign y20273 = ~1'b0 ;
  assign y20274 = ~n47587 ;
  assign y20275 = ~n47592 ;
  assign y20276 = n47593 ;
  assign y20277 = n47595 ;
  assign y20278 = n47596 ;
  assign y20279 = ~n47598 ;
  assign y20280 = ~n47599 ;
  assign y20281 = ~n47600 ;
  assign y20282 = ~n47603 ;
  assign y20283 = ~1'b0 ;
  assign y20284 = ~n47604 ;
  assign y20285 = ~n47606 ;
  assign y20286 = ~1'b0 ;
  assign y20287 = n47607 ;
  assign y20288 = n47610 ;
  assign y20289 = ~n47613 ;
  assign y20290 = ~n47614 ;
  assign y20291 = ~n47619 ;
  assign y20292 = ~n47626 ;
  assign y20293 = ~n47635 ;
  assign y20294 = ~1'b0 ;
  assign y20295 = ~1'b0 ;
  assign y20296 = ~n47636 ;
  assign y20297 = ~n47640 ;
  assign y20298 = n47643 ;
  assign y20299 = n47644 ;
  assign y20300 = ~1'b0 ;
  assign y20301 = ~n47645 ;
  assign y20302 = ~n47647 ;
  assign y20303 = n10424 ;
  assign y20304 = n47648 ;
  assign y20305 = n47649 ;
  assign y20306 = ~n47651 ;
  assign y20307 = n47654 ;
  assign y20308 = ~1'b0 ;
  assign y20309 = n47657 ;
  assign y20310 = n47658 ;
  assign y20311 = n47662 ;
  assign y20312 = ~1'b0 ;
  assign y20313 = ~n47664 ;
  assign y20314 = ~n47671 ;
  assign y20315 = n47673 ;
  assign y20316 = n47674 ;
  assign y20317 = ~n47676 ;
  assign y20318 = ~1'b0 ;
  assign y20319 = ~1'b0 ;
  assign y20320 = ~1'b0 ;
  assign y20321 = n47678 ;
  assign y20322 = ~n1048 ;
  assign y20323 = ~n47680 ;
  assign y20324 = n47681 ;
  assign y20325 = n47689 ;
  assign y20326 = n47693 ;
  assign y20327 = ~n47695 ;
  assign y20328 = n47696 ;
  assign y20329 = ~n47697 ;
  assign y20330 = n47700 ;
  assign y20331 = n47701 ;
  assign y20332 = ~n47703 ;
  assign y20333 = ~n47704 ;
  assign y20334 = n47705 ;
  assign y20335 = n47707 ;
  assign y20336 = ~n28270 ;
  assign y20337 = n47708 ;
  assign y20338 = ~1'b0 ;
  assign y20339 = n47711 ;
  assign y20340 = n47715 ;
  assign y20341 = n47716 ;
  assign y20342 = ~n47717 ;
  assign y20343 = n47733 ;
  assign y20344 = ~n47736 ;
  assign y20345 = n47738 ;
  assign y20346 = n47740 ;
  assign y20347 = ~n47742 ;
  assign y20348 = n47744 ;
  assign y20349 = ~1'b0 ;
  assign y20350 = ~1'b0 ;
  assign y20351 = ~n47746 ;
  assign y20352 = n47748 ;
  assign y20353 = n47749 ;
  assign y20354 = ~n47750 ;
  assign y20355 = n47753 ;
  assign y20356 = n47757 ;
  assign y20357 = n47760 ;
  assign y20358 = n47764 ;
  assign y20359 = ~n1341 ;
  assign y20360 = ~n47765 ;
  assign y20361 = ~1'b0 ;
  assign y20362 = ~1'b0 ;
  assign y20363 = n47767 ;
  assign y20364 = ~n47769 ;
  assign y20365 = ~n47770 ;
  assign y20366 = ~n47771 ;
  assign y20367 = ~n47772 ;
  assign y20368 = n47781 ;
  assign y20369 = n47782 ;
  assign y20370 = n47784 ;
  assign y20371 = ~1'b0 ;
  assign y20372 = n47786 ;
  assign y20373 = ~n47789 ;
  assign y20374 = ~n47791 ;
  assign y20375 = 1'b0 ;
  assign y20376 = ~1'b0 ;
  assign y20377 = ~n47792 ;
  assign y20378 = n47793 ;
  assign y20379 = n47794 ;
  assign y20380 = ~n47796 ;
  assign y20381 = n47798 ;
  assign y20382 = n47801 ;
  assign y20383 = n47803 ;
  assign y20384 = ~n47807 ;
  assign y20385 = ~1'b0 ;
  assign y20386 = n47809 ;
  assign y20387 = n47811 ;
  assign y20388 = n47812 ;
  assign y20389 = ~n47816 ;
  assign y20390 = ~n47819 ;
  assign y20391 = ~n47825 ;
  assign y20392 = n47828 ;
  assign y20393 = ~1'b0 ;
  assign y20394 = ~1'b0 ;
  assign y20395 = n47829 ;
  assign y20396 = ~n47830 ;
  assign y20397 = n47833 ;
  assign y20398 = ~n47837 ;
  assign y20399 = n47842 ;
  assign y20400 = n47849 ;
  assign y20401 = ~n47850 ;
  assign y20402 = ~n47857 ;
  assign y20403 = ~n47859 ;
  assign y20404 = n47862 ;
  assign y20405 = ~n47867 ;
  assign y20406 = 1'b0 ;
  assign y20407 = ~n47870 ;
  assign y20408 = ~n47871 ;
  assign y20409 = ~n47873 ;
  assign y20410 = n47874 ;
  assign y20411 = ~n47877 ;
  assign y20412 = n47880 ;
  assign y20413 = ~n47881 ;
  assign y20414 = ~n47883 ;
  assign y20415 = ~1'b0 ;
  assign y20416 = ~1'b0 ;
  assign y20417 = n47884 ;
  assign y20418 = n47885 ;
  assign y20419 = n47886 ;
  assign y20420 = 1'b0 ;
  assign y20421 = ~n47891 ;
  assign y20422 = ~n47893 ;
  assign y20423 = ~n47896 ;
  assign y20424 = n47898 ;
  assign y20425 = n47907 ;
  assign y20426 = n47909 ;
  assign y20427 = n47910 ;
  assign y20428 = n47912 ;
  assign y20429 = ~n47914 ;
  assign y20430 = ~n47915 ;
  assign y20431 = n47916 ;
  assign y20432 = n47918 ;
  assign y20433 = ~1'b0 ;
  assign y20434 = ~n47919 ;
  assign y20435 = ~1'b0 ;
  assign y20436 = ~n47922 ;
  assign y20437 = ~n47924 ;
  assign y20438 = ~n47926 ;
  assign y20439 = n22778 ;
  assign y20440 = ~n47931 ;
  assign y20441 = ~n47935 ;
  assign y20442 = ~n47936 ;
  assign y20443 = ~n47939 ;
  assign y20444 = ~1'b0 ;
  assign y20445 = ~n47942 ;
  assign y20446 = ~n47944 ;
  assign y20447 = n47946 ;
  assign y20448 = ~n47948 ;
  assign y20449 = ~1'b0 ;
  assign y20450 = ~n47950 ;
  assign y20451 = n1433 ;
  assign y20452 = n47951 ;
  assign y20453 = ~n47952 ;
  assign y20454 = ~1'b0 ;
  assign y20455 = ~1'b0 ;
  assign y20456 = ~1'b0 ;
  assign y20457 = ~n47954 ;
  assign y20458 = ~1'b0 ;
  assign y20459 = ~n47957 ;
  assign y20460 = n47958 ;
  assign y20461 = ~n47964 ;
  assign y20462 = ~1'b0 ;
  assign y20463 = n47966 ;
  assign y20464 = n47969 ;
  assign y20465 = n47971 ;
  assign y20466 = n32334 ;
  assign y20467 = n47975 ;
  assign y20468 = ~1'b0 ;
  assign y20469 = ~1'b0 ;
  assign y20470 = ~n47977 ;
  assign y20471 = ~1'b0 ;
  assign y20472 = n47979 ;
  assign y20473 = n47985 ;
  assign y20474 = n47986 ;
  assign y20475 = ~n47987 ;
  assign y20476 = ~1'b0 ;
  assign y20477 = ~1'b0 ;
  assign y20478 = n47989 ;
  assign y20479 = ~1'b0 ;
  assign y20480 = 1'b0 ;
  assign y20481 = ~1'b0 ;
  assign y20482 = ~n47990 ;
  assign y20483 = n47991 ;
  assign y20484 = n47994 ;
  assign y20485 = ~n47997 ;
  assign y20486 = n47998 ;
  assign y20487 = n48004 ;
  assign y20488 = ~1'b0 ;
  assign y20489 = ~n48006 ;
  assign y20490 = ~n48007 ;
  assign y20491 = ~1'b0 ;
  assign y20492 = n48009 ;
  assign y20493 = n48010 ;
  assign y20494 = ~n48012 ;
  assign y20495 = ~n48013 ;
  assign y20496 = 1'b0 ;
  assign y20497 = ~n48015 ;
  assign y20498 = ~1'b0 ;
  assign y20499 = ~n48017 ;
  assign y20500 = n48018 ;
  assign y20501 = ~1'b0 ;
  assign y20502 = ~n48023 ;
  assign y20503 = n48025 ;
  assign y20504 = ~n48033 ;
  assign y20505 = ~n48035 ;
  assign y20506 = ~n48037 ;
  assign y20507 = n48039 ;
  assign y20508 = ~n48040 ;
  assign y20509 = ~n48041 ;
  assign y20510 = ~n48051 ;
  assign y20511 = n48056 ;
  assign y20512 = n48059 ;
  assign y20513 = n48062 ;
  assign y20514 = ~1'b0 ;
  assign y20515 = ~n48065 ;
  assign y20516 = n48068 ;
  assign y20517 = n48069 ;
  assign y20518 = ~n48070 ;
  assign y20519 = n48073 ;
  assign y20520 = ~1'b0 ;
  assign y20521 = n48078 ;
  assign y20522 = n48080 ;
  assign y20523 = ~n48082 ;
  assign y20524 = ~n48083 ;
  assign y20525 = ~n48085 ;
  assign y20526 = n48088 ;
  assign y20527 = ~n48089 ;
  assign y20528 = ~n48090 ;
  assign y20529 = n48094 ;
  assign y20530 = n48095 ;
  assign y20531 = n48098 ;
  assign y20532 = ~1'b0 ;
  assign y20533 = ~n24721 ;
  assign y20534 = n48102 ;
  assign y20535 = ~1'b0 ;
  assign y20536 = n48103 ;
  assign y20537 = ~n48109 ;
  assign y20538 = ~n48113 ;
  assign y20539 = n48115 ;
  assign y20540 = ~1'b0 ;
  assign y20541 = ~n48116 ;
  assign y20542 = ~1'b0 ;
  assign y20543 = ~1'b0 ;
  assign y20544 = n48119 ;
  assign y20545 = ~n48121 ;
  assign y20546 = n48126 ;
  assign y20547 = ~n48132 ;
  assign y20548 = n48133 ;
  assign y20549 = ~n48141 ;
  assign y20550 = n48143 ;
  assign y20551 = n48144 ;
  assign y20552 = n48147 ;
  assign y20553 = n48148 ;
  assign y20554 = n48149 ;
  assign y20555 = n48152 ;
  assign y20556 = ~n48155 ;
  assign y20557 = ~n48157 ;
  assign y20558 = ~n48158 ;
  assign y20559 = ~1'b0 ;
  assign y20560 = ~1'b0 ;
  assign y20561 = ~n48160 ;
  assign y20562 = ~n48161 ;
  assign y20563 = n48164 ;
  assign y20564 = ~1'b0 ;
  assign y20565 = ~n48166 ;
  assign y20566 = ~n48167 ;
  assign y20567 = n48168 ;
  assign y20568 = n48169 ;
  assign y20569 = ~n48170 ;
  assign y20570 = ~n48172 ;
  assign y20571 = n48174 ;
  assign y20572 = ~1'b0 ;
  assign y20573 = n48176 ;
  assign y20574 = ~n48181 ;
  assign y20575 = ~1'b0 ;
  assign y20576 = ~1'b0 ;
  assign y20577 = ~n33566 ;
  assign y20578 = ~n48182 ;
  assign y20579 = n48184 ;
  assign y20580 = n48185 ;
  assign y20581 = ~n3014 ;
  assign y20582 = n48187 ;
  assign y20583 = n48188 ;
  assign y20584 = ~1'b0 ;
  assign y20585 = ~1'b0 ;
  assign y20586 = ~1'b0 ;
  assign y20587 = ~1'b0 ;
  assign y20588 = n48189 ;
  assign y20589 = n8107 ;
  assign y20590 = n48192 ;
  assign y20591 = ~1'b0 ;
  assign y20592 = ~1'b0 ;
  assign y20593 = ~n48195 ;
  assign y20594 = n48198 ;
  assign y20595 = ~n48199 ;
  assign y20596 = ~n48201 ;
  assign y20597 = ~n48204 ;
  assign y20598 = ~n48207 ;
  assign y20599 = ~n48208 ;
  assign y20600 = n48209 ;
  assign y20601 = n48211 ;
  assign y20602 = ~n48215 ;
  assign y20603 = ~1'b0 ;
  assign y20604 = n48217 ;
  assign y20605 = ~n4686 ;
  assign y20606 = 1'b0 ;
  assign y20607 = ~n48219 ;
  assign y20608 = ~n24259 ;
  assign y20609 = ~n48221 ;
  assign y20610 = ~1'b0 ;
  assign y20611 = n48222 ;
  assign y20612 = ~1'b0 ;
  assign y20613 = ~1'b0 ;
  assign y20614 = n48223 ;
  assign y20615 = ~n48225 ;
  assign y20616 = n48226 ;
  assign y20617 = ~n48227 ;
  assign y20618 = ~n829 ;
  assign y20619 = n48228 ;
  assign y20620 = n48229 ;
  assign y20621 = n48230 ;
  assign y20622 = ~1'b0 ;
  assign y20623 = ~1'b0 ;
  assign y20624 = n48231 ;
  assign y20625 = ~n48232 ;
  assign y20626 = ~n48233 ;
  assign y20627 = n48234 ;
  assign y20628 = n48235 ;
  assign y20629 = n48236 ;
  assign y20630 = n48239 ;
  assign y20631 = ~1'b0 ;
  assign y20632 = ~1'b0 ;
  assign y20633 = n48240 ;
  assign y20634 = n48241 ;
  assign y20635 = ~n48245 ;
  assign y20636 = n48247 ;
  assign y20637 = n28534 ;
  assign y20638 = ~n48249 ;
  assign y20639 = ~n48252 ;
  assign y20640 = n48253 ;
  assign y20641 = n48254 ;
  assign y20642 = ~1'b0 ;
  assign y20643 = ~1'b0 ;
  assign y20644 = n48263 ;
  assign y20645 = ~n48264 ;
  assign y20646 = ~n48268 ;
  assign y20647 = ~n48270 ;
  assign y20648 = ~n48273 ;
  assign y20649 = ~n48276 ;
  assign y20650 = n48278 ;
  assign y20651 = n48279 ;
  assign y20652 = n48280 ;
  assign y20653 = ~n48281 ;
  assign y20654 = ~1'b0 ;
  assign y20655 = ~n48283 ;
  assign y20656 = ~n48285 ;
  assign y20657 = ~1'b0 ;
  assign y20658 = ~n48287 ;
  assign y20659 = ~1'b0 ;
  assign y20660 = n48288 ;
  assign y20661 = n48290 ;
  assign y20662 = n48292 ;
  assign y20663 = n48294 ;
  assign y20664 = n48296 ;
  assign y20665 = n48298 ;
  assign y20666 = ~1'b0 ;
  assign y20667 = ~1'b0 ;
  assign y20668 = ~n48299 ;
  assign y20669 = ~n48303 ;
  assign y20670 = n48305 ;
  assign y20671 = n48307 ;
  assign y20672 = n48308 ;
  assign y20673 = ~1'b0 ;
  assign y20674 = n48312 ;
  assign y20675 = n48315 ;
  assign y20676 = ~n6944 ;
  assign y20677 = ~n48316 ;
  assign y20678 = 1'b0 ;
  assign y20679 = ~n48317 ;
  assign y20680 = n48319 ;
  assign y20681 = ~n48324 ;
  assign y20682 = n48327 ;
  assign y20683 = n48328 ;
  assign y20684 = ~n48330 ;
  assign y20685 = ~n48333 ;
  assign y20686 = n48334 ;
  assign y20687 = ~n48335 ;
  assign y20688 = ~1'b0 ;
  assign y20689 = n1261 ;
  assign y20690 = ~n48337 ;
  assign y20691 = ~n48341 ;
  assign y20692 = n48343 ;
  assign y20693 = n48347 ;
  assign y20694 = n48348 ;
  assign y20695 = n48349 ;
  assign y20696 = ~n48350 ;
  assign y20697 = ~n48351 ;
  assign y20698 = n48353 ;
  assign y20699 = ~n48354 ;
  assign y20700 = ~1'b0 ;
  assign y20701 = n48356 ;
  assign y20702 = n3790 ;
  assign y20703 = ~n5446 ;
  assign y20704 = ~n48358 ;
  assign y20705 = ~n48360 ;
  assign y20706 = ~1'b0 ;
  assign y20707 = ~n48364 ;
  assign y20708 = ~n48366 ;
  assign y20709 = ~1'b0 ;
  assign y20710 = ~n48370 ;
  assign y20711 = ~n48371 ;
  assign y20712 = ~n48374 ;
  assign y20713 = n48375 ;
  assign y20714 = n48377 ;
  assign y20715 = n48384 ;
  assign y20716 = ~n48388 ;
  assign y20717 = ~n48389 ;
  assign y20718 = n48391 ;
  assign y20719 = ~1'b0 ;
  assign y20720 = ~n48397 ;
  assign y20721 = n48398 ;
  assign y20722 = ~n35733 ;
  assign y20723 = n48400 ;
  assign y20724 = ~n48403 ;
  assign y20725 = ~1'b0 ;
  assign y20726 = n48404 ;
  assign y20727 = n48405 ;
  assign y20728 = n48406 ;
  assign y20729 = n48412 ;
  assign y20730 = n48415 ;
  assign y20731 = n48417 ;
  assign y20732 = ~1'b0 ;
  assign y20733 = ~n48421 ;
  assign y20734 = n48423 ;
  assign y20735 = ~n48424 ;
  assign y20736 = ~n48426 ;
  assign y20737 = n48427 ;
  assign y20738 = n48428 ;
  assign y20739 = n48433 ;
  assign y20740 = 1'b0 ;
  assign y20741 = ~1'b0 ;
  assign y20742 = ~1'b0 ;
  assign y20743 = n48436 ;
  assign y20744 = n48440 ;
  assign y20745 = ~1'b0 ;
  assign y20746 = n48443 ;
  assign y20747 = ~1'b0 ;
  assign y20748 = ~n48444 ;
  assign y20749 = n48446 ;
  assign y20750 = n48455 ;
  assign y20751 = n48458 ;
  assign y20752 = ~1'b0 ;
  assign y20753 = ~n48461 ;
  assign y20754 = ~n48463 ;
  assign y20755 = ~1'b0 ;
  assign y20756 = ~1'b0 ;
  assign y20757 = n48464 ;
  assign y20758 = n48465 ;
  assign y20759 = ~n48466 ;
  assign y20760 = ~n48467 ;
  assign y20761 = n48468 ;
  assign y20762 = n48469 ;
  assign y20763 = ~n48470 ;
  assign y20764 = ~1'b0 ;
  assign y20765 = ~n48473 ;
  assign y20766 = ~1'b0 ;
  assign y20767 = ~n48477 ;
  assign y20768 = ~n48480 ;
  assign y20769 = n48481 ;
  assign y20770 = n48482 ;
  assign y20771 = n48485 ;
  assign y20772 = ~n48486 ;
  assign y20773 = n48489 ;
  assign y20774 = n48491 ;
  assign y20775 = ~1'b0 ;
  assign y20776 = ~n48493 ;
  assign y20777 = n48494 ;
  assign y20778 = n48496 ;
  assign y20779 = ~n48498 ;
  assign y20780 = n48502 ;
  assign y20781 = ~n48503 ;
  assign y20782 = ~n48504 ;
  assign y20783 = ~n48506 ;
  assign y20784 = ~1'b0 ;
  assign y20785 = n48508 ;
  assign y20786 = n48509 ;
  assign y20787 = ~n48515 ;
  assign y20788 = ~1'b0 ;
  assign y20789 = n48519 ;
  assign y20790 = ~n48520 ;
  assign y20791 = n48523 ;
  assign y20792 = n48526 ;
  assign y20793 = ~n48529 ;
  assign y20794 = ~1'b0 ;
  assign y20795 = n48532 ;
  assign y20796 = n48533 ;
  assign y20797 = n48535 ;
  assign y20798 = ~1'b0 ;
  assign y20799 = ~n48536 ;
  assign y20800 = ~n48537 ;
  assign y20801 = n48542 ;
  assign y20802 = n48543 ;
  assign y20803 = ~1'b0 ;
  assign y20804 = ~1'b0 ;
  assign y20805 = ~n48545 ;
  assign y20806 = ~n48547 ;
  assign y20807 = n48548 ;
  assign y20808 = ~1'b0 ;
  assign y20809 = ~n30928 ;
  assign y20810 = ~1'b0 ;
  assign y20811 = ~n48549 ;
  assign y20812 = n48551 ;
  assign y20813 = n48553 ;
  assign y20814 = n48556 ;
  assign y20815 = n48557 ;
  assign y20816 = ~1'b0 ;
  assign y20817 = 1'b0 ;
  assign y20818 = ~1'b0 ;
  assign y20819 = ~1'b0 ;
  assign y20820 = 1'b0 ;
  assign y20821 = ~n48564 ;
  assign y20822 = ~n48567 ;
  assign y20823 = n48568 ;
  assign y20824 = n48571 ;
  assign y20825 = ~n48572 ;
  assign y20826 = ~n48578 ;
  assign y20827 = ~n48579 ;
  assign y20828 = ~n48581 ;
  assign y20829 = ~n48583 ;
  assign y20830 = n1680 ;
  assign y20831 = ~n48584 ;
  assign y20832 = n48586 ;
  assign y20833 = n48588 ;
  assign y20834 = n48589 ;
  assign y20835 = ~n48590 ;
  assign y20836 = ~n48591 ;
  assign y20837 = ~n48592 ;
  assign y20838 = ~n48595 ;
  assign y20839 = ~n48597 ;
  assign y20840 = ~n48600 ;
  assign y20841 = n48606 ;
  assign y20842 = n48607 ;
  assign y20843 = ~1'b0 ;
  assign y20844 = ~n48608 ;
  assign y20845 = ~n11472 ;
  assign y20846 = n48612 ;
  assign y20847 = ~n48613 ;
  assign y20848 = ~1'b0 ;
  assign y20849 = ~n48614 ;
  assign y20850 = n48620 ;
  assign y20851 = ~n48622 ;
  assign y20852 = ~n48625 ;
  assign y20853 = ~1'b0 ;
  assign y20854 = ~n22715 ;
  assign y20855 = ~n48626 ;
  assign y20856 = ~n48627 ;
  assign y20857 = n48628 ;
  assign y20858 = n48629 ;
  assign y20859 = ~n48631 ;
  assign y20860 = ~n48634 ;
  assign y20861 = ~n48636 ;
  assign y20862 = n48638 ;
  assign y20863 = ~1'b0 ;
  assign y20864 = ~n48642 ;
  assign y20865 = ~n15542 ;
  assign y20866 = ~n48643 ;
  assign y20867 = n48645 ;
  assign y20868 = ~1'b0 ;
  assign y20869 = ~n48649 ;
  assign y20870 = ~1'b0 ;
  assign y20871 = n48651 ;
  assign y20872 = ~n48652 ;
  assign y20873 = ~n48655 ;
  assign y20874 = ~n48658 ;
  assign y20875 = n3070 ;
  assign y20876 = ~n48659 ;
  assign y20877 = ~n48662 ;
  assign y20878 = n48667 ;
  assign y20879 = n48671 ;
  assign y20880 = ~1'b0 ;
  assign y20881 = ~1'b0 ;
  assign y20882 = ~n48673 ;
  assign y20883 = ~1'b0 ;
  assign y20884 = ~n48674 ;
  assign y20885 = n48676 ;
  assign y20886 = ~1'b0 ;
  assign y20887 = n48677 ;
  assign y20888 = ~n48679 ;
  assign y20889 = n48680 ;
  assign y20890 = ~n48682 ;
  assign y20891 = ~1'b0 ;
  assign y20892 = ~1'b0 ;
  assign y20893 = n48686 ;
  assign y20894 = ~1'b0 ;
  assign y20895 = n48688 ;
  assign y20896 = n48691 ;
  assign y20897 = n48693 ;
  assign y20898 = n48699 ;
  assign y20899 = n48700 ;
  assign y20900 = n48701 ;
  assign y20901 = ~n48704 ;
  assign y20902 = n48709 ;
  assign y20903 = ~n48716 ;
  assign y20904 = ~1'b0 ;
  assign y20905 = ~n48718 ;
  assign y20906 = ~n48719 ;
  assign y20907 = n48721 ;
  assign y20908 = n48723 ;
  assign y20909 = ~n48724 ;
  assign y20910 = ~n48727 ;
  assign y20911 = n48730 ;
  assign y20912 = ~n48731 ;
  assign y20913 = ~1'b0 ;
  assign y20914 = n48734 ;
  assign y20915 = ~n48735 ;
  assign y20916 = ~n48737 ;
  assign y20917 = ~n48739 ;
  assign y20918 = ~n48743 ;
  assign y20919 = ~n48744 ;
  assign y20920 = ~n48745 ;
  assign y20921 = n48746 ;
  assign y20922 = ~n21536 ;
  assign y20923 = n48749 ;
  assign y20924 = ~n48750 ;
  assign y20925 = n48752 ;
  assign y20926 = ~1'b0 ;
  assign y20927 = n48753 ;
  assign y20928 = ~n48757 ;
  assign y20929 = n48759 ;
  assign y20930 = ~n48763 ;
  assign y20931 = ~1'b0 ;
  assign y20932 = ~1'b0 ;
  assign y20933 = n48767 ;
  assign y20934 = n48774 ;
  assign y20935 = ~1'b0 ;
  assign y20936 = ~1'b0 ;
  assign y20937 = ~n48776 ;
  assign y20938 = n48777 ;
  assign y20939 = ~1'b0 ;
  assign y20940 = n48780 ;
  assign y20941 = n48783 ;
  assign y20942 = ~n48786 ;
  assign y20943 = ~1'b0 ;
  assign y20944 = ~n48793 ;
  assign y20945 = ~n48798 ;
  assign y20946 = n48799 ;
  assign y20947 = n48804 ;
  assign y20948 = n48809 ;
  assign y20949 = ~1'b0 ;
  assign y20950 = ~n48812 ;
  assign y20951 = ~n48814 ;
  assign y20952 = ~n48815 ;
  assign y20953 = ~n48816 ;
  assign y20954 = ~n48817 ;
  assign y20955 = n48820 ;
  assign y20956 = n48822 ;
  assign y20957 = ~n48823 ;
  assign y20958 = n48824 ;
  assign y20959 = ~1'b0 ;
  assign y20960 = ~n48826 ;
  assign y20961 = ~1'b0 ;
  assign y20962 = ~1'b0 ;
  assign y20963 = ~n48830 ;
  assign y20964 = n48832 ;
  assign y20965 = ~1'b0 ;
  assign y20966 = ~n48834 ;
  assign y20967 = n48838 ;
  assign y20968 = 1'b0 ;
  assign y20969 = 1'b0 ;
  assign y20970 = n48839 ;
  assign y20971 = n11434 ;
  assign y20972 = ~1'b0 ;
  assign y20973 = ~n48843 ;
  assign y20974 = ~n48845 ;
  assign y20975 = ~n48849 ;
  assign y20976 = n48850 ;
  assign y20977 = ~n48851 ;
  assign y20978 = ~n48852 ;
  assign y20979 = ~n48855 ;
  assign y20980 = ~n48857 ;
  assign y20981 = ~1'b0 ;
  assign y20982 = ~n48858 ;
  assign y20983 = ~1'b0 ;
  assign y20984 = ~n48859 ;
  assign y20985 = ~1'b0 ;
  assign y20986 = ~1'b0 ;
  assign y20987 = n48861 ;
  assign y20988 = n48863 ;
  assign y20989 = n48864 ;
  assign y20990 = ~n48869 ;
  assign y20991 = ~1'b0 ;
  assign y20992 = ~1'b0 ;
  assign y20993 = ~n48871 ;
  assign y20994 = n48872 ;
  assign y20995 = n48874 ;
  assign y20996 = n48877 ;
  assign y20997 = ~n48880 ;
  assign y20998 = ~n48881 ;
  assign y20999 = ~1'b0 ;
  assign y21000 = ~1'b0 ;
  assign y21001 = n48883 ;
  assign y21002 = ~n48885 ;
  assign y21003 = ~n48886 ;
  assign y21004 = ~1'b0 ;
  assign y21005 = n48887 ;
  assign y21006 = ~n48890 ;
  assign y21007 = ~n48891 ;
  assign y21008 = n48896 ;
  assign y21009 = ~n48898 ;
  assign y21010 = n48902 ;
  assign y21011 = ~n48907 ;
  assign y21012 = ~n48914 ;
  assign y21013 = ~1'b0 ;
  assign y21014 = ~1'b0 ;
  assign y21015 = ~n41786 ;
  assign y21016 = n48918 ;
  assign y21017 = ~n48919 ;
  assign y21018 = ~1'b0 ;
  assign y21019 = ~n48924 ;
  assign y21020 = ~n48927 ;
  assign y21021 = ~n48930 ;
  assign y21022 = n48931 ;
  assign y21023 = ~n10583 ;
  assign y21024 = ~1'b0 ;
  assign y21025 = ~1'b0 ;
  assign y21026 = n48937 ;
  assign y21027 = ~n48938 ;
  assign y21028 = ~n48939 ;
  assign y21029 = n48944 ;
  assign y21030 = n48945 ;
  assign y21031 = ~1'b0 ;
  assign y21032 = ~1'b0 ;
  assign y21033 = n48948 ;
  assign y21034 = ~n48950 ;
  assign y21035 = n48951 ;
  assign y21036 = ~n48953 ;
  assign y21037 = n647 ;
  assign y21038 = n48954 ;
  assign y21039 = n48955 ;
  assign y21040 = ~n48958 ;
  assign y21041 = n48961 ;
  assign y21042 = ~1'b0 ;
  assign y21043 = ~1'b0 ;
  assign y21044 = ~n48964 ;
  assign y21045 = n48966 ;
  assign y21046 = n48971 ;
  assign y21047 = n48976 ;
  assign y21048 = ~n48977 ;
  assign y21049 = n48978 ;
  assign y21050 = ~n48979 ;
  assign y21051 = n48982 ;
  assign y21052 = ~1'b0 ;
  assign y21053 = n48986 ;
  assign y21054 = n48988 ;
  assign y21055 = ~1'b0 ;
  assign y21056 = ~n48990 ;
  assign y21057 = ~n48993 ;
  assign y21058 = n48994 ;
  assign y21059 = n48995 ;
  assign y21060 = n48996 ;
  assign y21061 = ~n48997 ;
  assign y21062 = ~1'b0 ;
  assign y21063 = ~1'b0 ;
  assign y21064 = ~n48999 ;
  assign y21065 = 1'b0 ;
  assign y21066 = ~n49001 ;
  assign y21067 = ~n49002 ;
  assign y21068 = n49003 ;
  assign y21069 = ~n49004 ;
  assign y21070 = ~n49006 ;
  assign y21071 = ~n49007 ;
  assign y21072 = ~n49008 ;
  assign y21073 = n49009 ;
  assign y21074 = ~1'b0 ;
  assign y21075 = n49012 ;
  assign y21076 = ~n49014 ;
  assign y21077 = ~n49016 ;
  assign y21078 = ~1'b0 ;
  assign y21079 = ~1'b0 ;
  assign y21080 = n49019 ;
  assign y21081 = n49021 ;
  assign y21082 = ~n49022 ;
  assign y21083 = n49025 ;
  assign y21084 = n49028 ;
  assign y21085 = ~1'b0 ;
  assign y21086 = n49030 ;
  assign y21087 = ~1'b0 ;
  assign y21088 = ~1'b0 ;
  assign y21089 = n49032 ;
  assign y21090 = n49033 ;
  assign y21091 = ~n49038 ;
  assign y21092 = n49040 ;
  assign y21093 = n49041 ;
  assign y21094 = ~n49044 ;
  assign y21095 = ~1'b0 ;
  assign y21096 = ~n49045 ;
  assign y21097 = n49047 ;
  assign y21098 = n49048 ;
  assign y21099 = ~n49052 ;
  assign y21100 = ~n49057 ;
  assign y21101 = n49061 ;
  assign y21102 = ~n49063 ;
  assign y21103 = n49064 ;
  assign y21104 = ~n49065 ;
  assign y21105 = ~n49066 ;
  assign y21106 = ~1'b0 ;
  assign y21107 = n49070 ;
  assign y21108 = n9100 ;
  assign y21109 = n27496 ;
  assign y21110 = ~1'b0 ;
  assign y21111 = ~n49072 ;
  assign y21112 = ~n49074 ;
  assign y21113 = n49080 ;
  assign y21114 = ~n49081 ;
  assign y21115 = n49083 ;
  assign y21116 = ~n49089 ;
  assign y21117 = n49091 ;
  assign y21118 = n49094 ;
  assign y21119 = ~1'b0 ;
  assign y21120 = ~n49096 ;
  assign y21121 = n49098 ;
  assign y21122 = ~1'b0 ;
  assign y21123 = ~n49104 ;
  assign y21124 = ~n49105 ;
  assign y21125 = n49109 ;
  assign y21126 = ~n49113 ;
  assign y21127 = n49116 ;
  assign y21128 = ~1'b0 ;
  assign y21129 = ~n49118 ;
  assign y21130 = n49119 ;
  assign y21131 = ~n19534 ;
  assign y21132 = ~n49120 ;
  assign y21133 = ~n49121 ;
  assign y21134 = n49124 ;
  assign y21135 = ~n49125 ;
  assign y21136 = ~n1088 ;
  assign y21137 = ~n49127 ;
  assign y21138 = ~1'b0 ;
  assign y21139 = n49129 ;
  assign y21140 = n49132 ;
  assign y21141 = ~n49135 ;
  assign y21142 = ~1'b0 ;
  assign y21143 = n49138 ;
  assign y21144 = ~1'b0 ;
  assign y21145 = n49139 ;
  assign y21146 = n49142 ;
  assign y21147 = n49143 ;
  assign y21148 = ~n49144 ;
  assign y21149 = n49146 ;
  assign y21150 = ~n49147 ;
  assign y21151 = ~1'b0 ;
  assign y21152 = n49149 ;
  assign y21153 = ~n49155 ;
  assign y21154 = ~1'b0 ;
  assign y21155 = n49159 ;
  assign y21156 = n49160 ;
  assign y21157 = ~n49162 ;
  assign y21158 = n49169 ;
  assign y21159 = ~1'b0 ;
  assign y21160 = n49171 ;
  assign y21161 = ~n49172 ;
  assign y21162 = ~1'b0 ;
  assign y21163 = n49173 ;
  assign y21164 = n49176 ;
  assign y21165 = ~1'b0 ;
  assign y21166 = ~1'b0 ;
  assign y21167 = ~n49177 ;
  assign y21168 = n4822 ;
  assign y21169 = n49178 ;
  assign y21170 = ~n49179 ;
  assign y21171 = ~1'b0 ;
  assign y21172 = ~1'b0 ;
  assign y21173 = n49181 ;
  assign y21174 = ~n49182 ;
  assign y21175 = ~n49184 ;
  assign y21176 = n49186 ;
  assign y21177 = n49190 ;
  assign y21178 = n49191 ;
  assign y21179 = n49192 ;
  assign y21180 = ~n49194 ;
  assign y21181 = ~n49197 ;
  assign y21182 = ~1'b0 ;
  assign y21183 = ~n49201 ;
  assign y21184 = n49203 ;
  assign y21185 = ~n49206 ;
  assign y21186 = n49209 ;
  assign y21187 = n49211 ;
  assign y21188 = n49212 ;
  assign y21189 = ~n49213 ;
  assign y21190 = ~n49215 ;
  assign y21191 = n49222 ;
  assign y21192 = n49223 ;
  assign y21193 = ~1'b0 ;
  assign y21194 = ~n49224 ;
  assign y21195 = ~1'b0 ;
  assign y21196 = n49225 ;
  assign y21197 = n49231 ;
  assign y21198 = ~n49233 ;
  assign y21199 = ~1'b0 ;
  assign y21200 = n49234 ;
  assign y21201 = n49235 ;
  assign y21202 = ~n49241 ;
  assign y21203 = n49243 ;
  assign y21204 = ~n10851 ;
  assign y21205 = ~1'b0 ;
  assign y21206 = ~n49244 ;
  assign y21207 = ~1'b0 ;
  assign y21208 = n49246 ;
  assign y21209 = ~1'b0 ;
  assign y21210 = ~1'b0 ;
  assign y21211 = n49247 ;
  assign y21212 = n49250 ;
  assign y21213 = n49252 ;
  assign y21214 = ~n49253 ;
  assign y21215 = n49254 ;
  assign y21216 = n49258 ;
  assign y21217 = n49261 ;
  assign y21218 = ~n49263 ;
  assign y21219 = n49264 ;
  assign y21220 = ~n34953 ;
  assign y21221 = ~n49271 ;
  assign y21222 = ~n49277 ;
  assign y21223 = n49278 ;
  assign y21224 = ~n49282 ;
  assign y21225 = n49286 ;
  assign y21226 = ~n49287 ;
  assign y21227 = n49294 ;
  assign y21228 = ~n49299 ;
  assign y21229 = ~n49302 ;
  assign y21230 = ~1'b0 ;
  assign y21231 = ~1'b0 ;
  assign y21232 = n49311 ;
  assign y21233 = n49312 ;
  assign y21234 = ~n49316 ;
  assign y21235 = ~n49320 ;
  assign y21236 = ~n9470 ;
  assign y21237 = ~n49323 ;
  assign y21238 = ~1'b0 ;
  assign y21239 = ~n49325 ;
  assign y21240 = ~1'b0 ;
  assign y21241 = ~n49330 ;
  assign y21242 = ~n49334 ;
  assign y21243 = 1'b0 ;
  assign y21244 = n49336 ;
  assign y21245 = n49343 ;
  assign y21246 = n49346 ;
  assign y21247 = ~n49347 ;
  assign y21248 = ~n49349 ;
  assign y21249 = n49351 ;
  assign y21250 = ~n49355 ;
  assign y21251 = n49357 ;
  assign y21252 = ~n49359 ;
  assign y21253 = ~1'b0 ;
  assign y21254 = ~n49361 ;
  assign y21255 = n49363 ;
  assign y21256 = ~n49364 ;
  assign y21257 = n49365 ;
  assign y21258 = n49367 ;
  assign y21259 = n49369 ;
  assign y21260 = n49375 ;
  assign y21261 = ~1'b0 ;
  assign y21262 = n49376 ;
  assign y21263 = n49377 ;
  assign y21264 = ~n49379 ;
  assign y21265 = n49382 ;
  assign y21266 = n49383 ;
  assign y21267 = n49384 ;
  assign y21268 = n49385 ;
  assign y21269 = ~n49386 ;
  assign y21270 = ~1'b0 ;
  assign y21271 = n49391 ;
  assign y21272 = ~n49397 ;
  assign y21273 = ~n49398 ;
  assign y21274 = n24748 ;
  assign y21275 = ~n49400 ;
  assign y21276 = ~1'b0 ;
  assign y21277 = ~n49405 ;
  assign y21278 = n49413 ;
  assign y21279 = ~n49416 ;
  assign y21280 = ~n49417 ;
  assign y21281 = n49418 ;
  assign y21282 = ~1'b0 ;
  assign y21283 = ~1'b0 ;
  assign y21284 = ~n49422 ;
  assign y21285 = ~1'b0 ;
  assign y21286 = ~n49427 ;
  assign y21287 = ~n49429 ;
  assign y21288 = ~n49431 ;
  assign y21289 = ~n49432 ;
  assign y21290 = n49433 ;
  assign y21291 = ~1'b0 ;
  assign y21292 = n49435 ;
  assign y21293 = n49438 ;
  assign y21294 = ~n49440 ;
  assign y21295 = ~n49442 ;
  assign y21296 = ~n49444 ;
  assign y21297 = ~n49446 ;
  assign y21298 = ~1'b0 ;
  assign y21299 = n49448 ;
  assign y21300 = ~n49453 ;
  assign y21301 = n49456 ;
  assign y21302 = ~n49457 ;
  assign y21303 = n49462 ;
  assign y21304 = n49465 ;
  assign y21305 = n49467 ;
  assign y21306 = n49469 ;
  assign y21307 = ~n49471 ;
  assign y21308 = n49473 ;
  assign y21309 = ~n49476 ;
  assign y21310 = ~n49480 ;
  assign y21311 = n49481 ;
  assign y21312 = n49482 ;
  assign y21313 = ~n49483 ;
  assign y21314 = ~n49487 ;
  assign y21315 = ~1'b0 ;
  assign y21316 = ~n49488 ;
  assign y21317 = ~n31956 ;
  assign y21318 = ~n49492 ;
  assign y21319 = ~n49493 ;
  assign y21320 = ~1'b0 ;
  assign y21321 = n49495 ;
  assign y21322 = ~n49497 ;
  assign y21323 = ~n49500 ;
  assign y21324 = ~n49501 ;
  assign y21325 = ~1'b0 ;
  assign y21326 = ~n49503 ;
  assign y21327 = n49504 ;
  assign y21328 = n49507 ;
  assign y21329 = ~1'b0 ;
  assign y21330 = ~1'b0 ;
  assign y21331 = ~1'b0 ;
  assign y21332 = ~n49510 ;
  assign y21333 = n49513 ;
  assign y21334 = ~n49514 ;
  assign y21335 = ~n49515 ;
  assign y21336 = ~n49520 ;
  assign y21337 = ~n49522 ;
  assign y21338 = n49523 ;
  assign y21339 = n49529 ;
endmodule
